ELF              ��4   he      4    (           � �B  B           B  ���  �        �W  �2  �                 �    UU���r#  VW�����_^�y  �    �i���f�f�f�f�f����=��t$�    ��tU���h���Ѓ��Í�&    f�Í�&    ��&    ����-�����������t(�    ��tU���Ph���҃��Í�&    �t& �Í�&    ��&    ��=�� ugU�����V��S���������9�s�v ����������9�r��'����    ��t��hx��Q~��������e�[^]�Í�&    ��&    ��    ��t'U���h��hx��~������	�����&    f���������t$�"  ��Ã��t$�"  ��Ã��t$�o&  ��Ã��t$�_&  ��Ã��t$�O&  ��Ã��t$�?&  ���UWVS���t$(�|$,�T$4�\$0�T$�F�D$�G�D$�~ ��   �G)Ѕ���   �T$�$    �[���F9�~4�O��)�9�~)�$Ћl$�l� ������v��L$���D$�,��$�$9F~*�D$�G+D$;$~�F��~܋O��)څ�~Ѻ    롃�[^_]�UWVS��8�l$L�|$P�D$T�D$�L$X�L$ �t$\�L$`�L$�\$d�\$$�T$h�T$(j�P!  ���     �@    �@    ��9�
�D$�9�}R�L$9��D$�9���   t$9�|�D$�9���   �t$�T$�9�|�D$�9��  �؃�,[^_]Ã�j��   �     �@    �h�x��)���P�L$$�H��C�C   �����j�����j�   �     �@    �h�x�L$ �H�T$)����P���; t�S��S�P�C�C�|$�-�������)�D$��j�*   �     �@    �p�x�T$ +T$(�P�L$$�H���; t�S��S�P�C�C�D$�D$���������j��  �     �@    �h�p�L$ �H)��T$$)�P���; t�S��S�P�C�C�������S��(�\$0�St�T$�Kx�L$�D$    �D$    �C|�D$���   �D$�Cu	�=`� u#��j �D$P�D$(P�sphL�j�,  ��H[�hL�j j j ��PjQR��  �� hL�j j j ���   ��Pj�sx�C|Ct��P�  �� hL�j j j j�C|��P�sx�st�  �� hL�j j j j�C|��P���   Cx��P�st�]  �� 9(��6  hL�h�   h�   h�   j�s|�Cx��P�Ct��P�"  �� ��hL�h�   h�   h�   �Cx��P�Ct��P�CP��  �Ct�Sx�H�L$8�J�L$<�� hL�j2j2jdjj��RC|��P�  �� hL�j2j2jdjj�Cx��P�C|Ct��P�  �� hL�j2j2jdjj�Cx��P�C|Ct��P�k  �� hL�j2j2jdjj�Cx��P�C|Ct��P�C  �K|Kt�A�Kx�Q�� RPh �hL���  ��������hL�h```�h   �j�s|�Cx��P�Ct��P�  �� �����S��j j j h��h��j��)  ��������+��i��  ��+��Ѓ� =�  v,����̉��%����������    ��������[�ÍL$����q�U��WVSQ���   j j j hL��E�Pj�N)  ���T��X���P�V  �`������n  �8�   �<�   �D�����j�  �     �@    �@    �����j j j j hI�j��(  ��j j j �E�PhV�j�(  ��   ��   ��j hb��'  ���$   �  ����jj S�B'  �ǉ$�  �ƃ�WPS��&  ��h �Vjjj j ��  ��S�l'  ��j hm��-'  �Ã�jj P��&  �ǉ$�4  �ƃ�WPS�w&  ���   ���   �$  0 �  �������u%ǅ@���    ǅ8���    ǅD���    �  ����h��Vh   h   j j �:  �� �ǅ<���    fǅl���  fǅn���  fǅp���  fǅr���  ��j j j ��l���P��<���j�J'  ��@����ǃ� ����   �uܻ    � �    �	��D����B;ppt/��9���   ��9�@���vօ�tً�D����    ���9�u���9�@���vQ���+	  ��D����    ���9�u��Bƀ�   ��D����    ���9�u��B��l����   ����   �    ƀ�   �    �ك�h�   �  �Í�l����   �����l����Ct��n����Cx��p����C|��r������   ƃ�   �(��$   �;  �     �@    �X����D��� t=��8�����H��@����`���8�����<�����<���9�T�����  �7�����D������,���@���������  �d��h���<����  �5    �   ��D����  ��D����H��4������t�H��t�J�P��t���t�
��u���D�����@�����@���9�t��P�"  ����8�����H��8����ድ8�����j�  ��8����     �@    ��4����H����D��� ��   ��p��@�����@���9���   ����   ��D����    � ��9�u��@�(��`��Wx�h��J9���   �G��  �5d��Ot��<���O|�Y�9�}�Z9���9�|�J9�E+�<����5�)У ��$���  ��8�����D����E����    �o�����D����a���ǅt���   �Gp��|�����P��x���j��p�����l����wl�#  �� �m  ǅt���   �G�  �d�+Ot����)��
  �������  ��9���������������D����    �6��9�u��v�Ft9�~�F|9�}��Fx9�<���~���   9�<���}�����@���������9��������������D���� ���(  �    ��9�@��������9��~�������  ���ۡ    ���    t���5    �\����    ���i  �    ;(��_  �(�    �    �K  ��D������t�Q��t�P�A��t���t���u���D�����9�t��Q�Q  ���    ��  �A��8����߉�@�����X�����S��!  ������   ��`���� u�(���t׋�d�������t �у�tǅt���   ������x����ǅt���   ������x����Pp��|�����R��x�����t�����p�����l����pl�c!  �� �^����5h��5d�hL�h0��5���hL�j j j jjj j �H  ��,j
��l���S�5����!  ��hL�h�   h�   h�   j j S��  ��j j j hL��u�j�!  �� ���������j ��P���Pjh-��u�j��   �� ��P��� t>�-��Q�d��P���    H£d��A�؋h��B���    H£h��=$� t3�(��d��h�+��    HӉQt+ ��    HAx�`���j j j j ��T���Pj�6   �� ��T��� ������,��-��t���S�������   �=$� t�$� hL�h�   h�   j@�X���P�5T�j j �  �� �    ��@�����@��� �u  �y�����D����@���ǅt���   �d�+Ot)�����ȉ�x����Wp��|�����RP��t�����p�����l����wl�&  �� �=,� �Q����-�� �C����,� �$� ǅt���   �(�����������|�����x�����t�����p�����l����pl�  �� �������D����H��4��������(�    ��   ����D����s�F��������V��D����@��D������    ��   ��tȋ�D����    ���9�u����r� �������D����    ���9�u��Bƀ�    ��9�������9��R�����t���D����    ���9�u��B���    u���D����    ���9�u��(�9B�������R�����D�������(����    ��9��8���9��0�������Q������ߋ�D����Bƀ�   �����f�f�f�f��UWVS��
  ��>  ���D$(�|$$�ƃ�)����ŋD$ ��	��t>��QW�t$,�  ����u	��[^_]Ð���/VR�D$,�P�  ����[^_]Ð��QW�t$,�R  ������&    ��    UWVS�P
  ��w=  ���t$ �|$$�T$(��   t*�B���t�v ���>�����u��[^_]Í�&    �t& ������R��WV�  ����tӉ>��t̉~��tĉ~��[^_]Í�&    �t& ���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���|$$�L$,�D$4�\$8�t$(�T$0�|$�L$��y��D$    �L$��y�1����ȁ�   ���	���% �  ���͉���	�k	ǅ�~u;s}p�D2��L$�D$�D$�D��$��&    �D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�  �ù;  ���t$j j j j Vj �  ��$��[^� f��`  �;  UWVS��,�|$@�t$D�D$�L$L�D$P�\$T�T$X�l$\��y|$H1���y�1�����������	�	E�T$�D$��~\;u}W�D$H��D$�D��D$�
f���9u~9�]������)�;\$OT$H��R��t$�L$ ��P�\$�X�����;t$u���,[^_]Í�&    �  �:  UWVS��,�t$@�l$D�D$�L$L�D$P�|$T��yt$H1���y�1��؉������� �  ��	�	G�T$�D$��~i;o}d�D$H��D$�D��D$��t& ���9o~C�G�_������)����;\$OT$H��R�t$�L$ ���P�\$�~�����;l$u���,[^_]Í�&    ��    UWVS�  ���9  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$�������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�@  ��g8  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�,����� 9t$h�_�����L[^_]Í�&    UWVS�p  �×6  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�\����� 9t$l�_�����L[^_]Í�&    UWVS�  ���4  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�)�����9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$Ë$�f��UWVS�������3  ���D$<�|$8�t$0�D$�G�D$�D$D���Ơ��D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������ ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ�P����� ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�N����� 9|$�b�����[^_]Í�&    f�UWVS�����÷0  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��U��E�]�Mfof ��������]�U��E�]�M�o� ��������]�U��E�]�M��~4fn�fop�f��fs�f��fs�f��fs�f��f ������]Ð������                U��01�WVS�k����Ò/  ��(���  �����9��  C��  P���  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p��x�1����  �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � �����p  ��t   �g�����&    �t& �����.  ǀ|      ��x�ǀx      �    �B    ��p�ǀ�     �    �B    ��h�ǀ�      �    �B    ǀp      ǀt      ǀh      ǀl      ǀ`      ǀd      Í�&    �UWVS�0�����W-  ���|$0� ��&    ���p  �   ��t   �  �w �  ��t܋�|  �t$�|$0����  �|$0��x  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s��x  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ���|  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$������p��B1ҋD$~Q��@�����   ��   �E��  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,��p��E$���~��h�Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ�������������|  ���K�����
  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~��h��N,��p��ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��D
  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS�P�����w)  ���D$ ����   �P���)փ� C��	  �N�A=����~   �y��p�1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o��x  ����   ��t�J+J�ʋO)�9�|W�R	  ��[^_]Í�&    �v ��h  ��l   ����� ���� t
f=��t<�u���`  ��d   뱍�&    ���x  롍�&    ���p  ��t   ��[^_]Í�&    �v �G9�|  tU9�ta���t�B�G��t���x��G1�)Q���wW��  ���4�����&    �t& �o�������&    ���|  룍�&    �ǃx      듍t& WVS�t$�������'  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS�������&  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��  �G�P�������   �P9���   �T$��  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ�h  ��l   %��� =�� tDf����t=���t8�C  1���[��^_]Í�&    �p���&  ����[^_]Í�&    �t& ���`  ��d   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ�����f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f�S�C�����j#  �� j j j �D$ P�t$8j��  �D$,��8[�f�S������:#  ��j j j j �t$(j�  ��([Í�&    f�S�������
#  �� j �D$P�t$8�t$8�t$8j�g  �D$,��8[Í�&    ��&    S�������"  �� j �D$P�t$8�t$8�t$8j�'  �D$,��8[Í�&    ��&    S�c����Ê"  �� j �D$P�t$8�t$8�t$8j��  �D$,��8[Í�&    ��&    S�#�����J"  �� j �D$P�t$4�t$<�t$8j�  �D$,��8[Í�&    ��&    S�������
"  ���t$�t$�t$�������[Í�&    �t& S�������!  ���t$�t$�t$�������[Í�&    �t& S�����ê!  ���t$�t$�t$� �����[Í�&    �t& S�S�����z!  ���t$�t$�������[Í�&    ��&    �S�#�����J!  ���t$�������1�[ÐS������*!  ��j �t$�������   ��u
����[Ív ��P������1҃���[�f�f�f�f�f��S�������   �� j j j �D$ P�t$8j�;   �D$,��8[�f�S�����ê   ��j �t$0�t$0�t$0�t$(j�   ��([�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��WVS�D$�L$���ƍT�N��������~&1���&    �t& �:����Z�����9�|�[^_Ív W1�VS�D$��������  �|$�t$��t@�������	~%��W�T���u��� QW�l�������[^_Ív ��0�T���u��ٍv �0   f���[^_�f�1�Í�&    ��    �P���{  �����  1�Í�&    �v S�3�����Z  �� j j j �D$ P�t$8j�����D$,��8[�f�1��f�f�f�f�f�f�������t6U��S������&    �v �Ѓ�����u��[]Í�&    ��&    ��
����  /taskbar.lef /dev/mouse0 /close.bmp /bg1.bmp          zR |�        m���    CD H     8   a���    CD H     T   U���    CD H     p   I���    CD H     �   =���    CD H     �   1���    CD H  8   �   %����    A�A�A�A�C(�A�A�A�A�h      ����
   A�A�A�A�CLvP^@[
A�A�A�A�ACLBPx@JLBPn@oLBPm@kLBPm@   p  l  P���r   A�C0E8B<E@EDCHELBPHA�A0�E4B8B<B@DDBHALAPH0E4B8B<B@JDBHCLJPH0E4B8B<B@BDGHCLCPH0E4B8B<B@BDGHMLCPH0Q4E8E<E@BDCHGLGPH0C4E8E<E@EDGHGLDP\0E4B8B<B@BDBHDLGPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPW0A4A8E<E@H0H4E8E<E@BDCHGLGPH0 4   �  N���z    A�CBB B$E(E,B0lvA�        ����       ,   ,  }����   D Gu Fupu|uxut�   \  8����    A�A�A�A�N c$A(A,D0H G
A�A�A�A�BC$D(A,G0H C
A�A�A�A�BC$A(A,D0H    \   �  D����    A�A�A�A�N n
A�A�A�A�LC$F(D,A0H YA�A�A�A�   @  t���?    Cy 8   X  �����    A�A�A�A�C$�A�A�A�A�8   �  P���.    A�A�NFB B$B(A,B0HC�A� H   �  D����    K�A�A�A�C@�DAHFLHPL@IA�A�A�A� H     �����    K�A�A�A�C@�DAHDLJPL@IA�A�A�A� <   h  \���b   A�A�A�A�NPL@�A�A�A�A�X   �  �����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X      ����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   `  t����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   �  �����    A�A�A�A�C(�A�A�A�A�   �  ����          �  ����           t���W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   $  ����s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�  D   |  �����   A�F�A�A�N<Z@J0�
A�A�A�A�M      �  �����       T   �  l����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `   0	  �����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   �	  @����    A�A�A�WA H��A�A�  �   �	  �����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0<   \
  ���   A�A�A�A�C �
C�A�A�A�A 8   �
  �����    A�A�A�A��
�A�A�A�P   0   �
  \���.    A�N(B,B0B4E8D<B@LA�  0     X���'    A�NBB B$B(D,B0HA�  0   @  T���2    A�N(B,E0D4D8D<B@LA�  0   t  `���2    A�N(B,E0D4D8D<B@LA�  0   �  l���2    A�N(B,E0D4D8D<B@LA�  0   �  x���2    A�N(B,E0D4D8D<B@LA�  (     ����%    A�NDDD HA�   (   <  ����%    A�NDDD HA�   (   h  ����%    A�NDDD HA�   $   �  ����!    A�NDD HA�      �  ����    A�ND HC� 8   �  ����E    A�NBD HL
C�DCA HEC�0     ����.    A�N(B,B0B4E8D<B@LA�  0   P  ����-    A�NBD D$D(D,B0HA�  (   �  ����!    A�A�A�[�A�A�,   �  ����M    A�A�A�G�A�A�   D   �  ����n    A�C�A�tEA HC
�A�A�D[�A�A�    (  ����          <  ����       0   P  ����.    A�N(B,B0B4E8D<B@LA�     �  ����           ����    ����                                                                      @  �                          �             �   �            �����   �           ���������   �          �������������   �         �����������������   �        ���������������������   �       �������������������������   �      �����������������������������   �     ���������������������������������   �    �������������������������������������   �   ���������������������   �   �   �   �   �   ���������   ���������   �����      �����   �    ���������   �      �   �     ���������   �����      ����   ���������   �          ���������   �       ����   �   �����                 1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                                                                                                                                                                                                                                                                                            <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              ��                           >        ���    src/gfx/sse2.asm NASM 2.14.02 ��     %  . @   l    '   �       src/gfx/sse2.asm      �!0==?LL==0/!$!0==?LL==0/!#!0==>=0K�KYKYKYMK>1/""u�                                               t�          ��          A�          I�          x�          �          �           �          @�     	     ��     
                                                                                                                             ��   �         �      (   x�      ;   ��      =    �      P   P�      f   ��    
 u   ��    
 �   Ё      �   ��    
             ���   �      �   �      �    �      �            ��  ��                  ��           ��#           ��,           ��5           ��F  �       W  �       r  \�       �  e�       �  p�     5           ���  ���    �  ��    	 �  ��    	 �  ��    
 �  ��    
 �  ��    
 �  ��    
 �  ��    
            ��           ��           ��#           ��-           ��4           ��             ��@   �      V  x�    
 b  `�.     t  ���    �  d�    	 �  h�    
 �  ��!     �  бM     �  ��    
 �  ��     �  ��     �  ��    
   @�.     P  ��    
   �     $  �2     /  ��    
 ;  ���    g   ��     n  p�    
 v  ��    	 �  p�-     �  �     �  �    
 �  ��.     �  e��     �  ���    �  ��     �  0�    
   @�    	    �n       ��    
 -  p�%     3  L�    
 ;  %�     B  $�    
 �  t�      G  ��     U  ��    	 _  (�    
 f  ���     �  P��     �   �      �  ��    
 �  -�    
 �  @�%     �  ��     �   �    
 �  P�2     �   �W      $�     ;  ��    
 <  ��&     *  �%     P  ��   	 c  ��.     r  5�     z  @��    �  `��     �  ��     �  ,�    
 �  @�b    �  ���       `�s     %  ��    
 7  ��     
 C  p��     i  �    p  %��    u  a�    	 }  ��    	 �  0�?     �  ��    
 �  E�     �  A�      �  ��z     �  �     �  �     �  �E     �  ��     	 �  ��     
 �  `�    	 �  .�
      ��2     $  8�r    =  P��     �  ��!     a  �'     m  ��    	 v   �      �  U�     �  Я2     �  �      g  а     �   ��     �  ���     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp graphics.cpp text.cpp font.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset_sse2.loop memset_sse2.ret bigzero allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns memory.c filesystem.c ipc.c syscall.c itoa.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos l_max_inuse syscall reverse frameCounter liballoc_init liballoc_unlock lastUptimeMilliseconds ReceiveMessage _Znwm lemon_read bgClipRects _Z12DrawGradientiiii10RGBAColourS_P7Surface memcpy l_inuse __TMC_END__ SendMessage __DTOR_END__ dragOffset lemon_open _Z12surfacecpy_tP7SurfaceS0_8Vector2i malloc __x86.get_pc_thunk.ax mouseSurface __dso_handle itoa currentUptimeMilliseconds lseek surface _ZdlPv drag liballoc_lock keymap_us active _Z18memset32_optimizedPvjm calloc memcpy_sse2_unaligned frameRate mouseData _Z16memcpy_optimizedPvS_m closeButtonSurface lemon_write _Z8DrawCharciihhhP7Surface _Z30RecalculateBackgroundClipRectsP4ListIP8Window_sE currentUptimeSeconds mouseSurfaceBuffer liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main testKey font_default _Z5floord bgSurface _ZdaPv _fini _Z15UpdateFrameRatev liballoc_free _Znam access _edata _end redrawWindowDecorations _Z14SplitRectangle4RectS_ lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close font_old memset_sse2 _ZdaPvm lemon_readdir memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                    t�t                     !         ���   �2                 '         A�A3                    -      2   I�I3  -                 5         x�x3  �                 ?         �B                    F         �B                    M          � B                   V         @�@B  h                  \         ���Q  �                  a      0       �Q  +                 j              �Q                     y              �Q                    �              R  B                  �              GR                    �              bR  p                  �              �R                    �              �R                                  �R  �	     ?         	              �\  �                               �d  �                  