ELF          >     @     @        D
         @ 8  @                   @       @     4�     4�                  8�     8�B     8�B     (      �                   8�     8�B     8�B                           �C  �� �             H��    UH���������  �7� H��   �i���f.�     �` C H=` C t�    H��t	�` C ��f��ff.�     @ �` C H��` C H��H��H��?H�H��t�    H��t�` C ���ff.�     @ �=��  uwUH��� H��ATA�`�B S�h�B H��`�B H��H��H9�s%f.�     H��H�}� A��H�r� H9�r��0����    H��t
�`�B �����[A\�B� ]��ff.�     @ �    H��tU�� C �`�B H������]����D  ����UH��H��   H�E�A�    A�    �    �    H�ƿ   �!  �E��� �E�    �pC �M  9E�������   �E� �E�    ��� 9E�}kH��`���H���  �E�Hc�H��`���A�    A�    �    H�ƿ   �G!  H�E�H�E�E��ƿpC ��  H� H9E�����t�E���E���E�����t�E��ƿpC ��  ��� �E��=������UH��H��   H�E�A�    A�    �    �    H�ƿ   �   �E܉�� �E�    ��� 9E���  �E� H��`���H����  �E�Hc�H��`���A�    A�    �    H�ƿ   �Z   H�E�H�E��E�    �pC ��  9E�����t)�E�ƿpC ��  H� H9E�����t�E���E����E�������   ��   �RC  H�E�H�E�H��`���H��h���H�PH�HH��p���H��x���H�PH�H H�U�H�M�H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�U؉��   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�E�H�ƿpC �F  ��� �E��c������UH��AVAUATSH��   H�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸� C A�    A�    H�ƿ   �  �Y  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H���c  H��P���H�E��@����H��X���H�    ����H!�H	�H��X���H��X�����H�       H	�H��X���H��P���H��X���H��H��H�й� C ��H��H���?  �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H���  H��`���H��h���H�    ����H!�H��H��h���H�E��@������H�� H��h�����H	�H��h���H��`���H��h���H��H��H�й� C ��H��H���  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H����  H��p���H�E��@������H��x���H�    ����H!�H	�H��x���H��x�����H�       H	�H��x���H��p���H��x���H��H��H�й� C ��H��H���  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H���  H�E�H�U�H�    ����H!�H��H�E�H�E��@������H�� H�U���H	�H�E�H�E�H�U�H��H��H�й� C ��H��H���  A�    A�*�2   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H���O  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A�� C D���H��H����  H�E����   ����H�E����   ����H�E�H��H��h� C A��   A��   ��   H���9  H���E�   �E�   H�E�H���   H�E�H��H���{
  H�E�H�E�H�U�H��� C A�    A�    H���   �P  H�e�[A\A]A^]�UH��H���   �� C ��  H��� H��� H��H��H��� H���� �H��� f�HH���2  H��H�E�H�E�H�H�HH�k� H�l� H�PH�HH�e� H�f� H�@ H�c� �M� �C� ��H�H����<  H�;� H�E؋PH�E؋@�u�h�   A�    A��   �щ¾    �    ��  H��A�    A�    �    �    �    �   �3  �`�A �b�A �]�  H�E�H�Eк   �    H����  H�H�E�H�Eк    �    H�����  H�E�H�H���<<  H�E�H�u�H�U�H�E�H�Ѻ   H���z�  H�Eȋ@��H��H��H�H��H��H�E�H�H�E����    ���    ��  ��;  H�� �m� �c� H�M�A�@C I�ȉщ¾    �    ��  �l�A A�    A�    �    �    H�ƿ   �!  �    �w�A ��  �E��E��   �C ���@  ��� ��� A�� C D��� �щ¾    �    ��  ��� ��t,�\� �R� A�� C D��� �щ¾    �    ��  �E�    ��� 9E�}%�E��ƿpC �1  H�E�H�E�H���`����E����4�  �E��   �C ���  �� ��� ���Љ�� ��� ��� ���)Љ�� ��� ����   ��� ��� ��� H�#� )щʉ��   ��� ��� H�� )щʉ��   H��� ���   ��yH��� ǀ�       H��� ���   ��yH��� ǀ�       �1� �������#  �� �����  �� �pC ��  ���E��}� ��  �E��ƿpC ��  H�E���� H�E����   9���  ��� H�E����   H�E��@���9���  ��� H�E����   9��  ��� H�E����   H�E��@���9��Z  �E��ƿpC �v  H�ƿpC �  H�E�H��� �U� H�E����   �P�>� 9�|LH�E��@����u>�"� H�E����   )� H�E����   )��ȉ�� ��� ��� ��   H�E�   H�E��@����t0��� H�E����   )ЉE��� H�E����   )ЉE��4��� H�E����   )Ѓ��E��� H�E����   )Ѓ��E��E�H�� H�E�H	�H�E�H�E�H�@|H�E�H�E�H�@tH���u��u��u���x�����p���H���  H��0�	�m�������� ����t��� ��t���  ��� ����  ��� ��������  ���  ���  H�'� H����  ��� H�� ���   9���  ��� H��� ���   H��� �@���9��h  �n� H��� ���   9��M  �S� H��� ���   H��� �@���9��"  �+� H��� ���   �P�� 9�|H�j� �@������   H�U� H����   H�E�   H�=� �@����t6��� H�&� ���   )ЉE��� H�� ���   )ЉE��:��� H��� ���   )Ѓ��E�v� H��� ���   )Ѓ��E�E�H�� H�E�H	�H�E�H��� H�@|H�E�H��� H�@tH���u��u��u���x�����p���H���  H��0H��@���H���Q  H�������  H��P���H=�  ��   H=� u�H�1� H����   H��X���H����   H��X���H��H��t0H��X�����H��t!H�E�   H��X������� �B H�H�E��H�E�   H��X����� �B H�H�E�H��� H�@|H�E�H��� H�@tH���u��u��u���x�����p���H���  H��0�(H��X���H��u�=����H��X���H��u�1�����������������5�� ��� h� C j A�    A��   �   �   ���r  H���E�    �}��E�    �}��E���E���&� �$� ������H�A� H�E�H�@H��H����  �5T� �J� A�� C D�F� �   �   ���  ����UH��H���}��u��}�u'�}���  u�pC �   � �B �pC ��@ �3  ���UH����  �   ����]�UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]ÐUH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H��H�}��u�U�H�E���H���   ��UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H���^0  H�E��ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �?  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H��H�}�H�E��@��tH�E��    H���2�������H��H��H�D$    H�t$A�    A�    �    �   �!  H�D$H���H��H��H�T$A�    A�    �    �   ��  �D$H���H��Hc�A�    A�    �    �    �   ��  H���H��H��Hc�A�    L�D$H��H�¿   �  �D$H���H��H��Hc�A�    L�D$H��H�¿   �h  �D$H���H��H��Hc�Hc�A�    L�D$H�¿   �:  H�D$H���H��H��Hc�A�    L�D$�!   �  �D$H���H��t�    �4�H��H9�u��ATUSH��H��@��tH��t�    H�,�H��H9�u�[]A\�I��A��H���>	  M��t�J��H�+H��H9�u���AUATUSH��H��H��H��H	�t�@  H��[]A\A]�I��A��L)�I��H���P  M��t�L�L�A��s<A��u"E��t��E �A��t�E��B�D%�fB�D#�릋E �E��B�D%�B�D#��H�E H�D��H�T�H�T�H�KH���H)�H)�D������a�������    ��H�t H�4��9�r��B���SH���(   �-  �@    �     �T$�P�T$�P�T$�P�T$�PH�X[��,�f���*�f/�����)��US�D$L�T$ ��x?��xDE��A����A	�E��A��E	�A��   �M�J��~\A;r}V��l�D�\����    ��    �9�t3��A9Z~*A�B������~�9�~���E��A9�tԃ�A9B���[]�SD����AQ����PA��E���J���H��[�H��A��I��H��H�� H��H�� �������H���AWAVAUATUSH��A��A��A��A��L��A�@
J�, �R���B>��I���f���*������D��    A�~�A��E����   D;{��   D��G�T7�G�L,��   �����A��L�{G�7D�ZF�| D�XL�sG�<D�ZF�\ ����L�sE�A9�t6���C��9�~)A��F�\ A��u�D�rB�|5 u�D�rB�|5 u���D)�D9�t��9s~E��~�CA9�}��D���H��[]A\A]A^A_�AWAVAUATUSH��HA��A��A��D�L$L��$�   D��D����A�����E  E���I  E���$  A;|$�  ���    f���A*��|$��f���*��l$�L$��f���*���f���*��\$ �\��^��D$(������f���*�E��f���A*��d$0�\��^��D$8f���*͋D$��f���*��T$�\��^D$�Y��X��D,��D$(�Y��XD$ �D,�AT�YL$@�XL$8�,���PE��E��D���   D����������H��A9�t��A9\$�m���H��H[]A\A]A^A_�A��    ����E�A�    ����AWAVAUATUSH��HA��A��A��D�L$L��$�   D��D����A�����D  ���J  E���$  A;t$�  ��    f���A*��|$��f���*��l$�L$��f���*���f���*��\$ �\��^��D$(������f���*�E��f���A*��d$0�\��^��D$8f���*͋D$��f���*��T$�\��^D$�Y��X��D,��D$(�Y��XD$ �D,�AT�YL$@�XL$8�,���PE��E���   D����D���
�����H��A9�t��A9\$�m���H��H[]A\A]A^A_�A�A�    ����A��    ����H��A��H��H�� H��H�� APA�Љ���E���H���AVAUATUSA��H�� �~ ~nA�֋G)Ѕ�~bH��I���    �uA�D$B�.��D)�9�N���Hc�����Hc�HuB�<3��D���Hc�I|$�������9]~A�D$D)�9��[]A\A]A^�ATUSA��H�� L�VH�_�~ ��   I�ӉՋG)Ѕ�~vA�    �T���F9�~2�WA��E)�A9�~$A���H�A��=����v�A���D�Hc҉���A��D9N~(A���G)�D9�~�F��~�W��D)���~չ    �[]A\�H��H��H�T$A�    A�    �    �   �  H�D$H���H��H��A�    L�D$0H�L$(H�T$ �   �  H���H��H���   HD���%  H���H��H���   HD��%  H���H���$  H���H�������H���H���$  H���H���t$  H���UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo% #@ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo% #@ f��fs�f��f H����H��]Ð�����������                AWAVAUATUSH��A��L�t$P�L$D�L$��H��@�B L�,A��H��   H�D$A���D$�L��t6@��y�A�)�AV�D$PD�L$D�D$�   �   D���6���H����I��A��L;l$tA�m �   �H��[]A\A]A^A_�AWAVAUATUSH��H���T$L�|$P�?@��t?��A��E��E��A��@��H��AWE��E�ƋT$������H���;��H��@��u�H��[]A\A]A^A_�UH��SH�}�H�u�H�U�H�M�L�E�L�M�H�E�L�E�H�M�H�U�H�u�H�}�L���i�[]�UH��H���}��E�H�A�    A�    �    �    H�ƿ   �������UH��H��H�}�H�u�H�E�%�  H��tH�	� �   H�5�� H�=�� �z  H�E�H�U�H���  H��H��A�    A�    �    H�¿   ����H�E�H� H��u�������    ��UH��H�}�H�u�    ]�UH��H��H�}�H�E�A�    A�    �    �    H�ƿ    �������UH��H�=:� ����UH��H��H�E�A�    A�    �    �    H�ƿ   �w���H�E��E��E���UH��H��0�}�H�u�H�U�H�U�H�E�A�    A�    �    H�ƿ   �2���H�E�H��H�E�H�H�E�Hi�@B H��H�E�H��    ��UH��H�}��u��    ]�UH��H�}��    ]�UH��    ]�UH��]�UH��H���   H��X���H��P�����L���H��@���H��`���H�»C H��H���  H��`���H�5U� H���  H��H��@���H��H���  H�5>� H���  H��H��P���H��H���y  H�5"� H���j  H��L�����H���  H�5� H���H  H�5�� H���9  H��H��X���H��H���$  H�5�� H���  H���_  H��`���H����  ���UH��H���   H��X���H��P�����L���H��@���H��`���H�ºC H��H���:  H��`���H�5I� H���Z  H��H��@���H��H���E  H�52� H���6  H��H��P���H��H���!  H�5� H���  H��L�����H���)  H�5�� H����  H�5�� H����  H��H��X���H��H����  H�5�� H���  H���  H��`���H���  ���UH��H�}�H�u�H�E�]ÐUH��H��H�}�H�E��     H�E��@    H�E�H��H����   H�E��@ H�E��@ H�E��@ H�E��@ H�E��@ ���UH��H��H�}�H�u�H�E��H�E��H�E��PH�E��PH�E�H��H�U�H��H��H���   H�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��P��ÐUH��H��H�}�H�E�H��H���(   ��ÐUH��H��H�}�H�E�H����  H�E��@ ��ÐUH��H��H�}�H�E�H����  ��ÐUH��H��H�}�H�u�H�E�H���  H�E��PH�E��PH�E��@��tH�E�H�ƿ   �U���H��H�E�� ����UH��H��H�}�H�u�H�U�H�E�H��H���]  H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���[  H�E��ÐUH��H��H�}��u�H�U�H�E�H��H���w  H�E���UH��H��H�}�H�E�H� H�U�H��H��H���  H�E���UH��H��H�}�H�u�H�U�H�E�H��H���  H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���  H�E��ÐUH��H��H�}��u�H�U�H�E�H��H���  H�E���UH��H��H�}�H�E�H� H�U�H��H��H���  H�E���UH��H�}��]ÐUH��H�}��]ÐUH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H������H�E�H� H�U�H�M�H��H���Z  H�E�H���T������UH��H��0H�}�H�u�H�E�H���E���H�E؋ H�U�H�M�H�Ή��A  H�E�H���������UH��H��H�}�H�u�H�E�H�U�H��H���u� ���UH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H������H�E�H� H�U�H�M�H��H����   H�E�H���r������UH��H��0H�}�H�u�H�E�H���c���H�E؋ H�U�H�M�H�Ή���   H�E�H���/������UH��H��H�}�H�u�H�E�H�U�H��H���s� ���UH��H�� H�}�H�u�H�U�H�U�H�E�H��H����   ���UH��H��@�}�H�u�H�U�H�U�H�E�H��H���"���H�U�H�M��E�H�Ή��T  H�E�H���������UH��H�� H�}�H�u�H�U�H�U�H�E�H��H���  ���UH��H��@�}�H�u�H�U�H�U�H�E�H��H������H�U�H�M��E�H�Ή��N  H�E�H���!������UH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=�� �@ѿ�H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H����  �TH�E�� ��t%H�E�� ��tH��    H��uH�=�� �Eп��u�H�E�A�    A�   �    �
   H���q  ��ÐUH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=� ��Ͽ�H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���   �TH�E�� ��t%H�E�� ��tH��    H��uH�=|� ��ο��u�H�E�A�    A�   �    �
   H���X   ���UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���\   H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��� H�E��E�    �E���~H��    H��uH�=�� �Ϳ��M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�� �DͿ��E��P�U�H��D�-H�U�H�E�H��H���Z  � 9E�����tE�E�    H�U�H�E�H��H���4  � �U�)�9E�����t�U�H�E���H���8  �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���  �E��ڋE����E�}� x!�E�H��D���H�E���H����  �m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�E� H�E��E�    �E���~H��    H��uH�=\� �̿��M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=B� �˿��E��P�U�H��D�-H�U�H�E�H��H���   � 9E�����tE�E�    H�U�H�E�H��H���   � �U�)�9E�����t�U�H�E���H���M  �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���  �E��ڋE����E�}� x!�E�H��D���H�E���H����   �m��ِ��UH��H�}�H�u�H�E��H�E�� 9�}H�E��H�E�]ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=O� �bʿ�H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ��ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=�� �ɿ�H�E�H���   H��u)H�E�H� H�U�H��H��H�������H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ���UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�sH�U�H�E�HЋU�H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�H;E�s"H�U�H�E�H�H�M�H�U�H�� �H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H;E�s4H�E�    H�E�H;E�sgH�U�H�E�H�H�M�H�U�H�� �H�E���H�E�    H�E�H;E�s3H�E�H+E�H�P�H�E�H�H�E�H+E�H�P�H�E�H���H�E���H�E�]�UH��H�}�H�E�    H�E�    H�U�H�E�H�� ��tH�E�H�E���H�E�]�UH��H��H�}�H�E��    H���|   fH~�H�E��E���UH��H��H�}�H�E��
   �    H����   ��UH��H��H�}�H�E��
   �    H���   ��UH��H��H�}�H�E��
   �    H����  ��UH��H�� H�}�H�u�H�U�H�E�H��H����  fH~�H�E��E���UH��H��H�}�H�u�H�U�H�E�H��H���  ��UH��H�� H�}�H�u�H�U�H�E�H��H���-  �}�H�E��U�H�E��U��m���UH��H��0H�}�H�u��U�H�E�� ��t"H�E�� �����La  ������uH�E��ԐH�E�� <+uH��� �:   H�5�� H�=�� �����E� H�E�� <-u	�E�H�E��}�
t@�}� tH��� �B   H�5�� H�=�� �T����U�H�M�H�E�H��H���   �   H�E�    H�E�� ��tGH�E�� </~<H�E�� <91H�U�H��H��H�H�H��H�E�� ����0H�H�H�E�H�E��H�}� tH�E�H�U�H��}� t	H�E�H���H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H��`H�}�H�u��U�H�E�����H�E�H�E��E�    H�E�H�PH�U�� ���E�E���_  ������t�փ}�-u�E�   H�E�H�PH�U�� ���E���}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��E�Hc�H�������    H��H�E؋E�Hc�H�������    H��H�ЉE�H�E�    �E�    �E����\  ������t�m�0�4�E���S\  ��������   �E���_  ��t�7   ��W   )E�E�;E�}r�}� xH�E�H9E�rH�E�H9E�u�E�;E�~	�E������*�E�   �E�Hc�H�E�H��H�EȋE�Hc�H�E�H�H�E�H�E�H�PH�U�� ���E��<�������}� y
H�E�������}� tH�E�H��H�E�H�}� t�}� t
H�E�H���H�E�H�U�H�H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H���C H����  %���]�UH��H��H�}�H�� ��   H�5� H�=S� �����UH��H���}��E���H���C H����  ���UH��H��   ��\���H��`���H�ºC H��H������H��`���H�5� H���.���H���x���H��`���H���������UH��H�� H�}�H�u�H�U�H�M�H�E�H��H����
  �E��}� tH���C �U���    �H�E���UH��H�� H�}�H�u�H�E�H�E�H���!	  H�E�H�}� u�    �!H�E�H�E�H��H�E��    H������H�E���UH��H��� ��   H�5ڽ H�=� ����UH��H��H�}�H�E��    �    H���c����    ��UH��H��H�}�H��� ��   H�5�� H�=�� �C���UH��H���}��,����E����<���UH��H���}��E����'���UH��H���}�H�I� ��   H�5-� H�=h� �����UH��H��H�}�H�)� ��   H�5� H�==� ����UH��H��H�}�H�� ��   H�5׼ H�=� ����UH��H��`H�}�H�u�H�U�H�M�L�E�H�E�    H�E�H�E�H�E�H;E�s|H�E�H+E�H��H�E�H�U�H�E�H�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���ЉE܃}� yH�U�H�E�H�H�E�뛃}� ~H�U�H�E�H�H��H�E��H�E��.H�E�H;E�tH�8� ��   H�5�� H�=f� �����    ��UH��H��`H�}�H�u�H�U�H�M�H�E�    H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�E�H��H�E�H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���Ѕ�����ufH�E�H�E�H�E�H�E�H�E�    H�E�H;E�sEH�U�H�E�H�� �E�H�U�H�E�H�H�M�H�U�H�� �H�U�H�E�H��EǈH�E�벐H�E��M���H�E��������UH��H���}�H��� �  H�5�� H�=�� �w���UH��H��H�}�H��� �  H�5�� H�=ʺ �L���UH��H��H�}�H��� �  H�5d� H�=�� �!���UH��}�u�E��}�E��E��}�ЉE�H�E�]�UH��H��H�}�H�u�H�b� �'  H�5� H�=J� �����UH��H��H�}�H�u�H�8� �+  H�5� H�=� ����UH��SH��HH�}�H�u��M� H�E�H�E�H�E�H�U�H�E�H�H�E�H�E�H�E�H�E�H��H�E�H�}� uOdH�%    H������f�   dH�%    H������f�@  dH�%    H�������@    H�E��@	���bH�E�H� H��H�dH�%    H������H��H�U�H�u�H�E�H���ӉE�}� tH�I� �;  H�5� H�=\� ����H�E�H+E�H��H[]�UH��H���   H��X���H��P���H��H���H��`���H�ºC H��H�������H��`���H�5/� H������H���O���H��`���H�������H��X���H��uH��� �@  H�5K� H�=� ����H��P���H��uH��� �A  H�5 � H�=� �����H��H���H��uH�Y� �B  H�5�� H�=�� ����H��P���� ��uH�,� �C  H�5ȷ H�=�� ����H��P����H��X����҉�   ��UH��H��H�}��u�H��� �H  H�5}� H�=�� �:���UH��H��pH�}�H�u�H�U��� H�E�f�E�  f�E�  �E�    H�E�    H�E�    H�E�H�E�H�E�H�E�H�E�H��    H�E�H�H�E�H�}� uNH�E�H� H�� H� H�M�H�U�H�u�H�}��ЉE�}� tH�;� �U  H�5Ƕ H�=8� ����H�E��H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� tH��� �Z  H�5y� H�=� �6���H�E�H+E�H��H�E�H�E�H;E�sH�E�H��    H�E�H��     H�E���UH��H�� H�}�H�u�H�U�H��� �e  H�5� H�=H� �����UH��H��P  H������H�=�� �zf  H��������   H������H�ºC H��H���
���H������H�5�� H���*���H��H������H��H���  H���_���H������H�������H��������H��tIH��`���H�ºC H��H������H�EH��H��`���H��H���5  H������H��`���H�������	� H��H������H��H���  ���UH��H��   H��X����ڒ H��H��X���H��H���  H�E�H�=�� �`e  H������tXH��`���H�ºC H��H�������H��`���H�5�� H������H��H�E�H��H���z  H���L���H��`���H�������H�E���UH��H��   H��X���H��P����/� H��H��P���H��X���H��H���  H�E�H�=�� �d  H������t|H��`���H�ºC H��H���B���H��`���H�5� H���b���H��H��X���H��H����  H�5� H���>���H��H�E�H��H���  H���v���H��`���H���	���H�E���UH��SH��8H�}�H�u�H�U�H�E�H��w
�  �   H�E�H�P�H�E�H!�H��t�  �~�.� H��H�U�H�E�H��H���P  H� H��H����  H�E�H�}� u�  �CH�E�H�P�H�E�H!�H��tH�y� ��  H�5� H�=.� ����H�E�H�U�H��    H��8[]�UH��H�� H�}�H�u�H�U�H�?� ��  H�5�� H�=ֲ �X���UH��H���}��u��}�u�}���  uH���C H���   ���UH����  �   ����]ÐUH��H��H�}�H�E��q  H���   ���UH��H�}��u�H�E��U�H�E�ǀ�	     H�E����	  =o  wH�E����	  �P�H�E�Hcҋ�H�E����	  �P�H�E�Hcҋ���1�i�e�lH�E����	  ��H�E����	  �H�E�Hc҉�H�E����	  �PH�E����	  �x����]ÐUH��H�}��E�    �E�߰�H�E؋��	  =o  �N  �E�    �}��   kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE�E����  H�E�Hcҋ��U���1E�����D����1�H�E؋U�Hc҉��E���E��   �}�n  kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE��E������H�E�Hcҋ��U���1E������D����1�H�E؋U�Hc҉��E��H�E؋��	  %   ���H�E؋ %���	ЉE�H�E؋�0  �U���1E�����D��1�H�E؉��	  H�E�ǀ�	      H�E؋��	  �HH�U؉��	  H�U�H����E�E���1E�E���%�V,�1E�E���%  ��1E�E���1E�E�]ÐUH��H�� H�}�H�u��U�H�U�H�E�H��H�������H�E��U��H�E���UH��H�}�H�E�H�     H�E�H�@    H�E�H�@    H�E�H�@    H�E�H�@     H�E��@(    �]�UH��H�}�H�E�H��?]�UH��H��H�}�H�U��   �������tH�l� �   H�5�� H�=�� �������UH��H�}�H�E��    ��]�UH��H��PH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH� � �   H�5į H�=� ����f���E�H�E��.   H����} H�E�H�E�H���p���H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� �����J  �������  �M��Q� �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   �� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�5�� H�=î �����H�E�H;E�sbH�E�H�E�� �����-I  ������uBH�E�� ����0�*��^E��M��X��E��M��\� �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E��~-� fW��E��E���UH��H��@H�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH��� �   H�5w� H�=�� ����f���E�H�EȾ.   H���{ H�E�H�E�H���#���H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� �����G  �������  �M��� �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   ��� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�5M� H�=v� ����H�E�H;E�sbH�E�H�E�� ������F  ������uBH�E�� ����0�*��^E��M��X��E��M��'� �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E�� � W��E��E���UH��H��pH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH��� �   H�5+� H�=T� �h������}�H�E��.   H���My H�E�H�E�H�������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sNH�E�� �����mE  ��������   �m��-�� ���}�H�E�� ����0�E��E��m����}�H�E��H�}� ��   �-�� �}�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�5� H�=>� �R���H�E�H;E�sVH�E�H�E�� �����D  ������u6H�E�� ����0�E��E��m����m����}��m��-� ���}�말����H�}� tH�E�H�U�H��}� t�m����}��m���UH��H��H�}�H�u�H�U�H�E�H��H���0  H�E���UH��}�H�E�   �E�H9E�vH���B �U�H���U�E�   �E�H+E�H��H�E�E�H+E�H�P�E��H�H!�H�E�H�E�H��H�E؋E�Hc�H�E�H�H�E؉�H��H��]�UH��H��@H�}�H�E�   H�E������_���H9E�����tG�E�    �E�H�U�H��H9�s#�E����3���H9E�����t�E��   �E���H�E�H���   H�E�H������H��?   H)�H��H�E�H�E�H�E�H�E�H��H�E�H�E�   ��H��H�E�H)�H��H�E�   ��H��H��H�H�P�H�E���H��H��H�E�H�U�H�E�H�H�E�H�H���ÐUH��H��H�}�H�u�H�E�H� H�U�H��H����   ��ÐUH��H��H�}�H�u�H�E�H� H�U�H��H���
  ��UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���  ��UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]�UH��H��0H�}�H�u�H�E�H������H�E�H� H�U�H�M�H��H���J
  H�E�H���S������UH��SH��xH�}�H�u�H�}� �D  H�E�H�E�H�E�H�PH�E�H��H���}
  H�U�H�E�H��H����
  H�E�H�}� uH��    H��uH�=ަ �I���H�E�� ����   H�E�H�@H9E�tH��    H��uH�=� ����H�E�H�PH�E�H��H���  H�E�H�P H�E�H�@H   H��H)�H�E�H�P H�E�H���  H�E�H� H�U�H�RH��   H�U�H�RH�� ���H��H��H���y� �    �   H�E�� ��tH��    H��uH�=ͦ �h���H�E�H���6  H�E�H�E�H�E�H%  ��H��H�E�H9�tH��    H��uH�=� �$���H�E؋@HH�H��H��H��H�E�H�H��H�E�H�E؋@H�������H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=� 貦��H�U�H�E�H��H���  H�E�H�@PH�����E�H�E؋@L��uH��    H��uH�=.� �i���H�E�H�ƿ   �����H��H���w
  H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H���e
  ����t�   ��    ��tH��    H��uH�=� �����H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H���F
  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���X	  H�E�H���  �   H�E�H���  ����H��x[]�UH��SH��   H��x���H��p���H��p��� uHǅp���   H��p��� �  ��  H��p���H���Y����E�}�~H��    H��uH�=w� �⤿��E�H�H��H��H��H��x���H�H��H�E�H�U�H�E�H��H���  H�E�H�@H���*  H�E�H�@H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=N� �a���H�E�H�U�H��H���  ����tH��    H��uH�=j� �-���H�E�H� H��t$H�E�H�U�H�H��H���K  ����t�   ��    ��tH��    H��uH�=w� �ڣ��H�E�H�H�E�H�PPH�E؋@L�PH�E؉PLH�E�H�@PH���$  H�E�H�PH�E�H��H���	  H�E�H��H���	  H��H�E�H�P��  H�E�H���@  �U�H��x�����H����	  H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=D� ����H�E�H�U�H��H���L  ����tH��    H��uH�=`� �뢿�H�E�H� H��t$H�E�H�U�H�H��H���	  ����t�   ��    ��tH��    H��uH�=m� 蘢��H�E�H�H�E�H�PPH�EЋ@L�PH�EЉPLH��x���H�PH�E�H��H���Z  H��x���H�PH�E�H��H���
  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H����  H�E�H����
  H�E�H�@PH��uH��    H��uH�=7� �ڡ��H�E�H�PH�E�H��H���M  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���  H�E�H���S  H�]�H�E�H���  �   H��p���H�  H% ���H�E�H�U�H��x���H��H���M
  H�E�H��x���H�PH�E�H��H���  H��x���H�PH�E�H��H����  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H���  H�E�H�@H��H�E�H����  H��H�Ĉ   []�UH��SH��hH�}�H�u�H�U�H�}� uH�U�H�E�H��H���!���H����  H�}� uH�U�H�E�H��H�������    �  H�E�H�E�H�E�H�PH�E�H��H���&  H�U�H�E�H��H���m  H�E�H�E�H����  H�}� uH��    H��uH�=�� �柿�H�E�� ����   H�E�H�E�H�E؋@H������H�E�H�E�H;E�w	H�]��  H�U�H�E�H��H���C���H�E�H�}� u
�    ��   H�U�H�M�H�E�H��H���z���H�U�H�E�H��H������H�]��   H�E�� ��tH��    H��uH�=O� �*���H�E�H�@H9E�tH��    H��uH�=�� ����H�E�H�@H9E�sH�]��WH�U�H�E�H��H������H�E�H�}� u�    �2H�E�H�PH�M�H�E�H��H������H�U�H�E�H��H�������H�]�H�E�H���   H��H��h[]�UH��H��`H�}�H�u�H�U�H�E�H�5E� H���>���H�E�H�������H�E�H�M�   H��H���:���H�E�H�U�H�M�H��H����  H�E�H������H�E�H���������UH��H��H�}�H�u�H�E�H�U�H�H�E��@ H�E�H���  ���UH��H��H�}�H�E��@��tH�E�H���  ��ÐUH��H�� H�}�H�u�H�E�H��H����  H�E�H�}� ��   H�E�H�@H9E�sH�E�H����  H�E���H�E�H�PH�E�H�@H�H9E�rH�E�H���  H�E��H�E�H�@H9E�rH�E�H�PH�E�H�@H�H9E�rH��    H��uH�=ܢ ��H�E���    ��UH��H��0H�}�H�u�H�E�H���)  H�E�H�E�H���7  H�E�H�}� uH�U�H�M�H�E�H��H���4  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���g	  H�E�H�E�H���  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���I	  ���UH��H��H�}�H�E��@����tH��    H��uH�=n� ���H�E�H� H�������H�E��@ ��ÐUH��H�}�H�E�H�     �]�UH��H�}�H�u�H�E�H�E�H�E�H�@H9E�r H�E�H�PH�E�H�@H�H9E�s�   ��    ]ÐUH��H�� H�}�H�u�H�E�H���  H������tH�E�H�U�H��H����
  �   H�E�H����
  H�E�H�E�H�HH�U�H�E�H��H���5  ��tAH�E�H���M  H������tH�E�H�U�H�M�H��H���J  �VH�E�H���  H�E��H�E�H���a  H������tH�E�H�U�H�M�H��H���_  �H�E�H���2  H�E��\�����UH��H��0H�}�H�u�H�E�H���
  H�E�H�E�H����  H�E�H�}� uH�U�H�M�H�E�H��H���0  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���c  H�E�H�E�H���F
  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���E  ���UH��H�� H�}�H�E�H���Z	  H�E�H�}� u�    �,H�E�H����	  H������tH�E�H����	  H�E���H�E���UH��SH��XH�}��u�H�E�H� �   H����t H�E�H�E�H�� H%  ��H�EЋE��������H�E�H�E�    H�}�   w
H�E�HE���H�}��� vH��    H��uH�=�� �䘿�H�E�H�ƿ�   �d���H�ø   H+E�H�M�H�U�H�4�U���H��H���  H�]�H�E�    H�E�    H�E�H�@H9E�sHH�E�H�PH�E�H�H�ƿ   �����H��H������H�]�H�E�H�U�H�H�E�H�E�H�E�HE��H�E�H�U�H�PPH�E�H��X[]�UH��H�� H�}�H�u�H�E�H���`  H������tH�E�H�U�H��H���]  �   H�E�H���2  H�E�H�E�H�HH�U�H�E�H��H����  ��tAH�E�H���  H������tH�E�H�U�H�M�H��H���f  �VH�E�H����  H�E��H�E�H����  H������tH�E�H�U�H�M�H��H���]  �H�E�H����  H�E��\�����UH��H��H�}�H�E��@��tH��    H��uH�=)� ����H�E�H� H������H�E��@���UH��SH��(H�}�H�u�H�E�%�  H��tH��    H��uH�=&� 豖��H�E�H� H�U�H��   H��H���$r H�E�H�E�H�ƿH   ����H��H�E�H��   H�E�H���   H���  H�]�H�E�H��([]�UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���  �UH�E�� ��t%H�E�� ��tH��    H��uH�=� �ؕ��H�u�H�E�A�    A�   �    �
   H���C  ��ÐUH��H�}�H�E�H� ]�UH��H��H�}�H�E�H���m  H�@��UH��H��H�}�H�E�H���O  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���-  H�E�H�}� tH�]�H�E�H����  H�X H�}� tH�]�H�E�H����  H�XH�E�H����  �@(������t8H�E�H����  ��tH�E�H���  �@(   �H�U�H�E�H��H����  H�E�H�������H��uH�E�H������H9E�t*H�E�H�������H9E�uH�E�H�������H��t�   ��    ��tH��    H��uH�=� �4���H�E�H���9  H�E�H�}� uH�E�H�U�H��rH�E�H���g���H9E�����tH�]�H�E�H����  H�X�EH�E�H���X���H9E�����tH��    H��uH�=7� 貓��H�]�H�E�H���  H�XH�}� tH�]�H�E�H���o  H�H�E�H���`  H�@    H�E�H���L  H�@    H�E�H���8  H�     H�E�H���%  H�@    H�E�H���  H�@     H�}� tH�U�H�E�H��H���5  �H��H[]�UH��H��H�}�H�E�H����  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H��� ���H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���H  H�X�EH�E�H�������H9E�����tH��    H��uH�=� �)���H�]�H�E�H���  H�XH�]�H�E�H����  H�H�E�H����  �X(H�E�H����  �X(H�]�H�E�H���  H�XH�}� tH�]�H�E�H���  H�H�]�H�E�H���  H�XH�}� tH�]�H�E�H���s  H�H�E�H���}���H������tH�]�H�E�H���c���H���B  H�X H�E�H���K���H��H�E�H���#  H�XH�E�H���)  H��H�E�H���  H�X H�E�H���
  H������tH�]�H�E�H����  H����  H�XH�E�H����  H�@    H�E�H���  H�@    H�E�H���  H�     H�E�H���  H�@    H�E�H���s  H�@     H�U�H�E�H��H����  H�U�H�E�H��H���  �H��H[]ÐUH��H�}�H�E�H� ]ÐUH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=Q� ����H�E�H�U�H�H�U�H�E�H��H���  H�U�H�E�H��H���  ���UH��H�}�H�u�H�U�H�E�H�PH�E�H�@H9���]�UH��H��H�}�H�E�H���  H�@��UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=� �Z���H�E�H������H������tH��    H��uH�=� �*���H�]�H�E�H���&  H�XH�]�H�E�H���  H�H�E�H���T  H�E�H�}� tH�]�H�E�H����  H�X H�]�H�E�H����  H�XH�]�H�E�H����  H�X H�]�H�E�H���  H�XH�U�H�E�H��H���  H�U�H�E�H��H���  H�U�H�E�H��H���  �H��8[]�UH��H��H�}�H�E�H���O  H�@�ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=A� ����H�E�H������H������tH��    H��uH�=a� �ԍ��H�]�H�E�H����  H�XH�]�H�E�H���  H�H�E�H���  H�E�H�]�H�E�H���  H�X H�]�H�E�H���  H�XH�]�H�E�H���q  H�X H�}� tH�]�H�E�H���V  H�XH�U�H�E�H��H����  H�U�H�E�H��H���B  H�U�H�E�H��H����  �H��8[]ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���=  H�E�H�}� tH�]�H�E�H����  H�X H�}� tH�]�H�E�H���  H�XH�E�H���  �@(������t8H�E�H����  ��tH�E�H���p  �@(   �H�U�H�E�H��H���  H�E�H������H��uH�E�H�������H9E�t*H�E�H���i���H9E�uH�E�H������H��t�   ��    ��tH��    H��uH�=�� �؋��H�E�H���I  H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���  H�X�EH�E�H��� ���H9E�����tH��    H��uH�=۔ �V���H�]�H�E�H���R  H�XH�}� tH�]�H�E�H���7  H�H�E�H���(  H�@    H�E�H���  H�@    H�E�H���   H�     H�E�H����  H�@    H�E�H����  H�@     H�}� tH�U�H�E�H��H����  �H��H[]�UH��H��H�}�H�E�H���  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H�������H�E�H�}� uH�E�H�U�H��rH�E�H���o���H9E�����tH�]�H�E�H���  H�X�EH�E�H������H9E�����tH��    H��uH�=�� �͉��H�]�H�E�H����  H�XH�]�H�E�H���  H�H�E�H���  �X(H�E�H���  �X(H�]�H�E�H���  H�XH�}� tH�]�H�E�H���i  H�H�]�H�E�H���V  H�XH�}� tH�]�H�E�H���;  H�H�E�H���}���H������tH�]�H�E�H���c���H���
  H�X H�E�H���K���H��H�E�H����  H�XH�E�H���9  H��H�E�H����  H�X H�E�H���  H������tH�]�H�E�H���   H���  H�XH�E�H���  H�@    H�E�H���v  H�@    H�E�H���b  H�     H�E�H���O  H�@    H�E�H���;  H�@     H�U�H�E�H��H���
  H�U�H�E�H��H���#  �H��H[]ÐUH��H�� H�}�H�u�H�U�M�H�E�H�M�H�U�   H���  H�E��U�PHH�E��@L    H�E�H�@P    H�E�H��XH����������UH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=�� �^���H�E�H�U�H�H�U�H�E�H��H���	  H�U�H�E�H��H����  ���UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=�� ���H�E�H���I���H������tH��    H��uH�=�� ���H�]�H�E�H���  H�XH�]�H�E�H���  H�H�E�H������H�E�H�}� tH�]�H�E�H���\  H�X H�]�H�E�H���H  H�XH�]�H�E�H���4  H�X H�]�H�E�H���   H�XH�U�H�E�H��H���  H�U�H�E�H��H���<  H�U�H�E�H��H���  �H��8[]ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=�� 躅��H�E�H���/���H������tH��    H��uH�=� 芅��H�]�H�E�H���b  H�XH�]�H�E�H���N  H�H�E�H���U  H�E�H�]�H�E�H���+  H�X H�]�H�E�H���  H�XH�]�H�E�H���  H�X H�}� tH�]�H�E�H����   H�XH�U�H�E�H��H���_  H�U�H�E�H��H���  H�U�H�E�H��H���]  �H��8[]ÐUH��H�� H�}��u�H�U�H�M�H�E��U�H�E�H�U�H�PH�E�H�U�H�PH�E�H��H���������UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�}��   H�E�H�]�UH��H��H�}�H�E�H�������H�@ ��UH��H��H�}�H�}� u�    �H�E�H�������@(�����ÐUH��SH��XH�}�H�u�H�E�H���}����@(������tH��    H��uH�=S� �n���H�E�H���s  H�E�H�}� �\  H�E�H������H9E�������   H�E�H������H������tH��    H��uH�=U� ����H�E�H���}���H��������@(��������   H�E�H���X���H�E�H�E�H���H���H��H�E�H��H���  H�E�H������H9E�����tH��    H��uH�=)� 脂��H�E�H���`����@(   H�E�H���M����@(   H�E�H�������H�E��  H�E�H������H9E�����tH��    H��uH�=� ����H�E�H���o���H������tH��    H��uH�=M� �聿�H�E�H���?���H�������@(������tzH�E�H������H�E�H�U�H�E�H��H���  H�E�H������H9E�����tH��    H��uH�=0� �s���H�E�H���O����@(   H�E�H���<����@(   H�E�H������H�E�H�E�H������H����  ��tH�E�H������H���  ��t�   ��    ��toH�E�H��������@(������t+H�E�H��������@(   H�U�H�E�H��H��������  H�E�H�������@(   H�E�H�������@(   �  H�E�H���j����@(�E�H�E�H�������H9E������  H�E�H������H���i�����tH�E�H������H����  ��t�   ��    ��tQH�E�H���x���H�E�H�U�H�E�H��H���h  H�E�H��������@(   H�E�H��������@(   H�E�H�E�H�E�H���E���H�����������tH��    H��uH�=�� ���H�U�H�E�H��H���R  H�E�H���d����@(   �]�H�E�H���N����X(H�E�H�������H���7����@(   �M  H�E�H������H9E�����tH��    H��uH�=�� ���H�E�H������H��������tH�E�H���Q���H���~  ��t�   ��    ��tQH�E�H���G���H�E�H�U�H�E�H��H���y  H�E�H�������@(   H�E�H���x����@(   H�E�H�E�H�E�H�������H����������tH��    H��uH�=)� �L~��H�U�H�E�H��H���  H�E�H�������@(   �]�H�E�H��������X(H�E�H���k���H��������@(   ��H��X[]�UH��H��H�}�H�E�H������H� ��UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H���  ����uH�E�H������H�E��Ԑ���UH��H��H�}�H�u�H�E�H���x  ��ÐUH��H��H�}�H�u�H�E�H���g  ��ÐUH��H�� H�}�H�u�H�E�H���	  H�E�H�}� uH�E�H���#  �@(   �  H�E�H���  �@(   H�E�H����  �@(��������  H�E�H���L	  H�E�H�}� tH�E�H����  �@(��t�   ��    ��tH��    H��uH�=�� �|��H�E�H�������H9E�uH�E�H������H����  ��t�   ��    ��tYH�E�H���L  �@(   H�E�H���9  �@(   H�E�H������H���  �@(   H�U�H�E�H��H��������  H�E�H������H9E�uH�E�H���%���H���U  ��t�   ��    ��tYH�E�H���  �@(   H�E�H���  �@(   H�E�H�������H���  �@(   H�U�H�E�H��H�������j  H�E�H������H9E�������   H�E�H�������H9E�����t;H�U�H�E�H��H���C  H�U�H�E�H��H����  H�E�H���  �@(   �&H�U�H�E�H��H���  H�E�H����   �@(   H�E�H����   �@(   �   H�E�H���N���H9E�����tH��    H��uH�=1� �z��H�E�H�������H9E�����t;H�U�H�E�H��H���"  H�U�H�E�H��H���o  H�E�H���G   �@(   �&H�U�H�E�H��H���G  H�E�H���   �@(   H�E�H���   �@(   ����UH��H�}��X   H�E�H�]�UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H����  ����uH�E�H���  H�E��Ԑ���UH��H��H�}�H�E�H������H�@ ��UH��H��H�}�H�}� u�    �H�E�H���^����@(�����ÐUH��SH��XH�}�H�u�H�E�H���5����@(������tH��    H��uH�=� �y��H�E�H���s  H�E�H�}� �\  H�E�H���+���H9E�������   H�E�H���e���H������tH��    H��uH�=� �x��H�E�H���5���H�������@(��������   H�E�H������H�E�H�E�H��� ���H��H�E�H��H���q  H�E�H������H9E�����tH��    H��uH�=�� �x��H�E�H�������@(   H�E�H�������@(   H�E�H������H�E��  H�E�H���v���H9E�����tH��    H��uH�=�� �w��H�E�H�������H������tH��    H��uH�=� �|w��H�E�H�������H���t����@(������tzH�E�H������H�E�H�U�H�E�H��H���   H�E�H�������H9E�����tH��    H��uH�=Ą �w��H�E�H�������@(   H�E�H��������@(   H�E�H���%���H�E�H�E�H������H���%  ��tH�E�H���R���H���  ��t�   ��    ��toH�E�H�������@(������t+H�E�H���x����@(   H�U�H�E�H��H��������  H�E�H���M����@(   H�E�H���:����@(   �  H�E�H���"����@(�E�H�E�H���T���H9E������  H�E�H���9���H���i�����tH�E�H���v���H���1  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���Z  H�E�H�������@(   H�E�H�������@(   H�E�H�E�H�E�H�������H�����������tH��    H��uH�=L� �/u��H�U�H�E�H��H���D
  H�E�H�������@(   �]�H�E�H�������X(H�E�H������H��������@(   �M  H�E�H���p���H9E�����tH��    H��uH�=#� �t��H�E�H���?���H��������tH�E�H�������H����  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���k	  H�E�H���C����@(   H�E�H���0����@(   H�E�H�E�H�E�H���Y���H����������tH��    H��uH�=�� ��s��H�U�H�E�H��H���
  H�E�H��������@(   �]�H�E�H�������X(H�E�H�������H�������@(   ��H��X[]�UH��H��H�}�H�E�H���w���H� ��UH��H�� H�}�H�u�H�E�H���[���H�E�H�}� uH�E�H�������@(   �  H�E�H�������@(   H�E�H��������@(��������  H�E�H�������H�E�H�}� tH�E�H�������@(��t�   ��    ��tH��    H��uH�=ׁ �r��H�E�H�������H9E�uH�E�H������H��������t�   ��    ��tYH�E�H���D����@(   H�E�H���1����@(   H�E�H������H�������@(   H�U�H�E�H��H��������  H�E�H������H9E�uH�E�H���T���H��������t�   ��    ��tYH�E�H�������@(   H�E�H�������@(   H�E�H������H�������@(   H�U�H�E�H��H�������j  H�E�H�������H9E�������   H�E�H�������H9E�����t;H�U�H�E�H��H���  H�U�H�E�H��H���  H�E�H��� ����@(   �&H�U�H�E�H��H���f  H�E�H��������@(   H�E�H��������@(   �   H�E�H���F���H9E�����tH��    H��uH�=M� �p��H�E�H�������H9E�����t;H�U�H�E�H��H����  H�U�H�E�H��H���-  H�E�H���?����@(   �&H�U�H�E�H��H���  H�E�H�������@(   H�E�H�������@(   ����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�&l H�E��E�    �E���~H��    H��uH�=� �o���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=� �Fo���E��P�U�H��D�-H�U�H�E�H��H���\���� 9E�����tE�E�    H�U�H�E�H��H���6���� �U�)�9E�����t�U�H�E���H�������E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H��跤���E��ڋE����E�}� x!�E�H��D���H�E���H��臤���m��ِ��UH��H��H�}�H�}� u�   �H�E�H���*����@(�����ÐUH��SH��8H�}�H�u�H�E�H���*���H�E�H�}� tH�E�H������H9E�t�   ��    ��tH��    H��uH�=~ ��m��H�E�H���)���H�E�H�E�H�������H�E�H�}� tH�]�H�E�H������H�H�]�H�E�H���p���H�XH�]�H�E�H���\���H�H�]�H�E�H���I���H�XH�]�H�E�H���5���H�H�}� uH�E�H�U�H��rH�E�H������H9E�����tH�]�H�E�H�������H�X�EH�E�H���~���H9E�����tH��    H��uH�=�} ��l��H�]�H�E�H������H�XH�U�H�E�H��H���'���H�U�H�E�H��H�������H��8[]�UH��SH��8H�}�H�u�H�E�H������H�E�H�}� tH�E�H�������H9E�t�   ��    ��tH��    H��uH�=�} �2l��H�E�H������H�E�H�E�H���'���H�E�H�}� tH�]�H�E�H�������H�H�]�H�E�H�������H�XH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H������H�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���W���H�X�EH�E�H�������H9E�����tH��    H��uH�=} �8k��H�]�H�E�H������H�XH�U�H�E�H��H������H�U�H�E�H��H���t����H��8[]�UH��H�}��    ]�UH��H�}��    ]�UH��SH��8H�}�H�u�H�E�H���8���H�E�H�}� tH�E�H���I���H9E�t�   ��    ��tH��    H��uH�=!{ �tj��H�E�H������H�E�H�E�H�������H�E�H�}� tH�]�H�E�H���I���H�H�]�H�E�H���6���H�XH�]�H�E�H���"���H�H�]�H�E�H������H�XH�]�H�E�H�������H�H�}� uH�E�H�U�H��rH�E�H������H9E�����tH�]�H�E�H������H�X�EH�E�H���D���H9E�����tH��    H��uH�=�z �zi��H�]�H�E�H���v���H�XH�U�H�E�H��H�������H�U�H�E�H��H��������H��8[]�UH��SH��8H�}�H�u�H�E�H������H�E�H�}� tH�E�H���T���H9E�t�   ��    ��tH��    H��uH�=Az ��h��H�E�H���m���H�E�H�E�H���5���H�E�H�}� tH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H������H�H�]�H�E�H���o���H�XH�]�H�E�H���[���H�H�}� uH�E�H�U�H��rH�E�H���|���H9E�����tH�]�H�E�H������H�X�EH�E�H������H9E�����tH��    H��uH�=�y ��g��H�]�H�E�H�������H�XH�U�H�E�H��H���I���H�U�H�E�H��H���6����H��8[]�UH��H��H�}�H�}� u�   �H�E�H���~����@(������UH��H�� �}��F H�E��E���H�U�H�E���H����  �E�}� t�    ��[ H�E���H���O ����UH��H�� �}��@F H�E��E���H�U�H�E���H���  �E�}� t�    ���Z H�E���H���&P ����UH��H�� �}���E H�E��E���H�U�H�E���H���5  �E�}� t�    ��jZ H�E���H���P ����UH��H�� �}��E H�E��E���H�U�H�E���H����  �E�}� t�    ��Z H�E���H���Q ����UH��H�� �}��>E H�E��E���H�U�H�E���H���  �E�}� t�    ��Y H�E���H���Q ����UH��H�� �}���D H�E��E���H�U�H�E���H���3  �E�}� t�    ��hY H�E���H���TS ����UH��H�� �}��D H�E��E���H�U�H�E���H����
  �E�}� t�    ��Y H�E���H���S ����UH��H�� �}��<D H�E��E���H�U�H�E���H���
  �E�}� t�    ��X H�E���H���0T ����UH��H�� �}���C H�E��E���H�U�H�E���H���1
  �E�}� t�    ��fX H�E���H���T ����UH��H�� �}��C H�E��E���H�U�H�E���H����	  �E�}� t�    ��X H�E���H���U ����UH��H�� �}��:C H�E��E���H�U�H�E���H���	  �E�}� t�    ��W H�E���H���U ����UH��H�� �}���B H�E��E���H�U�H�E���H���/	  �E�}� t�    ��E����!
  ����UH��H�� �}��B H�E��E���H�U�H�E���H����  �E�}� t�    ��E���������UH��H�� �}���B H�E��M�H�U�H�E���H���B �E�}� t�    ���V H�E���H���lK ����UH��H�� �}��B H�E��M�H�U�H�E���H���JB �E�}� t�    ��V H�E���H����K ����UH��H�� �}��/B H�E��M�H�U�H�E���H����A �E�}� t�    ��,V H�E���H���LL ����UH��H�� �}���A H�E��M�H�U�H�E���H���A �E�}� t�    ���U H�E���H����L ����UH��H�� �}��A H�E��M�H�U�H�E���H���QA �E�}� t�    ��U H�E���H���bM ����UH��H�� �}��6A H�E��M�H�U�H�E���H����@ �E�}� t�    ��3U H�E���H���O ����UH��H�� �}���@ H�E��M�H�U�H�E���H���@ �E�}� t�    ���T H�E���H���O ����UH��H�� �}��@ H�E��M�H�U�H�E���H���X@ �E�}� t�    ��T H�E���H���P ����UH��H�� �}��=@ H�E��M�H�U�H�E���H���@ �E�}� t�    ��:T H�E���H���P ����UH��H�� �}���? H�E��M�H�U�H�E���H���? �E�}� t�    ���S H�E���H����P ����UH��H�� �}��? H�E��M�H�U�H�E���H���_? �E�}� t�    ��S H�E���H���ZQ ����UH��H�� �}��D? H�E��M�H�U�H�E���H���? �E�}� t�    ��E�����  ����UH��H��  H������H������H������H��H����  H������H�5=s H����  H������H������H������H��H���  ��t
�   �X  H������H�5�r H���  H������H������H������H��H����  ��t
�   �  H������H�5�r H���`  H������H������H������H��H���  ��t
�   ��  H������H�5�r H���  H������H������H������H��H���N  ��t
�   �  H������H�5Er H����  H������H������H������H��H���
  ��t
�   �H  H������H�5r H���  H������H������H������H��H����  ��t
�   �  H�� ���H�5�q H���P  H�� ���H�����H������H��H���  ��t
�   ��  H�����H�5�q H���  H�����H�����H������H��H���>  ��t
�   �|  H�� ���H�5Mq H����  H�� ���H��(���H������H��H����  ��t
�	   �8  H��0���H�5q H���  H��0���H��8���H������H��H���  ��t
�
   ��   H��@���H�5�p H���@  H��@���H��H���H������H��H���r  ��t
�   �   H��P���H�5�p H����  H��P���H��X���H������H��H���.  ��t�   �oH��`���H�ºC H��H���Ԇ��H��`���H�5@p H������H��H������H��H���߆��H�5,p H���І��H������H��`���H��譆���    ��UH��H���}�H�u�H��p �  H�5�o H�=p �Ɂ��UH��H�� �}��: H�E��E���H�U�H�E���H����   �E�}� t�E���O H�E���H���M ��UH��H�� �}��.: H�E��E���H�U�H�E���H���y   �E�}� t�E���N H�E���H����M ��UH��H���}�H��o �  H�50o H�=Qo �����UH��H���}�H��o �$  H�5o H�='o �Ӏ��UH��H��`H�}���H�U��E��E��E��E���x H�E��@��t�U�H�E���    ��   H�E�H�E�H�E�H��H�E�H�E�H�E�H�E�H��H�E�f�E�  f�E�  �E�    H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� t�E��]H�U�H�E�H9�tH��n �>   H�5em H�=�m ����H�U�H�E�H9�tH��n �?   H�59m H�=um �����    ��UH��}��}�v�}�t�}�v�}��   w�   ��    ]�UH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�PH�E�H�� ��tH�E�H�@H�PH�E�H�P�Ԑ]�UH��H�}�H��H��H��H�E�H�U�H�E�H�PH�E�H9�t�    �LH�E�    H�E�H�@H9E�s1H�E�H�H�E�H��H�M�H�E�H�� 8�t�    �H�E����   ]�UH��ATSH���   H��H��H��H�� ���H�����H�E�    H��@ C H� H�U�H��H�H� H���F  H��@ C H� H�U�H��H�H�H�����H��H������H������    �=   H����  H�E�H�}����   H�� ���H�ºC H��H��蒂��H�� ���H�5fm H��貂��H��H�����H����  I��H�����H����  H��H�E�L��H���.  H�U�H�E�H��H��H���  H�5+m H���W���H��衂��H�� ���H���4����GH�U�H������    H���  H�E�H�U�H�� ���H�����H�E�H��H��������tH�E��H�E�����H������H���   [A\]�UH���[b ������tRH�=Kb �K ������t=�1 H�0H�=b �  H�="b �K H�VJ H�5�a H����@ H���|��H��a ]�UH��H�� ����H�E�H�E�H����  H��H��@ C H� H9�������   H�E�H����  H�E�    H��@ C H� H�U�H��H�H� H��t+H��@ C H� H�U�H��H�H�E�H��H���  H�E��H�E�    H�U�H�E�H��H���
	  H�E�H���@  H��H��@ C H�����UH��SH��HH��H��H��H��H��H�u�H�}�H�U��ȈE�����H�E�H�E�H����  H��H��@ C H� H9�����tH�� �>   H�5*k H�=Kk �o{��H�U�H�E�H��H������H�E�H�}��t&�}� ��   H�]�H�U�H�E�H��H���  H��fH�E�H����  H� H������tH�� �F   H�5�j H�=�j ��z��H�]�H�E�H���  H�H�E�    H�U�H�E�H��H����  H�E�H���  H��H��@ C H��H��H[]�UH��SH��(H��H��H��H�E�H�U��f���H�E�H�E�H����  H��H��@ C H� H9�����tH��~ �Q   H�5�i H�=j �?z��H�U�H�E�H��H���f���H�E�H�}��uH��    H��uH�=j �S��H�E�H����  H��vH�E�H���  H� H��t�   ��    ��tH�a~ �W   H�5mi H�=j �y��H�E�H���}  H�P�H�E�H��H���"  H��H�U�H�E�H��H���  H��H���l  H�E�H���  H�E�H���  H�     H�E�H���  H��H��@ C H��H��([]�UH��H��@H�}�H�U�H�E�H��H���|���H�U�H�E�H��H���:���H�E�H�}��u
�    �   H��@ C H� H�U�H��H�H�H�E�H��H���-���H�Eк    �=   H���E  H�E�H�}��uH�E} �i   H�5?h H�=�h �x��H�E�H���c  H��H�E�H��H���UH��SH��8H�}�H�U�H�E�H��H������H�Eк    �=   H����  H�E�H�}��uH��| �q   H�5�g H�=�h �x���S���H�U�H�Eо    H���3  H�u�H��H��H��H�й   H��H��������    H��8[]�UH��ATSH��  H������H������������H������H�����H��H�������H������    �=   H���  H�E�H�}����   H�� ���H�ºC H��H����{��H�� ���H�5�g H����{��H��H�����H���	  I��H�����H���	  H��H�E�L��H���g  H�U�H�E�H��H��H����  H�5�g H���{��H����{��H�� ���H���m{��H���C �   �������   H������H������H�����H�5�g H�Ǹ    �tO  ������tH�%{ ��   H�5f H�=Zg �Vv��H�����H��uH��z ��   H�5�e H�=[g �+v���v��������� ��D��H�����H������H�E�H��H���d���H�u�H�E�D��H��H��H��������    H��  [A\]�UH��H�� H�}�����H�U�H�E�H��H������H�U�H�E�H��H��������    ��UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H�}��H�U؈E�H�E�H�E�H�E�H�@H9E�s#H�E�H�H�E�H�� 8E�uH�E��H�E���H������]ÐUH��H�}�H�E�H� ]ÐUH��H�}�H�E�H�@]�UH��H�� H�}�H��H��H��H�E�H�U�H�U�H�E�H��H���S  H�E���UH��H��0H�}�H�u�H�U�H�U�H�E�H�H�E�H�@H9�vH��    H��uH�=�e ��M��H�E�H�H�E�H�H�U�H�E�H��H���.  H�E�H�U���UH��SH��H�}�H�u�H�]�H�E�H���-  H�H�E�H�@    H�E�H�@    H�E�H�@    �H��[]�UH��H�� H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H�U�H�RH��H��蒣����ÐUH��H�}�H�E�H�@]�UH��H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H�@    �]�UH��H�� H�}�H�u�H�E�H�@H�PH�E�H��H���[  H�E�H�PH�E�H�@H��H�H�ƿ   �8u��H�U�H�H�H�E�H�E�H�@H�PH�E�H�PH�E��ÐUH��SH��(H�}�H�u�H�E�H�@H�PH�E�H��H����  H�E�H���   H��H�E�H�PH�E�H�@H��H�H�ƿ   �t��H�H�E�H�E�H�@H�PH�E�H�PH�E�H��([]ÐUH��H�}�H�u�H�E�H�@H�U�H��H�]ÐUH��H�}�H�E�H�PH�E�H�@H��H��H�]ÐUH��H�}�H�E�H�@]�UH��H�}�H�E�H� ]�UH��H�� H�}�H�u�H�E�H�������H�E�H�E�H�������H��H�E�H�H�E�H������H��H�E�H����UH��H�� H�}�H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��H�H���a���H�E�H�E���UH��H��0H�}�H�u�H�E�H���}s��H�M�H�U�H�E�H�0H�@H��H���H  H�E�H���Ct�����UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H�}�H�E�H� ]ÐUH��SH��8H�}�H�u�H�E�H�@H9E���   H�E�H�H�E�H�E�H�U�H��H��H��觠��H�E�H�E�    H�E�H�@H9E�sHH�E�H�@H�U�H��H�H���X���H��H�E�H��    H�E�H�H�ƿ   �dr��H�H�E��H�E�    H�E�H�@H9E�sH�E���H�E�H�U�H�RH��H������H�E�H�U�H�PH�E�H�U�H�P��H��8[]�UH��H��PI��H��L��L��H��H�u�H�}�H�U�H�M�H�E�H�E�H�E�    H�E�H9E���  H�U�H�E�H�� �E�}�`v�}�zv�}�@v �}�Zw�E���H�E���H������q  �}�/v �}�9w�E���H�E���H����~���K  �}� uH�E��    H����~���/  �E��H�=�` � H������t�E���H�E���H���~����   �}�\uH�E�H�5�` H���>x����   �}�"uH�E�H�5p` H��� x���   �}�'uH�E�H�5U` H���x���   �}�
uH�E�H�5:` H����w���   �}�	uH�E�H�5` H����w���fH�E�H�5` H���w��H�E�H�M��   H��H��蹔���E�E�H�U�H�M�H�E�H��H���*   H�E�H���q��H�E��}   H���}��H�E��4������UH��H��@H�}�H�u�H�U�H�U�H�E�H��H���Fp��H�E؋ H�U�H�M�H�Ή��Zu��H�E�H���p����ÐUH��H��H�}�H�u�H���B H�PH�E�H�H�E��@H    H�E��@L    H�E�H�U�H�PPH�E�H��XH���6   H�E�H�@    H�E�H�@�   H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�@0    H�E�H�@8    H�E��@@    H�E��@D    H�E�H��H�=2R ��  ���UH��H���   H��H���H���B H�PH��H���H�H��H���H�P0H��H���H�@8H9�tFH��`���H�ºC H��H����p��H��`���H�5�q H���q��H���Wq��H��`���H����p��H��H���H�@H��t�I  H��H��H���H�@H��H������H��H���H��H�=cQ �   H��X���H��X���H��H�=FQ ��   ���UH��H��H�}�H�E�H�������H�E��p   H���Kg���ÐUH��H��H�}�H�E�H�@PH��tH�E�H�@PH�U�H�������ÐUH��H���   H��(���H�� ���H�����H�����H�����H��uH�7� �W   H�5�p H�=�p �)k��H��(���H���u  ������t
������%  H��(����@L����   H��(���H� H��(H� H�����H��8���H�� ���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��  H��8���H��uH��(����@D����H��(����PDH��8���H�����H��    �y  H��(����@@��tVH��(���H�@(H��tFH��@���H�»C H��H����m��H��@���H�5�o H���n��H���_n��H��@���H����m��H��(����@@    H��(���H�PH��(���H�@(H9��  H��(���H���
  �E��}� t�E���  H��(���H���  �E�}� t�E��  H��(���H���4  H��(���H� H��(H� H��(���H�RH��(���H�qH��0���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��8  H��0���H��u1H��(����@D����H��(����PDH�����H�     �    ��   H��0���H��(���H�P H��0���H��(���H�P(H��(���H�PH��(���H�@(H9�rH��� ��   H�5�m H�=Un �h��H��(���H�P(H��(���H�@H)�H��H�E�H�����H�E�H��H���C   H� H�E�H��(���H�PH��(���H�@H�H�U�H�� ���H��H���x��H��(���H�PH�E�H�H��(���H�PH�����H�U�H��    �ÐUH��H��   H�����H�����H�����H�� ���H�����H��uH��� ��   H�5m H�=%m �g��H�����H����  ������t
������Q  H������@L����   H�����H�P0H�����H�@8H9�tH�1� ��   H�5�l H�=m �g��H�����H� H��0H� H�����H�� ���H�����H������ЉE��}� t!H������@D����H������PD�E��  H�� ���H��uH��� ��   H�5l H�=�l �f��H�� ���H�� ���H��    �e  H�����H�PH�����H�@H9�u@H�����H���2  �E�}� t�E��*  H�����H���&
  �E��}� t�E��
  H������@@��uVH�����H�@(H��tFH��0���H�»C H��H���i��H��0���H�5~k H����i��H���(j��H��0���H���i��H������@@   H�����H�PH�����H�@H9�rH��� ��   H�5�j H�=�k �xe��H�����H�PH�����H�@H)�H��H�E�H�����H�E�H��H���<  H� H��(����E� H������@L��u@H��(���H������
   H���
 H�E�H�}� tH�E�H��H+����H��(����E�H��(���H��uH�͆ ��   H�55j H�=)k �d��H�����H���d	  H��(���H�����H�HH�����H�@H�H�����H��H���u��H�����H�P0H�����H�@8H9�trH�����H�PH�����H��0H��H���7  H�H�����H�P0H�����H�PH��(���H�H�E�H�����H�P8H�E�H��H���W���H�H�����H�P8�6H�����H�PH�����H�P0H�����H�PH��(���H�H�����H�P8H�����H�P(H�����H�HH��(���H�H�E�H�E�H��H���ޓ��H�H�����H�P(H�����H�PH��(���H�H�����H�P�}� tH�����H���  ������t������H��(���H�� ���H��    �ÐUH��H��H�}����E�H�E�H�@H��uH�� ��   H�5Uh H�=Oi ��b��H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��E���ÐUH��H��H�}��u�H�E�H�P0H�E�H�@8H9�tH��� ��   H�5�g H�=�h �fb��H�E��U�PL�    ��UH��H�}�H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�P0H�E�H�P8�]ÐUH��H�� H�}�H�E�H�P8H�E�H�@0H9�tH�E�H����  �E��}� t�E��+H�E�H���  �E��}� t�E��H�E�H���_����    ��UH��H�� H�}�H�u�H�E�H� H��8H� H�U�H�}�H�Ѻ   �    �ЉE��}� t�E��)H�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H��    ��UH��H��@H�}�H�uЉU�H�E�H����  �E��}� t�E���   �}�ueH�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� ��   H�E؋@D����H�E؉PD�E��|�}� t%�}�tH��� �  H�5�e H�=]g �y`��H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� tH�E؋@D����H�E؉PD�E��H�E�H��������    �ÐUH��H�� H�}�H�E�@H��t�    �_H�E�H� H��H� H�U�H�JHH�U�H��H���ЉE��}� t�E��/H�E�@H��uH�� �%  H�5(e H�=�f �_���    �ÐUH��H��H�}�H�E��@L��t�    �aH�E�H� H�� H� H�U�H�JLH�U�H��H���Ѕ�����t������/H�E��@L��uH�r� �/  H�5�d H�=Wf �+_���    �ÐUH��H��0H�}�H�E�H��������E��}� t�E���  H�E�H�P0H�E�H�@8H9�u
�    �  H�E؋@H��u\H�E�H� H��8H� H�U�H�R0H��H�U�H�R H��H)�H�U�H�}�H�Ѻ   �ЉE��}� t�E��S  H�E�H�P0H�E�H�P �_H�E؋@H��tH��� �B  H�5�c H�=�e �H^��H�E�H�P H�E�H�@0H9�tH�k� �C  H�5�c H�=�e �^��H�E�H�P H�E�H�@8H9���   H�E�H� H��0H� H�U�H�J8H�U�H�R H)�I��H�U�H�JH�U�H�R H�4H�U�H�}�H��L���ЉE�}� tH�E؋@D����H�E؉PD�E��`H�E�H��uH�� �M  H�5�b H�=vc �j]��H�E�H�P H�E�H�H�E�H�P H�E�H�P0H�E�H�H�E�H�P0�#����    �ÐUH��H���   H��8���H��8���H��������E��}� t�E���   H��8����@H����   H��8���H�@H��H��8���H�@ H)�H��H�E�H��8���H� H��8H� H��H���H�u�H��8���H�Ѻ   �ЉE�}� ttH��8����@D����H��8����PDH��P���H�ºC H��H����`��H��P���H�5�c H���a��H�E��H���^  H���>a��H��P���H����`���E���    ��    ��UH��H�� H�}�H�E�H��������E��}� t�E��   H�E�@H��u4H�E�H�PH�E�H�@(H9�tH�	~ �m  H�5!a H�=Lc �[��H�E�H�P0H�E�H�@8H9�tH��} �o  H�5�` H�=aa �r[��H�E�H�@    H�E�H�@     H�E�H�@(    �    ��UH��H�� H�}�H�E�H�@H��uH�~} �x  H�5�` H�=�b �[��H�E�H�@H��u-�  H��H�E�H�@H��H������H�E�H�E�H�U�H�P���ÐUH��H�� H�}��u�H�U�H�E�H�U�H��H������H����B H�PH�E�H�H�E��U�Pp��ÐUH��H�}�H�E��@p]ÐUH��H��   H��X���H��X���H�P0H��X���H�@8H9�tFH��`���H�ºC H��H���^��H��`���H�5�a H����^��H���"_��H��`���H���^��H��X����@p��� �E��}� t�E���    �ÐUH��H�� H�}�H�u�H�E�@pH�U�H�Ѻ   �    ��� �E��}� uH�E��    �    ��}�-  uH�E��    �    ��E���UH��H��   H��X���H��P���H��    H��u6H��{ ��  H�5�^ H�=?a �?Z��H��P����    �    �   H��X����@p���2���E��}� uH��P����    �    �h�}�"  uH��P����    �    �KH��`���H�ºC H��H���=]��H��`���H�5�` H���]]��H���]��H��`���H���:]��������ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u�����
 �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u����
 �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u��U�H�M�H�E�@pH�MЋU�H�u����
 �E��}� t�E���    �ÐUH��H�}��]ÐUH��H���   H��8���H��< H�E�H�E�H���  H��H���H�E�H����  H��@���H��@���H��H���H��H����  ����   H��H���H���  H�E�H�E�H��������E�}� tFH��P���H�ºC H��H���e[��H��P���H�5Y_ H���[��H����[��H��P���H���b[��H��H���H���q  �]������UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���������UH��H��H�}�H�E�H�������ÐUH��H��H�}�H�u��[
 H��H�E�H��H���a  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��p  H������H������H�������+   H�����  H�����E�H������� <ru�}� t�E�   �   �E�   �   H������� <wu�}� t	�E�   ��E�   �M�  �oH������H�ºC H��H����Y��H������H�5�] H����Y��H��H������� ����H���+  H�5�] H����Y��H���Z��H������H���Y��H������H������� ����   H������� <+u
H��������H������� <bu
H�������H������� <eu�M� @  H�������H��P���H�ºC H��H����X��H��P���H�56] H���Y��H��H������H��H���Y��H�5] H����X��H���=Y��H��P���H����X��H�������(���H�������M�H��������H���H �E�}� tH���C �U��    �.�� H��H�U�H������H��H���q  H��tH����    ��UH��H��H�}�H�u�� H��H�E�H��H����  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��   ��\���H��P���H��`���H�ºC H��H���W��H��`���H�5\ H����W��H�5\ H���W��H���X��H��`���H���W��� H��H�U�H��\���H��H���  H��tH����    ��UH��H�� H�}�H�}� t
H�E�H����    H�E��E�    H�E�H���g���������t�E�����H�E�H� H��H� H�U�H���Ѕ�����t�E�����H�E�H�������E���UH��H��0H�}�H�u��U�H�}� t
H�E�H����    H�E��U�H�M�H�E�H��H�������E�}� tH���C �U��������    ��UH��H��0H�}�H�}� t
H�E�H����    H�E�H�U�H�E�H��H��������E�}� tH���C �U�H�������H�E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���*���������t�������    ��UH��H��H�}�H�E�H��������UH��H��@H�}�H�uЉU�H�M�H�}� t
H�E�H����    H�E��}�u1H�E��   H�������E�}� ��   H���C �U��������}�u-H�E��   H��������E��}� tZH���C �U��������L�}�u-H�E��   H�������E�}� t'H���C �U�������H���C �   �������    ��UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E��    �    H������H�E�@<�����H�E�P<���UH��H�� �}�H�u�H�}� t
H�E�H����    H�E��E���H�E���H�������E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���
������UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H���'��H�E�H�E�H���  D� H�E�H������H�������I��H�E�H�ƿx   �Q��H��L��D��H������H��H��8[A\A]]�UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H���~��H�E�H�E�H���  D� H�E�H������H������I��H�E�H�ƿx   �oP��H��L��D��H���u���H��H��8[A\A]]�UH��H���}��u��}���   �}���  ��   H�=s3 ��   �    �    H�=}3 � ���H�q H�5j3 H���@ H����M���    �   H�=�3 �����H�> H�5�3 H���@ H���M���    �   H�=4 ����H� H�54 H���@ H���\M��H�=f4 �����H�� H�5S4 H�=�����6M�����UH����  �   �����]ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@ �]�UH��SH��(H�}�H�u�H�E�H��uH��    H��uH�=�U �6&��H�E�H���3  H�E�H�U�H�E�H��H���+  �@��tH��    H��uH�=�U ��%��H�U�H�E�H��H����  H� H������tH��    H��uH�=V �%��H�U�H�E�H��H���  H�@H������tH��    H��uH�=!V �|%��H�E�H�@H��uH�E�H���  H��H�E�H��HH�E�H�XH�U�H�E�H��H���T  H�XH�E�H���t  H��H�E�H�PH�E�H��H���*  H�H�E�H�U�H�PH�U�H�E�H��H���  �@H�U�H�E�H��H���3  H�E�H��([]�UH��H�� H�}�H�u�H�U�H�E�H��H����  �@����tH��    H��uH�=�U �$��H�U�H�E�H��H����  H�E��ÐUH��SH��8H�}�H�u�H�E�H��uH��    H��uH�=�U �8$��H�U�H�E�H��H���=  �@����tH��    H��uH�=�U � $��H�U�H�E�H��H���  H���-  H�E�H�U�H�E�H��H����  H�@H�E�H�E�H��u9H�E�H�PH�E�H9�tH��    H��uH�=�U �#��H�E�H�U�H�P�pH�E�H���  H��H�E�H��H���~  H�PH�E�H9�����tH��    H��uH�=�U �:#��H�]�H�E�H���3  H��H�E�H��H���0  H�XH�}� ueH�E�H� H���  H��H�E�H9�����tH��    H��uH�=�U ��"��H�E�H���  H�E�H�E�H����  H��H�E�H��   H�U�H�E�H��H���  H� H���  H��H�E�H9�����tH��    H��uH�=�U �_"��H�U�H�E�H��H���d  H���  H�E�H�E�H���|  H��H�U�H�E�H��H���6  H�H�E�H���  H��H�E�H9�����tH��    H��uH�=�U ��!��H�U�H�E�H��H����  H�     H�U�H�E�H��H����  H�@    H�U�H�E�H��H���  �@ H�E�H��8[]�UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]�UH��H��H�}��u�H�U�H�E�H��H���  H�E���UH��H�� H�}�H�E�H� H���(  H��H�E�H��H���g  H�E��ÐUH��H�� H�}�H�E��    H���C  H�E��ÐUH��H��H�}�H�u�H�U�H�E�H��H���w  ����UH��H��H�}�H�E�H�H�E�H��H���r  H�H�E�H�H�E���UH��H�}�H�E�H� ]ÐUH��H��H�}����E�H�U�H�E�H��H���\  H�E���UH��H��H�}�H�u�H�}� t-H�E�H� H� H�U�H����H�M�H�E��p   H��H���\  ����UH��H�}�H�E�]�UH��H�}�H�E�]ÐUH��H��H�}�H�u�H�E�H���O  H��H�E�H��H���X  ��UH��H�}�H�E�H� ]ÐUH��H�}�H�u�H�E�H�U�H��]�UH��H��0H�}�H�u�H�E�H���H��H�E؋ H�U�H�M�H�Ή��  H�E�H����H����ÐUH��H�}�H�u�H�E�H�H�E�H� H9���]�UH��H��H�}�H�u�H�E�H���   H��H�E�H��H���   ��UH��H��0H�}�H�u�H�E�H���~G��H�E�� ��H�U�H�M�H�Ή��v   H�E�H���FH����ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���   ���UH��H��H�}�H�E�H���  �ÐUH��H�}�H�u�X   H�E�H�]�UH��H��@�}�H�u�H�U�H�U�H�E�H��H���"G��H�U�H�M��E�H�Ή��Y  H�E�H���G�����UH��SH��hH�}�H�u�H�U�H�}� �  H�}� �  vH�U�H�E�H��H���u����  H�E�H�E�H�E�H%  ��H�E�H�E�H�U�H��H���Ӂ������tH��    H��uH�=�Y �r��H�E��@HH�H��H��H��H�E�H�H��H�E�H�E��@H���r��H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=�Y � ��H�U�H�E�H��H����~��H�E�H�@PH�����E�H�E��@L��uH��    H��uH�=�Y ���H�E�H�ƿ   �7E��H��H���ŀ��H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H��賀������t�   ��    ��tH��    H��uH�=�Y �B��H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H��蔀��H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H����}����H��h[]�UH��H�}�H�E�]�UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=m\ �@���u�H�E�A�    A�   �    �
   H���   ���UH��H��0H�}�u�U��M�D�E�D�ȈEԃ}� y=�E��؉E��M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ   H���VN��H���3�M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��E H�E��E�    �E���~H��    H��uH�=�a �)���E���}���Hc�H�E�H���E��H�M�H��T��E���}��E��}� t맀}� t2�E���~H��    H��uH�=�a �����E��P�U�H��D�-H�U�H�E�H��H����N��� 9E�����tE�E�    H�U�H�E�H��H���N��� �U�)�9E�����t�U�H�E���H���rO���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���;O���E��ڋE����E�}� x!�E�H��D���H�E���H���O���m��ِ��UH��H��H�}�H����B H�PH�E�H�H�E�H���x�����ÐUH��H��H�}�H�E�H������H�E��x   H���:���ÐUH��H��H�}�H�� ��   H�5�a H�=%b ��>��UH��H�� H�}�H�u�H��    H��u3H�ڈ ��   H�5�a H�=b �?��H���C �   ������4H�U�H�E�H��H������E��}� tH���C �U���������    ��UH��H�� �}�H�u��U�H�M�H�e� ��   H�51a H�=ka �&>��UH��H�R� ��   H�5a H�=Ha �>��UH��H��H�}�H�/� ��   H�5�` H�=a ��=��UH��H�� H�}�H�u�H�U�H�� ��   H�5�` H�=�` �=��UH��H��H�}�H�u�H�݇ ��   H�5�` H�=�` �v=�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���$  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L�����UH��H���   H��(���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��X C H� H��0���H��(���H��H���  ��L�����L�����UH��H�}��u�H�U�}���   �E�H��    H��^ �H�H��^ H���H�E��H�E���]H�E��H�E�f��NH�U�H�E�H��AH�U�H�E�H��4H�U�H�E�H��'H�U�H�E�H��H�E�H�U�H��H�E��H�E����]�UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��� �p  H�5=] H�=w] �2:��UH��H���   H��(���H�� ���H�����H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�����H�� ���H��(���H����  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L����ÐUH��H�}�H�E�H� � ]�UH��H�}�H�E��@�PH�E��PH�E�H� H�HH�U�H�
� ]�UH��H��   H�����H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�Hǅ0���    Hǅ8���    H�����H��0���ǅ���   ǅ���0   H�EH�� ���H��P���H��(���H�����H�� ���H��0���H��H���7  ��L�����L�����UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���c3  H�U�H�M�H�E�H��H���9  H�M�H�U�H�u�H�E�H��H���9  H�E��ÐUH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H������H�E�H��tH�E�H� �U��҉�H�������H�E�H��t�E���    ��UH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H���#���H�E�H��tH�E�@�PH�E�PH�E�H��t�E���    ��UH��H��@H�}�H�u�H�U�H�}� t
H�E�H����    H�E�H�E�    H�E�    H�E�H�E�H�U�H�M�H�E�H��H���P$  ���UH��H��H�}�H�u�H��X C H� H�U�H�M�H��H���8�����UH��H��H�}�H�u�H�2� ��  H�5�X H�=�X �5��UH��SH��   H�}�H�u�H��x���H��p���H�}� u
�    �   H�M�H��p���H�H�VH�H�QH�FH�AH�E�H�P�H�M�H�E�H��H���3  H�U�H�M�H�E�H��H����=  H�M�H��x���H�u�H�E�H��H����=  H�]�H�E�H��H�E�H�E�H�PH�E�H��H�������H� H��  H�E�H�Ĉ   []�UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���1  H�U�H�M�H�E�H��H���D  H�M�H�U�H�u�H�E�H��H���"D  H�U�H�E�H��  H�E���UH��H�� H�}�H�u�H�U�H��~ ��  H�5W H�=UW �4��UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�O~ ��  H�5�V H�=DW �3��UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��} ��  H�5+V H�=�V � 3��UH��H�� H�}�H�u�H�U�H��} ��  H�5�U H�=�V ��2��UH��H�� H�}�H�u�H�U�H��} ��  H�5�U H�=fV �2��UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�1} ��  H�5MU H�=�U �B2��UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��| ��  H�5�T H�=vU ��1��UH��H�� H�}�H�u�H�U�H�M�H��| ��  H�5�T H�=?U �1��UH��H�� H�}�H�u�H�U�H�M�H�s| ��  H�5gT H�=U �\1��UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�| ��  H�5�S H�=�T ��0��UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��{ ��  H�5wS H�=T �l0��UH��H��H�}�H�u�H�t{ ��  H�5HS H�=�S �=0��UH��H��H�}�H�u�H�U{ ��  H�5S H�=�S �0��UH��H�� H�}�H�U�H�E�H�Ѻ   �   H���u  H�E�H�}�t�������E�����UH��H��0H�}�H�u�H�U�H�}� uH��z ��  H�5�R H�=]S �/��H�E�    H�E�H��H9E�uH�U�H�E�H��  H�E��oH�E�H���L����E�}��u"H�}� tH�U�H�E�H��  H�E��?�    �8H�U�H�E�HЋU��}�
uH�E�H�PH�E�H��  H�E��
H�E��o�����UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���  H������t�������   ��UH��H���}�H�u�H�U��E�H�։�������UH��H��H�}�H�u�H�E�H���@��H��H�U�H�E�H�Ѻ   H���  H������t�������   ��UH��H��H�}�H�u�H�U�H�E�H��H��������UH��H��H�}�H�E�H���	  ��UH��H��H�}�H�E�H���������UH��H��P C H� H���]	  ]�UH��H��P C H� H������]�UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���?  H������t�������E���UH��H���}�H�u�H�U��E�H�։�������UH��H���}�H��X C H��E�H�։��s�����UH��H���}��E����������UH��H��@H�}�H��X C H� H��tH��X C H� H����    H�E�H�E�    H�E�H���Z>��H�E�H�E�H;E�sQH�E�H+E�H��H�M�H�E�H�4H�M�H�E�H������������t������NH�E�H��u������>H�E�HE��H�U�H�E�H�Ѻ   H�5 P H���d���������t�������   ��UH��H��H�}�H�Vw �f  H�5O H�=�O �,��UH��H�� H�}��u�H�U�H�+w �g  H�5�N H�={O ��+��UH��H���}�H�u�H�w �h  H�5�N H�=MO �+��UH��H��H�}�H�u�H��v �i  H�5}N H�=O �r+��UH��H��H�}��u�H��v �j  H�5ON H�=�N �D+��UH��H��H�}�H��v �k  H�5$N H�=�N �+��UH��H�uv �l  H�5N H�=�N ��*��UH��H���}�H�u�H�Pv �m  H�5�M H�=tN ��*��UH��H���}�H�-v �n  H�5�M H�=JN �*��UH��H���}�H�u�H�v �o  H�5{M H�=N �p*��UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���  ��UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���!  ��UH��H��H�}�H�u�H��u �z  H�5�L H�="M ��)��UH��H��H�}�H�u�H�]u �  H�5�L H�=�L �)��UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�H���C � �E�H�}� t-H�E�� ��t"H��H C H� H�U�H�5M H�Ǹ    �����E�����  H��H��H C H� H�5�L H�Ǹ    �������UH��SH���   H�����H�����H�����H����� t
H����� uH���C �   H�������^  H�E�    H�E�    H�����H� H��tH�����H� H�E�H�����H� H�E�H�}� u��  �   H���WX��H�E�H�E�   H�����H�M�H�E�H��H���d���H������tH��������   H�E�H���9��H�E�H�U�H�E�H�� 
H�E�H�PH�E�H��  H�� ���H�ºC H��H���T,��H�� ���H�5�K H���t,��H��H�E�H�PH�M�H�E�H��H������H�U�H�E�H��H��H��蔲��H���,��H�� ���H���,��H�����H�U�H�H�����H�U�H�H�E�H��H���   []�UH��H�� H�}�H�u��U�H�M�H��r ��  H�5J H�=OJ �
'��UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���   ��L�����L�����UH��H��pH�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�E�H���%  H�U�H�M�H�E�H��H���<  H�M�H�U�H�u�H�E�H��H���<  H�E�H���%  H�U�H�E�H��  H�U�H�E�H�H�E���UH��H��   H��X���H��`���H�ºC H��H���*��H��`���H�5qI H���5*��H���*��H��`���H���*�����UH��H��   H��X���H��`���H�ºC H��H���)��H��`���H�5FI H����)��H���$*��H��`���H���)�����UH��H��   H��X���H��`���H�ºC H��H���_)��H��`���H�5I H���)��H����)��H��`���H���\)�����UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�H�U�H�E�H�Ѻ   �   H�������H������t�������E�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H������������tHH������H�ºC H��H����'��H������H�5�G H����'��H���9(��H������H����'���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H������������tHH��@���H�ºC H��H����&��H��@���H�5�F H���'��H���N'��H��@���H����&���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H���R���������tHH������H�ºC H��H���%��H������H�5�E H���%��H����%��H������H���%���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H���g���������tHH��@���H�ºC H��H���$��H��@���H�5�D H����$��H���%��H��@���H���$���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H�� H�}��u�H�U�H�gk �b  H�5�B H�=�B ���UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� ����譓��������tbH�� ���H��� ����茓��������t
H�� �����H�����H���+��������`�����������  H�����H��������H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� ����跐����tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H�ºC H��H����!��H�� ���H�5-B H���"��H���P"��H�� ���H����!��H�� ����T  H�� ���� <muSH������H�ºC H��H���!��H������H�5�A H���!��H����!��H������H���!��H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H�8A �H�H�,A H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H�A �H�H�A H����E�
   H�E�    H�����H��������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���m����E�륀}�0uHH�����H���g���H�����H���D����E׀}�xu!H�����H���@���H�����H�������E׀}�/~2�}�9,H�����H������H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H�������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H������H�E�H��H���E׃�AH�H�H�E�H�����H���]����E��;����}�/~S�}�7MH�����H���N���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H�������E�뭐����H�}� ��  H�U؋M�H�E���H���L����  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���n����E��H�}� �/  H�UȋM�H�E���H�������  H�E�    H�����H���-����E��}�0uHH�����H���)���H�����H�������E��}�xu!H�����H������H�����H��������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H���e���H�E�H��H���E���AH�H�H�E�H�����H���'����E��C���H�}� ��  H�U��M�H�E���H���p�����  H�E�H�E�H�����H��������E��E�    �}� t�E���������u�   ��    ��tPH�����H������H�}� t�E�Hc�H�E�H��E��H�����H���|����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H���'����E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H�������H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H���%��ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H���0����E��}� te�E�;E�}]H�����H���$����E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H��������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H�������E��}�0uHH�����H������H�����H���^����E��}�xu!H�����H���Z���H�����H���7����E��}�/~2�}�9,H�����H���-���H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H�������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H������H�E�H��H���E���AH�H�H�E�H�����H�������E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E���UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� ��������������tbH�� ���H��� �����ͅ��������t
H�� �����H�����H����������衅����������  H�����H���B�����H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� �����������tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H�ºC H��H���'��H�� ���H�5n4 H���G��H�����H�� ���H���$��H�� ����T  H�� ���� <muSH������H�ºC H��H������H������H�5*4 H������H���0��H������H������H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H��: �H�H��: H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H��: �H�H��: H����E�
   H�E�    H�����H�������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H�������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���H����E�륀}�0uHH�����H������H�����H�������E׀}�xu!H�����H���i���H�����H��������E׀}�/~2�}�9,H�����H���<���H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H�������H�E�H��H���E׃�AH�H�H�E�H�����H���8����E��;����}�/~S�}�7MH�����H���w���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H��������E�뭐����H�}� ��  H�U؋M�H�E���H�������  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H�������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���I����E��H�}� �/  H�UȋM�H�E���H��������  H�E�    H�����H�������E��}�0uHH�����H���R���H�����H��������E��}�xu!H�����H���+���H�����H�������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H�������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H������H�E�H��H���E���AH�H�H�E�H�����H�������E��C���H�}� ��  H�U��M�H�E���H��������  H�E�H�E�H�����H�������E��E�    �}� t�E����H}����u�   ��    ��tPH�����H�������H�}� t�E�Hc�H�E�H��E��H�����H���W����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H�������E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H���(���H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H������ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H�������E��}� te�E�;E�}]H�����H���M����E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H�������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H���`����E��}�0uHH�����H������H�����H���9����E��}�xu!H�����H������H�����H�������E��}�/~2�}�9,H�����H���V���H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H�������H�E�H��H���E���AH�H�H�E�H�����H���Z����E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H��H�}����E�H�E�H�H�E�H�Ѻ   �   H���l���H�E�H�@H�PH�E�H�P���UH��SH��H�}�H�u�H�E�H�H�E�H�����H��H�E�H�ٺ   H������H�E�H������H��H�E�H�@H�H�E�H�P�H��[]ÐUH��H�� H�}�H�u�H�U�H�E�H�H�u�H�E�H�Ѻ   H������H�E�H�PH�E�H�H�E�H�P��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H�}����E�H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]�UH��H�}�H�u�H�E�    H�U�H�E�H�� ��t>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�밐]ÐUH��H�}�H�u�H�U�H�E�    H�E�H;E�s>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�븐]ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�PH�E�H�@    �]�UH��H�}����E�H�E�H�PH�E�H�@H9�sH�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]ÐUH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���e���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E�H�     H�E�H�@    H�E�H�@    �]�UH��H��0H�}�H�E�H�PH�E�H�@H9���   H�E�   H�E�H�@H�H�E�H�U�H�E�H��H���c0��H� H�E�H�E�H���'!��H�E�H�E�H��uH��K ��   H�5�" H�=�" �����H�E�H�PH�E�H�H�E�H��H���A��H�E�H� H������H�U�H�E�H�H�E�H�U�H�PH�E�H�PH�E�H�@H9�rH�+K ��   H�5\" H�=�" �Q�����ÐUH��H��H�}����E�H�E�H�������H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P���UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���k���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E��@]�UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=
$ ��־�H��x���� <%uH�E��%   H����  H��x����  H�E�H���1���H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�# �K־��H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�# �־��u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�# �վ��*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�# �qվ������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�# �&վ�������E���tH��    H��uH�=#$ ��Ծ��E���tH��    H��uH�=a$ ��Ծ�H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=�$ �Ծ�H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=0$ ��Ӿ�돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=6$ �Ӿ�H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=D$ �gӾ�H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H���������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�# �Ҿ�H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�# �MҾ��H�U�H�E�H��H���"  H�E�H�U�H��H��H����  H�E�H��������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=�# ��Ѿ�H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�# �Ѿ��N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�# �7Ѿ�H�U�H�E�H��H���$���H��x���� ���M�H�U�H�E�H���<  H�E�H������H��x���H�E�H���x����g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�= ��Ͼ�H��x���� <%uH�E��%   H����  H��x����  H�E�H���;���H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=� �UϾ��H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=� �Ͼ��u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=� ��ξ��*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=  �{ξ������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�= �0ξ�������E���tH��    H��uH�=- �ξ��E���tH��    H��uH�=k ��;�H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=� �;�H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=: ��̾�돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=@ �̾�H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=N �q̾�H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H���������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=� ��˾�H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=� �W˾��H�U�H�E�H��H���,  H�E�H�U�H��H��H����  H�E�H��������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=� ��ʾ�H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=� �ʾ��N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=� �Aʾ�H�U�H�E�H��H���.���H��x���� ���M�H�U�H�E�H���p  H�E�H������H��x���H�E�H�������g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���I  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�= ��Ⱦ�H��x���� <%uH�E��%   H���  H��x����  H�E�H���E���H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=� �_Ⱦ��H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=  �Ⱦ��u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�= ��Ǿ��*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=
 �Ǿ������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�= �:Ǿ�������E���tH��    H��uH�=7 �Ǿ��E���tH��    H��uH�=u ��ƾ�H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=� �ƾ�H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=D �ƾ�돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=J �ž�H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=X �{ž�H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���	  H�E�H�U�H��H��H����	  H�E�H���������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=� ��ľ�H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=� �aľ��H�U�H�E�H��H���6	  H�E�H�U�H��H��H����  H�E�H�������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=� ��þ�H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=� �þ��N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=� �Kþ�H�U�H�E�H��H���8���H��x���� ���M�H�U�H�E�H���  H�E�H������H��x���H�E�H�������g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���}  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=( �����H��x���� <%uH�E��%   H���P  H��x����  H�E�H���O���H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=� �i����H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=
 �%����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�= ������*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�= ���������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�= �D���������E���tH��    H��uH�=A �����E���tH��    H��uH�= �����H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=� 輿��H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=N ����돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=T �Ǿ��H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=b 腾��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H���������   �E�    H��x���� </~H��x���� <9~H��    H��uH�= �ڽ��H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=� �k����H�U�H�E�H��H���@  H�E�H�U�H��H��H����  H�E�H�������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=� �꼾�H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=� 襼���N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=� �U���H�U�H�E�H��H���B���H��x���� ���M�H�U�H�E�H����  H�E�H������H��x���H�E�H�������g������UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H��������ÐUH��H��H�}����E�H�E�H� �U��H���0�����ÐUH��SH��H�}�H�u�H�E�H���#���H�E��@H�E�H���c�����H�E�H�ƿ   �������H��[]�UH��H��H�}�H�u�H�U�H�E�H��H���  H�E��ÐUH��SH��H�}�H�u�H�E�H������H�E��@H�E�H��������H�E�H�ƿ   �c�����H��[]�UH��SH��(  H��������H��������������������������E��3�   ��H��    H��, �H�H��, H���H������H�XH������H������H��H���G���������H������H� ������H������I��H����  H������H�������  H������H�XH������H�����H��H�������������H������H� ������H�����I��H���c  H�����H���B����  H������H�XH������H��0���H��H������������H������H� ������H��0���I��H���#  H��0���H��������C  H�������@��tH�
* �*   H�5� H�=� ����H�������@��tH��) �+   H�5p H�=v �e���H�������@��tH��) �,   H�5B H�=[ �7���H�������@��tH��) �-   H�5 H�=C �
��������� tH�Y) �.   H�5� H�=6 �����H������H��H���r�����tH�#) �/   H�5� H�=, ����H������H�H���C � ��藎  H��H��������  ������ tH��( �3   H�5e H�=� �Z���H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ºC H��H���r���H��P���H�5n H������H����������H���Ԗ��H�5s H���o���H������H��P���H���L���H��' �;   H�5�  H�=A �~����H��(  []�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���p�����ÐUH��H��H�}����E�H�E�H� �U��H��������ÐUH��SH��(  H��������H��������������������������E��3�   ��H��    H�z) �H�H�n) H���H������H�XH������H������H��H������������H������H� ������H������I��H���   H������H���y����  H������H�XH������H�����H��H������������H������H� ������H�����I��H���=,  H�����H�������  H������H�XH������H��0���H��H���[���������H������H� ������H��0���I��H���3  H��0���H�������C  H�������@��tH��% �*   H�5t�  H�=i	 �i���H�������@��tH��% �+   H�5F�  H�=L	 �;���H�������@��tH��% �,   H�5�  H�=1	 ����H�������@��tH�o% �-   H�5��  H�=	 ����������� tH�G% �.   H�5��  H�=	 ����H������H��H���H�����tH�% �/   H�5��  H�=	 ����H������H�H���C � ���m�  H��H���4����  ������ tH��$ �3   H�5;�  H�=� �0���H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ºC H��H���H���H��P���H�5D H���h���H����������H��誒��H�5I H���E���H������H��P���H���"���H��# �;   H�5_�  H�= �T����H��(  []�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H��������ÐUH��H��H�}����E�H�E�H� �U��H���8�����ÐUH��SH��(  H��������H��������������������������E��3�   ��H��    H� & �H�H�& H���H������H�XH������H������H��H�������������H������H� ������H������I��H���0  H������H���O����  H������H�XH������H�����H��H������������H������H� ������H�����I��H���<  H�����H��������  H������H�XH������H��0���H��H���1���������H������H� ������H��0���I��H���kC  H��0���H�������C  H�������@��tH��! �*   H�5J�  H�=? �?���H�������@��tH��! �+   H�5�  H�=" ����H�������@��tH��! �,   H�5��  H�= �����H�������@��tH�U! �-   H�5��  H�=� ���������� tH�-! �.   H�5��  H�=� ����H������H��H��������tH��  �/   H�5c�  H�=� �X���H������H�H���C � ���C�  H��H�������  ������ tH��  �3   H�5�  H�=Z ����H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ºC H��H������H��P���H�5 H���>���H����������H��耎��H�5 H������H���e���H��P���H�������H�� �;   H�55�  H�=� �*����H��(  []�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���D�����ÐUH��H��H�}����E�H�E�H� �U��H���z�����ÐUH��SH��(  H��������H��������������������������E��3�   ��H��    H��" �H�H��" H���H������H�XH������H������H��H�������������H������H� ������H������I��H���g@  H������H���%����  H������H�XH������H�����H��H���h���������H������H� ������H�����I��H����K  H�����H��������  H������H�XH������H��0���H��H������������H������H� ������H��0���I��H���ES  H��0���H���c����C  H�������@��tH�� �*   H�5 �  H�= ����H�������@��tH�� �+   H�5��  H�=�  �����H�������@��tH�� �,   H�5��  H�=�  ����H�������@��tH�[ �-   H�5��  H�=�  ���������� tH�3 �.   H�5o�  H�=�  �d���H������H��H���������tH�� �/   H�59�  H�=�  �.���H������H�H���C � ����  H��H�������  ������ tH�� �3   H�5��  H�=0  �����H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ºC H��H�������H��P���H�5��  H������H����������H���V���H�5��  H�������H���;���H��P���H�������H�� �;   H�5�  H�=��  � ����H��(  []�UH��SH��(H�}�H�u�H�E��@��t$H�E��@��tH�U�H�E�H��H���Q  �   H�E��@��tAH�E��@����t2H�E�H�������E�H�E�H��������H�E�H�ƿ   ������KH�E��@����t<H�E��@��t0H�E�H��������E�H�E�H��������H�E�H�ƿ   �6����H�E�H�PH�E�H��H��H���P  �H��([]�UH��H��H�}�H�E��@����tH��    H��uH�=� �K���H�E���UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=� �ר��H��x����@��tH��    H��uH�=� 讨��H��x����@��tH��    H��uH�= 腨��H��x����@��tH��    H��uH�=J �]���H�E�H�5� H���0���H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���dO  �  H��x����@��tH��    H��uH�= �Ƨ��H��x����@��tH��    H��uH�=R 蝧��H��x����@��tH��    H��uH�=� �t����}� tH��    H��uH�=� �T���H��x���H��H���]�����tH��    H��uH�= �#����E�    H��x����@��9E�}H�E��    H�������E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H���P����?  H��x����@��tH��    H��uH�=� 脦��H��x����@��tH��    H��uH�=  �[����}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH� H�E�H�U�H�E�H��H����L��H�E�H���aW���E�H��x���H��H���������t!H��x���H��H���>���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H��������E�뽋E�E�H��x����@9E���  H�E��    H�������E��֋E�E�H��x����@9E�}H�E��    H���~����E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H���,����E�뵃}�tH��    H��uH�=u �h���H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�� H�E�H�U�H�E�H��H����K  H�E�H���$L  �E�H��x���H��H��������t!H��x���H��H���U���� 9E�~�   ��    ��tH��x���H��H���+���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H��������E�뱋ẺE�H��x����@9E���   H�E��    H�������E��֋ẺE�H��x����@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���/����E��H��    H��uH�=  �q�������ÐUH��SH��H�}�H�u�H�E�H� H��H���b�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��� �����tH�E�H� H��H���M������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���	I  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���(�����tH�E�H� H��H���u������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���I  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���P�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���YG  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���������t&H�E�H� H��H���&���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���x�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����G  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H���O���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���E  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���)�����t&H�E�H� H��H���v���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���5F  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�� �H�H�� H���H�E��@��tH��    H��uH�=��  �圾�H�E��@��tH��    H��uH�=$�  远���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=��  �뛾�H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H���������t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���g�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���>C  �W  H�E��@��tH��    H��uH�=�  �ߚ��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���P����}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  �J���H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=��  �䙾�H�E��@��tH��    H��uH�=#�  辙��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�  �F���H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=�  �����H�E��@��tH��    H��uH�=O�  躘��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=��  �����H�E��@��tH��    H��uH�=+�  �֗��H�E�H��H��������tH��    H��uH�=]�  託���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���c@  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���9>  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����=  �   �}� tH��    H��uH�=G�  �2���H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���>  �H��    H��uH�=5�  谕�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5O�  H���F����H��    H��uH�=9�  �D������UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=��  �Ӕ��H��x����@��tH��    H��uH�=��  誔��H��x����@��tH��    H��uH�=�  联��H��x����@��tH��    H��uH�=F�  �Y���H�E�H�5��  H��薹��H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���o=  �  H��x����@��tH��    H��uH�=�  ���H��x����@��tH��    H��uH�=N�  虓��H��x����@��tH��    H��uH�=��  �p����}� tH��    H��uH�=��  �P���H��x���H��H���Y�����tH��    H��uH�=�  �����E�    H��x����@��9E�}H�E��    H�������E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H��謷���?  H��x����@��tH��    H��uH�=��  耒��H��x����@��tH��    H��uH�=��  �W����}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��  H�E�H�U�H�E�H��H����8��H�E�H���]C���E�H��x���H��H��������t!H��x���H��H���:���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���6����E�뽋E�E�H��x����@9E���  H�E��    H�������E��֋E�E�H��x����@9E�}H�E��    H���ڵ���E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H��舵���E�뵃}�tH��    H��uH�=q�  �d���H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH���  H�E�H�U�H�E�H��H����7  H�E�H��� 8  �E�H��x���H��H��������t!H��x���H��H���Q���� 9E�~�   ��    ��tH��x���H��H���'���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���=����E�뱋ẺE�H��x����@9E���   H�E��    H�������E��֋ẺE�H��x����@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H��苳���E��H��    H��uH�=
�  �m�������ÐUH��SH��H�}�H�u�H�E�H� H��H���^�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���I������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���7  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��腵����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���$�����tH�E�H� H��H���q������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���37  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��讴����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���L�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���d5  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���ճ����t&H�E�H� H��H���"���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���t�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���5  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���������t'H�E�H� H��H���K���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��蜲����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���3  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���%�����t&H�E�H� H��H���r���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���ı����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����3  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�4�  �H�H�(�  H���H�E��@��tH��    H��uH�=��  �ሾ�H�E��@��tH��    H��uH�= �  軈���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=��  �燾�H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H���������t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���c�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H����0  �W  H�E��@��tH��    H��uH�=�  �ۆ��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H��謫���}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  �F���H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=��  �����H�E��@��tH��    H��uH�=�  躅��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�  �B���H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=�  �܄��H�E��@��tH��    H��uH�=K�  趄��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=��  �����H�E��@��tH��    H��uH�='�  �҃��H�E�H��H���ޫ����tH��    H��uH�=Y�  褃���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���.  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���D,  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����+  �   �}� tH��    H��uH�=C�  �.���H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���=,  �H��    H��uH�=1�  謁�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5K�  H��謦���H��    H��uH�=5�  �@������UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=��  �π��H��x����@��tH��    H��uH�=��  覀��H��x����@��tH��    H��uH�=
�  �}���H��x����@��tH��    H��uH�=B�  �U���H�E�H�5��  H���>���H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���+  �  H��x����@��tH��    H��uH�=�  ���H��x����@��tH��    H��uH�=J�  ���H��x����@��tH��    H��uH�=��  �l���}� tH��    H��uH�=��  �L��H��x���H��H���U�����tH��    H��uH�= �  ����E�    H��x����@��9E�}H�E��    H��豢���E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H���j����?  H��x����@��tH��    H��uH�=��  �|~��H��x����@��tH��    H��uH�=��  �S~���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��  H�E�H�U�H�E�H��H����$��H�E�H���Y/���E�H��x���H��H��������t!H��x���H��H���6���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H��������E�뽋E�E�H��x����@9E���  H�E��    H���Ġ���E��֋E�E�H��x����@9E�}H�E��    H��蘠���E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H���F����E�뵃}�tH��    H��uH�=m�  �`|��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH���  H�E�H�U�H�E�H��H����#  H�E�H���$  �E�H��x���H��H��� �����t!H��x���H��H���M���� 9E�~�   ��    ��tH��x���H��H���#���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H��������E�뱋ẺE�H��x����@9E���   H�E��    H���˞���E��֋ẺE�H��x����@9E�}H�E��    H��蟞���E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���I����E��H��    H��uH�=�  �iz������ÐUH��SH��H�}�H�u�H�E�H� H��H���Z�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���E������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���$  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��聡����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��� �����tH�E�H� H��H���m������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����$  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��誠����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���H�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���#  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���џ����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���p�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���!#  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���������t'H�E�H� H��H���G���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��蘞����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���R!  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���!�����t&H�E�H� H��H���n���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���q!  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H���  �H�H���  H���H�E��@��tH��    H��uH�=��  ��t��H�E��@��tH��    H��uH�=�  �t���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=��  ��s��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��輛����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���_�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���z  �W  H�E��@��tH��    H��uH�=�  ��r��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���j����}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  �Br��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=��  ��q��H�E��@��tH��    H��uH�=�  �q��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�  �>q��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=�  ��p��H�E��@��tH��    H��uH�=G�  �p��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=��  ��o��H�E��@��tH��    H��uH�=#�  ��o��H�E�H��H���ڗ����tH��    H��uH�=U�  �o���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���p  �   �}� tH��    H��uH�=?�  �*n��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H����  �H��    H��uH�=-�  �m�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5G�  H���T����H��    H��uH�=1�  �<m�����UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=��  ��l��H��x����@��tH��    H��uH�=��  �l��H��x����@��tH��    H��uH�=�  �yl��H��x����@��tH��    H��uH�=>�  �Ql��H�E�H�5��  H��趓��H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���  �  H��x����@��tH��    H��uH�=�  �k��H��x����@��tH��    H��uH�=F�  �k��H��x����@��tH��    H��uH�=}�  �hk���}� tH��    H��uH�=��  �Hk��H��x���H��H���Q�����tH��    H��uH�=��  �k���E�    H��x����@��9E�}H�E��    H�������E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H���ґ���?  H��x����@��tH��    H��uH�=��  �xj��H��x����@��tH��    H��uH�=��  �Oj���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH� �  H�E�H�U�H�E�H��H������H�E�H���U���E�H��x���H��H��������t!H��x���H��H���2���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���\����E�뽋E�E�H��x����@9E���  H�E��    H���,����E��֋E�E�H��x����@9E�}H�E��    H��� ����E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H��讏���E�뵃}�tH��    H��uH�=i�  �\h��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH���  H�E�H�U�H�E�H��H����  H�E�H���  �E�H��x���H��H���������t!H��x���H��H���I���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���c����E�뱋ẺE�H��x����@9E���   H�E��    H���3����E��֋ẺE�H��x����@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H��豍���E��H��    H��uH�=�  �ef������ÐUH��SH��H�}�H�u�H�E�H� H��H���V�����t'H�E�H� H��H��裼��� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���A������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���P  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���}�����t&H�E�H� H��H���ʻ��� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���i������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���o  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��覌����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���D�����tH�E�H� H��H��葺�����   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���͋����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���l�����tH�E�H� H��H��蹹�����   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���������t'H�E�H� H��H���C���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��蔊����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H����  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H���j���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��載����tH�E�H� H��H���	������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�4�  �H�H�(�  H���H�E��@��tH��    H��uH�=޾  ��`��H�E��@��tH��    H��uH�=�  �`���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=��  ��_��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��踇����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���[�����tH�E�H��H��諵�����   H�E��PH�u�H�E�A��A�ȉѺ
   H���  �W  H�E��@��tH��    H��uH�=�  ��^��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���҅���}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=ӽ  �>^��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=ݽ  ��]��H�E��@��tH��    H��uH�=�  �]��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  �:]��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=	�  ��\��H�E��@��tH��    H��uH�=C�  �\��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=�  ��[��H�E��@��tH��    H��uH�=�  ��[��H�E�H��H���փ����tH��    H��uH�=Q�  �[���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���=	  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �   �}� tH��    H��uH�=;�  �&Z��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���y  �H��    H��uH�=)�  �Y�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5C�  H���̀���H��    H��uH�=-�  �8Y�����UH��H�� H�}�H�u�H�E�H�������E�H�E�H��������H�E�H�E�H���������H�E�����UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�E�H��������E�H�E�H���������H�E�H�E�H��������H�E�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H����ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�@H��    H�E�HЋ ��tH�E�H�@H�PH�E�H�P�͐]ÐUH��H�}�H�E�H�@]�UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H����  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���A  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����	  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���-  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H����
  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���6  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���"  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���+  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���~  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���   H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���s  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�֚  H�E��E�    �E���~H��    H��uH�=�  �CQ���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=ƺ  ��P���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H�������� �U�)�9E�����t�U�H�E���H���s���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����r���E��ڋE����E�}� x!�E�H��D���H�E���H���r���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�.�  H�E��E�    �E���~H��    H��uH�=@�  �O���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  �)O���E��P�U�H��D�-H�U�H�E�H��H���?���� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���Yq���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���"q���E��ڋE����E�}� x!�E�H��D���H�E���H����p���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  ��M���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�  �M���E��P�U�H��D�-H�U�H�E�H��H��蠂��� 9E�����tE�E�    H�U�H�E�H��H���z���� �U�)�9E�����t�U�H�E���H���o���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���o���E��ڋE����E�}� x!�E�H��D���H�E���H���So���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=��  �TL���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=׵  ��K���E��P�U�H��D�-H�U�H�E�H��H�������� 9E�����tE�E�    H�U�H�E�H��H���Ҁ��� �U�)�9E�����t�U�H�E���H���n���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����m���E��ڋE����E�}� x!�E�H��D���H�E���H���m���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�?�  H�E��E�    �E���~H��    H��uH�=Q�  �J���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=/�  �:J���E��P�U�H��D�-H�U�H�E�H��H���P��� 9E�����tE�E�    H�U�H�E�H��H���*��� �U�)�9E�����t�U�H�E���H����n���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���n���E��ڋE����E�}� x!�E�H��D���H�E���H���cn���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  �I���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �H���E��P�U�H��D�-H�U�H�E�H��H���}��� 9E�����tE�E�    H�U�H�E�H��H���}��� �U�)�9E�����t�U�H�E���H���"m���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����l���E��ڋE����E�}� x!�E�H��D���H�E���H���l���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=�  �]G���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�  ��F���E��P�U�H��D�-H�U�H�E�H��H���	|��� 9E�����tE�E�    H�U�H�E�H��H����{��� �U�)�9E�����t�U�H�E���H���k���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���Lk���E��ڋE����E�}� x!�E�H��D���H�E���H���k���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�P�  H�E��E�    �E���~H��    H��uH�=b�  �E���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=@�  �KE���E��P�U�H��D�-H�U�H�E�H��H���az��� 9E�����tE�E�    H�U�H�E�H��H���;z��� �U�)�9E�����t�U�H�E���H����i���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���i���E��ڋE����E�}� x!�E�H��D���H�E���H���ti���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  �D���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �C���E��P�U�H��D�-H�U�H�E�H��H���x��� 9E�����tE�E�    H�U�H�E�H��H���x��� �U�)�9E�����t�U�H�E���H����f���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���f���E��ڋE����E�}� x!�E�H��D���H�E���H���f���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H� �  H�E��E�    �E���~H��    H��uH�=�  �mB���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  ��A���E��P�U�H��D�-H�U�H�E�H��H���w��� 9E�����tE�E�    H�U�H�E�H��H����v��� �U�)�9E�����t�U�H�E���H���Me���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���e���E��ڋE����E�}� x!�E�H��D���H�E���H����d���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�Y�  H�E��E�    �E���~H��    H��uH�=k�  ��@���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=Q�  �\@���E��P�U�H��D�-H�U�H�E�H��H���ru��� 9E�����tE�E�    H�U�H�E�H��H���Lu��� �U�)�9E�����t�U�H�E���H���c���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���wc���E��ڋE����E�}� x!�E�H��D���H�E���H���Gc���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=˨  �&?���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �>���E��P�U�H��D�-H�U�H�E�H��H����s��� 9E�����tE�E�    H�U�H�E�H��H���s��� �U�)�9E�����t�U�H�E���H���b���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����a���E��ڋE����E�}� x!�E�H��D���H�E���H���a���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=#�  �~=���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  �=���E��P�U�H��D�-H�U�H�E�H��H���"r��� 9E�����tE�E�    H�U�H�E�H��H����q��� �U�)�9E�����t�U�H�E���H����c���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���c���E��ڋE����E�}� x!�E�H��D���H�E���H���cc���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�i�  H�E��E�    �E���~H��    H��uH�={�  ��;���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=Y�  �d;���E��P�U�H��D�-H�U�H�E�H��H���zp��� 9E�����tE�E�    H�U�H�E�H��H���Tp��� �U�)�9E�����t�U�H�E���H���"b���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����a���E��ڋE����E�}� x!�E�H��D���H�E���H���a���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�  H�E��E�    �E���~H��    H��uH�=ԣ  �/:���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=��  ��9���E��P�U�H��D�-H�U�H�E�H��H����n��� 9E�����tE�E�    H�U�H�E�H��H���n��� �U�)�9E�����t�U�H�E���H���`���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���L`���E��ڋE����E�}� x!�E�H��D���H�E���H���`���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�"�  H�E��E�    �E���~H��    H��uH�=4�  �8���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  �8���E��P�U�H��D�-H�U�H�E�H��H���3m��� 9E�����tE�E�    H�U�H�E�H��H���m��� �U�)�9E�����t�U�H�E���H����^���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���^���E��ڋE����E�}� x!�E�H��D���H�E���H���t^���m��ِ��UH��H�}�H�u�H�E�H�E�H�E�H�E�H�E�� ��tH�E�H�PH�U��H�E�H�HH�M����H�E��  H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E�H;E�sH�E�H�PH�U��  H�E���H�E�]�UH��H��H�}�H�u�H�E�H���[n��H��H�E�H�H�E�H��H�������H�E���UH��H��@H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H���n��HE�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E��  H�E���UH��H�}�H�u�H�U�H�E�    H�E�H;E�sIH�U�H�E�H�� �E�H�U�H�E�H�� �E��E�:E�s�������E�:E�v�   �H�E�뭸    ]�UH��H�}�H�u�H�E�    H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H��H�}�H�u�H�U�H�E�H��H���k�����UH��H�}�H�u�H�U�H�E�    H�E�H;E�r�    �\H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H�� H�}�H�u�H�U�H�=�  �g   H�5��  H�=��  �^Z��UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s)H�U�H�E�H�� �U�8�uH�U�H�E�H��H�E��͸    ]�UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E��ă}� uH�U�H�E�H���    ]�UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H���N���H��t�   ��    ��tH�E��H�E����UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t=H�U�H�E�H�� ��H�E���H�������H������tH�U�H�E�H��H�E�뱸    ��UH��H�� H�}�u�H�E�H���?j��H�E�H�E�    H�E�H;E�w8H�E�H+E�H��H�E�H�� ��9E�uH�E�H+E�H��H�E�H��H�E�뾸    ��UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H������H��u�   ��    ��tH�E��H�E����UH��H�}�H�u�H�E�    H�U�H�E�H�� ����   �E�H�E�    H�U�H�E�H�� ��tGH�U�H�E�H�� ��t-H�U�H�E�H�H�E�H��H�M�H�E�H�� 8�t�E� ��H�E�맀}� tH�U�H�E�H��H�E��h����    ]�UH��H��0H�}�H�u�H�U�H�E�H��uH�ܫ  ��   H�50�  H�=e�  ��V��H�}� t
H�E�H�E��#H�E�H� H��tH�E�H� H�E��
�    �   H�E�� ��t$H�E�� ��H�E���H������H��t�   ��    ��tH�E���H�E�H�E�H�E�� ��t$H�E�� ��H�E���H���R���H��u�   ��    ��tH�E���H�E�� ��tH�E��  H�E�H�U�H��H��H�E�H�     H�E���UH��H��H�}�H�u�H�M�H�E�H��< H��H��������UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E���H�U�H�E�H�]�UH��H��H�}�H�u�H�@�  ��   H�5��  H�=Ħ  �PU��UH��H��H�}�H�u�H��  ��   H�5\�  H�=��  �!U��UH��H��H�}�H�u�H��  ��   H�5-�  H�=f�  ��T��UH��H�� H�}�H�u��U�H�ǩ  ��   H�5��  H�=4�  ��T��UH��H�� H�}�H�u��U�H���  ��   H�5ɥ  H�=�  �T��UH��H�� H�}�H�u��U�H�s�  ��   H�5��  H�=Х  �\T��UH��H�� H�}�H�u��U�H�I�  ��   H�5e�  H�=��  �*T��UH��H��H�}�H�u�H�#�  ��   H�56�  H�=o�  ��S��UH��H�� H�}�H�u�H�U�H���  ��   H�5�  H�=<�  ��S��UH��H�� H�}�H�u�H�U�H�̨  ��   H�5Ф  H�=	�  �S��UH��H�� H�}�H�u�H�U�H���  ��   H�5��  H�=֤  �bS��UH��H��H�}�H�u�H�{�  ��   H�5n�  H�=��  �3S��UH��H�� H�}�H�u�H�U�H�O�  ��   H�5;�  H�=t�  � S��UH��H��H�}�H�u�H�(�  ��   H�5�  H�=E�  ��R��UH��H��H�}�H�u�H��  ��   H�5ݣ  H�=�  �R��UH��H�� H�}�H�u�H�U�H�֧  ��   H�5��  H�=�  �oR��UH��H�� H�}�H�u�H�U�H���  ��   H�5w�  H�=��  �<R��UH��H�� H�}�H�u�H�U�H���  ��   H�5D�  H�=}�  �	R��UH��H��H�}��u�H�Z�  ��   H�5�  H�=O�  ��Q��UH��H��H�}�H�u�H�3�  ��   H�5�  H�= �  �Q��UH��H��H�}�H�u�H��  ��   H�5��  H�=�  �}Q��UH��H��H�}��u�H��  ��   H�5��  H�=â  �OQ��UH��H��H�}�H�u�H���  ��   H�5[�  H�=��  � Q��UH��H��H�}�H�u�H���  ��   H�5,�  H�=e�  ��P��UH��H�� H�}�H�u�H�U�H�k�  ��   H�5��  H�=2�  �P��UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s6H�E�H��    H�E�HЋ 9E�uH�E�H��    H�E�H��H�E����    ]�UH��H��H�}�H��  �  H�5h�  H�=��  �-P��UH��H�� H�}��u�H�U�H���  �  H�56�  H�=o�  ��O��UH��}�E�-�  ��C�  ��H��    H���  �H�H�y�  H���H�Q�  H�E���   H�`�  H�E���   H�h�  H�E���   H�t�  H�E���   H���  H�E��   H���  H�E��   H���  H�E��   H���  H�E��   H���  H�E��sH���  H�E��fH�ҡ  H�E��YH��  H�E��LH��  H�E��?H� �  H�E��2H�4�  H�E��%H�;�  H�E��H�I�  H�E��H�^�  H�E�H�E�]�UH��H��0�}�H�u�H�U؋E������H�E�H�U�H�M�H�E�H��H������H�E�H���`��H9E�����t�   ��    ��UH��H�� H�}�H�u�H�U�H�U�H�M�H�E�H��H����^��H��H�E�H���UH��H�� H�}�H�u�H�E�H���_��H�E�H�E�H�PH�M�H�E�H��H���^��H�U�H�E�H���UH��H��0�}�H�u�H�U�H�M�H�u�H�U��E�H�H�M�A�    I��H�ƿ   �vK���E�Hc�H�E�H�H�E�H� H���u�������    ��UH��H��0�}�H�u�H�U�H�M�H�u�H�U��E�H�H�M�A�    I��H�ƿ   �K���E����u�������E�Hc�H�E�H��    ��UH��H��0�}�H�u��U�H�M�H�u��E�Hc�H�U��E�H�A�    I��H�ƿ   �J��H�E�H�E�H�}��u������H�E�H�U�H��    ��UH��H��0H�}�u�H�U�H�U�H�E�A�    A�    �    H�ƿ   �MJ���E���u�������U�H�E؉�    ��UH��H���}��E�H�A�    A�    �    �    H�ƿ   ��I���    ��UH��H�� H�}�u�H�U��M�H�E��H���K����E���t�E��������    ��   ��UH��H����2 ������t-H�=�2 �J  ������tH�=�2 �u  H�=�2 �s  ��4 ������t<H�=�4 �  ������t'H�=�2 �d  H��H�=�2 �q  H�=`4 �'  �d4 ������tDH�=T4 ��  ������t/H�=g2 �  H�E�H�E�H��H�= 4 �  H�=4 ��  H�=4 ��  �ÐUH��H�� H�}�H�u�H�U�H�E�H��H���I��������tH���  �   H�5a�  H�=��  �J��H�E��ÐUH��H�� H�}�H�u�H�U�H�E�H�U�H��H���DI��������tH���  �!   H�5�  H�=\�  �HJ�����UH��H�}�H�E��     �]ÐUH��H��H�}�H�E�H����   H�E�H�ƿ   �L�����UH��H�}�H�E�]�UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H���   H�E�H�������H��H�E�H�ƿ�  ��K��H��H���   �H��[]�UH��H�}�H�E�]�UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H����   H�E�H�������H�H�E�H�ƿ   �VK��H��H����   �H��[]�UH��H�}�H�E�]�UH��H�}�H�E��  �]�UH��H�}�H�E�H�Ƹ    �9   H��H���H��]ÐUH��ATSH��H�}�H�u�H�E�H�U�H�H�E�H��H���r���H�E�H��H���n   H�E�H�@     H�E�H��(�   I��H��xL���i   I�� H����H��[A\]ÐUH��H�}�H�E�H�     �]�UH��H�}�H�u�H�E�H�U�H��]�UH��H��H�}�H�E�H���N   H�}�:   ���UH��H��H�}�H�E�H������H�E�H�@    H�E�H��H���$   ���UH��H�}�]ÐUH��H�}�H�E�H�     �]�UH��H��H�}�H�E�H���   H�}�������UH��H�}�H�E�H�     �]�UH��H�}�H����B H�PH�E�H��]ÐUH��H��H�}�H�E�H�������H�E��   H����B����UH���f0 ������tJH�=V0 �  ������t5H�=10 ��  H�=50 ��  H�y H�50 H����A H����F��H��/ ]�UH��H�}��u�H�U�U�H�E��    ]�UH��H��/ ]�UH��H�}����E�ЈE�H����B H�PH�E�H�H�E��U�PH�E��U��P	�]ÐUH��H�}�H�E��     H�E��@    �]�UH��H�}�H�E�� ]�UH��H�}�H�E��@]ÐUH��H�� H�}�H�u�H�E�H� � �E�H�E� ����   �E���x�U�H�E�P�-  �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    �   �E�%�   =�   t/�E�%�   =�   tH���  �'   H�5��  H�=��  �E���   �q�E�%�   =�   tH���  �,   H�5]�  H�=Λ  ��D��H�E�@�����E���?	�H�E�PH�E� �P�H�E�H�E�H� H�PH�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�E�H� � �E��}�vH���  �>   H�5Ӛ  H�=l�  �XD��H�E�H� �U��H�E�H� H�PH�E�H�H�E�H� H�PH�E�H��    ��UH��H��H�}�H�E��    �   H���X���H��h�B H�PH�E�H���ÐUH��H��H�}�H��h�B H�PH�E�H�H�E�H���<�����ÐUH��H��H�}�H�E�H������H�E��   H���/?���ÐUH��SH��XH�}�H�u�H�U�H�M�H�E�� f��tH�L�  �W   H�5ƙ  H�=��  �KC��H�E�H�PH� H�E�H�U�H�E�H�������H�E�H���  ��tH�E�H���  ��t�   ��    ����   H�U�H�E�H��H�������E�}� t�E��   H�E�H������������t�H�U�H�E�H�H�E�H���o���������t�    �MH�E�H�H�E�H���L����H�E�H� H�PH�E�H��@���H�E�H������������t�   ��    H��X[]ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH��  �s   H�5{�  H�=T�  � B��H�E�H�PH� H�E�H�U�H�E�H���x���H�E�H���F  ��tH�E�H���v  ��t�   ��    ����   H�U�H�E�H��H���s����E��}� t�E��   H�E�H���4���������t�H�U�H�E�H�H�E�H���$���������t�    �OH�E�H��������H�E�H� �H�E�H� H�PH�E�H��>���H�E�H�������������t�   ��    �ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH�w�  ��   H�53�  H�=�  �@��H�E�H�PH� H�E�H�U�H�E�H���0���H�E�H�     H�E�H����  ��ttH�U�H�E�H��H���D����E��}� t�E��tH�E�H������������t�H�U�H�E�H�H�E�H�������������t�    �8H�E�H� H�PH�E�H��|���H�E�H������������t�   ��    ��UH��H��`H�}�H�u�H�U�H�M�H�E�� f��tH�3�  ��   H�5�  H�=��  �?��H�E�H�PH� H�E�H�U�H�E�H���V  ��tH�E�H���f  ��t�   ��    ����   H�E�H� � �E؋E؅�u
�    �   H�E�H�E�H�E�H��H�E�H�U�H�M�H�E�H��H���x����E��}�tY�}� t�E��pH�U�H�E�H9�tH�d�  ��   H�5P�  H�=8�  ��>��H�E�H� H�PH�E�H�H�U�H�E�H��"��������H�U�H�E�H� H9�t�   ��    ��UH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}��   ]ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t2��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ºC H��H����A��H��`���H�5H�  H����A��H���6B��H��`���H����A���    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t ��T���/v��T���9w�   �[�    �T��T���vFH��`���H�ºC H��H���A��H��`���H�5ޔ  H���2A��H���|A��H��`���H���A���    ��UH��H��   H��X�����T�����T���wH��X���H���:�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���fv��T���@v��T���Fw�   �[�    �T��T���vFH��`���H�ºC H��H���4@��H��`���H�5P�  H���T@��H���@��H��`���H���1@���    ��UH��H��   H��X�����T�����T���wH��X���H���\�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ºC H��H���V?��H��`���H�5  H���v?��H����?��H��`���H���S?���    ��UH��H��   H��X�����T�����T���wH��X���H���~�����t�   ��    ���r  ��T���!�W  ��T���"�J  ��T���#�=  ��T���$�0  ��T���%�#  ��T���&�  ��T���'�	  ��T���(��   ��T���)��   ��T���*��   ��T���+��   ��T���,��   ��T���-��   ��T���.��   ��T���/��   ��T���:��   ��T���;��   ��T���<t~��T���=tu��T���>tl��T���?tc��T���@tZ��T���[tQ��T���\tH��T���]t?��T���^t6��T���_t-��T���`t$��T���{t��T���|t��T���}t	��T���~u�   �[�    �T��T���vFH��`���H�ºC H��H���F=��H��`���H�5�  H���f=��H���=��H��`���H���C=���    ��UH��H��   H��X�����T�����T���wH��X���H���n�����t�   ��    ��t ��T��� v��T���~w�   �[�    �T��T���vFH��`���H�ºC H��H���<��H��`���H�5��  H���<��H����<��H��`���H���<���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T��� t	��T���	u�   �n�    �g��T���vYH��`���H�ºC H��H����;��H��`���H�5.�  H����;��H��T�����H���	<��H���)<��H��`���H���;���    �ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��tD��T��� t-��T���	t$��T���
t��T���t��T���t	��T���u�   �[�    �T��T���vFH��`���H�ºC H��H����:��H��`���H�5��  H��� ;��H���J;��H��`���H����:���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���v��T���~w�   �[�    �T��T���vFH��`���H�ºC H��H���&:��H��`���H�5"�  H���F:��H���:��H��`���H���#:���    ��UH��H��   H��X�����T�����T���wH��X���H���N�����t�   ��    ��t ��T���`v��T���zw�   �[�    �T��T���vFH��`���H�ºC H��H���l9��H��`���H�5h�  H���9��H����9��H��`���H���i9���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ºC H��H���8��H��`���H�5��  H����8��H���9��H��`���H���8���    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t��T���@v��T���Zw��T����� �U��T���vFH��`���H�ºC H��H����7��H��`���H�5G�  H���8��H���e8��H��`���H����7����T�����UH��H��   H��X�����T�����T���wH��X���H���"�����t�   ��    ��t��T���`v��T���zw��T����� �U��T���vFH��`���H�ºC H��H���C7��H��`���H�5ߍ  H���c7��H���7��H��`���H���@7����T�����UH��H�� ]ÐUH��H��H�}�H�u�H�E�H���F1����ÐUH��H��H�}�H�u�H�E�H���&1���W1���UH��H�� H�}��E�    H�E�H�pH�U���   ��������u�
��uH�=��  ��0�����UH��H�}�H�E�H���    ��]�UH��H��   H��`���H�»C H��H���5��H��`���H�5b�  H���5��H��H�EH��H���   H����5��H��`���H���m5�����UH��H�� H�}�H�E�H�E�H�E�H������H�E�� ������tH�E�H���D����    ��   ��UH��H��H�}�H�E�H�E�H�E��   �H�E�H���������UH��H��H�}�H�u�H�U�H�E�H��H���   H�E���UH��H��0H�}�H�u�H�E�H����2��H�E�H� H�U�H�M�H��H���   H�E�H���3�����UH��H��`H�}�H�u�H�U�H�E�H�5V�  H���_8��H�E�H���2��H�E�H�M�   H��H����V��H�E�H�U�H�M�H��H���   H�E�H���63��H�E�H���*3�����UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���Z   �UH�E�� ��t%H�E�� ��tH��    H��uH�=�  �	��H�u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���   H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�s�  H�E��E�    �E���~H��    H��uH�=��  �E���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �����E��P�U�H��D�-H�U�H�E�H��H����<��� 9E�����tE�E�    H�U�H�E�H��H����<��� �U�)�9E�����t�U�H�E���H����<���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���<���E��ڋE����E�}� x!�E�H��D���H�E���H���`<���m��ِ��D  H�9�  H���t3UH��S�P�B H��D  ��H��H�H���u�H��[]�f.�     ��J���         r close.bmp /shell.lef /dev/mouse0               0123456789abcdef       ../sysdeps/lemon/generic/lemon.cpp !(size & 0xFFF) libc panic!          sys_anon_allocate        0123456789abcdef  In function  , file  : 
 __ensure( ) failed  ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!        0123456789abcdef       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    ../options/ansi/generic/stdlib-stubs.cpp *string != '+' !negative !"Not implemented" mlibc: srandom() is a no-op i == j !"decode_wtranscode() errors are not handled" mlibc: Broken mbtowc() called wc mbs max_size *mbs MLIBC_DEBUG_MALLOC mlibc (PID ?): free() on    mlibc (PID ?): malloc() returns  mlibc (PID ?): realloc() on   returns  !(reinterpret_cast<uintptr_t>(p) & (align - 1)) ../options/internal/include/mlibc/strtofp.hpp   !"hex numbers in strtofp are unsupported"       ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:348: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:365: Assertion 'fra->type == frame_type::large' failed!       ../subprojects/frigg/include/frg/slab.hpp:366: Assertion 'address == fra->address' failed! 0x   ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       strtofp strtofp strtofp strtol rand_r abort     at_quick_exit   quick_exit system mktemp        bsearch abs labs llabs ldiv lldiv mblen mbtowc wctomb   mbstowcs        wcstombs lock   posix_memalign  strtod_l              $@       �           A               �                   �@                            @        0123456789abcdef       ../options/internal/include/mlibc/charcode.hpp nseq.it == nseq.end wseq.it == wseq.end alnum alpha blank cntrl digit graph lower print punct space upper xdigit mlibc: wctype(" ") is not supported     ../options/ansi/generic/ctype-stubs.cpp !"Not implemented"      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       promote iswctype        towlower        towupper                ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"  0123456789abcdef  mlibc: environment string "     " does not contain an equals sign (=)   ../options/ansi/generic/environment.cpp environ == vector.data() !vector.back() ../options/ansi/generic/environment.cpp:84: Assertion 'k != size_t(-1)' failed! vector.size() >= 2 && !vector.back() s != size_t(-1)    !"Environment strings need to contain an equals sign" mlibc: environment variable " " contains an equals sign %s=%s     asprintf(&string, "%s=%s", name, value) > 0 string      ../subprojects/frigg/include/frg/string.hpp:72: Assertion 'from + size <= _length' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{     ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed! lock     assign_variable unassign_variable getenv putenv setenv           0123456789abcdef       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    mlibc warning: File is not flushed before destruction   ../options/ansi/generic/file-io.cpp max_size    mlibc: Cannot read-write to same pipe-like stream __offset < __valid_limit __dirty_begin == __dirty_end io_size > 0 && "io_write() is expected to always write at least one byte" __offset < __buffer_size chunk __offset       __dirty_begin == __dirty_end && "update_bufmode() must only be called before performing I/O"    whence == SEEK_SET || whence == SEEK_END _type != stream_type::unknown  _bufmode != buffer_mode::unknown        _type == stream_type::pipe_like __io_offset == __dirty_begin hit io_seek() error  __offset == __valid_limit __buffer_size       mlibc warning: File is not flushed before closing       Library function fails due to missing sysdep    mlibc: sys_isatty() failed while determining whether stream is interactive      mlibc warning: Failed to flush file before exit() Illegal fopen() mode ' ' Illegal fopen() flag '       [31mmlibc: fdopen() ignores the file mode [39m        ../subprojects/frigg/include/frg/list.hpp:104: Assertion 'element' failed!      ../subprojects/frigg/include/frg/list.hpp:106: Assertion '!h(borrow).in_list' failed!   ../subprojects/frigg/include/frg/list.hpp:107: Assertion '!h(borrow).next' failed!      ../subprojects/frigg/include/frg/list.hpp:108: Assertion '!h(borrow).previous' failed!  ../subprojects/frigg/include/frg/list.hpp:79: Assertion 'h(ptr).in_list' failed!        ../subprojects/frigg/include/frg/list.hpp:164: Assertion 'it._current' failed!  ../subprojects/frigg/include/frg/list.hpp:165: Assertion 'h(it._current).in_list' failed!       ../subprojects/frigg/include/frg/list.hpp:170: Assertion '_back == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:173: Assertion 'h(traits::decay(next)).previous == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:179: Assertion 'traits::decay(_front) == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:183: Assertion 'traits::decay(h(previous).next) == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:188: Assertion 'traits::decay(erased) == it._current' failed! ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/slab.hpp:471: Assertion 'slb->contains(pointer)' failed!       ../subprojects/frigg/include/frg/slab.hpp:475: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:482: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:485: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed! lock read write unget update_bufmode seek     _init_type      _init_bufmode   _write_back _reset      _ensure_allocation              determine_bufmode               ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"  0123456789abcdef  ../options/ansi/generic/stdio-stubs.cpp new_buffer count < limit !"Not implemented"     Library function fails due to missing sysdep    a���o���~�������������������    Functionality is not implemented max_size > 0 
 %s:  %s
 returns:       mlibc: File locking (flockfile) is a no-op      mlibc: File locking (funlockfile) is a no-op    mlibc: File locking (ftrylockfile) is a no-op   mlibc: fread() I/O errors are not handled       mlibc: fwrite() I/O errors are not handled do_scanf: ' not implemented! do_scanf: m not implemented!    �������������������������������������������������������������������������������������a������������������������������������������������������������������������������������پ�����������'���������������r��������������������������������������������E������������������������������������������������������� �����������������������"���\�����������������������������������../subprojects/frigg/include/frg/formatting.hpp:200: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:213: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:217: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:221: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:225: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:229: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:235: Assertion '!opts.always_sign' failed!      ../subprojects/frigg/include/frg/formatting.hpp:236: Assertion '!opts.plus_becomes_space' failed!       ../subprojects/frigg/include/frg/formatting.hpp:240: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:247: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:254: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:258: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:262: Assertion '*s >= '0' && *s <= '9'' failed! ../subprojects/frigg/include/frg/formatting.hpp:266: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:275: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:279: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:286: Assertion '*s' failed! 0���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u�������u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���d���u�������u�������u���u���u���u�������u���u������u���u���u���u���u������?���a���a�������a���a���a���a���a���a���a���B�������a���a���a���a�������a���a���a���a���'�����������a���a�������a�������a���a���?���!opts.fill_zeros !opts.left_justify !opts.alt_conversion opts.minimum_width == 0    szmod == frg::printf_size_mod::default_size !opts.precision     [31mmlibc: Unknown printf terminator ' '[39m !"Illegal printf terminator"     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/optional.hpp:97: Assertion '_non_null' failed! ../subprojects/frigg/include/frg/formatting.hpp:299: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:300: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:301: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:302: Assertion 'opts.minimum_width == 0' failed! 0x     ../subprojects/frigg/include/frg/formatting.hpp:307: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:308: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:309: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:310: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:311: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:317: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:318: Assertion '!opts.alt_conversion' failed! (null)    ../subprojects/frigg/include/frg/formatting.hpp:341: Assertion 'szmod == printf_size_mod::long_size' failed!    (   n   u   l   l   )           ../subprojects/frigg/include/frg/formatting.hpp:364: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/formatting.hpp:374: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:375: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:384: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:396: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:413: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:419: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:420: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:432: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:437: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:438: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:454: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:455: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:456: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:470: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:477: Assertion '!"Unexpected printf terminal"' failed! %f       ../subprojects/frigg/include/frg/formatting.hpp:494: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{      ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! remove rename    renameat        tmpfile tmpnam  freopen setbuf scanf    operator() vscanf       operator()      operator()      vsscanf fwprintf        fwscanf vfwprintf       vfwscanf        swprintf        swscanf vswprintf       vswscanf        wprintf wscanf  vwprintf        vwscanf fgets fgetwc fgetws fputwc fputws fwide getwc   getwchar putwc  putwchar        ungetwc fgetpos fsetpos lock    getdelim        operator() expand       fgets_unlocked  ����������������������������������������������������������������������������������������������=�����������������������������������`�����������=���������=��������������������Y���Y���Y���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u���u�������u���u���u���u���u���u���u���u���u���u�����������Y���Y���Y���u�������u���u���u�������������������u���u�������u�������u���u�����������������������������������������������������������������������������������R�����������������������������������������������R�������������������R������������������S���R�����������������������R�����������R������������)���)���)���)���)���)���)���)���)���)���)���)���)���)���)���)�������)���)���)���)���)���)���)���)���)���)���K����������������)�������)���)���)���n�����������K���)���)���K���)�������)���)�������b�����������������������������������������������]�������������������]�����������������������c�����������������������F�����������^����������������������������� ����������� �����������������������������������b�����������������������������������]��������������]�����������������c�����������������F��������^���+��/��/��/��/��/��/��/��/��/��/��/���'��/��/��/��/���'��/��/��/��/��/���)��/��/��/��/��/���,��/��/���*��../options/ansi/generic/string-stubs.cpp !"Not implemented" m   Functionality is not implemented        Operation would block (EAGAIN) Access denied (EACCESS) Bad file descriptor (EBADF) File exists already (EEXIST) Access violation (EFAULT) Operation interrupted (EINTR) Invalid argument (EINVAL) I/O error (EIO)       Resource is directory (EISDIR)  No such file or directory (ENOENT) Out of memory (ENOMEM)       Expected directory instead of file (ENOTDIR)    Operation not implemented (ENOSYS)      Operation not permitted (EFAULT) Broken pipe (EPIPE) Seek not possible (ESPIPE) No such device or address (ENXIO) Unknown error code (?)    �\���]���]���]���\���]���\���]���]���]���]���]���]���]���]���]���]���\���\���]���]���]���]���\���\���\���]��]���]���]���]���]���]���]���]���]���]���]���]���]���]��]���]���]���]��&]���]���]���]��@]���]��3]���]���]���]���]���]��t]���]���]���]��M]��Z]���]���]���]���]��g]��    strxfrm strtok_r wcstod wcstof  wcstold wcstol  wcstoll wcstoul wcstoull wcscpy wcsncpy wmemcpy wmemmove wcscat wcsncat wcscmp  wcscoll wcsncmp wcsxfrm wmemcmp wcschr  wcscspn wcspbrk wcsrchr wcsspn wcsstr wcstok wcslen     wmemset         ../options/internal/generic/allocator.cpp       !mlibc::sys_anon_allocate(length, &ptr) !mlibc::sys_anon_free((void *)address, length) map unmap                 0123456789abcdef       ../options/internal/generic/charcode.cpp        (uc & 0b1100'0000) == 0b1000'0000 || (uc & 0b1111'1000) == 0b1111'1000  (uc & 0b1100'0000) == 0b1000'0000       wc <= 0x7F && "utf8_charcode cannot encode multibyte chars yet" !st.__progress cps.it == cps.end        encode_wtranscode       operator()              decode_wtranscode_length        operator()      decode_wtranscode decode         0123456789abcdef       mlibc: charset::is_alpha() is not implemented for the full Unicode charset      mlibc: charset::is_digit() is not implemented for the full Unicode charset      mlibc: charset::is_xdigit() is not implemented for the full Unicode charset     mlibc: charset::is_alnum() is not implemented for the full Unicode charset      mlibc: charset::is_punct() is not implemented for the full Unicode charset      mlibc: charset::is_graph() is not implemented for the full Unicode charset      mlibc: charset::is_blank() is not implemented for the full Unicode charset      mlibc: charset::is_space() is not implemented for the full Unicode charset      mlibc: charset::is_print() is not implemented for the full Unicode charset      mlibc: charset::to_lower() is not implemented for the full Unicode charset      mlibc: charset::to_upper() is not implemented for the full Unicode charset      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!  0123456789abcdef      0123456789abcdef      __cxa_guard_acquire contention  mlibc: Pure virtual function called from IP  0x ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!              zR x�        ̍��I    A�CD     <   ����2    A�Cm      \   �{��   A�C    |   �|���   A�C� $   �   G~���   A�CN�����   �   ����	   A�C      �   ����-    A�Ch         ����    A�CL         ����"    A�C]      @  ����-   A�C(    `  ����"    A�C]       �  �����    A�CE��      �  @����    A�C�     �  ы��>    A�Cy      �  ����-    A�Ch        ϋ��    A�CP      $  u���:    D u    <  ����0    D k    T  ����,    Dg    l  Ï��.    D i    �  ُ��.    D i    �  ���/    D j    �  ���(    D c    �  ���       (   �  ���S    B�A�A �d
ABA8     @����    B�B�A �A(�D0Y
(A ABBA     H  ���>    A�|      d  ���           x  ����    A�A��A      �  ~���"    A�HG PA     �  |���&    Da H   �  ����'   B�B�B �B(�A0�A8�D@8A0A(B BBB   X   $  e����   B�B�B �B(�A0�A8�D��T�a�W
8A0A(B BBBA   X   �  �����   B�B�B �B(�A0�A8�D��T�a�W
8A0A(B BBBA      �  ޔ��(    DS P  8   �  ����    B�B�B �A(�A0�|(A BBB  ,   4  :����    B�A�A ��AB         d  ����1    D l    |  ɕ��+    Df    �  ܕ��    DU    �  ޕ��    DU    �  ����    DI    �  ֕��    DI    �  ̕��    DI      ��    DI P   $  �����    B�B�B �B(�A0�A8�DPMXF`aPa8A0A(B BBB   P   x  ���p    B�B�B �B(�A0�A8�DPlXB``PI8A0A(B BBB       �  ���>    A�CA�x   �  <���6    A�Cq        R����    A�C�     ,  ����    A�CN      L  ����6    A�Cq      l  Ɨ��    A�C      �  ����;    A�Cv      �  ח��c    A�C^     �  ���    A�CM      �  ���    A�CJ        ����    A�CF       (  ���    A�CB          L  ���    A�CM      l  ԙ��\    A�CW     �  ����    A�C�     �  ����    A�CZ      �  I���   A�C    �  5���   A�C    	  D���#    A�C^      ,	  H���    A�CV      L	  D���V    A�CQ     l	  z���)    A�Cd      �	  ����    A�CF      �	  p���)    A�Cd      �	  z���(    A�Cc      �	  ����,    A�Cg      
  ����)    A�Cd      ,
  ����    A�CF      L
  ����)    A�Cd      l
  ����(    A�Cc      �
  ����,    A�Cg      �
  ����    A�CF      �
  ����    A�CF      �
  z���4    A�Co        ����E    A�C@     ,  ����C    A�C~      L  ֚��&    A�Ca      l  ܚ��4    A�Co      �  ���E    A�C@     �  ���C    A�C~      �  8���&    A�Ca      �  >���*    A�Ce        H���J    A�CE     ,  r���*    A�Ce      L  |���J    A�CE     l  �����    A�C�     �  W����    A�C�     �  Ԝ���    A�C�     �  �����    A�C�     �  ���U    A�CP       6���U    A�CP     ,  k����   A�C�    L  ����   A�C�    l  i���(    A�Cc      �  r����    A�C�     �  ����    A�C�     �  ����F    A�CA     �  ����Z    A�CU       �����    A�C�     ,  ����<    A�Cw      L  ����     A�C[      l  �����    A�C�     �  D����   A�C�    �  ����6    A�Cq      �  
���Q    A�CL     �  ;���    A�CN        .���B    A�C}      ,  P���    A�CQ      L  ����-    A�Ch      l  ����$    A�C_      �  ����$    A�C_      �  ����$    A�C_      �  ����3    A�Cn      �  ʢ��%    A�C`        Ϣ��9    A�Ct      ,  ���J   A�CE    L  ���+    A�Cf      l  ���G   A�CB    �  D���+    A�Cf      �  O���    A�CU      �  I���+    A�C      �  X���"    A�C]        Z���Z    A�CU     (  ����I    A�CD     H  ����V    A�CQ     h  ���#    A�C      �  ����)    A�Cd      �  ���+    A�C      �  ���    A�C      �  ���    A�C      �  	���*    A�C        ���+    A�C      0  &���+    A�C      L  5����    A�C�     l  ����   A�C    �  ���*    A�C      �  ����+    A�C      �  ���+    A�C      �  ���&    A�Ca         ���/    A�C        -���/    A�C       8  @���   A�CE��      \   ���1   A�C,    |  1���.    A�C      �  C���=   A�C8    �  `���3    A�C      �  w����    A�C�     �  S����    A�C�       ׭���    A�C�      4  �����    A�CE��      X  2���3    A�C      t  ���M   A�CH    �  K���L   A�CG    �  w���   A�C    �  t���)    A�Cd      �  }���    A�Cz       ܹ���    A�C�     4  ����)    A�Cd      T  ĺ��(    A�Cc      t  ̺��0    A�Ck      �  ܺ��+    A�Cf      �  ���E    A�C@      �  ���h   A�CE�^      �  P����   A�CH��        ����#   A�CE�     @  ����}    A�Cx     `  8���2    A�Cm      �  J���'    A�Cb      �  R����    A�C�     �  �����    A�C�     �  ����O    A�CJ        ����    A�CQ         ����I    A�CD     @  �����    A�C�     `  �����    A�C�     �  V���X    A�CS      �  ����D   A�CE�:     �  �����    A�C�     �  ����L    A�CG        �����    A�CE��      (  &����    A�C�     H  ����    A�CL      h  ����    A�CY      �  ����    A�CY       �  ����a   A�CE�W     �  ����    A�CY       �  �����   A�CE��       8���    A�CL      0  *���j    A�Ce     P  t���(    A�Cc      p  |���    A�CY       �  z���7   A�CE�-     �  ����    A�CY       �  ����7   A�CE�-      �  ����a   A�CE�W       ����    A�CY       <  �����   A�CE��     `  D���d    A�C_     �  ����j    A�Ce      �  ����7   A�CE�-      �  ����7   A�CE�-     �  ����K    A�CF       %���W    A�CR     (  \���    A�CQ      H  R���    A�CY      h  P���1    A�Cl       �  b����   A�CE��     �  ���    A�CX      �  ����H    A�CC     �  &���    A�CZ        &���    A�CZ      ,  &���V   A�CQ    L  \���    A�CQ      l  R���H    A�CC     �  z���    A�CY      �  x���1    A�Cl       �  �����   A�CE��     �  )���    A�CX        &���V   A�CQ    0  \����   A�C�    P  ����1    A�Cl       p  �����   A�CE��      �  r����   A�CE��     �  ����    A�CJ      �  ����    A�CJ       �  �����   A�CE��        H����   A�CE��     @  ����1    A�Cl      `  ]���/    A�Cj       �  l���    A�CP          �  � ��   A�C    �  ���0    A�Ck      �  Q���V    A�CQ       ����V    A�CQ     $  ����V    A�CQ     D  ����V    A�CQ     d  )���V    A�CQ     �  _���V    A�CQ     �  ����V    A�CQ     �  ����V    A�CQ     �  ���V    A�CQ        7���V    A�CQ     $   m���V    A�CQ     D   ����K    A�CF     d   ����J    A�CE     �   ����S    A�CN     �   +���S    A�CN     �   ^���S    A�CN     �   ����S    A�CN     !  ����S    A�CN     $!  ����S    A�CN     D!  *���S    A�CN     d!  ]���S    A�CN     �!  ����S    A�CN     �!  ����S    A�CN     �!  ����S    A�CN     �!  )���H    A�CC     "  Q����   A�C�    $"  ����.    A�C      @"  ���Q    A�CL     `"  =���Q    A�CL     �"  n���*    A�C      �"  |���*    A�C      �"  ����R    A�CM      �"  ����    A�Cz         �"  ���*    A�Ce       #  3����   A�CJ���   @#  ����o    A�Cj     `#   ���    A�C�      �#  � ��?   A�CE�5      �#  ���r   A�CE�h     �#  ���    A�C�      �#  ����    A�CE��       $  G���   A�CJ���   0$  ��>    A�Cy      P$  \��S    A�CN     p$  ���    A�CL      �$  ���    A�CM      �$  t��6    A�Cq      �$  ���r    A�Cm      �$  ���P    A�CE�F      %  ��C    A�C~      4%  ,��    A�CM      T%  ��4    A�Co      t%  2��w    A�Cr      �%  ����    A�CE�{      �%  ���!    A�C\      �%  ���%    A�C`      �%  ���    A�CM      &  ���    A�CL      8&  ���O    A�CJ     X&  ��I    A�CD     x&  /��I    A�CD     �&  X��*    A�Ce      �&  b��    A�CL       �&  T���    A�CE��      �&  -	��   A�C    '  ��N    A�CI     <'  B���    A�C�     \'  ����    A�C�     |'  ���+    A�Cf      �'  ���/    A�Cj      �'  ����   A�C�    �'  Z���   A�C�    �'  ��m    A�Ch     (  P��T    A�CO     <(  ���?    A�Cz      \(  ���h    A�Cc     |(  ���n    A�Ci     �(  :��   A�C    �(  4��    A�Cz     �(  ����    A�C|     �(  ����   A�C�    )  ���    A�C    <)  ����    A�C�     \)  r��u    A�Cp     |)  ���E    A�C@     �)  ���    A�CL      �)  ����    A�C�     �)  Z��h    A�Cc     �)  ����    A�C�     *  v��U    A�CP     <*  ���U    A�CP     \*  ���E    A�C@     |*  ��    A�CF      �*  ����    A�C�     �*  ���4    A�Co      �*  ���    A�CU      �*  ���*    A�Ce      +  ���    A�CZ      <+  ���    A�CL      \+  ���E   A�C@    |+  � ��*    A�Ce      �+  � ��    A�CZ      �+  � ��    A�CL      �+  � ���    A�C�     �+  d!���    A�C|     ,  �!��f    A�Ca     <,  "��]    A�CX     \,  H"��I    A�CD     |,  q"��    A�CU      �,  k"���    A�C�     �,  4#��R    A�CM     �,  f#��B    A�C}      �,  �#��5    A�Cp      -  �%��"    A�C]      <-  �%��*    A�Ce       \-  �%���   A�CE��     �-  N'��a    A�C\      �-  �'���   A�CE��     �-  K*��+    A�Cf      �-  V*��(    A�Cc      .  ^*��3    A�Cn      $.  r*��#    A�C^      D.  v*��(    A�Cc      d.  ~*��2    A�Cm      �.  �*��    A�CL      �.  �*��*    A�Ce      �.  �*��G    A�CB     �.  �!��    A�CI      /  �*��    A�CI   $   $/  �!���    A�CI���v      L/  �!��    A�CI   $   l/  �!���    A�CI���v      �/  *��    A�CI      �/   *��0    A�Ck      �/  *��    A�CL      �/  *��    A�CU      0  �)��C    A�C~      40   *��"    A�C]      T0  "*��0    A�Ck      t0  2*��G    A�CB     �0  Z*��1    A�Cl      �0  k*��    A�CU      �0  f*��    A�CU      �0  `*��J    A�CE      1  �*��<   A�CE�2     81  �,��    A�CI      X1  �,���    A�C�     x1  -���    A�C�     �1  �-���   A�C�    �1  �.��-    A�Ch      �1  /��+    A�Cf      �1  ����    A�C�      2  � ��    A�CP          <2  �i��&    A�Ca      \2  �i��H    A�CC      |2  j��e    A�CE�[      �2  Hj��M    A�CH     �2  vj��&    A�Ca      �2  |j��<    A�Cw       3  �j��g    A�Cb      3  �j��c    A�C^     @3  $k��6    A�Cq      `3  :k��Q    A�CL     �3  lk��S    A�CN     �3  �k��O    A�CJ     �3  �k��.    A�Ci      �3  �k��	   A�C     4  �l��L    A�CG      4  �l��S    A�CN     @4  (m��O    A�CJ     `4  �,��+    A�C      |4  �,���    A�C�     �4  -��5    A�C      �4  7-��#    A�C      �4  >-��+    A�C      �4  M-��3    A�C      5  d-��2    A�Cm      ,5  v-���    A�C�     L5  
.���    A�C�     l5  �.���    A�C�     �5  5/���    A�C�     �5  �/��x    A�C      �5  0���    A�C�     �5  �0���    A�C�     6  H1��    A�CO      (6  <1��0    A�Ck      H6  L1���    A�C�     h6  2��}    A�Cx     �6  b2��b    A�C]     �6  �2��[    A�CV     �6  �2��`    A�C[     �6  3��/    A�Cj      7  .3��/    A�C       $7  A3���    A�CH��      H7  �3���    A�C�     h7  j4��3    A�C      �7  �4��x    A�C      �7  �4��x    A�C      �7  95��3    A�C      �7  P5��3    A�C      �7  g5��x    A�C      8  �5��x    A�C      ,8  6��7    A�C      H8  :6��7    A�C      d8  U6��x    A�C      �8  �6��x    A�C      �8  7��/    A�C      �8   7��/    A�C      �8  37��D    A�C      �8  W7���    A�C�     9  8��K    A�CF     49  78��"    A�C]      T9  98��P    A�CK     t9  i8��%    A�C`      �9  n8��    A�CU      �9  h8��    A�CU      �9  b8��    A�CS      �9  Z8��    A�CS      :  R8��I    A�CD     4:  {8��"    A�C]      T:  }8��$    A�C_      t:  �8��    A�CR      �:  x8���    A�C�     �:  59��+    A�C      �:  D9��2    A�C      �:  Z9��.    A�C      ;  l9��/    A�C      $;  9��.    A�C      @;  �9��+    A�C      \;  �9��#    A�C      x;  �9��.    A�C      �;  �9��*    A�C      �;  �9��.    A�C      �;  �9��2    A�Cm      �;  �9��2    A�Cm      <  �9��/    A�C      (<  :��/    A�C      D<  #:��    A�CQ      d<  :��    A�CO      �<  :��    A�CO      �<  :��z    A�Cu      �<  [:���   A�CH��     �<  �;��6    A�C      =  <���    A�C�     $=  �<���    A�C�     D=  =��[    A�CV     d=  Q=��[    A�CV     �=  �=��[    A�CV     �=  �=��    A�CQ      �=  �=��    A�CO      �=  �=��    A�CO      >  �=��D    A�C      $>  �=��;   A�C6    D>  �?��;   A�C6    d>  �A��2    A�C      �>  8c��    A�CM      �>  �A���   A�C�    �>  
c��*    A�Ce      �>  c���   A�C�     ?  TO���   A�C�     ?  �i��*    A�Ce      @?  �i���   A�C�    `?  Vp��*    A�Ce      �?  `p���   A�C�    �?  w��*    A�Ce      �?  w���   A�C�    �?  �}��    A�CK       @  �}��1    A�Cl       @  �}��)    A�Cd       @@  �}��N    A�CE�D      d@  �}��)    A�Cd       �@  ~��N    A�CE�D       �@  ,~���   A�CH��     �@  ց��1    A�Cl      �@  ���)    A�Cd       A  ����   A�CH��     0A  ����1    A�Cl      PA  ����)    A�Cd       pA  �����   A�CH��     �A  b���1    A�Cl      �A  t���)    A�Cd       �A  ~����   A�CH��      �A  (����    A�CE��      B   ���;    A�Cv      <B  ����   A�C�     \B  ֔���    A�CE��       �B  �����    A�CE��       �B  >����    A�CE��       �B  �����    A�CE��       �B  �����    A�CE��       C  \����    A�CE��       4C  ����   A�CE��     XC  ����d    A�C_     xC  ����   A�C�     �C  �����    A�CE��       �C  T����    A�CE��       �C  ����    A�CE��       D  �����    A�CE��       (D  n����    A�CE��       LD  $����    A�CE��       pD  ֫���   A�CE��     �D  g���d    A�C_     �D  �����   A�C�     �D  f����    A�CE��       �D  ����    A�CE��       E  λ���    A�CE��       @E  �����    A�CE��       dE  6����    A�CE��       �E  ����    A�CE��       �E  �����   A�CE��     �E  /���d    A�C_     �E  s����   A�C�     F  .����    A�CE��       4F  �����    A�CE��       XF  �����    A�CE��       |F  L����    A�CE��       �F  �����    A�CE��       �F  �����    A�CE��       �F  f����   A�CE��     G  ����d    A�C_     ,G  ;���J    A�CE     LG  e���    A�CL      lG  V���J    A�CE     �G  ����W    A�CR     �G  ����Y    A�CT     �G  ����    A�CM      �G  �����    A�C�     H  c���U    A�CP     ,H  ����W    A�CR     LH  ����W    A�CR     lH  ����    A�C�     �H  ����U    A�CP     �H  ����W    A�CR     �H  ����W    A�CR     �H  (����    A�C�     I  ����U    A�CP     ,I  ����W    A�CR     LI  ���W    A�CR     lI  J����    A�C�     �I  ����U    A�CP     �I  ����W    A�CR     �I  5����   A�C�    �I  �����   A�C�    J  E����   A�C�    ,J  �����   A�C�    LJ  L����   A�C�    lJ  �����   A�C�    �J  \����   A�C�    �J  �����   A�C�    �J  c����   A�C�    �J  �����   A�C�    K  s����   A�C�    ,K  �����   A�C�    LK  z����   A�C�    lK  ����   A�C�    �K  �����   A�C�    �K  	����   A�C�    �K  ����S    A�CN     �K  �����    A�C�     L  +���;    A�Cv      ,L  F����    A�C}     LL  ����r    A�Cm     lL  ����r    A�Cm     �L  L���%    A�C`      �L  Q����    A�C�     �L  ����3    A�C      �L  ����Y    A�CT     M  ���i    A�Cd     (M  Q���m    A�Ch     HM  ����n    A�Ci     hM  ����p    A�Ck     �M  <���m    A�Ch     �M  �����    A�C�     �M  ���*   A�C%    �M  &���,    A�Cg      N  2���\    A�CW     (N  n���/    A�C      DN  ����/    A�C      `N  ����/    A�C      |N  ����2    A�C      �N  ����2    A�C      �N  ����2    A�C      �N  ����2    A�C      �N  ����/    A�C      O  ���3    A�C      $O  )���3    A�C      @O  @���3    A�C      \O  W���/    A�C      xO  j���3    A�C      �O  ����/    A�C      �O  ����/    A�C      �O  ����3    A�C      �O  ����3    A�C      P  ����3    A�C       P  ����.    A�C      <P  ����/    A�C      XP  ���/    A�C      tP  $���.    A�C      �P  6���/    A�C      �P  I���/    A�C      �P  \���3    A�C      �P  s���f    A�Ca     Q  ����+    A�C       Q  ����2    A�C      <Q  ����@   A�C;    \Q  ����]    A�CX     |Q  ; ��7    A�Cr      �Q  R ��H    A�CC     �Q  z ��f    A�Ca     �Q  � ��a    A�C\     �Q  ��g    A�Cb     R  H��W    A�CR     <R  ��:    A�Cu      \R  ���C    A�C~      |R  T��    A�CP      �R  ����    A�C�     �R  p��Q    A�CL     �R  ���R    A�CM     �R  ���,    A�Cg      S  ���    A�CI      <S  ���    A�CI       \S  ���P    A�CE�F      �S  ���    A�CI      �S  ���    A�CI       �S  ���P    A�CE�F      �S  ��    A�CI      T  ���    A�CM      $T  ���%    A�C`       DT  ���{    A�CG��o    hT  D��    A�CQ      �T  :��    A�CU      �T  4��$    A�C_      �T  8��7    A�Cr      �T  O��
    A�CE      U  :��    A�CQ      (U  0��$    A�C_       HU  4��    A�CQ          lU  ��=    A�Cx      �U   ��     A�C[      �U   ��    A�CK      �U  ��    A�CL      �U  ���   A�C�    V  l��|    A�Cw     ,V  f��    A�CX      LV  d��+    A�Cf      lV  o��g    A�Cb     �V  ���    A�CZ      �V  ���    A�CH      �V  (��7    A�Cr      �V  @��-    A�Ch      W  N��+    A�Cf       ,W  Z��K   A�CE�A     PW  ���G   A�CB    pW  ���   A�C    �W  ���X   A�CS    �W  �	��    A�CZ      �W  �	��    A�CZ      �W  �	��    A�CZ      X  �	��    A�CZ       0X  �	��    A�CZ          TX  �	��    A�CJ      tX  �	���    A�C�     �X  n
���    A�C�     �X  ���    A�C�     �X  ����    A�C�     �X  ���   A�C    Y  t���    A�C�     4Y  ���    A�C�     TY  ����    A�C�     tY  z���    A�C�     �Y  ���    A�C�     �Y  ����    A�C�     �Y  H���    A�C�     �Y  ����    A�C�     Z  x��    A�CH      4Z  f��    A�CZ      TZ  f��!    A�C          tZ  h��J    A�CE     �Z  ���    A�CU      �Z  ���f    A�Ca     �Z  ���J    A�CE     �Z  ���.    A�Ci      [  
��)    A�Cd      4[  ��E    A�C@     T[  8��}    A�Cx     t[  ����    A�C�     �[  ��W    A�CR     �[  K���   A�C�         7@     PJ@     4�@     ��������        ��������        ��A     	�A     A�A     �B     �B     A+B     fIB     �|B     q~B     �B     �B                     �@     B�@      �@     ��@     �@     ��@     L�@     ��@                                     ��A     ��A     ��A     ��A     ��A     ��A                     ��A     ��A     ��A     6�A     ~�A     ��A                                     ��A     ��A     ��A     ��A                                                                    1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `  �C     C     C     �C     GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             ]@     �      L@     I       �@     2       �@     -       �@            @     "       *@     -      X@     "       z@     �       H@     �       �@     -                       ,    D       @"@     �                       ,    �       N$@     >                       ,    �       �$@     �                      �   �'       y&@           �(@            �(@     \        )@     �       �)@            �)@     #       �)@            �)@     V       J*@     )       t*@            �*@     )       �*@     (       �*@     ,       �*@     )       (+@            4+@     )       ^+@     (       �+@     ,       �+@            �+@            �+@     4       �+@     E       C,@     C       �,@     &       �,@     4       �,@     E       %-@     C       h-@     &       �-@     *       �-@     J       .@     *       ,.@     J       v.@     �       G/@     �       �/@     �       �0@     �       Q1@     U       �1@     U       �1@     �      �3@     �      95@     (       b5@     �       6@     �                       ,    \E       �6@     �                      �   �G       N8@           fJ@             �J@     �       4K@     �      �(@            �(@     \        )@     �       �)@            M@     6       :M@     Q       �M@            �M@     B       �M@            �)@     #       �)@            �)@     V       �M@     M      CP@     L      �R@           �*@     )       (+@            4+@     )       �+@     ,       �T@     )       �T@            TU@     �       RV@     )       |V@     (       �V@     0       �V@     +       �+@            �+@            �,@     4       �,@     E       h-@     &       �V@     E       DW@     h      �Z@     �      \_@     #      .@     *       a@     }       �a@     2       .b@     '       Vb@     �       c@     �       �c@     O       *d@            @d@     I       �d@     �       ~e@     �       :f@     X       �f@     D      �g@     �       �h@     L       i@     �       �/@     �       �i@     �       Rj@            cj@            �j@            �j@     a      m@             m@     �      �o@            �o@     j       (p@     (       Pp@            np@     7      �q@            �q@     7      �r@     a      ]u@            |u@     �      x@     d       lx@     j       �x@     7      z@     7      F{@     K       �{@     W       �{@            �{@            |@     1       N|@     �      �@            .�@     H       v�@            ��@            ��@     V      �@            "�@     H       j�@            ��@     1       ��@     �      }�@            ��@     V      ��@     �      ��@     1       ʑ@     �      j�@     �      
�@            �@            (�@     �      Ȗ@     �      h�@     1       95@     (       6@     �                       \   ��       ��@           �(@     \       �)@            ��@           ��@     0       �)@     #       �)@            �@     R       4�@            �*@     )       (+@            4+@     )       �+@     ,       �+@            �+@            �,@     4       �,@     E       h-@     &       .@     *       �/@     �                       �   ��       ��@     3	      :M@     Q       �M@            �M@     B       �M@            �(@            �(@     \        )@     �       �)@            M@     6       �@     *       �)@     #       �)@            �)@     V       �@     R       �@     S       �*@     )       (+@            4+@     )       d�@            v�@            ��@     6       �+@     ,       ��@     r       4�@            0�@     P       ��@     C       Ĳ@            ֲ@     4       
�@     w       ��@     �       �@     !       *�@     %       P�@            b�@            s�@     O       ´@     I       �+@            �+@            �,@     4       �,@     E       �@     I       h-@     &       T�@     *       ~�@            �T@            TU@     �       RV@     )       ��@     �       .@     *       ��@           DW@     h      |V@     (       �/@     �       6@     �       ��@     N       �a@     2       .b@     '       Vb@     �       c@     �       �c@     O       *d@            @d@     I       �d@     �       �Z@     �      ,.@     J       Rj@            �h@     L       cj@            �j@            �j@     a      m@             m@     �      �o@            �o@     j       (p@     (       Pp@            np@     7      �q@            �q@     7      ~e@     �       :f@     X       �f@     D      �g@     �       i@     �       �0@     �       �{@            �{@            |@     1       N|@     �      �@            .�@     H       v�@            ��@            ��@     V      �@            ]u@            "�@     H       j�@            �r@     a      |u@     �      x@     d       lx@     j       �x@     7      z@     7      F{@     K       �1@     U       ��@     1       ʑ@     �      j�@     �      
�@            �@            }�@            ��@     1       (�@     �      Ȗ@     �      ��@     �      ��@     V      �3@     �      h�@     1       95@     (                           /                      �   �      �@     g       �(@            �(@     \        )@     �       �)@            :M@     Q       �M@            �M@     B       �M@            �)@     #       �)@            �)@     V       J�@     "       l�@     *       ��@     �      �*@     )       (+@            4+@     )       �+@     ,       �T@            TU@     �       RV@     )       2�@     a       ��@     �      J*@     )       t*@            �*@     )       �*@     ,       s�@     +       �V@     +       ��@     (       |V@     (       ��@     3       ��@     #       �@     (       F�@     2       x�@            ��@     *       ��@     G       ��@            �+@            �+@            	�@            �@     0       H�@            Z�@            �,@     4       �,@     E       h-@     &       DW@     h      �+@     4       �+@     E       �,@     &       t�@     C       �Z@     �      ��@     "       ��@     0       
�@     G       R�@     1       ��@            ��@            .@     *       �a@     2       .b@     '       Vb@     �       c@     �       �c@     O       *d@            @d@     I       �d@     �       �-@     *       ��@     J       ~e@     �       :f@     X       �f@     D      �g@     �       �h@     L       i@     �       �@     <      >�@            �/@     �       Rj@            cj@            �j@            �j@     a      m@             m@     �      �o@            �o@     j       (p@     (       Pp@            np@     7      �q@            �q@     7      v.@     �       L�@     �       �r@     a      ]u@            |u@     �      x@     d       lx@     j       �x@     7      z@     7      F{@     K       �{@            �{@            |@     1       N|@     �      �@            .�@     H       v�@            ��@            ��@     V      �@            "�@     H       j�@            ��@     �       ��@     1       ��@     �      }�@            ��@     V      ��@     1       ʑ@     �      j�@     �      
�@            �@            (�@     �      Ȗ@     �      �3@     �      ��@     �      h�@     1       95@     (       6@     �       �@     -       B�@     +                       �   ��      n�@     	;      :M@     Q       �M@            �M@     B       �M@            �(@            �(@     \        )@     �       �)@            M@     6       �@     *       x"A     &       �"A     H       �"A     e       L#A     M       �#A     &       �#A     <       �#A     g       d$A     c       �$A     6       �$A     Q       P%A     S       �%A     O       �%A     .       "&A     	      ,'A     L       x'A     S       �'A     O       �)@     #       �)@            (A            �)@     V       �V@     +       .(A     *       X(A     �      $/A     *       N/A     �      s�@     +       6A     *       D6A     �      �T@            TU@     �       |V@     (       �*@     )       (+@            4+@     )       ��@     6       �+@     ,       =A     *       :=A     �      �+@            �+@            DA            DA     1       HDA     )       rDA     N       �DA     )       �DA     N       8EA     �      IA     1       8IA     )       bIA     �      0MA     1       bMA     )       �MA     �      �Z@     �      �,@     4       �,@     E       �@     I       h-@     &       ZQA     1       �QA     )       �QA     �      �UA     �       ��@            �VA     ;       �VA     �      �]A     �       p^A     �       F_A     �        `A     �       �`A     �       �aA     �       �bA     �      [jA     d       ��@     *       �jA     �      �qA     �       trA     �       JsA     �       $tA     �       �tA     �       �uA     �       �vA     �      _~A     d       �~A     �      ��A     �       x�A     �       N�A     �       (�A     �       ��A     �       ؉A     �       ��A     �      c�A     d       �a@     2       .b@     '       @d@     I       ~e@     �       :f@     X       �c@     O       �f@     D      �g@     �       �h@     L       �d@     �       i@     �       .@     *       ��@           ǒA     �      ��A     �       |�A     �       R�A     �       ,�A     �       �A     �       ܝA     �       ��A     �      g�A     d       ˦A     J       �A            &�A     J       p�A     W       �@     R       v�@            ȧA     Y       "�A            4�A     �       ӨA     U       (�A     W       
�@     G       �A     W       ֩A     �       u�A     U       ʪA     W       !�A     W       x�A     �       �A     U       l�A     W       Rj@            Pp@            �q@            �r@     a      ]u@            |u@     �      �o@            x@     d       *d@            lx@     j       (p@     (       cj@            �x@     7      �j@            z@     7      �o@     j       np@     7      �q@     7      F{@     K       �/@     �       6@     �       ��@     N       ìA     W       �A     �       ��A     U       �A     W       e�A     �      �A     �      ��A     �      T�A     �      ��@     J       ��A     �      ��A     �      L�A     �      �A     �      ��A     �      ;�A     �      �A     �      ��A     �      �@            j�@            ��@     1       ��@     �      }�@            "�@     H       ��@            v�@            ��@     V      �{@            m@            .�@     H       �{@            ��@     V      ,.@     J       *�A     �      ��A     �      z�A     �      �A     �      95@     (       L�@     �       h�@     1       (�@     �      Ȗ@     �      �@            
�@            �@            |@     1       ʑ@     �      j�@     �      �0@     �       ��@     �       �1@     U       �3@     �      ��@     �                      ,    �]      ��A     �                      ,    p      ��A                           |   t      ��A     �      �(@            4�A            J�A     ,       v�A            ��A            ��A     P       ��A            ��A            ��A     P       N�A            \�A            n�A     %       ��A     {       �A            &�A            @�A     $       d�A     7       ��A     
       ��A            ��A     $       ��A                            L   ˓      ��A     �       ��A     =       �A             0�A            @�A            R�A     �      ��A     |       X�A     7       ��A     -       ��A     +       ��A     K      6�A     G      ~�A           ��A     X      ��A            
�A            *�A            J�A            j�A                            �   U�      ��A     s      �(@            �(@     \        )@     �       �)@            �)@     #       �)@            �)@     V       �*@     )       (+@            4+@     )       �+@     ,       ^+@     (       �+@            �+@            �,@     4       �,@     E       h-@     &       %-@     C       .@     *       ,.@     J       �/@     �       �0@     �       �1@     U       �3@     �      95@     (       6@     �                       ,    ��      ��A     A                       �   ��      @�A     B      �(@            �(@     \        )@     �       �)@            M@     6       �)@     #       �)@            �)@     V       J*@     )       t*@            �*@     )       ��A     )       �*@     ,       �+@            �+@            �+@     4       �+@     E       ��A     E       �,@     &       �-@     *       ��A     }       v.@     �       m�A     �       �A     W       c�A     �      95@     (       b5@     �                                       @       �	  #  a                   �  5   �  m  H   �  �  [   �  �  n   �  �  	�   �  �  J  �   int �   �  �  �n   -  u   4  �   ,  )     <   3  O   �  b     4�   �  P  h  �    �  �   bpp 	�   �  �   
 �    �  �n   	�  J  i	  �
  (	�  x 	�    y 		�   h  	�   �  	�   �  	�   �  	
�   ݨ  		�  �  	

�     
�     	  �  '  x 	�    y �    +  	  '     r  r �    g �   b �   a �    o	  8  "�  �  �  #�   @  $�   �D  %�   �  &�   
 �  �  n    �  �  '~  ()�   �    *�    h  +
�   �  ,
�     -�   bpp .�   }  /�   @  0�   �  1
�   �  2
�   g  3�    (
  4�   $ �   5�  E  6  �  
h  
�  |B  /  x �    y �   h  �   �  �      �   {  /  �  �   l,  �  tD  �  (  �    �  ?  n   _ D  �  I @�    �      	\  �  #	\  �  &	\    )	\   �  ,	\  (�  -	\  0
  2�   8�  5�   < 
�  Q  8"K  �  K�  
�  �  L�  �  M�  (D	  Y  =  �    z  �   msg �   �  �   V  �     F	  
  �  �q  
�  G  ��  8  ��   }  ��   �  ��   s
  [   |  A"�  
�  �   �  \   �h   w  �  �  �.  �  �P   A  X  
  h  .  �  �    �  m:  
@  P  �  h   �  �\  
b  h  �  �  �   �   h   �  �"�  
�  �   PH-  V J�   @  Kn   pos Ln   �  NS  �
  OS   ��  P_  (G Q�  0P  S�  8�  T�  @�p  U�  H W  �S  q  ��   ѷ  �h   �  �-  �  �k  
q  n   �  �  n   �  n    
5   �  �  
�  �  �   �  :�   �  L�  x N�   y O�   c  Q�  p   w1  M   y�   �  y�    z�  ]  z�     |�  �	  (�    [    h  [   �  	�   ݨ  
�  �  H   �  5   !  5   
  h    �  =  q  (Q,	  �  S�      T�     V,	  E  W�  �  X2	     Z�     
�  
�   �  \�  G  [   ��	  \   �
  pmoc�  stib�	  ltuoH  tolp �	  �E	    ��  5  ��   �  �H   �  ��   �
  �[   �  ��   T	  �   4  ��	  
�	  
  h   d  �.
  �  �h   o  ��	   /  �
    $H
  
N
  �  +�
  �  -;
   �  .;
  �  /h   �  D�
  n�  F;
   W   G;
   �  I�
  �  @<>  h  >�   �  ?�  �  A�  �  B�  �  C�     E�  (  F�  0  G�  8 }
  I�
  �
   s�  �  u�	   h  v�	  @  x�  >  z�  V  {�   �  }K  2  �#�  
�  �  .  �"�  
�  /  �  � �  
�  ]	  ��  �   �	   �  �	    �	  �  �	  	  �	   ,  �  (�  �  0�  �	  8{  �  @O  !�	  HS  "�  P  $.
  XR   )1  h  +�	  �f  ,�	  �  -�	  ��  .�	  �\  0�	  ��  1�	  ��  3�	  � 	  4�	  ��  6  �@  7�  �:  8h  ��  <�  �P  =�  ��  >�  ��  @�
  ��
  B.
  �    Ch  ��  E�  � �   �  
�  �  Xm  �
  o�     p.
  	  qU  �  r�  P �  $%  
  �  0\h  �  ^�   �
  _�  �  `  �  a�	    b.
   	  d>  0�  e�	  p  f�	  x�  g�  ��  i�	  ��  k�  ��  l�	  �:  m�	  �A  o8	  �b  q�	  �f  rb  � �  th    �  u�      w�   �  x�   �  zh    �  |z  ( *  F#u  
{  �  A�  �
  C�   8  D�  #  E�	    F�	     [   ��  �     bmysO  cinu=  sijs�    bg�  5gib&  snawk  ahoj�    bgX  sijs�    bg{  5gib  snaw^
  ahojH  BODA4   EBDA9
  CBDA�  1tal�  2tal   nmra R
  �  #   `)�  
�  �   
�	  
�  
h    �)�  
�  �   
  8HU  >  J�	   V  K�	  }	  M�	  �
  N�	  f  P�    Q�   �  R�  (�  S�  0 �  U�  #  �$o  
u  4	  �  �)�  
�  �  �   �  n    !]  �  	 �B     v  �B�  ,  C�   �  D?  pos E'  �   F�  � l  "fb I
�  	� C     !�   JP  	� C     !�	  K�  	� C     �   R  n    !y  MB  	C     !�  N'  	 �B     !�  O�  	C     !  P�  	C     !<  Q'  	C     !0  S�  	(�B     !  U�  	C     !�  W�  	 C     !�  X	�  	(C     !�  sr  	)�B     !q  t�  	@C     !o  v�   	hC     #�    $�  
  |  �     $�  8  �  �    �    $�  !n  �  �     $�  *I  �  �    (   $&  ;�
  �  �    (   %�  L�  (    !    [    %:  P�  (  :  E    [    $|  Z0  Z  j    [   (   %�  dX  �   �  �     %   h`  (  �  �    [    %\  }  (  �  �     %  �N  (  �  �     &*  ��   &�  ��  'num �[   (T (   
Z    
�  #y  �  &�  	�   &�  
�  'obj (  )    w  }  �   (T (   
.  �  !�  wZ  	pC     !   x(  	�C     *&  h  +N  7@            �,�  �  �  -�  #  -  �    .�       �@     -       �)  /�  �h 0�  �@     >       �e  1�  ��   �l1p  ��   �h 2!  �  H@     �       ��  3�  #  �X4pos P[   �T5_�  S�  �h6�@     8       7i U[   �d  8�  �  z@     �       �  3�  #  �H4obj *(  �@5"O  +�  �X 9e  )  3  -�  �   :  �  V  X@     "       �_  /)  �h 8�  ~  *@     -      ��  3�  #  �H4pos h[   �D5_�  n�  �h7obj r(  �X;P@     	       �  5yu  j(  �P 6d@     8       7i p[   �d  8�    @     "       �7  3�  #  �h4pos L[   �d 2j  V  �@            �c  3�  #  �h ,g  q  {  -�  #   :c  �  �  �@     -       ��  /q  �h <�  ��   
@     �	      ��  5�
  ��  �H5l  ��  �@5?  ��   ��5�   ��  ��5�  ��  ��5�  ��   ��6@     u      =msg eY  ��~;�@     7       �  =i �   �l6�@            =win (  ��  ;�@     
        =i )�   �h6@     �      =win *(  ��66@     �       >	  3Y  ��~>�  5�   �d>�  6�   �`   ;<@     �       a  >	  SY  ��~>�  U�   �\>�  V�   �X ;q@     �       �  >I  jY  ��~ 6v@     &       =i ��   �T6�@            =j ��   �P    
�  ?Q  �f  G@     �      �  4win �(  ��5�  �'  �� ?�  �%  e@     �      ��  5n  ��   �L6�@     �      7j �
�   �l6�@     �      5�  ��  �k5�  �?  ��~5�  ��  �X;�@     D       �  7i ��   �d 6O@     �       7win �(  �P    ?c  z�  ]@           ��  5n  {�   �T6�@     �       7i ~
�   �l6�@     �       5�  	�  �k6�@     }       7j ��   �d6�@     e       5�  �?  ��~5�  ��  �X     
?  �  9  �  �  -�  �   :�    �  �@     2       ��  /�  �h @�  Q  '  L@     I       �=  4l 0=  �h4r E=  �` A3   N    �  @"@     0#@     �  src/gfx/sse2.asm NASM 2.14.02 �@"@              �      H  %  �  N$@     >       z  �  �  �  �  N   �  �  �  int �  �  B   	  N$@     >       �  q   �`  &q   �X  5q   �P  Dq   �H�  Sq   �@   bq   ��  Y	   v  �  �  �  �$@     �      ,  �  �  �@   �  �  E  6  int Z     Z   �  �  �    -   �  �  @   �  �  �@   �  �     4�   �  �   r  	-�  	D  +�  F  	�  ,�  K  
�  =	I  Z   %  �   
�  9s  Z   D  �  Z    
,  0m  Z   h  Z   �  �   �  (�  f   �  "�  b  ?  �  `   
w  �  Z   �  �   4    
�  �  Z   �  4   �   �  *  Z     std  c  �  h  q  j  �  c  �  �    4  :  x   �  q    R  X  x   T c  v c    �  �  �  q  j  �  c  �  ,  �  �  �  �   �  �  �  �  �  �   T c  v c   m  2  �  q  �j  T Z   �  �    �  �>  q  �j  T Z   �  �    6  ��  j  6  �?  j   l  c      h  F  z  �  frg 	Q  �  �  o   �  �  
 �   .  
7f   !�    "�  {*  #�  |Z   $�  ~;      z   %�      z  Z     &)    ?  E  �   &)  a  Z  e  �  �   &)  �  z  �  �  �   &)  �  �  �  �  �   &)  *�  �  �  �  �   &)  0x  �  �  �  �   &(  8  �    �  Z    '�  =O  �    )  �  �   'c  Q�  c  B  H  �   'c  T�  c  a  g  �   'm  X�  c  �  �  �   'R  \+  �  �  �  �   'R  `[  �  �  �  �   '!  d�  �  �  �  �   $f  �  �  �  �   (�  ��   (�  �c  T Z    �  )p  J�  
,  �  5  *�  *�   +�  	��A     �   `  +�  	p�B     �  �  ,a   -Z   ,  -�  ,�    ,Z   Z   .:  �  .�    �  |  +:  	��A     />  /P  0  H�  r&@            �1  CZ   g&@            �2  X&@            �X  3ѷ  =�  �h 2%  F&@            ��  3ѷ  9�  �h3  9'Z   �d �   -   4D  �%@     c       �  3  0Z   �\31  0'�  �P3�  03�  �H50  1�   �h5�  1�   �` 4h  �%@     ;       �?  5\  )�   �`6pid ,	f   �l 7x  �%@            �4�  `%@     6       ��  8msg  `  �h 2�  M%@            ��  3ѷ  �   �h3@  *4   �` �   4�  �$@     �       �	  3@  4   �h3ѷ  ,�  �`9  	  	��A      :�   	  ;@    	  4�  �$@     6       �N	  3x  Z   �l i	  J   q     �  &  �  �             �  �  �<   �  �  E  6  std  �  �  �   q  �  �  �  �  �  {   �   �   	�   �  q  {   �   �   	�   
T �  v �    a   �  J  q  �  �  �  �  ,  �       	�   �  �  �   4  :  	�   
T �  v �   �   2  �|  q  ��  
T "  �  !    �  ��  q  ��  
T "  �  '    6  ��  �  6  �?  �   l  �    n   �   F  �   J  �  �  �  �  �  �  int "  frg 	�  �  :  o   C  �  	 o  .  	7�   %  "  ,�  �   �  hex  �  �  �  {�  �  |"  �  ~;  �  �  	�    �    �  	�  	"    !)        	
   !)  a     +  	
  ":   !)  �  @  K  	
  "   !)  �  `  k  	
  "   !)  *�  �  �  	
  "!   !)  0x  �  �  	
  "'   !(  8  �  �  	
  	"   #�  =O  -  �  �  	
  "�   #c  Q�  �      	3   #c  T�  �  '  -  	
   #m  X�  �  F  L  	3   #R  \+    e  k  	3   #R  `[  9  �  �  	
   #!  d�  ?  �  �  	
   f  �  �  �  	
   $�  ��   $�  ��  
T "   �  �*  2�  �*  3Z(      	E   	   6C  �  )  4  	E  "o   $   <o   $�  ="  $�)  >�  $�   ?�  $�'  @�  $�#  A�  $<  B�  $�  C�  %�*  E&  �  �  	E  	"   &�*  >  �  	E  "�    �  'p  J9  (�-  N�!  $  
P   
T �  "�  "�  "�  ""  ""  ""  "�   (!  Na!  f  
P �	  
T �  "^  "�  "�  ""  ""  ""  "�   (�'  x<+  �  
P   
T �  "�  "�  ""  ""  ""  "�   ()  x  �  
P �	  
T �  "^  "�  ""  ""  ""  "�   (�  ��+    
T �  
F   "�  "�  "�   )4  ��)  
T �  
F �	  "�  "�  "^    �  
9  �  B  �  [	  �)  E#  t    	t  "�   q,  �	�  q,  �#  �  �  	  "t   *q,  _   �  �  	  "�   +�  	~-  �  �  �  	  "�   p,  �*      	  	"   )  "	�  �  $  /  	  "9   �$  'a&  C  N  	  "�   �$  1�  b  m  	  "�   ,�)  >t   ,ܨ  ?d  ,7&  @
0   �,)  A�  ��   	  �  �  �  
T �  	  "�   -c.  	�*  �  �  
T �  	  "�      �  H`*    	  	  	t   !�#  M�"  .	  9	  	t  "�   ,.  Q�   .U(  �  /].  <   � �  c  �)  E�&  |	  �	  	B  "�   q,  �	�
  q,  �&  �	  �	  	M  "B   *q,  N"  �	  �	  	M  "X   +�  	�   ^  �	  �	  	M  "X   p,  �"  	
  
  	M  	"   )  "	�(  ^  ,
  7
  	M  "9   �$  'r  K
  V
  	M  "�   �$  1�,  j
  u
  	M  "�   ,�)  >B   ,ܨ  ?d  ,7&  @
0   �,)  A�  ��   	6-  ^  �
  �
  
T �  	M  "�   -c.  	�$  ^  �
  
T �  	M  "�    �	  �  H�#  �	    !  	B   !�#  M�  6  A  	B  "�   ,.  Q�   .U(  �  /].  <   � 0�  
i    �  
T "  "  "   (`)  �@%  �  
F   "�  "�  "�   (`)  �O'  �  
F   "�  "�  "�   (f  �v,  �  
F �	  "�  "�  "^   (f  ��  %  
F �	  "�  "�  "^   1N#  3�  O  
T �  
F   "|  "�   1�  3�%  y  
T �  
F   "�  "�   1�  3,  �  
T �  
F �	  "|  "^   2   3n$  
T �  
F �	  "�  "^    3H  	�A     �  �  �  �  3a  	x�B     �  �  �  
  4)  5"  4�  5�  4�  �  4"  "  �  E  6:  \  6�  �  �  |  3G  	�A     'r  
6  <&  
�  7<&  

9(  �  �  	6    �  
'%  �  	6  "�    P(  
  7P(  
6"  �  �  	<    �  
�'  	  	<  "�    8D  
+�  S  8�  
,�  [	   �  �  [	  B  �	  M  4�
  4�	  9�  t  :<    S  t      4�  4  ;�  ;�  </  �  6@     �       ��  =�  �  �h>s '�  �d <7
  �  b5@     �       �  =�  S  �h>s '�  �d ?c  95@     (       �O  
T "  >a   �h>b #  �` @�  �3@     �      �{  
P   
T �  A��  N�  ��A�   N$�  ��A�'  N1�  ��A3(  N?"  ��Ah  O"  ��A�)  O"  ��A�D  O#�  ��B4  P�  �XBݨ  S{  ��Ck T"  ��D�4@     E       8  Ci a"  �l D�4@     -       [  Ci d"  �h E5@     0       Ci f"  �d  9�  �  :<    @$  �1@     �      ��  
P �	  
T �  A��  N^  ��A�   N$�  ��A�'  N1�  ��A3(  N?"  ��Ah  O"  ��A�)  O"  ��A�D  O#�  ��B4  P�  �XBݨ  S{  ��Ck T"  ��D�2@     E       t  Ci a"  �l D:3@     -       �  Ci d"  �h Eg3@     0       Ci f"  �d  @f  �1@     U       �I  
P   
T �  A��  x�  �hA�   x!�  �dA3(  x-"  �`Ah  x8"  �\A�)  y"  �XA�D  y�  �TFGi$  {	�    @�  Q1@     U       ��  
P �	  
T �  A��  x^  �hA�   x!�  �dA3(  x-"  �`Ah  x8"  �\A�)  y"  �XA�D  y�  �TFGi$  {	�    @�  �0@     �       �2  
T �  
F   A�  ��  �l>fo �/�  �`A��  �6�  �X <N  Q  �/@     �       �m  =�  �  �h>str 1�  �` @  G/@     �       ��  
T �  
F �	  A�  ��  �l>fo �/�  �`A��  �6^  �X <V
  �  v.@     �       ��  =�  S  �h>str 1�  �` @�  ,.@     J       �P  
F   A�  �!�  �L>fo �8�  �@A��  �?�  �� @�  .@     *       ��  
F   A�  � �  �h>fo �7�  �`A��  �>�  �X @�  �-@     J       ��  
F �	  A�  �!�  �L>fo �8�  �@A��  �?^  �� @�  �-@     *       �A  
F �	  A�  � �  �h>fo �7�  �`A��  �>^  �X <	  `  h-@     &       �|  =�  z  �hA/&  M�  �` 4�  @%  %-@     C       ��  
T �  
F   H�  3|  �HH��  3!�  �@ 4�  @O  �,@     E       �  
T �  
F   H�  3�  �HH��  3!�  �@ I�  *  @  J�  �  K�)  t   L  �  c  �,@     4       �t  M*  �hM3  �` <!  �  �,@     &       ��  =�  H  �hA/&  M�  �` @y  C,@     C       ��  
T �  
F �	  H�  3|  �HH��  3!^  �@ @�  �+@     E       �C  
T �  
F �	  H�  3�  �HH��  3!^  �@ I�	  Q  g  J�  S  K�)  B   LC  �  �  �+@     4       ��  MQ  �hMZ  �` I�  �  �  J�    J  )   L�  6.  �  �+@            ��  M�  �h I�  �     J�     L�  9*  #  �+@            �,  M�  �h <  K  �+@     ,       �`  =�  �  �hN9  �  <�  �  ^+@     (       ��  
T �  =�  �  �hA�  �  �d <�  �  4+@     )       ��  
T �  =�  �  �hA�  �  �` I�  �    J�  �  J  )   L�  *$  (  (+@            �1  M�  �h <�  P  �*@     )       �]  =�  z  �` <
  |  �*@     ,       ��  =�  S  �hN9  �  <�
  �  �*@     (       ��  
T �  =�  S  �hA�  �  �d <�
  �  �*@     )       �  
T �  =�  S  �hA�  �  �` I�	  #  6  J�  S  J  )   L  v(  Y  t*@            �b  M#  �h <  �  J*@     )       ��  =�  H  �` Ik  �  �  J�    K�  *!   O�  %'  �  �)@     V       ��  M�  �hM�  �` I�  �    J�    J  )   O�  g  *  �)@            �3  M�  �h I�  A  K  J�     O3    n  �)@     #       �w  MA  �h PA'  �'@           ��  A�*   �  ��~Az�  7�  ��~Aػ  J�  ��~A�%  �  ��~ P�,  y&@           �5  A�*   �  ��~Az�  7�  ��~Aػ  J�  ��~A�%  �  ��~ Q�  2F  Y  J�  K  J  )   O5  .  |  �)@            ��  MF  �h 4�  Q�  2�  �  J�  K  "�   O�  �  �   )@     �       ��  M�  �hM�  �` I�  �  �  J�  K   O�  K    �(@     \       �#  M�  �h R.  ^    �(@            �f  A@  #0   �h>p /  �` i	  J   �     �  �.  �  �6@     �      �  �  �9   �  |.   -   8@     <       ��   s  �   �Xlen !	-   �h"8@     &       i "-   �`  �   �  	�   m	 a  i7@     �       �a  
� a  �Hsrc 'h  �@
@  3-   ���.  t  �X�.  t  �P�7@     4       A  i -   �h �7@     E       i -   �`  a  s  h  �   ! a  7@     Z       �  
� c  �Hsrc <n  �@
@  H-   ���.  t  �`�.  t  �X/7@     4       i -   �h  �	 a  �6@     F       ��  
� a  �Xc �  �T
@  (-   �H�.  t  �`�6@     )       i -   �h  int  �Z   �  e�  T~  �            �  @�>  5   fint 5   @Q  M   S   �  S   @�o  M   �  k   �  "�  �   �  �   �  �   �  �  �  "�  ��   "3  ~   �   "  4�   �   "�  ��   �   "�:  	  g  A$G  1  Or  5    /rem 5    "%G  	  A_S  e  Or  �    /rem �    "`S  =  AQD  �  Or  �   /rem �   �  "RD  q  hfrg �  iN�  �	�  On <   pOm <   �P�v  �   ߰�jmsb �      �P73  �   ���N�  ;]  '  -  �   @  u  A  L  �  �     �  w�  �   d  j  �   k_st >�   l|  ?5   �	 B�  �  Qo   �  m�   �  n.  7�   7%  5   ,�  %�   %�  Rhex  S�  3  o�  {>  p�  |5   �  ~;    "  �   C�    2  �  5     )    S  Y  �   )  a  n  y  �  �   )  �  �  �  �  �   )  �  �  �  �  �   )  *�  �  �  �  �   )  0x  �  �  �     (  8      �  5    &�  =O    2  =  �  �   &c  Q�  �  V  \     &c  T�  �  u  {  �   &m  X�  �  �  �     &R  \+  �  �  �     &R  `[    �  �  �   &!  d�    �  �  �   f  �      �   �  ��   �  ��  T 5    �  �*  2  �*  3Z(  Y  _       	   6C  8  w  �     �      <�   �  =5   �)  >�  �   ?�  �'  @�  �#  A�  <  B�  �  C�  q�*  E&  �       5    r�*  >       =X    8  Dp  J�  8qK  N�Y  r  P    T �   2#  �   �  5   5   5   S    8�2  x ;  �  P    T �   2#  �   5   5   5   S    s�R  ��>  T �   F    �   8  2#    B�  

�  Q�  
�  �  
�  �)  
E#       #  �   q,  �
	�  q,  
�#  A  L  !#  #   ,q,  
_   `  k  !#  ,#   -�  
	~-  2#  �  �  !#  ,#   p,  
�*  �  �  !#  5     )  
"	�  2#  �  �  !#  �   �$  
'a&  �  �  !#  S    �$  
1�      !#  �   3�)  
>#   3ܨ  
?�"  37&  
@
�   �3)  
A�  � �3  
	#t  2#  e  p  T   !#     Tc.  
	�*  2#  �  T �  !#  �        �  
H`*     �  �  #   �#  
M�"  �  �  #  �   3.  
Q�   4U(  �  t].  �   � U�  BE3  		  u��  
	   Dd^  	  E<	  V4j  �    F)	  7G  5   i	  %�   Rred %h^   �o  0!
  �o  �F  �	  �	  6!   ,�o  �D  �	  �	  6!  A!   -�  �z  G!  �	  �	  6!  A!   tl     �    pU    �I     �D  !   [r  "D	  ( i	  q  %r
  �Q  '!=  �  T
  T f  e#   W�  '1Q  �  T �  N#    dV  5  Xh 8<  6!  �
  N#   pl  =�n  N#  �
  N#   �p  B�^  N#  �
  N#   lU  Ef|  N#  �
  N#   �I  I�  N#     N#   �D  LE  N#    N#    <3  Pfm  N#  2  8  �#   9�E  U�L  �  S  N#   9�_  Z�M  �  n  N#    c  djw  �  �  �#   , c  gar  �  �  �#  �#   -�  i
J  �#  �  �  �#  �#    ��  op  N#  �  �  �#   �D  |+G  �    �#  N#   ��  ��z    -  �#  N#  N#   5>  ��@  B  R  �#  N#  N#   �F  �4\  g  r  �#  N#   '�  Dj  �  �  �#  N#   O  $d  �  �  �#  N#  N#   �U  D�6  �  �  �#  N#  N#   �  x�E  �  �  �#  N#    q  �nq       �#  N#   �9  1y  6  A  �#  N#   '�=  Ӏ  V  a  �#  N#   '�z  #�8  v  �  �#  N#   0L  0Nx  �  �  �  �#   0L  9�/  �  �  �  �#  N#    �#  �#   :?3  �   D 	  T �  ;�P  �Z  A &
   r
  v�5  ��  (��  (�  (�-  (��
  (��
  (�  Gr
   'Z|  �@  h  s  �#  �   '�F  �V�  �  �  �#  N#   :�R  ��  T �  ;�P  �Z  L �  A &
   .H  5T  Xh 8�4  6!  �  e#   pl  =&i  e#    e#   �p  B�Z  e#    e#   lU  EP  e#  6  e#   �I  I�f  e#  P  e#   �D  L}S  e#  j  e#    <3  PO]  e#  �  �  �#   9�E  U�g  �  �  e#   9�_  Z)?  �  �  e#    c  d8  �  �  �#   , c  g~u  �  �  �#  �#   -�  i'O  �#      �#  �#    ��  oAs  e#  2  8  �#   �D  |�k  M  X  �#  e#   ��  ��0  m  }  �#  e#  e#   5>  ��A  �  �  �#  e#  e#   �F  �X  �  �  �#  e#   '�  �1  �  �  �#  e#   O  
e  �    �#  e#  e#   �U  DxT    .  �#  e#  e#   �  xfC  D  O  �#  e#    q  �{l  e  p  �#  e#   �9  E}  �  �  �#  e#   '�=  �9  �  �  �#  e#   '�z  #�`  �  �  �#  e#   0L  0�_  �  �  �  �#   0L  9�a  �    %  �#  e#    �#  �#   :?3  �   D Y  T f  ;�P  �Z  XA &
   �  w�~  �(�8  (�X  (�}  (�  (�  (�j  G�   'Z|  �<R  �  �  �#  �   '�F  �/L  �  �  �#  e#   :�R  ��  T f  ;�P  �Z  XL �  A &
    E"  V4j  �    F  /�  Y  xclz �3  5   Q  �    T �    y��  �$"  7 Q  5   ��  %�   %ʃ  %QS   g  �U  H�	a  �U  ���  �  �  N#  g  �   �    ,�U  ���  �  �  N#  Y#   -�  �
`D  _#  �  	  N#  Y#    ��  ��b  �  !  ,  N#     �U  ��   WS  ��   p ��   �=  �   �  �U  ��	  G�   �U  �Pc  �  �  e#  �   �   5    ,�U  �z  �  �  e#  p#   -�  �4  v#  �  �  e#  p#   �  �<   H�D  ��   L$H  �|#  P�B  �  X f  %\  �	�  %\  �/  ?  E  |#   ,%\  �l5  Y  d  |#  �$   -�  ��h  �$  |  �  |#  �$   �E  �|#      �R  �	�  T�  ��v  �  �  �#  Y#  Y#    �.   �	  �.  �R�  �  �  �#   �E  �	R!   �o  �e#  �e  �   "1|  �  u  ��=  <  G  C#  �#   Yu  (�t  \  g  C#  �#   z�  *�K  �#  �  �  C#  �#   &�  ��o    �  �  C#  �    0�  L�g    �  �  C#    �    �  ~��  �  �  C#     �I  �Ճ       C#    �    &WV  1	e;  �   9  ?  C#   {C  >
$                         @       H�v  @ �   H�`  A �    �~  H�U  �   �  �    �.  W�N  �   �  �    HQC  j<   1zz  l�   |  oK>  �  �  �    1́  |�   1]C  �   |�D  ��    I�~  ��<  N#  4  ?  C#  �    I��  &q  e#  X  c  C#  5    IFS  %n^  N#  |  �  C#  �    '4  7:k  �  �  C#   ']  >�J  �  �  C#  N#   �[  �
�#   �1  �R!  "�U  �'  L  ��  �=  �	�    eu  �`$  (4sz  "  4tZ  R!   Y  }4^  V  �B  X�;  K  V  8#  C#   0�  [kt    p  {  8#  �    �I  _p3  �  �  8#    �    �  c"u  �  �  8#     0V  g�c    �  �  8#    �    ~ZD  lC#   4sz  "  4tZ  R!   J�v  �+i	  J�D  �7Y  J�D  �7	  Smv  �  �~  �  V  \  p$   �~  e/  q  �  p$  	  "   �~  GZ  �  �  p$  "   Y�~  !�b  �  �  p$  {$   �~  #�.  �  �  p$  �$   �~  (�Y  �    p$  5    &�  - R  �$    %  p$  4   �~  2J�  :  @  p$   |  8�Y  U  [  p$   &f3  >C  �  t  z  p$   &Gc  B=K  �  �  �  p$  "   �1  G	"   e3  H�  4tZ  R!   4  �  
i  �  �  T 5   �  �   8`)  �zZ    F    ]  8  2#   8`)  �O'  ;  F    �  8  2#   ZV  3��  e  T   F    >  2#   Z�  3�%  �  T �  F    �>  2#   Wvo  
j  �?  T �   �?  �?    �  �/  )7�  �  )>  �  )An  �  )1c    �  �  �   �  ��   o E  �6  �std  �  �  �  1q  �  "�  �   �  �  /  S  Y  �    �  q  /  q  w  �   T �  [v �      �  �  1q  �  "�  �   �  ,  �  �  �  �    �  �  �  �  �  �   T �  [v �   �  2  �0  1q  ��  T 5   \�  ]�    �  �]  1q  ��  T 5   \�  ]    ^6  ��  �  ^6  �?  �   l  �  )  "  �  )F  �  �  <�  	@�A     Z   �  =�  <�  	��B     �  �  �  �  <   K5   3  K�  �  3  5   5   8     _:    _�  =  �  X  =F  |  Q  c  �<�  	R�A     Dr  &!  <&  �  �<&  
9(  �  �  &!   C�  '%  �  &!  �    `D  +�  �  `�  ,�  �  7\z  5      %�   %σ  %�=  %�^  %mS   �1  b   /it �   /end �  ac  7�  �  T   Z   �"   C Z    fT  �   /it �"   /end F  ac  �3  �  �   �   �"   C Q   �z  	
�:  �  �   T �  �  C    p  	
�B  D  �   T D  �  C   ,R  	
ׁ  �D   !  T �D  �  C   U�  �  6	  6.	  i	  6!  !
  i	  6  #Q  �!  #Q  C|  s!  y!  "   ,#Q  �B  �!  �!  "  "   -�   k  "  �!  �!  "  "   �~  �A  �!  �!  "   |  �  �!  �!  "   3̀  5     R!  R!  "  �!  R!  H  l"  �map vU  �   @"  K"  l"  �    C]   �f  ["  l"  �   �     "   �"  �z  �    F�  �   �:  �       �   Q  =�"  b   S   �"  !�    E�"  �G  r"   F�"  <�"  
        ��Q3  ��  	�C     �  #     !#  �     '  8#  Y  C#  �  N#  a  �  f  e#    f    |#  r
  �#    r
  N#  �  �#  	  �#  �  �#  T  �  e#  Y  �#  �  "  "  Y  �   
$  !�    �#  )�{  ?  )�7  m  )f  {  )]f  �  b=Y  �   �b�N  �   �Vn  �     )�7    �  p$  !�    4  p$  �  K4  4  �    6]  6o  �9w  PJ@            ���  !J@     /       ��$  �  �5   �lp  �5   �h 	�  %  6@     �       �1%  �  '#  �hs 
'S   �d .�  95@     (       �n%  T 5   a �  �hb #�  �` �  h�@     1       ��%  "O  Ze#  �h 	p  �%  Ȗ@     �      ��%  �  �#  ��n e#  ��u e#  �Xv e#  �Pw e#  �H 	O  &  (�@     �      �e&  �  �#  ��n �e#  ��u �e#  �Xv �e#  �Pw �e#  �H .3
  �@            ��&  T f  "O  'e#  �h .T
  
�@            ��&  T �  "O  'N#  �h 	   �&  j�@     �      �/'  �  �#  ��n N#  ��u N#  �Xv N#  �Pw N#  �H 	�  N'  ʑ@     �      ��'  �  �#  ��n �N#  ��u �N#  �Xv �N#  �Pw �N#  �H S  ��@     1       ��'  "O  ZN#  �h 0  ��@     �      ��(  P    T �   ��  N2#  ���   N$�   ���'  N1�  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#S   ��~4  P�  �Xݨ  S�(  ��
k T5   ��#�@     E       �(  
i a5   �l #8�@     -       �(  
i d5   �h e�@     0       
i f5   �d  S   �(  !�    	R  )  ��@     V      �S)  �  �#  �Xn �N#  �Ptl  �N#  �h�R  �N#  �` �  }�@            �~)  q,  =e#  �h 	.  �)  ��@     �      �{*  �  �#  ��n xe#  ��tl  {e#  �Ps �e#  �XTr  �D	  ��#��@     �       *  x �e#  �H #��@     z       0*  x �e#  �@ #K�@     Q       W*  .\  �e#  �� ��@     Q       .\  �e#  ��  �  ��@     1       ��*  "O  Ue#  �h P  j�@            ��*  q,  Le#  �h 	�  �*  "�@     H       �+  �  �#  �X"O  #e#  �P_�  $e#  �h .�  �@            �H+  q,  8e#  �h 	�  g+  ��@     V      ��+  �  �#  �Xn �e#  �Ptl  �e#  �h�R  �e#  �` 	�  �+  ��@            ��+  �  �#  �h"O  e#  �` 	A  �+  v�@            �,  �  �#  �h"O  N#  �` 	a  6,  .�@     H       �c,  �  �#  �X"O  #N#  �P_�  $N#  �h �
  �@            ��,  q,  =N#  �h 	�  �,  N|@     �      ��-  �  �#  ��n xN#  ��tl  {N#  �Ps �N#  �XTr  �D	  ��#}@     �       -  x �N#  �H #9~@     z       @-  x �N#  �@ #�@     Q       g-  .\  �N#  �� .�@     Q       .\  �N#  ��  8  |@     1       ��-  "O  UN#  �h    �{@            ��-  q,  LN#  �h .
  �{@            �.  q,  8N#  �h r  �{@     W       ��.  P    T �   ��  x2#  �h�   x!�   �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yS   �P��i$  {	�     �  �.  �.  �  T#  +�B  �g  +�=  �%�   +�U  �6�    *�.  �[  �.  F{@     K       � /  �.  �h�.  �d�.  �X�.  �P 	-  ?/  z@     7      �z/  �  �#  �Htl  �N#  �@"O  �"N#  ��*L  �N#  �X 	  �/  �x@     7      ��/  �  �#  �Htl  �N#  �@"O  �!N#  ��M�  �N#  �X 	�  �/  lx@     j       �0  �  �#  �h"O  |N#  �` y  0  K0  �  k#  +�=  ��   +�U  �)�   +$w  �65    *0  �X  n0  x@     d       ��0  0  �h&0  �`20  �X>0  �T 	�  �0  |u@     �      �1  �  �#  ��"O  e#  ���/   e#  ��tl  e#  �X�  e#  �PpU  e#  �H 6  ]u@            �91  q,  Ie#  �h 	  X1  �r@     a      ��1  �  �#  ��"O  De#  ��.\  D$e#  ��M�  Ee#  �X*L  Fe#  �Ptl  Ze#  �H 	}  �1  �q@     7      �2  �  �#  �Htl  �e#  �@"O  �"e#  ��*L  �e#  �X   �q@            �=2  q,  Ee#  �h 	X  \2  np@     7      ��2  �  �#  �Htl  �e#  �@"O  �!e#  ��M�  �e#  �X   Pp@            ��2  q,  Be#  �h 2�  �2  (p@     (       �3  �  �#  �ha �!Y#  �`b �1Y#  �X 	8  '3  �o@     j       �C3  �  �#  �h"O  |e#  �` 2j  b3  �o@            �o3  �  �#  �h 	�  �3   m@     �      ��3  �  �#  ��"O  N#  ���/   N#  ��tl  N#  �X�  N#  �PpU  N#  �H �
  m@            �4  q,  IN#  �h 	�  84  �j@     a      ��4  �  �#  ��"O  DN#  ��.\  D$N#  ��M�  EN#  �X*L  FN#  �Ptl  ZN#  �H �
  �j@            ��4  q,  EN#  �h �
  cj@            ��4  q,  BN#  �h 2  5  Rj@            �5  �  �#  �h �  �i@     �       �q5  T �   F    �  ��   �hfo �/8  �`��  �62#  �X 	�  �5  �/@     �       ��5  �  '#  �hstr 
1�  �` 	c  �5  i@     �       �6  �  I#  �H@  %8�   �@WS  +�   �Xfra -N#  �P 	%  '6  �h@     L       �46  �  v$  �h 	s  S6  �g@     �       ��6  �  �#  �X"O  �N#  �P_�  �N#  �h 	?  �6  �f@     D      �U7  �  I#  ���  45   ��WS  
�   �@�1  �   ���f  	�   �Xslb e#  ����  |#  �Pag@     ^       off �   �Hwg@     >       �  |#  ��   	  t7  :f@     X       ��7  �  �#  �X_�  pe#  �h 	�  �7  ~e@     �       �8  �  �#  �H"O  e#  �@B>  e#  �h`w  e#  �`�e@     I       M�  e#  �X  	�  -8  �d@     �       �Z8  �  �#  �X"O  �e#  �P_�  �e#  �h 2	  y8  @d@     I       ��8  �  T#  �Xp �  �P
adr �	�   �h +  �8  �8  �  �#   5�8  �c  �8  *d@            ��8  �8  �h 	@  9  �c@     O       �9  �  v$  �h 	r  19  c@     �       ��9  �  �#  �H"O  N#  �@B>  N#  �h`w  N#  �`�c@     I       M�  N#  �X  	  �9  Vb@     �       ��9  �  I#  �XWS  �6�   �P_�  �N#  �h �  �9  �9  �  v$    <    *�9  a4   :  .b@     '       �):  �9  �h �  7:  M:  �  v$  +�1  "   *):  S�  p:  �a@     2       ��:  7:  �h@:  �` �  a@     }       ��:  F    �  � ]  ��fo �78  ����  �>2#  ��   .@     *       �$;  F    �  � �  �hfo �78  �`��  �>2#  �X 	�  C;  \_@     #      �<  �  I#  ��ѷ  L/  ��q  L?�   ��WS  V�   �XCx  X4  ��fra YN#  �P#)`@     �       �;  slb _e#  �H�1  `
�   �@ku  e	  �� �`@     �       ku  s	  ��  	�  -<  �Z@     �      �@=  �  I#  ��~p �1�   ��~#�Z@     �      �<  �  �5   �\bkt �#  �P`v  4  ���  |#  ��#d[@     *      �<  slb 	e#  �H �\@     �      slb 	e#  �@Cx  #4  ��  �^@     �       @  :�   ��fra ;N#  ��Cx  =4  ��~  	�  _=  DW@     h      �>  �  I#  ��~ѷ  ~+  ��~WS  ��   �XCx  �4  ��fra �N#  �Pslb �e#  �Hbkt ��#  �@�1  �	�   ��`v  �4  ��H  ��  ���  �|#  ��   ;  �V@     E       �c>  T   F    �  3>  �H��  3!2#  �@ 	�  �>  h-@     &       ��>  �  #  �h/&  
M�  �` �  e  �,@     E       ��>  T �  F    �  3�>  �H��  3!2#  �@ -  �>  ?  �  '#  +�)  
#   5�>  �  5?  �,@     4       �F?  �>  �h?  �` "  T?  g?  �  �    <    5F?  6.  �?  �+@            ��?  T?  �h   �?  �?  �  �   5�?  9*  �?  �+@            ��?  �?  �h �   .�  �V@     +       �@  T �   a �?  �hb #�?  �` 	�  9@  �V@     0       �f@  �  >#  �hѷ  g  �`j  g)�   �X 	V  �@  |V@     (       ��@  �  >#  �h@  [�   �` 	�  �@  RV@     )       ��@  �  >#  �hѷ  c  �` �  TU@     �       �mA  @  W0�   ��
tc Y�   �`
e b�   �X
f c�   �P
ip d�   �H
is e�   �@�U@     :       
i [�   �l  .�  �T@            ��A  idx H6�   ��
tc J�   �h
s O5   �d
ip P�   �X
is Q�   �P
f R�   �H 	F  B  �T@     )       �B  T   �  '#  �h�  
  �` 	�  >B  �+@     ,       �SB  �  '#  �h>�  �  	p  yB  4+@     )       ��B  T �  �  '#  �h�  
�  �` �  �B  �B  �  '#    <    5�B  *$  �B  (+@            ��B  �B  �h 	�  C  �*@     )       �C  �  #  �` M   =C  �   �R@           ��C  T �  str 	
�  ���;  	
#C  ��Lret 	1�T@        D  	�B     �'  	�  ��JC  	�  �`
dot 	�  ��
end 	�  ���Q  	�  ��
tmp 	�  �XM�  
d 	"�  �@  Z    D  !�    �C  i	  �   CP@     L      ��D  T D  str 	
�  ���;  	
#C  ��Lret 	1[R@        D  	�B     �'  	�  �[JC  	D  �l
dot 	�  �P
end 	�  �H�Q  	�  �@
tmp 	�  �`M�  
d 	"D  �\  J  �   �M@     M      ��E  T �D  str 	
�  ���;  	
#C  ��Lret 	1P@        D  	�B     �'  	�  �WJC  	�D  �h
dot 	�  �H
end 	�  �@�Q  	�  ��
tmp 	�  �`M�  
d 	"�D  �X  �  �E  �E  �  �  +�  *�   *�E  %'  F  �)@     V       �F  �E  �h�E  �` �   F  3F  �  �    <    *F  g  VF  �)@            �_F   F  �h >  mF  wF  �  �   *_F    �F  �)@     #       ��F  mF  �h $�~  ��D  �I@     3       �
G  �2  �*�  �h�;  �EC  �`loc �V�   �X  G  	HB      Z   G  !�    
G  $ �  �5   %I@     �       ��G  out ��G  �H)�  �'�   �@@  �5�   ��p �  �X  �G  	8B        Z   �G  !�    �G  $�  ~  OH@     �       �H  ptr ~  ��~@  ~!�   ��~�2    �h $L  u  �G@     �       �KH  @  u�   ��~�2  v  �h ��  j�F@     �       �}H  ptr j  ��} $�_  d�   |F@     3       ��H  �^  dM   �h��  d<L  �`�1  dN�   �X  G  	(B      $�1  L�   ?E@     =      �J  wcs L�"  ��mbs L+�  ���t  L7�   ��cc MJ  �hst Nr"  �P  O   �@�1  Pb   ��  G  	B     #�E@     N       �I  @  S
�   ���E@     H       e T�  �d  �E@            e Y
�  �`CF@     7       n ]
�   �X    !  $>  G5   E@     .       �pJ  �.  GM   �hwc G"Q  �d  �J  	B      Z   �J  !�    pJ  $�p  >5   �C@     1      ��J  wc > �"  ��~mbs >;�  ��~�1  >G�   ��~  �J  	B      $J  /5   �B@           ��K  mbs /�  ���p  /#�   ��cc 0J  �Xwc 1
Q  �P  2   �@�1  3b   ��  �K  	B     wC@     Z       e :
�  �T  Z   �K  !�    �K  $�1  *	�  �B@     /       �L  �   *�  �h�  *+�  �`  �K  	�B      $�1  &e  ~B@     /       �iL  �   &�   �h�  &�   �`  yL  	�B      Z   yL  !�    iL  �div  1  XB@     &       ��L  �    5   �\�   5   �Xr !1  �h $G  �  -B@     +       �M  �   �  �h  �K  	�B      $G  �   B@     +       �_M  �   �   �h  yL  	�B      �abs 5   �A@     *       ��M  �   5   �l  �M  	�B      Z   �M  !�    �M  N�f  ��@@           ��N  V �  ����  ��   ��@  �-�   ���K  �	O  ���@@     �       i  �   �h�@@     �       u 	  �PA@     �       j �   �`&A@     �       v 
  �H9s  
M   �@w  	
M   ��jA@     V       k 
�   �X|A@     =       yu  
S   ��       �5   O  ]  ]   �N  3]  �  �?@     �       ��O  key �]  ��V �,]  ����  �9�   ��@  �G�   ���K  �	O  ��
i �	�   �h
j �	�   �`   D  	�B     @@     |       
k �
�   �Xkz  ��  �P
res �5   �L  wu  �M   �?@     +       �5P  >M   �h  �J  	�B      �`  �5   �?@     +       �zP  �^  ��  �h  �J  	�B      ?�v  �e?@     *       ��P  x  �5   �l  �P  	�B      Z   �P  !�   
 �P  ?gS  �P?@            ��P  x  �5   �l ?�v  �6?@            �,Q  x  �5   �l �v  �5   ?@     +       �qQ  >x  �sQ  �h  �Q  	�B      �qQ  Z   �Q  !�    yQ  #  �5   �>@     )       ��Q  >x  �sQ  �h ?�B  ��>@     #       ��Q    �K  	�B      f  �  i>@     V       �BR  ��  ��   �X@  �#�   �P
ptr �  �h w  �   >@     I       ��R  [/  ��   �X@  �.�   �P
ptr �  �`
ret �5   �l N��  ��=@     Z       ��R  >�   ��~ N+|  ��=@     "       ��R  s ��   �l 	P  �5   y=@     +       �3S  >�"  �h  �J  	�B      ��R  �5   _=@            �Tf  �?  4=@     +       ��S  �^  �4�  �hend �NC  �`V �W5   �\ �Q  [�   �:@     G      �jT  �2  [.�  ���;  [FC  ��V [R5   ���t  ]�   �P
s _jT  �h
acc `�   ��
c a5   �d}~  b�   �H
neg c5   �`
any c5   �\�Q  c5   �D r   �2  V�  �:@     +       ��T  �^  V*�  �hend VDC  �`V VM5   �\ Yw  0�   x9@     J      �AU  �^  0$�  �Xend 0>C  �PV 0G5   �L  �J  	�B     �'  ;�  �oJC  G�   �` �1  -�  ?9@     9       ��U  �^  -,�  �hend -FC  �` 2w  *D  9@     %       ��U  �^  *%�  �hend *?C  �` +w  '�D  �8@     3       �V  �^  '&�  �hend '@C  �` �Q  $�  �8@     $       �6V  �^  $�  �h �=  !�   �8@     $       �hV  �^  !�  �h �=  5   {8@     $       ��V  �^  �  �h �9  �D  N8@     -       ��V  �^  �  �h 2�!  �V  �M@            ��V  �  	"  �h 	�!  W  �M@     B       �7W  �  	"  �h  yL  	1B      .7  �M@            �`W  x )�   �h v	  nW  xW  �  <!   5`W  1~  �W  :M@     Q       ��W  nW  �h 	_  �W  M@     6       ��W  �  &  �`c 63�  �\�>  78  �h c�  2�W  X  �  &    <    *�W  .  4X  �)@            �=X  �W  �h   c  2TX  cX  �  &  =X   *CX  �  �X   )@     �       ��X  TX  �h]X  �` E  �X  �X  �  &   *�X  K  �X  �(@     \       ��X  �X  �h �.  ^    �(@            �Y  @  #�   �hp /  �` 2L  >Y  4K@     �      �Z  �  �  �H��0   Z  �P
res 3�   �X_K@     N      
y -�   �\#_K@     {       �Y  
kk #5   �loK@     e       
y $�   �d  �K@     {       
kk (5   �h�K@     e       
y )�   �`    �   Z  !�    Z  2-  ?Z  �J@     �       �YZ  �  �  �hs �   �d   gZ  qZ  �  �   *YZ  /  �Z  fJ@             ��Z  gZ  �h d�    "df    " �   �  �  ^�  �  �
          �K  3�  e6   �  6   L�  	
N   �  �  �  �N   �  E  6  �  �  �  
6   �  �  int �   3  �    �   	�z  �    	F�  �   	�:  6    
std  h  �  m  q  o  �  h  �  �    9  ?  }   �  q    W  ]  }   T h  v h    �   �  �  q  o  �  h  �  ,  �  �  �  �   �  �  �  �  �  �   T h  v h   r  2  �  q  �o  T �   �  �
    �  �C  q  �o  T �   �  �
    6  ��  o  6  �?  o   l  h      m  F    �  frg 	2
  �  �  o   �  �   �  .  7G
   %  �   ,�  �   �  hex  �  I  �  {T  �  |�    �  ~;  2  8  g
   !�    H  g
  �     ")    i  o  r
   ")  a  �  �  r
  #�   ")  �  �  �  r
  #}
   ")  �  �  �  r
  #�
   ")  *�  �  �  r
  #�
   ")  0x      r
  #�
   "(  8  $  /  r
  �    $�  =O  �
  H  S  r
  #�   $c  Q�  h  l  r  �
   $c  T�  h  �  �  r
   $m  X�  h  �  �  �
   $R  \+  }
  �  �  �
   $R  `[  �
  �  �  r
   $!  d�  �
      r
    f  �  !  '  r
   	�  �   	�  �h  T �    �  �*  2   �*  3Z(  o  u  �
   	   6C  N  �  �  �
  #�   	   <�   	�  =�   	�)  >�  	�   ?h  	�'  @h  	�#  Ah  	<  Bh  	�  Ch  %�*  E&    �
  �     &p  J�  �  "o�  ׈  C  I  �
   "o�  ��  ^  i  �
  #A
   "o�  �  ~  �  �
  #A
  #\    $�  �  A
  �  �  �
   $�  #��  �
  �  �  �
  #\    $@  '	7�  \   �  �  �
   $
�  +p�  h  	    �
  #!   $�  3�  h  -  8  �
  #!   $��  7	
�  \   Q  a  �
  #L
  #\    $Ĉ  ?	ȉ  \   z  �  �
  #L
   $R�  G�  !  �  �  �
  #\   #\    	з  XA
   	o Y	\   '�  L
   !  �  
�  �  �  �  �	   �)  E#      X  #   q,  �	j	   q,  �#  >  I  c  #X   (q,  _   ]  h  c  #n   )�  	~-  t  �  �  c  #n    p,  �*  �  �  c  �    )  "	�  t  �  �  c  #�    �$  'a&  �  �  c  #L
    �$  1�   	  	  c  #A
   *�)  >X   *ܨ  ?z  *7&  @
\   �*)  Ah  �+c.  	�*  t  ^	  T A
  c  #A
      �  H`*    �	  �	  X   "�#  M�"  �	  �	  X  #A
   *.  Q   'U(    ,].  N   � -�  .`)  �O'  �	  F   #A
  #N  #t   /�  3�%  %
  T A
  F   #Z  #t   u�  \!!   0�  	�B     S
  A
  �  L
  0�  	��B       g
  �  r
  1�   2�   1I  2�  1�  I  1�   �   N  �
  3:  �  3�  #  �  !  �
  �  �
  1S
  |  0�  	�B     4r  �  <&  U  5<&  
9(  3  9  �   !�  '%  I  �  #A
    6D  +�  �  6�  ,�  �	  \z  �   �  �   σ  �=  �^  mS   �1  �  7it A
   7end A
  8c  7�  h  �  �  �   C S
   �  >  7it �   7end �  8c  օ  h  0  6  �   C 6    � qp  +w�  r��  u  _  �  #�
  #�    f�  #�   9� �  +w�  0K�  u  �  �  #L
  #�    :(�  "��  h  #p      �  6   =   �  >  1p  ;P  <6   ���   A�  ��  ]�  ��  u�  ^�  U�  �  �  	��  
��  )�  ��    =��  �  X    c  1j	  1  >L
  �  ?N    @C  @U  A�  �  �/@     �       ��  B�  i  �hCstr 1A
  �` D�	  .@     *       �  F   E�  � A
  �hCfo �7N  �`E��  �>t  �X A�	  >  h-@     &       �Z  B�  ^  �hE/&  MA
  �` 1G
  D�	  �,@     E       ��  T A
  F   F�  3Z  �HF��  3!t  �@ G*  �  �  H�  i  I�)  X   J�  �  �  �,@     4       �  K�  �hK�  �` G8    #  H�  m
  H  �    J  6.  F  �+@            �O  K  �h G  ]  g  H�  m
   JO  9*  �  �+@            ��  K]  �h A�  �  �+@     ,       ��  B�  i  �hL�  �  AC	  �  4+@     )       �	  T A
  B�  i  �hE�  A
  �` G�    *  H�  i  H  �    J	  *$  M  (+@            �V  K  �h Ao	  u  �*@     )       ��  B�  ^  �` M�  �  4�@            ��  B�  �
  �XE�  +%!  �@Ne�@     G       Oi .\   �h  GI  �  �  H�  �
  Pcs  A
   J�  ~�  "  �@     R       �3  K�  �hK�  �` G  A  T  H�  x
  H  �    Q3  g  w  �)@            ��  KA  �h GT  �  �  H�  x
   Q�    �  �)@     #       ��  K�  �h R��  #)   |�@     *       �  L)   �lS    	`B      >S
    ?N      R:�  )   R�@     *       �W  L)   �lS    	PB      R �  �   �@     Q       ��  Tnc �   �\Ucc �  �hUcp p  �`N�@     &       Ue 
u  �d  |  �  R�  
�   ��@     Q       �D  Tnc 
�   �\Ucc �  �hUcp p  �`NĤ@     &       Ue 
u  �d  RΈ  �   ��@     .       ��  L)   �lLB   �`S    	@B      VЈ  �
B   ��@     �      ��  Ccs �A
  ��|Os �%
  ��} V�  ��   q�@     H       �7  Cnc �)   �\Occ ��  �hOcp �p  �`N��@     %       Oe �
u  �d  V��  ��   �@     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N2�@     %       Oe �
u  �d  V�  ��   ˟@     S       �  Cnc �)   �\Occ ��  �hOcp �p  �`Nߟ@     %       Oe �
u  �d  VU�  ��   x�@     S       �{  Cnc �)   �\Occ ��  �hOcp �p  �`N��@     %       Oe �
u  �d  V��  ��   %�@     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N9�@     %       Oe �
u  �d  V��  ��   Ҟ@     S       �S  Cnc �)   �\Occ ��  �hOcp �p  �`N�@     %       Oe �
u  �d  V��  ��   �@     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N��@     %       Oe �
u  �d  VD�  ��   ,�@     S       �+  Cnc �)   �\Occ ��  �hOcp �p  �`N@�@     %       Oe �
u  �d  V�  ��   ٝ@     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N�@     %       Oe �
u  �d  Vև  ��   ��@     S       �  Cnc �)   �\Occ ��  �hOcp �p  �`N��@     %       Oe �
u  �d  V;�  ��   3�@     S       �o  Cnc �)   �\Occ ��  �hOcp �p  �`NG�@     %       Oe �
u  �d  V��  x�   ��@     S       ��  Cnc x)   �\Occ y�  �hOcp zp  �`N��@     %       Oe {
u  �d  VC�  l�   ��@     J       �G  Cnc l�   �\Occ m�  �hOcp np  �`N��@     (       Oe o
u  �d  V��  d�   K�@     K       ��  Cnc d�   �\Occ e�  �hOcp fp  �`N_�@     (       Oe g
u  �d  V�  \�   ��@     V       �  Cnc \�   �\Occ ]�  �hOcp ^p  �`N	�@     (       Oe _
u  �d  V��  T�   ��@     V       ��  Cnc T�   �\Occ U�  �hOcp Vp  �`N��@     (       Oe W
u  �d  V]�  L�   I�@     V       ��  Cnc L�   �\Occ M�  �hOcp Np  �`N]�@     (       Oe O
u  �d  Vm�  D�   �@     V       �c  Cnc D�   �\Occ E�  �hOcp Fp  �`N�@     (       Oe G
u  �d  VJ�  <�   ��@     V       ��  Cnc <�   �\Occ =�  �hOcp >p  �`N��@     (       Oe ?
u  �d  VM�  4�   G�@     V       �;  Cnc 4�   �\Occ 5�  �hOcp 6p  �`N[�@     (       Oe 7
u  �d  V��  ,�   �@     V       ��  Cnc ,�   �\Occ -�  �hOcp .p  �`N�@     (       Oe /
u  �d  V�  $�   ��@     V       �  Cnc $�   �\Occ %�  �hOcp &p  �`N��@     (       Oe '
u  �d  V��  �   E�@     V       �  Cnc �   �\Occ �  �hOcp p  �`NY�@     (       Oe 
u  �d  Ve�  �   �@     V       ��  Cnc �   �\Occ �  �hOcp p  �`N�@     (       Oe 
u  �d  Vg�  �   ��@     V       �W  Cnc �   �\Occ �  �hOcp p  �`N��@     (       Oe 
u  �d  W�  ��@     0       ��  Cc "*p  �l A�  �  ��@           �8  B�  �  ��Cnc 0L
  ��Cwc 0-�  ��Ouc 1{   �oX  7�  �PX�1  8�  �@Ost 9�   ��S  H  	8B     N%�@     .       Oe ;u  �h  >S
  H  ?N    8  Y   2^  q  H�  �
  H  �    QM  .  �  �)@            ��  K^  �h G[  �  �  H�  �
   Q�  K  �  �(@     \       ��  K�  �h i	  J   �T   P  ^�  �  �            �T  1�>  5   _int 5   1Q  M   
X   M   �  X   1�o  M   �  ��   p   �  `�  �  �  �   I @'    M       	p   �  #	p   �  &	p     )	p    �  ,	p   (�  -	p   0
  25   8�  55   < Q  8"�   1�  K?  
'  1�  L?  1�  M?  E  a6  �  i  �  �  �  �  ��     4�  �  bstd  �  �  $  -q  �  �  �  �  �  �  �  �  �   �  q  �      �   T �  Iv �    �  �  �  -q  �  �  �  �  ,  C  g  m  �   �  �  C  �  �  �   T �  Iv �   )  2  ��  -q  ��  T 5   J�  K�%    �  ��  -q  ��  T 5   J�  K�%    ��  `  �U  a5  T �D   ��  `<  �U  aM   T �'   L6  ��  �  L6  �?  �  -�  j>   �  !�  `  �  T �D  �D   5+�  =�  �  T M   �'  �'   -�  j>(  M��  !�  �  T �'  �'    l  �  .  �  
$  .F  6  
�  cfrg '$  >E3  	  d��     ?d^  	  @J  N4j  �    A7  BG  5   w  /�   Ored /h^   �o  0/  �o  �F  �  �  1$   )�o  �D  �  �  1$  <$   *�  �z  B$  �  �  1$  <$   tl  �    �  �   pU  �   �I   �   �D  !�    [r  "R  ( w  q  %�  �Q  '!=  �  b  T t  (   M�  '1Q  �  T �  �'    dV  5	  Ph 8<  1$  �  �'   pl  =�n  �'  �  �'   �p  B�^  �'  �  �'   lU  Ef|  �'  �  �'   �I  I�  �'    �'   �D  LE  �'  (  �'   <3  Pfm  �'  @  F  /(   8�E  U�L  �  a  �'   8�_  Z�M  �  |  �'    c  djw  �  �  /(   ) c  gar  �  �  /(  :(   *�  i
J  @(  �  �  /(  :(   ��  op  �'  �  �  /(   �D  |+G      /(  �'   ��  ��z  +  ;  /(  �'  �'   5>  ��@  P  `  /(  �'  �'   �F  �4\  u  �  /(  �'    �  Dj  �  �  /(  �'   O  $d  �  �  /(  �'  �'   �U  D�6  �  �  /(  �'  �'   �  x�E      /(  �'    q  �nq  #  .  /(  �'   �9  1y  D  O  /(  �'    �=  Ӏ  d  o  /(  �'    �z  #�8  �  �  /(  �'   0L  0Nx  �  �  �  /(   0L  9�/  �  �  �  /(  �'  �%  F(  F(   2?3  ��    D 	  T �  9�P  �T  A 4   �  Q�5  ��	  !��  !�  !�;  !��  !��  !�(  C�    Z|  �@  v	  �	  W(  �    �F  �V�  �	  �	  W(  �'   2�R  ��  T �  9�P  �T  L �  A 4   .H  5b  Ph 8�4  1$  �	  (   pl  =&i  (  
  (   �p  B�Z  (  *
  (   lU  EP  (  D
  (   �I  I�f  (  ^
  (   �D  L}S  (  x
  (   <3  PO]  (  �
  �
  b(   8�E  U�g  �  �
  (   8�_  Z)?  �  �
  (    c  d8  �
  �
  b(   ) c  g~u  �
    b(  m(   *�  i'O  s(    (  b(  m(   ��  oAs  (  @  F  b(   �D  |�k  [  f  b(  (   ��  ��0  {  �  b(  (  (   5>  ��A  �  �  b(  (  (   �F  �X  �  �  b(  (    �  �1  �  �  b(  (   O  
e      b(  (  (   �U  DxT  ,  <  b(  (  (   �  xfC  R  ]  b(  (    q  �{l  s  ~  b(  (   �9  E}  �  �  b(  (    �=  �9  �  �  b(  (    �z  #�`  �  �  b(  (   0L  0�_  �  �  �  b(   0L  9�a  �    3  b(  (  �%  y(  y(   2?3  ��    D g  T t  9�P  �T  XA 4   �	  e�~  �!�F  !�f  !��  !�
  !�*
  !�x
  C�	    Z|  �<R  �  �  (  �    �F  �/L  �  �  (  (   2�R  ��  T t  9�P  �T  XL �  A 4    @0  N4j  �    A  /�  g  fclz �3  5   _  �    T �    g��  �$0  B Q  5   ��  /�   /ʃ  /QS   u  �U  H�	o  �U  ���  �  �  �'  u  �  p    )�U  ���  �  �  �'  (   *�  �
`D  (      �'  (   ��  ��b  �  /  :  �'  �    �U  ��   WS  ��  p �|   �=  �A!   �  �U  ��	'  C�   �U  �Pc  �  �  (  �  p   5    )�U  �z  �  �  (  (   *�  �4  (  �  �  (  (   �  �<   H�D  ��   L$H  �$(  P�B  �A!  X t  %\  �	�  %\  �/  M  S  $(   )%\  �l5  g  r  $(  4)   *�  ��h  :)  �  �  $(  4)   �E  �$(    ,  �R  �	�  R�  ��v  �  �  L(  (  (    �.   �	)  �.  �R�  �    �(   �E  �	M$   �o  �(  �e  �)   1|  �N!  u  ��=  J  U  �'  �(   Su  (�t  j  u  �'  �(   h�  *�K  �(  �  �  �'  �(   �  ��o  �   �  �  �'  p    0�  L�g  �   �  �  �'  �   p    �  ~��  �    �'  �    �I  �Ճ    .  �'  �   p    WV  1	e;  p   G  M  �'   iC  >�(                         @       D�v  @ �   D�`  A �    �~  H�U  p   �  �    �.  W�N  p   �  p    DQC  j<   -zz  l|   |  oK>  �     �    -́  ||   -]C  |   j�D  �|    E�~  ��<  �'  B  M  �'  �   E��  &q  (  f  q  �'  5    EFS  %n^  �'  �  �  �'  p     4  7:k  �  �  �'    ]  >�J  �  �  �'  �'   �[  �
�(   �1  �M$  �U  �[!  L  ��  �=  �	p    eu  �)  (+sz  %  +tZ  M$   g  k4^  V  �B  X�;  Y  d  �'  �'   0�  [kt  �   ~  �  �'  p    �I  _p3  �  �  �'  �   p    �  c"u  �  �  �'  �    0V  g�c  �   �  �  �'  �   p    lZD  l�'   +sz  %  +tZ  M$   >�    To   $  m�   P  n.  7�%   B%  5   ,u  /�   /�  Ohex  :�  �  o�  {�  p�  |5   �  ~;  �  �  �%   F�    �  �%  5     )    �  �  �%   )  a      �%     )  �  !  ,  �%  �%   )  �  A  L  �%  �%   )  *�  a  l  �%  �%   )  0x  �  �  �%  �%   (  8  �  �  �%  5    �  =O  �%  �  �  �%  u   c  Q�  �  �  �  �%   c  T�  �      �%   m  X�  �  '  -  �%   R  \+  �%  F  L  �%   R  `[  �%  e  k  �%   !  d�  �%  �  �  �%   f  �  �  �  �%   �  ��   �  ��  T 5    u  �*  2�  �*  3Z(  �  �  �%   	   6C  �  
    �%  P      <P   �  =5   �)  >u  �   ?�  �'  @�  �#  A�  <  B�  �  C�  q�*  E&  �  �  �%  5    r�*  >  �  �%  �R    �  ?p  Jm  5�-  N�!    P �  T �   �'  �   �  5   5   5   X    5�'  x<+  B  P �  T �   �'  �   5   5   5   X    s�  ��+  T �   F �  �   �  �'    :�    o�  ׈  �  �  &   o�  ��  �  �  &  {%   o�  �  �  �  &  {%  p    �  �  {%  �  �  &   �  #��  &      &  p    @  '	7�  p   6  <  &   
�  +p�  �  U  `  &  m   �  3�  �  y  �  &  m   ��  7	
�  p   �  �  &  X   p    Ĉ  ?	ȉ  p   �  �  &  X    R�  G�  m  �  �  &  p   p    з  X{%   o Y	p   +�  X    m  Qj�  u   j�  "��  F  V  $&  /&  p    2ܨ  &/&   2@  '	p    #  >�  	
z  T�  	�  �  	�  �)  	E#  �  �  e'  Q&   q,  �		7  q,  	�#  �  �  p'  e'   )q,  	_        p'  {'   *�  		~-  �'  #  .  p'  {'   p,  	�*  B  M  p'  5    )  	"	�  �'  e  p  p'  z   �$  	'a&  �  �  p'  X    �$  	1�  �  �  p'  {%   3�)  	>e'   3ܨ  	?�'  37&  	@
p   �3)  	A�  �d�  		u�  �'      T #  p'  #   Rc.  		�*  �'  +  T {%  p'  {%    �  �  	H`*  �  T  Z  e'   �#  	M�"  o  z  e'  {%   3.  	QQ&   +U(  Q&  t].  �   � u�  :<�   
<!  Ɍ  
�A�  �  �  �'  5   Ɍ  
��  �  �  �'  �'   Ɍ  
$ď      �'  �'   ��  
�Ќ  #  .  �'  5    �  
+
n�  �'  G  R  �'  �   �  
�R�  �'  k  v  �'  �'   �  
�J�  �'  �  �  �'  �'   p�  
4��  �'  �  �  �'  �'   p�  
8��  �'  �  �  �'  �'   Gpop 
��  M   �    �'   �  
D��      �'   �  
J��  _'  5  ;  �'   �  
Nٕ  �'  T  Z  �'   @  
R	@�  p   s  y  �'   ��  
V��  �  �  �  �'   ݱ  
Z��  _'  �  �  �'   ݱ  
^��  �'  �  �  �'   Gend 
b�  _'  �  �  �'   Gend 
f7�  �'        �'   *  
j�  �'  -   3   �'   *  
m�  �'  L   R   �'   �  
q��  �'  k   q   �'   �  
tJ�  �'  �   �   �'   �  
x�  �'  �   �   �'  p    �  
{P�  �'  �   �   �'  p    T�  
��  �   �   �'  p    C  
�5   �  
�_'  @  
�	p   [�  
�	p   T M   +H  5   �  H�v  �+w  H�D  �7g  H�D  �7	  :mv  �"  �~  �  �!  �!  )   �~  e/  �!  �!  )    %   �~  GZ  �!  �!  )  %   S�~  !�b  �!  �!  )  ")   �~  #�.  
"  "  )  ()   �~  (�Y  *"  5"  )  5    �  - R  .)  N"  Y"  )  h!   �~  2J�  n"  t"  )   |  8�Y  �"  �"  )   f3  >C  �  �"  �"  )   Gc  B=K  �  �"  �"  )  �$   �1  G	�$   e3  H�  +tZ  M$   h!  �  
i  �%  !#  T 5   �%  �%   5`)  �@%  H#  F �  �   �  �'   ;N#  8��  w#  T �   F �  �?  �  �'   ;`)  ��  �#  F �  #  �  �'   5`)  �O'  �#  F �  {%  �  �'   ;e�  3ˑ  �#  T #  F �  rE  �'   ;�  3�%  $  T {%  F �  �E  �'   u�  \!m   6  6<  
w  1$  /  w  6"  #Q  �$  #Q  C|  n$  t$  �$   )#Q  �B  �$  �$  �$  	%   *�   k  %  �$  �$  �$  	%   �~  �A  �$  �$  �$   |  �  �$  �$  �$   3̀  5     M$  
M$  �$  �$  M$  H  f%  vmap vU  �  :%  E%  f%  p    F]   �f  U%  f%  �  p     
%  <)  	�B     
_   {%  <B  	��B     
�  �%  
u  �%  <   75   �  7u  u  
�  5   
5   
�  �%  U:  �  U�  �  �  
m  &  
  &  _   |  
#  $&  
5&  w<�  	�B     ?r  �&  <&  �&  x<&  
9(  s&  y&  �&   F�  '%  �&  �&  {%    VD  +�  �  V�  ,�  �   
Q&  @"'  y%�  *'  WR�  O�&  $   WT�  <�&  $  {%  �   z  -{z�  ('�'  |��  p   $    A�&  %M   :'  &�     <�&  	�C     }�  _'  	@ C     
M   
�  e'  
�  p'  7  �  %X   �'  &�    
5  �'  
g  �'  
�  �'  <!  7�  �  M   S   7M   
S   
<!  �'  ~&  �   
�  �'  o  �  
t  (  '  t  
,  $(  
�  /(  	  �  �'  
�  L(  
	  W(  
�	  b(  b  �	  (  
g  (  
�  %  0  g  %|   �(  &�    �(  .�{  M  .�7  {  .f  �  .]f  �  X=Y  �   �X�N      Vn       .�7    %�  )  &�    
h!  )  �"  7h!  h!  �  ,  6<  6N  '�"  95@     (       ��)  T 5   a �%  �hb #�%  �` �
  h�@     1       ��)  "O  Z(  �h �  �3@     �      ��*  P �  T �   ��  N�'  ���   N$�   ���'  N1�  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P{%  �Xݨ  S�*  ��k T5   ��#�4@     E       �*  i a5   �l #�4@     -       �*  i d5   �h 5@     0       i f5   �d  %X   �*  &�    `  +  ��@     V      �E+  �  5(  �Xn ��'  �Ptl  ��'  �h�R  ��'  �` <  d+  ��@     �      �B,  �  h(  ��,n x(  ��	tl  {(  �Ps �(  �X	Tr  �R  ��#��@     �       �+  x �(  �H #��@     z       �+  x �(  �@ #K�@     Q       ,  	.\  �(  �� ��@     Q       	.\  �(  ��  ~  a,  Ȗ@     �      ��,  �  h(  ��,n (  ��u (  �Xv (  �Pw (  �H ]  �,  (�@     �      �-  �  h(  ��,n �(  ��u �(  �Xv �(  �Pw �(  �H �
  ��@     1       �9-  "O  U(  �h �	  }�@            �d-  q,  =(  �h 'A  �@            ��-  T t  "O  '(  �h 'b  
�@            ��-  T �  "O  '�'  �h .  �-  j�@     �      �..  �  5(  ��,n �'  ��u �'  �Xv �'  �Pw �'  �H   M.  ʑ@     �      ��.  �  5(  ��,n ��'  ��u ��'  �Xv ��'  �Pw ��'  �H a  ��@     1       ��.  "O  Z�'  �h   �1@     U       �R/  P �  T �   ��  x�'  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �TY�i$  {	�     �  `/  �/  �  �'  $�B  �u  $�=  �%�  $�U  �6p    "R/  �[  �/  F{@     K       ��/  `/  �hi/  �du/  �X�/  �P ;  �/  z@     7      �,0  �  5(  �Htl  ��'  �@"O  �"�'  ��*L  ��'  �X   K0  �x@     7      ��0  �  5(  �Htl  ��'  �@"O  �!�'  ��M�  ��'  �X �  �0  lx@     j       ��0  �  5(  �h"O  |�'  �` �  �0  �0  �  (  $�=  ��  $�U  �)p   $$w  �65    "�0  �X   1  x@     d       �A1  �0  �h�0  �`�0  �X�0  �T �  `1  |u@     �      ��1  �  h(  ��"O  (  ���/   (  ��	tl  (  �X	�  (  �P	pU  (  �H   �1  �r@     a      �?2  �  h(  ��"O  D(  ��.\  D$(  ��	M�  E(  �X	*L  F(  �P	tl  Z(  �H ^
  j�@            �j2  q,  L(  �h �  �2  "�@     H       ��2  �  h(  �X"O  #(  �P	_�  $(  �h D
  ]u@            ��2  q,  I(  �h '�	  �@            �3  q,  8(  �h �  +3  ��@     V      �c3  �  h(  �Xn �(  �Ptl  �(  �h�R  �(  �` �  �3  ��@            ��3  �  h(  �h"O  (  �` O  �3  v�@            ��3  �  5(  �h"O  �'  �` o  �3  .�@     H       �'4  �  5(  �X"O  #�'  �P	_�  $�'  �h �  �@            �R4  q,  =�'  �h �  q4  N|@     �      �O5  �  5(  ��,n x�'  ��	tl  {�'  �Ps ��'  �X	Tr  �R  ��#}@     �       �4  x ��'  �H #9~@     z       5  x ��'  �@ #�@     Q       +5  	.\  ��'  �� .�@     Q       	.\  ��'  ��  F  |@     1       �z5  "O  U�'  �h   �{@            ��5  q,  L�'  �h '�  �{@            ��5  q,  8�'  �h B  �0@     �       �'6  T �   F �  �  ��   �lfo �/�  �`��  �6�'  �X q  F6  i@     �       ��6  �  �'  �H@  %8p   �@	WS  +�  �Xfra -�'  �P �	  �6  �g@     �       ��6  �  ](  �X"O  ��'  �P	_�  ��'  �h M  �6  �f@     D      ��7  �  �'  ���  45   ��	WS  
�  �@	�1  �   ��	�f  	p   �Xslb (  ��	��  $(  �Pag@     ^       off p   �Hwg@     >       	�  $(  ��   (  �7  :f@     X       ��7  �  h(  �X_�  p(  �h �  �7  ~e@     �       �]8  �  h(  �H"O  (  �@	B>  (  �h	`w  (  �`�e@     I       	M�  (  �X  �  |8  �q@     7      ��8  �  h(  �Htl  �(  �@"O  �"(  ��*L  �(  �X *
  �q@            ��8  q,  E(  �h f  9  np@     7      �<9  �  h(  �Htl  �(  �@"O  �!(  ��M�  �(  �X 
  Pp@            �g9  q,  B(  �h �  �9  (p@     (       ��9  �  R(  �ha �!(  �`b �1(  �X F  �9  �o@     j       ��9  �  h(  �h"O  |(  �` x
  :  �o@            �:  �  h(  �h �  3:   m@     �      ��:  �  5(  ��"O  �'  ���/   �'  ��	tl  �'  �X	�  �'  �P	pU  �'  �H �  m@            ��:  q,  I�'  �h �  �:  �j@     a      �=;  �  5(  ��"O  D�'  ��.\  D$�'  ��	M�  E�'  �X	*L  F�'  �P	tl  Z�'  �H �  �j@            �h;  q,  E�'  �h �  cj@            ��;  q,  B�'  �h Y"  �;  �h@     L       ��;  �  )  �h (  �;  Rj@            ��;  �  5(  �h !#  ,.@     J       �<<  F �  �  �!�   �Lfo �8�  �@��  �?�'  �� �  [<  �Z@     �      �n=  �  �'  ��~p �1p   ��~#�Z@     �      (=  �  �5   �\bkt �(  �P	`v  h!  ��	�  $(  ��#d[@     *      �<  slb 	(  �H �\@     �      slb 	(  �@	Cx  #h!  ��  �^@     �       	@  :�   ��fra ;�'  ��	Cx  =h!  ��~  �  �=  �d@     �       ��=  �  �(  �X"O  �(  �P	_�  �(  �h   �=  @d@     I       �>  �  �'  �Xp ��   �Padr �	�   �h 9  >  >  �  *(   (>  �c  =>  *d@            �F>  >  �h t"  e>  �c@     O       �r>  �  )  �h �  �>  c@     �       ��>  �  5(  �H"O  �'  �@	B>  �'  �h	`w  �'  �`�c@     I       	M�  �'  �X  )  ?  Vb@     �       �<?  �  �'  �XWS  �6�  �P	_�  ��'  �h "  J?  ]?  �  )    <    "<?  a4  �?  .b@     '       ��?  J?  �h �!  �?  �?  �  )  $�1  %   "�?  S�  �?  �a@     2       ��?  �?  �h�?  �` �   H#  ��@     N       �B@  T �   F �  �  8�?  �H,fo 8-�  �@��  84�'  �� p  a@  6@     �       �{@  �  v'  �hs 	'X   �d �  �@  �/@     �       ��@  �  v'  �hstr 	1{%  �` d  �@  |V@     (       ��@  �  �'  �h@  [p   �` �  A  DW@     h      ��A  �  �'  ��~ѷ  ~+�   ��~	WS  ��   �X	Cx  �h!  ��fra ��'  �Pslb �(  �Hbkt ��(  �@	�1  �	p   ��	`v  �h!  ��	H  ��  ��	�  �$(  �� w#  ��@           �iB  F �  ��  '#  ��,fo <�  ����  C�'  ��p iB  �`��@     �      i p   �hҶ@     �      c 	i  �_   
p  �#  .@     *       ��B  F �  �  � {%  �hfo �7�  �`��  �>�'  �X �   �B  ��@     �       �\C  �  �'  ��\�  
�4p   ��c�  
�	p   �H��  
�_'  �@#ٵ@     ^       <C  i 
�p   �X 7�@            i 
�p   �P  �  {C  RV@     )       ��C  �  �'  �hѷ  c�   �` �  TU@     �       �'D  @  W0p   ��tc Y�   �`e b�   �Xf c�   �Pip d�   �His e�   �@�U@     :       i [�   �l  '�  �T@            ��D  idx H6�   ��tc J�   �hs O5   �dip P�   �Xis Q�   �Pf R�   �H 5  'l  ~�@            ��D  T �D  x *�D  �h �  �D  �D  �  &  Zs  {%  $p *p    (�D  c�  E  T�@     *       �7E  �D  �h�D  �`�D  �X Z  VE  h-@     &       �rE  �  k'  �h/&  	M{%  �` u  �#  �@     I       ��E  T #  F �  �  3rE  �H��  3!�'  �@ �%  �#  �,@     E       �F  T {%  F �  �  3�E  �H��  3!�'  �@ �   F  6F  �  v'  $�)  	e'   (F  �  YF  �,@     4       �jF   F  �h)F  �` �  xF  �F  �  �%    <    (jF  6.  �F  �+@            ��F  xF  �h �  �F  �F  �  �%   (�F  9*  �F  �+@            ��F  �F  �h �  G  ´@     I       �6G  �  �'  �Xkz  
�M   �h �  s�@     O       ��G  T M   x �'  �Xy �'  �Pyu  M   �h '�  b�@            ��G  T �'  x *�'  �h Z  �G  P�@            ��G  �  �'  �h R   �G  *�@     %       �
H  �  �'  �h �   )H  �@     !       �EH  �  �'  �h�  
{p   �` v  dH  ��@     �       ��H  �  �'  �Hkz  
�#�'  �@ѷ  
�_'  �X R  �H  
�@     w       ��H  �  �'  �Xkz  
�(�'  �Pѷ  
�_'  �h   �H  ֲ@     4       �$I  �  �'  �X޲@            i 
Ep   �h    CI  Ĳ@            �PI  �  �'  �h   ^I   ~I  �  �'    <   Y�i 
�p     "PI  ɐ  �I  ��@     C       ��I  ^I  �X�pI  �I  �qI   �pI  ��@            �qI  �h  �  �I   �I  �  �'  $C  
�(5   "�I  ��  "J  0�@     P       �3J  �I  �X�I  �P <  RJ  4�@            ��J  �  &  �X�  +%m  �@e�@     G       i .p   �h  �  �J  ��@     r       ��J  �  &  �X^�  G&p   �P@  G3p   �H M  �J  �+@     ,       �K  �  v'  �h�z  �  �  2K  ��@     6       �NK  T #  �  v'  �h�  	#  �P   mK  v�@            �zK  �  &  �h �  �K  d�@            ��K  �  &  �h   �K  4+@     )       ��K  T {%  �  v'  �h�  	{%  �` .  �K  	L  �  v'    <    (�K  *$  ,L  (+@            �5L  �K  �h <  TL  �*@     )       �aL  �  k'  �` �  �L  �@     S       ��L  �  &  �Xc 7X   �TX�  7#p   �H!�@     9       i 8p   �h  �  �L  �L  �  &  Zcs  {%   (�L  ~�  M  �@     R       �M  �L  �h�L  �` L  -M  CM  �  �%  $�  *�%   "M  %'  fM  �)@     V       �wM  -M  �h6M  �` �  �M  �M  �  �%    <    "wM  g  �M  �)@            ��M  �M  �h �  �M  �M  �  �%   "�M    �M  �)@     #       �N  �M  �h =��  �5   ��@     >       �:N  �  �{%  �X =��  x5   ��@     �      ��N  �  x{%  ��}q  x*{%  ��}7�  x55   ��}|�  y$  ��~s z	p   �X�^  �M   ��}4  �N  	0+B      %_   �N  &�    �N  =ҕ  m5   �@     �       �DO  �^  m{%  ��|�  n$  �@s o	p   �X4  �N  	)+B      =��  bM   G�@     �       ��O  �  b{%  ��k c�   �h|�  g$  �@s h	p   �`4  �N  	"+B      �&  ի@     r      �P  �  O)$  �@Ɍ  P�'  �X4  P  	+B     k S�   �P %_   P  &�    P  �&  ��@     ?      ��P  �  <'$  ���^  <9{%  ��7�  <F�  ��Ɍ  =�'  �X4  �P  	 +B     k @�   �P %_   �P  &�    �P  �&  ɩ@     �       ��P  Ɍ  .�'  �`�@     P       i 5p   �h  '  Z�@     o       �.Q  Ɍ  ).�  	�C      '  ��@     �      ��Q  �  ,$  ��}ا@     o      i p   �X�@     <      |�  $  ��~s 
p   �P   1  �Q  �Q  �  *&  [ݨ  "/&  [@  "(p    (�Q  ��  �Q  �@     *       �R  �Q  �h�Q  �`�Q  �X �  5R  M@     6       �_R  �  �%  �`c 63P  �\�>  7�  �h \}  2pR  �R  �  �%    <    "_R  .  �R  �)@            ��R  pR  �h �  \�  2�R  �R  �  �%  �R   "�R  �  �R   )@     �       �	S  �R  �h�R  �` �  S  !S  �  �%   "	S  K  DS  �(@     \       �MS  S  �h �.  ^  �   �(@            ��S  @  #p   �hp /�   �` �$  �S  �M@            ��S  �  %  �h �$  �S  �M@     B       ��S  �  %  �h4  T  	�*B      %_   T  &�    �S  'E  �M@            �:T  x )�   �h �  HT  RT  �  7$   (:T  1~  uT  :M@     Q       �~T  HT  �h i	  J  ]�  A!  "]t  A!  " p    �%  �  ��  �  �~  �>  	3   	�C     int Q  P   	�C     V   �  �o  P   	�C      �u   ?&  x�  G�  �  �          5  7�>  5   yint 5   7Q  M   S   !�  S   7�o  M   �  �|   k   !�  |   z!�  !�  !�  !�  !�  �   !�  !�  �  �|     4�   �   �  �   I @l    M       	k   �  #	k   �  &	k     )	k    �  ,	k   (�  -	k   0
  25   8�  55   < Q  8"�   7�  K�  l  7�  L�  7�  M�  �  �   !E  {6  |std  �  �  7  4q  �  �  �  �  �  �    	  �   �  q  �  !  '  �   T �  [v �    �  �  �  4q  �  �  �  �  ,  V  z  �  �   �  �  V  �  �  �   T �  [v �   <  2  ��  4q  ��  T 5   \�  .�'    �  �  4q  ��  T 5   \�  .�'    ]k�  l]��  ~��  `>  �U  a�  T �0   -�  j>*  ��  `k  �U  a5   T �'   A�  `�  �U  a�0  T T   i�  [�  �U  \�c  T �c   �  [�  �U  \�b  T �b   ^6  ��  �  ^6  �?  �  -�  j>x  ��  !Q�  �    T T  T   Ay�  �&  <  T �b  �U   -�  j>�  U�  �  �'  i  T �'  �V   -�  j>W  A��  '  �  T �c  �V   -�  j>�   !l  �  5  �  7  5F  I  �  }frg 	�'  B�  �  _o   �  ~�   
  .  7�'   <%  5   ,/  #�   #�  `hex  a�  �  ��  {�  ��  |5   �  ~;  k  q  �'   C�    �  �'  5     )    �  �  �'   )  a  �  �  �'  �   )  �  �  �  �'  �'   )  �  �    �'  �'   )  *�    (  �'  �'   )  0x  =  H  �'  �'   (  8  ]  h  �'  5    '�  =O  �'  �  �  �'  /   'c  Q�  �  �  �  �'   'c  T�  �  �  �  �'   'm  X�  �  �  �  �'   'R  \+  �'      �'   'R  `[  �'  !  '  �'   '!  d�   (  @  F  �'   f  �  Z  `  �'   �  �<   �  ��  T 5    /  �*  2p  �*  3Z(  �  �  (   	   6C  �  �  �  (  
      <
   �  =5   �)  >/  �   ?�  �'  @�  �#  A�  <  B�  �  C�  ��*  E&  K  V  (  5    ��*  >  d  (  �t    �  Dp  Jn	  6��  Nc�  �  P �	  T 5   m1  5   �  5   5   5   S    6�-  N�!  	  P �	  T �   m1  �   �  5   5   5   S    6ۮ  x��  B	  P �	  T 5   m1  5   5   5   5   S    ���  ��  T 5   F �	  5   �  m1    B�  	
n	  _�  	w	  �  	�  �)  	E#  �	  �	  Q1  T(   q,  �		U  q,  	�#  �	  �	  \1  Q1   /q,  	_   �	  �	  \1  g1   0�  		~-  m1  
  "
  \1  g1   p,  	�*  6
  A
  \1  5    )  	"	�  m1  Y
  d
  \1  n	   �$  	'a&  x
  �
  \1  S    �$  	1�  �
  �
  \1  �'   �)  	>Q1   ܨ  	?�0  7&  	@
k   �)  	A�  �/�  		`�  m1  �
    T S   \1  S    �  		��  m1  #  .  T 5   \1  5    Mc.  		�*  m1  I  T �'  \1  �'    �	  �  	H`*  �	  r  x  Q1   �#  	M�"  �  �  Q1  �'   .  	QT(   U(  T(  b].  |   � �  	�  �)  	E�&  �  �  �1  �(   q,  �		3  q,  	�&      �1  �1   /q,  	N"  &  1  �1  �1   0�  		�   �1  I  T  �1  �1   p,  	�"  h  s  �1  5    )  	"	�(  �1  �  �  �1  n	   �$  	'r  �  �  �1  S    �$  	1�,  �  �  �1  �'   �)  	>�1   ܨ  	?�0  7&  	@
k   �)  	A�  �Mc.  		�$  �1  '  T �'  �1  �'    �  �  	H�#  �  P  V  �1   �#  	M�  k  v  �1  �'   .  	Q�(   U(  �(  b].  |   � BE3  	�  ���  �   Dd^  	�  E�  N4j  �    O�  <G  5     #�   `red #h^   �o  0�  �o  �F  "  (  �/   /�o  �D  <  G  �/  �/   0�  �z  �/  _  j  �/  �/   tl  �    �  �   pU  �   �I   �   �D  !�    [r  "�  (   q  %
  �Q  '!=  �  �  T �  �2   c�  '1Q  �  T *  �2    dV  5�  dh 8<  �/  0  �2   pl  =�n  �2  J  �2   �p  B�^  �2  d  �2   lU  Ef|  �2  ~  �2   �I  I�  �2  �  �2   �D  LE  �2  �  �2   <3  Pfm  �2  �  �  �2   F�E  U�L  �  �  �2   F�_  Z�M  �    �2    c  djw       �2   / c  gar  4  ?  �2  �2   0�  i
J  �2  W  b  �2  �2   ��  op  �2  z  �  �2   �D  |+G  �  �  �2  �2   ��  ��z  �  �  �2  �2  �2   5>  ��@  �  �  �2  �2  �2   �F  �4\  �  
  �2  �2   $�  Dj    *  �2  �2   O  $d  @  P  �2  �2  �2   �U  D�6  f  v  �2  �2  �2   �  x�E  �  �  �2  �2    q  �nq  �  �  �2  �2   �9  1y  �  �  �2  �2   $�=  Ӏ  �  �  �2  �2   $�z  #�8      �2  �2   (L  0Nx  �  3  9  �2   (L  9�/  �  S  m  �2  �2  �'  �2  �2   G?3  ��    D �  T *  =�P  �u  A �   
  P�5  �Z  )��  )��  )��  )�J  )�d  )��  >
   $Z|  �@       3  3   $�F  �V�     +  3  �2   G�R  �3  T *  =�P  �u  L 3  A �   .H  5�  dh 8�4  �/  �  �2   pl  =&i  �2  �  �2   �p  B�Z  �2  �  �2   lU  EP  �2  �  �2   �I  I�f  �2  �  �2   �D  L}S  �2    �2   <3  PO]  �2       3   F�E  U�g  �  ;  �2   F�_  Z)?  �  V  �2    c  d8  j  p  3   / c  g~u  �  �  3  &3   0�  i'O  ,3  �  �  3  &3   ��  oAs  �2  �  �  3   �D  |�k  �  �  3  �2   ��  ��0      3  �2  �2   5>  ��A  *  :  3  �2  �2   �F  �X  O  Z  3  �2   $�  �1  o  z  3  �2   O  
e  �  �  3  �2  �2   �U  DxT  �  �  3  �2  �2   �  xfC  �  �  3  �2    q  �{l  �    3  �2   �9  E}    )  3  �2   $�=  �9  >  I  3  �2   $�z  #�`  ^  i  3  �2   (L  0�_  �  �  �  3   (L  9�a  �  �  �  3  �2  �'  23  23   G?3  ��    D �  T �  =�P  �u  XA �   Z  e�~  �)��  )��  )�  )��  )��  )�  >Z   $Z|  �<R  L  W  83  3   $�F  �/L  l  w  83  �2   G�R  �3  T �  =�P  �u  XL 3  A �    E�  N4j  �    O�  /�  �  fclz �3  5   �  |    T |    ���  �$�  < Q  5   �%  #�   #ʃ  #QS      �U  H�	�  �U  ���  K  `  �2     �   k    /�U  ���  t    �2  �2   0�  �
`D  �2  �  �  �2  �2   ��  ��b  �  �  �  �2  �    �U  �%   WS  ��   p �w   �=  �\#   *  �U  ��	�  >*   �U  �Pc  &  ;  �2  �   k   5    /�U  �z  O  Z  �2  �2   0�  �4  �2  r  }  �2  �2   �  �<   H�D  ��   L$H  ��2  P�B  �\#  X �  %\  �	.  %\  �/  �  �  �2   /%\  �l5  �  �  �2  4   0�  ��h  4       �2  4   �E  ��2    �  �R  �	e  M�  ��v  �  T  3  �2  �2    �.   �	�  �.  �R�  �  �  C3   �E  �	�/   �o  ��2  �e  ��   1|  �i#  u  ��=  �  �  ~1  I3   gu  (�t  �     ~1  O3   ��  *�K  U3    %  ~1  O3   '�  ��o  �   >  I  ~1  k    (�  L�g  �   c  s  ~1  �   k    �  ~��  �  �  ~1  �    �I  �Ճ  �  �  ~1  �   k    'WV  1	e;  k   �  �  ~1   �C  >k3                         @       Q�v  @ �   Q�`  A �    �~  H�U  k   >  �    �.  W�N  k   X  k    QQC  j<   4zz  lw   |  oK>  �  �  �    4́  |w   4]C  w   ��D  �w    H�~  ��<  �2  �  �  ~1  �    H��  &q  �2  �  �  ~1  5    HFS  %n^  �2    #  ~1  k    $4  7:k  8  >  ~1   $]  >�J  S  ^  ~1  �2   �[  �
I3   �1  ��/  �U  �v#  L  �x  �=  �	k    eu  ��3  (sz  d0  tZ  �/   �  �4^  V�  �B  X�;  �  �  s1  ~1   (�  [kt  �       s1  k    �I  _p3  .  >  s1  �   k    �  c"u  T  _  s1  �    (V  g�c  �   y  �  s1  �   k    �ZD  l~1   sz  d0  tZ  �/   D;�  �"  B�  ֚  9  c�  T�  �  �  �0   ˷  $�0  �  �   �  &�0  ��     �  �  )�  �0  u�  �0   ���  R�"   S�v   E>  hh %ҧ  	1  n  y  1  y   S�  "6   �  *	�   R�"   hh -	1�  	1  �  �  /1  y   �  2�  �  �  /1  y   R  5��  y  �  �  :1   
�  9��  �        :1  E1   �  <��  �  4   ?   :1  E1   j�  @�  K1  W   ]   /1   j�  D(�  �  u   �   /1  5    ^�  Ky    �  I�  N.�  �  �   �   1  y   ��  S-�  �   �   1   j�  V��  �  �   �   1  �    S˷  !4�  p�  g}�  �  !  $!  1  �    �F  x��  �  <!  L!  1  �  �    ��  ���  �  d!  j!  1   *  �s�  y  �!  �!  1   �  ��  y  �!  �!  1   �  ���  �   �!  �!  1   K�  �A�  �   �!  �!  1   »  �A�  �   �!  "  1  �   ķ  �g�  "  )"  1  �  1   ݱ  �נ  �  A"  G"  1   iend ���  �  _"  e"  1   )  ��    �  �y  T L)  �  �"    Ӝ  �"  �  ��  �0  �"  �"  �0  �0   T L)  H �  =�P  �u  X v�  
#  R�"   fget 
��  �0  
#  1   Tag �  T �"   ��  \#  m�  9�  �0  B#  �0   T L)  )�  �0  u�  �0   T�v  �+  T�D  �7�  T�D  �7�  amv  %  �~  �  �#  �#  �3   �~  e/  �#  �#  �3  �  ^0   �~  GZ  �#  �#  �3  ^0   g�~  !�b  $  $  �3  �3   �~  #�.  %$  0$  �3  �3   �~  (�Y  E$  P$  �3  5    '�  - R   4  i$  t$  �3  �#   �~  2J�  �$  �$  �3   |  8�Y  �$  �$  �3   'f3  >C  �  �$  �$  �3   'Gc  B=K  �  �$  �$  �3  M0   �1  G	M0   e3  H�  tZ  �/   �#  y�  ��  �  

i  �'  H%  T 5   �'  �'   6`)  ���  o%  F �	  5   �  m1   6f  ��  �%  F �  �'  �  �1   6`)  �O'  �%  F �	  �'  �  m1   ݻ  
�  �0  �%  Tag �  T �"  1   I�  3w�  &  T S   F �	  ,(  m1   I�  3�  ;&  T 5   F �	  �'  m1   I   3n$  e&  T �'  F �  nQ  �1   I�  3�%  �&  T �'  F �	  nQ  m1   A��  4  �&  T |-  H  �  J�  �&  .�'  .�b   KU  �'  �&  8�b   Aʣ  4  #'  T |-  H  �  J�  '  .�'  .�c   KU  �'  '  8�c   6��  i�  N'  T L)  H  �  KU  �0   vo  

j  Y  t'  T |   Y  Y   cʳ  
	
��  Y  T |   Y  Y    2�  	@+B     Z   �'  2�  	��B     <  �'  /  �'  <   85   �  8/  /  �  5   5   �  (  j:  �  j�  �  !�  Z   !|  2|	  	R+B     Dr  j/  <&  �(  k<&  
9(  v(  |(  j/   C�  '%  �(  j/  �'    P(  �(  kP(  6"  �(  �(  p/   C�  �'  �(  p/  �'    lD  +�  �	  l�  ,�  �  <�  5   
!)  #&�   #�  #i�   <��  5   L)  #&�   #Ȼ  #ب  #��   m}�  pL)  C-  >�   �w�  `4   }�  0ݥ  �)  �)  �0  )4   /}�  ��  �)  �)  �0  q4   0�  �  �0  �)  �)  �0  q4   ��  @Ҧ  L)  �)  �)  �0  5    C�  LU�  *  *  �0   �G #Ƙ  5   L)  /*  5*  �0   ��  V��  5   M*  b*  �0  M   k   G4   �  �G�  5   z*  �*  �0  �'  k   G4   K�  ���  �*  �*  �0  S    ��  �V�  5   �*  �*  �0  !)   ��  ��  �*  �*  �0   ��  ��  5   +  	+  �0   ��  ��  5   !+  ,+  �0  M4   H��  ?�  5   E+  U+  �0  �  5    ?ٷ  2�  5   L)  v+  �+  �0  ;4   ?v�  3�  5   L)  �+  �+  �0  A4   ?��  4��  5   L)  �+  �+  �0  M   k   G4   ?�  5j�  5   L)  ,  ,  �0  �'  k   G4   ?��  6D�  5   L)  :,  O,  �0  �  5   M4   (�  �  5   i,  o,  �0   (�  )c�  5   �,  �,  �0   (��  3�  5   �,  �,  �0   (��  U��  5   �,  �,  �0   (f  fT�  5   �,  �,  �0   ��  w�  -  -  �0   �U  B�(  H�  C!)  L?�  D%)4  Pl�  H(%  X L)  Et-  N��  $�   �  !9  ��  'Z-   OH-  mw�  xKL)  d/  >L)   nw�  |�  �-  �-  4  4   nw�  ��  �-  �-  4  #4   $w�  ��  �-  �-  4  5   )4   �fd ���  5   	.  .  4   �G �*�  5   |-  1.  7.  4   @ٷ  �6�  5   |-  Y.  d.  4  ;4   @v�  �4�  5   |-  �.  �.  4  A4   @��  �k�  5   |-  �.  �.  4  M   k   G4   @�  �'�  5   |-  �.  �.  4  �'  k   G4   @��  ��  5   |-  !/  6/  4  �  5   M4   �_fd \5   p�v�  Ů  |-  X/  4  5     |-   T(  �(  9�  9�    �/  �    9�  #Q  H0  #Q  C|  �/  �/  M0   /#Q  �B  �/  �/  M0  X0   0�   k  ^0  �/  0  M0  X0   �~  �A  0  0  M0   |  �  30  90  M0   ̀  5     �/  �/  M0  H0  �/  H  �0  imap vU  �   �0  �0  �0  k    C]   �f  �0  �0  �   k     d0  L)  �0  �  �0  %S   �0  &|    9M-  �  �"  �0  L)  �"  �"  J  9  1  9  2f-  	�C     �  /1  �   :1  �   �  �	  Q1  �	  \1  U  �	  �  s1  �  ~1  �  �1  �  �1  3  �  E%2  K&�  �|-  K��  �|-  K�  �|-  P;�  �	2  �;�  ��1  �1  \2   ���  �2  \2  5     K4�  ��1   ���1  2�1  	 C     2�1  	�C     2�1  	 C     �1  \2  22  	xC     Ux  �	H C     U�  �	P C     U�  �	X C     *  �2  �  *  �  �2  �  �  �  �2  
  �2  �  
  �2  3  3  �  3  Z  3  �  Z  �2  �  83  e  d0  �  �  %w   k3  &|    [3  5�{  �  5�7    5f    5]f  X  o=Y  f   �o�N  �   �Vn  �     5�7  �  %e  �3  &|    �c  .d  �b  �b  �#  �3  %  8�#  �#  .  �  |-  4  8|-  d/  /4  �;4  �0   �(  !)  k   �  �5   `4  � f4  �Y�  S4  C-  �&  �   9�  9�  ���  4�@            ���  A�@     �       ��4  	�  w5   �l	p  w5   �h VE/  K�4  5  �  4    <     �4  3�  '5  B�@     +       �05  �4  �h  �4  �  S5  �@     -       �\5  �4  �h d
  {5  6@     �       ��5  �  b1  �hs 	'S   �d ""%  95@     (       ��5  T 5   a 
�'  �hb 
#�'  �` ;  h�@     1       ��5  "O  Z�2  �h �  ��@     �      �)7  P �	  T 5   ��  Nm1  ���   N$5   ���'  N1�  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#S   ��4  P�'  �Xݨ  S)7  ��k T5   ��e�@     E       �6  i a5   �l ��@     -       	7  i d5   �h ��@     0       i f5   �d  %S   97  &|    �  �3@     �      �e8  P �	  T �   ��  Nm1  ���   N$�   ���'  N1�  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#S   ��4  P�'  �Xݨ  S)7  ��k T5   ���4@     E       "8  i a5   �l �4@     -       E8  i d5   �h 5@     0       i f5   �d    �8  Ȗ@     �      ��8  �  !3  ��3n �2  ��
u �2  �X
v �2  �P
w �2  �H �  �8  (�@     �      �19  �  !3  ��3n ��2  ��
u ��2  �X
v ��2  �P
w ��2  �H "�  �@            �c9  T �  "O  '�2  �h "�  
�@            ��9  T *  "O  '�2  �h �  �9  j�@     �      ��9  �  �2  ��3n �2  ��
u �2  �X
v �2  �P
w �2  �H �  :  ʑ@     �      �a:  �  �2  ��3n ��2  ��
u ��2  �X
v ��2  �P
w ��2  �H �  ��@     1       ��:  "O  Z�2  �h �  �:  ��@     V      ��:  �  �2  �Xn ��2  �Ptl  ��2  �h�R  ��2  �` �  }�@            �;  q,  =�2  �h �  -;  ��@     �      �<  �  !3  ��3n x�2  ��tl  {�2  �P
s ��2  �XTr  ��  ����@     �       �;  
x ��2  �H ��@     z       �;  
x ��2  �@ K�@     Q       �;  .\  ��2  �� ��@     Q       .\  ��2  ��     ��@     1       �6<  "O  U�2  �h 	  ��@     �       ��<  P �	  T 5   ��  xm1  �X�   x!5   �T3(  x-5   �Ph  x85   �L�)  y5   �H�D  yS   �D�@     ;       i$  {	�   �l  �  j�@            �=  q,  L�2  �h I  %=  "�@     H       �R=  �  !3  �X	"O  #�2  �P_�  $�2  �h "g  �@            �}=  q,  8�2  �h :  �=  ��@     V      ��=  �  !3  �Xn ��2  �Ptl  ��2  �h�R  ��2  �` )  �=  ��@            �>  �  !3  �h	"O  �2  �` �  />  v�@            �L>  �  �2  �h	"O  �2  �` �  k>  .�@     H       ��>  �  �2  �X	"O  #�2  �P_�  $�2  �h 0  �@            ��>  q,  =�2  �h v  �>  N|@     �      ��?  �  �2  ��3n x�2  ��tl  {�2  �P
s ��2  �XTr  ��  ��}@     �       Q?  
x ��2  �H 9~@     z       u?  
x ��2  �@ �@     Q       �?  .\  ��2  �� .�@     Q       .\  ��2  ��  �  |@     1       ��?  "O  U�2  �h �  �{@            �@  q,  L�2  �h "  �{@            �A@  q,  8�2  �h 7  O@  }@  �  �2  *�B  �   *�=  �%�   *�U  �6k     A@  �[  �@  F{@     K       ��@  O@  �hX@  �dd@  �Xp@  �P �  �@  z@     7      �A  �  �2  �Htl  ��2  �@"O  �"�2  ��*L  ��2  �X �  :A  �x@     7      �uA  �  �2  �Htl  ��2  �@"O  �!�2  ��M�  ��2  �X �  �A  lx@     j       ��A  �  �2  �h"O  |�2  �`   �A  �A  �  �2  *�=  ��   *�U  �)k   *$w  �65     �A  �X  B  x@     d       �0B  �A  �h�A  �`�A  �X�A  �T z  OB  |u@     �      ��B  �  !3  ��	"O  �2  ��	�/   �2  ��tl  �2  �X�  �2  �PpU  �2  �H �  ]u@            ��B  q,  I�2  �h �  �B  �r@     a      �YC  �  !3  ��	"O  D�2  ��	.\  D$�2  ��M�  E�2  �X*L  F�2  �Ptl  Z�2  �H B	  L�@     �       ��C  T 5   F �	  �  �5   �lfo �/�  �`��  �6m1  �X �  �C  v.@     �       ��C  �  �1  �hstr 	1�'  �`   
D  �q@     7      �ED  �  !3  �Htl  ��2  �@"O  �"�2  ��*L  ��2  �X �  �q@            �pD  q,  E�2  �h �  �D  np@     7      ��D  �  !3  �Htl  ��2  �@"O  �!�2  ��M�  ��2  �X �  Pp@            ��D  q,  B�2  �h 1@  E  (p@     (       �;E  �  3  �ha �!�2  �`b �1�2  �X �  ZE  �o@     j       �vE  �  !3  �h"O  |�2  �` 1  �E  �o@            ��E  �  !3  �h *  �E   m@     �      �!F  �  �2  ��	"O  �2  ��	�/   �2  ��tl  �2  �X�  �2  �PpU  �2  �H ~  m@            �LF  q,  I�2  �h P  kF  �j@     a      ��F  �  �2  ��	"O  D�2  ��	.\  D$�2  ��M�  E�2  �X*L  F�2  �Ptl  Z�2  �H d  �j@            ��F  q,  E�2  �h J  cj@            �!G  q,  B�2  �h 1�  @G  Rj@            �MG  �  �2  �h �
  lG  �/@     �       ��G  �  b1  �hstr 	1�'  �` "�"  >�@            ��G  p 
%1  �h �  �G  �@     <      �sH  �  �1  ��	ѷ  �1�   ��	@  �Ak   ��WS  �|   �X
slb ��2  �P
bkt �C3  �H�1  �	k   �@`v  ��#  ��H  ��  ���  ��2  �� �  �H  i@     �       ��H  �  �1  �H	@  %8k   �@WS  +�   �X
fra -�2  �P t$  �H  �h@     L       ��H  �  �3  �h   I  �g@     �       �GI  �  3  �X	"O  ��2  �P_�  ��2  �h �  fI  �f@     D      �J  �  �1  ��	�  45   ��WS  
�   �@�1  |   ���f  	k   �X
slb �2  ����  �2  �Pag@     ^       
off k   �Hwg@     >       �  �2  ��   �  ;J  :f@     X       �WJ  �  !3  �X_�  p�2  �h Z  vJ  ~e@     �       ��J  �  !3  �H	"O  �2  �@B>  �2  �h`w  �2  �`�e@     I       M�  �2  �X  H%  ��@     J       �&K  F �	  �  �5   �Lfo �/�  �@��  �6m1  �� o%  �-@     *       �vK  F �  �  � �'  �hfo �7�  �`��  �>�1  �X W  �K  �d@     �       ��K  �  >3  �X	"O  ��2  �P_�  ��2  �h 1�  �K  @d@     I       �
L  �  �2  �Xp ��   �Padr �	|   �h �  L  "L  �  �2   ,
L  �c  EL  *d@            �NL  L  �h �$  mL  �c@     O       �zL  �  �3  �h 
  �L  c@     �       ��L  �  �2  �H	"O  �2  �@B>  �2  �h`w  �2  �`�c@     I       M�  �2  �X  �  M  Vb@     �       �DM  �  �1  �X	WS  �6�   �P_�  ��2  �h 0$  RM  eM  �  �3    <     DM  a4  �M  .b@     '       ��M  RM  �h �#  �M  �M  �  �3  *�1  ^0    �M  S�  �M  �a@     2       ��M  �M  �h�M  �` �%  .@     *       �9N  F �	  �  � �'  �hfo �7�  �`��  �>m1  �X 1�"  XN  ��@            �rN  �  �0  �hx �0  �` �%  ��@            ��N  Tag �  T �"  p 
1  �h   �N  R�@     1       ��N  �  y1  �h	ѷ  _�   �`	@  _(k   �X �%  
�@     G       �AO  T S   F �	  	�  3,(  �H	��  3!m1  �@ �  `O  ��@     0       �|O  �  51  �hptr -y  �` 1�  �O  ��@     "       ��O  �  @1  �h�  9$E1  �` %  �O  �Z@     �      ��P  �  �1  ��~p �1k   ��~�Z@     �      �P  �  �5   �\
bkt C3  �P`v  �#  ���  �2  ��d[@     *      oP  
slb 	�2  �H �\@     �      
slb 	�2  �@Cx  #�#  ��  �^@     �       @  :|   ��
fra ;�2  ��Cx  =�#  ��~  &  t�@     C       �3Q  T 5   F �	  	�  3�'  �H	��  3!m1  �@ V  RQ  �,@     &       �nQ  �  �1  �h/&  	M�'  �` �'  ;&  �+@     E       ��Q  T �'  F �  	�  3nQ  �H	��  3!�1  �@ �  �Q  �Q  �  �1  *�)  	�1   ,�Q  �  R  �+@     4       �R  �Q  �h�Q  �` s  5R  DW@     h      ��R  �  �1  ��~	ѷ  ~+�   ��~WS  �|   �XCx  ��#  ��
fra ��2  �P
slb ��2  �H
bkt �C3  �@�1  �	k   ��`v  ��#  ��H  ��  ���  ��2  �� x  S  h-@     &       �$S  �  W1  �h/&  	M�'  �` e&  �,@     E       �nS  T �'  F �	  	�  3nQ  �H	��  3!m1  �@ �	  |S  �S  �  b1  *�)  	Q1   ,nS  �  �S  �,@     4       ��S  |S  �h�S  �` �  �S  �S  �  51  *_�  2y   ,�S  ݙ  T  Z�@            �T  �S  �h�S  �` �0  "�  H�@            �TT  T T  x *T  �h W  sT  �@     0       ��T  �  1  �hptr %y  �` "(#  	�@            ��T  К  �0  �h q  �T  �T  �  �'    <    ,�T  6.  �T  �+@            �U  �T  �h W  U  U  �  �'   ,U  9*  BU  �+@            �KU  U  �h �  �&  ��@     �       ��U  T |-  H  �  J�  �U  .�'  .�b   C  KU  ��p+�U  �'  �&   ѷ  �   �H@�  +�'  ����  +�&  �� <  "  ��@            �V  T �b  x .�U  �h �&  +�@     �       ��V  T |-  H  �  J�  XV  .�'  .�c   C  KU  ��p+{V  �'  '   ѷ  �   �H@�  +�'  ����  +'  �� i  "H  ��@            ��V  T �'  x .�V  �h �  "u  �@            �W  T �c  x .�V  �h #'  ��@     G       �aW  T L)  H  �  C  KU  �hѷ  (�0  �` �
  �W  ��@     *       ��W  T S   �  b1  �h�  	S   �d 1�  �W  x�@            ��W  �  @1  �h ?   �W  F�@     2       ��W  �  51  �h    X  �@     (       �6X  �  @1  �h�  <$E1  �` G"  UX  ��@     #       �bX  �  1  �X )"  �X  ��@     3       ��X  �  1  �X �  �X  |V@     (       ��X  �  y1  �h	@  [k   �`   �X  ��@     (       �Y  T 5   �  b1  �h�  	5   �d �   "N'  �V@     +       �OY  T |   a 
Y  �hb 
#Y  �` "t'  s�@     +       ��Y  T |   a 
	Y  �hb 
	#Y  �` s  �Y  �*@     ,       ��Y  �  �1  �hLn	  �    �Y  �*@     )       �Z  T �'  �  �1  �h�  	�'  �` T  Z  #Z  �  �1    <    ,Z  v(  FZ  t*@            �OZ  Z  �h 8  nZ  J*@     )       �{Z  �  �1  �` �!  �Z  ��@     �      ��Z  �  1  ��it ��  ���  ��   �H��  �y  �Pz�  ��   �X �   [  2�@     a       �[  �  1  �Xptr N&y  �P >  >[  RV@     )       �[[  �  y1  �h	ѷ  c�   �` >  TU@     �       ��[  @  W0k   ��tc Y|   �`e b|   �Xf c|   �Pip d|   �His e|   �@�U@     :       i [�   �l  "$  �T@            �Z\  idx H6�   ��tc J|   �hs O5   �dip P|   �Xis Q|   �Pf R|   �H A
  y\  �+@     ,       ��\  �  b1  �hLn	  �  .  �\  4+@     )       ��\  T �'  �  b1  �h�  	�'  �` "
  �\  �\  �  b1    <    ,�\  *$  ]  (+@            �]  �\  �h Z  <]  �*@     )       �I]  �  W1  �` !  h]  ��@     �      ��]  �  1  �Hkz  g#�   �@u�  iy  �X �  �]  �]  �  �0   ,�]  l�  �]  l�@     *       ��]  �]  �h �   �]  �]  �  1   ,�]  �  ^  J�@     "       �^  �]  �h   )^  ?^  �  �'  *�  *�'    ^  %'  b^  �)@     V       �s^  )^  �h2^  �` H  �^  �^  �  �'    <     s^  g  �^  �)@            ��^  �^  �h �  �^  �^  �  �'    �^    �^  �)@     #       �_  �^  �h q��  t��@     5       �D_  	Q t�  �Xz�  u�0  �h -��  n5   ��@     B       ��_  3c n5   �\	Q n�  �Pz�  o�0  �h q��  hT�@     R       ��_  	Q h�  �Xz�  i�0  �h -��  N5   k�@     �       ��`  	Q N�  �H	ݨ  N$M   �@	)  N05   ��	@  N=k   ��z�  P�0  �h��@     1       o`  
e R
5   �d ��@     -       �`  
e W
5   �` �@     -       
e \
5   �\  -��  J5   Q�@            ��`  	Q J�  �h -��  D5   �@     I       �,a  	Q D�  �Xz�  E�0  �h -��  :�   ��@     ]       ��a  	Q :�  �Hz�  ;�0  �hֲ  <�  �X��@     1       
e =	5   �d  -��  15   E�@     f       �$b  	Q 1�  �X	�  1!�   �P	s�  1-5   �Lz�  2�0  �hr�@     2       
e 3	5   �d  -�  &5   ��@     �       �vb  	Q &�  �Xz�  '�0  �`
e (5   �l -x�  �  '�@     �       �tc  3fd 5   ��~	)  "�'  ��~eI�  #r7�  �b  �b  �3  5    s�   c  ��@     *       �c  �b  �  Lc  �h	��  #�0  �` ta�  )4  @c  �@            �Rc  �  Lc  �h�3   u��  ��@            �L�0  �h   -��  ��  ��@     E      ��d  	@�  ��'  ��}	)  �+�'  ��}   �5   �l��  ��  �k
fd 5   ��}PI�  �d  r7�  d  d  �3  5    s�  3d  ,�@     *       �Pd  �c  �  d  �h	��  �0  �` ta�  )4  sd  v�@            ��d  �  d  �h�3   u��  V�@            �L�0  �h  e�@     7       
e 	5   �d  -�  �5   �@            ��d  	Q ��  �h -�  �5   ��@     4       �?e  	Q ��  �Xz�  �4  �h �1  Me  �e  �  b2    <   Wvit ��0  X��  1  Xױ  �  X�  �  Wve �5      �?e  �e  ��@     �       �@f  Me  ��~w_e  �e  :`e  :le  :ue  :~e  ��e  :�e    Y_e  �@     �       ;`e  �`;le  �h;ue  ��~;~e  ��~Y�e  k�@     [       ;�e  �\   �1  Nf  Xf  �  b2   �@f  xf  ��@            ��f  Nf  �h �.  �f  ��@     E       ��f  �  4  �X	�  ��  �P	s�  �(5   �L	ͨ  �7M4  �@��@     '       
e �	5   �l  �.  g  L�@     U       ��g  �  4  �X	ݨ  �#�'  �P	�1  �2k   �H	ִ  �DG4  �@
s �
�   �`d�@     (       
e �	5   �l  �.  �g  ��@     U       �h  �  4  �X	ݨ  �M   �P	�1  �+k   �H	ִ  �=G4  �@
s �
�   �`�@     (       
e �	5   �l  d.  0h  �@     �       ��h  �  4  ��~	)  �-A4  ��~+  �h  	�HB     ]�@     �       
e �	5   �l  %Z   �h  &|    �h  7.  �h  ��@     h       ��h  �  4  �X	�U  �*;4  �P�  ��  �`
e �5   �l .  i   �@     �       �>i  �  4  ��~s�@            
e �	5   �l  1�-  ]i  ��@            �ji  �  4  �h �-  xi   �i  �  4  �fd �5   �@�  �!)4    ji  c�  �i  ��@     E       ��i  xi  �h�i  �d�i  �X �,  �i  2�@     u       �(j  �  �0  �X+  8j  	�HB     
ptr |�   �h %Z   8j  &|    (j  �,  \j  j�@     �       ��j  �  �0  �X+  �j  	�HB     v�@            
e g	5   �l  %Z   �j  &|    �j  �,  �j  J�@            �Uk  �  �0  ��~\�@             k  
e V
5   �l ��@     �       ͨ  Z	�  ��~(�  [�   �`��@     �       
e \5   �\   �,  tk  V�@     �      �@l  �  �0  �H+  Pl  	�HB     b�@            �k  
e 4	5   �l ��@     Z       �k  ͨ  =	�  �X��@     J       
e >
5   �h  ~�@     �       �  H
k   �P~�@     i       
e I
5   �d   %Z   Pl  &|    @l  o,  tl  ��@     �       ��l  �  �0  �h+  �l  	�HB      %Z   �l  &|    �l  O,  �l  T�@            �m  �  �0  �X+  m  	�HB     r�@     0       
e #	5   �l  %Z   m  &|   
 m  ,+  <m  :�@           �n  �  �0  �H	�  �  �@	s�  +5   ��ͨ  	�  �P+  'n  	�HB     M�@            �m  
e 	5   �l p�@     e       �m  (�  �   �`��@     D       
e 
5   �\   �@     @       
e 
5   �X  %Z   'n  &|    n  	+  Kn  ��@     n       ��n  �  �0  �Xֲ  � M4  �P(�  ��  �`��@     3       e �	5   �l  �*  �n  d�@     h       �o  �  �0  �X��@            �n  e �5   �l ��@            e �
5   �h  1�*  "o  $�@     ?       �/o  �  �0  �h �*  No  ��@     T       �}o  �  �0  �h)  �/!)  �d+  �o  	�HB      %Z   �o  &|    }o  �*  �o  b�@     m       ��o  �  �0  �hc � S   �d+  �o  	zHB      %Z   �o  &|    �o  b*  p  ��@     �      �-q  �  �0  ��~ݨ  �&�'  ��~�1  �5k   ��}ִ  �GG4  ��}+  �o  	tHB     ��  �|   ��~һ  ��  �o!�@     �       �p  �  �
k   ��~[�@     Y       e �
5   �h  �@             �p  e �
5   �d 5�@             q  e �
5   �` T�@     @       nl �M   �X  5*  Lq  ��@     �      �xr  �  �0  ��~ݨ  VM   ��~�1  V.k   ��~ִ  V@G4  ��~+  'n  	oHB     ��  �|   �X��@     �       �q  �  \
k   ��~��@     Y       e ]
5   �l  ��@           �  x
k   ��~��@             4r  e q
5   �h ϼ@             Wr  e s
5   �d ��@     a       e y
5   �`   �)  �r  κ@     /       ��r  �  �0  �h �)  �r   �r  �  �0    <   W�it H�     �r  ��  �r  ��@     +       ��r  �r  �h  �r  ˾  "s  ��@     �       �Zs  �r  ��~w�r  :s  :�r   Y�r  ݹ@     �       ;�r  ��~  n)  hs   ~s  �  �0  *@�  0%)4    Zs  ?�  �s  �@     �       ��s  hs  �hqs  �` 10  �s  �M@            ��s  �  S0  �h 0  �s  �M@     B       �t  �  S0  �h+  'n  	jHB      "�  �M@            �Ft  x )|   �h   Tt  ^t  �  �/   ,Ft  1~  �t  :M@     Q       ��t  Tt  �h V9  2�t  �t  �  (    <     �t  .  �t  �)@            ��t  �t  �h p  VV  2�t   u  �  (  �t    �t  �  #u   )@     �       �4u  �t  �h�t  �` �  Bu  Lu  �  (    4u  K  ou  �(@     \       �xu  Bu  �h �.  ^  �   �(@            ��u  @  #k   �hp /�   �` !i	  !J  ZL)  %  "Z*  \#  "Z�  \#  " �   Y1  t�  ��  �  0"          *�  E�>  5   uint 
5   EQ  M   X   FM   +�  
X   E�o  M   $2�  (|   v=�  �   -�   �   1�     +�  
�   w�  �   J>�   �    J��   �   J��   �   J�   �    +�  
�   x$9�  cp   $�  ��   
�   $�    +�  I @�    M       	�   �  #	�   �  &	�     )	�    �  ,	�   (�  -	�   0
  25   8�  55   < $Q  8"  $�  9�   
�  E�  K�  �  F�  E�  L�  E�  M�  +�  
�  +�  +�  +�  $��  �  $�  ��   $_�  /  $  4  
0  +�  K3�  e�   $��  �  +E  y6  zstd  `  �  �  =q  g  $�  `  .�  �  �  �  �  u   .�  q  �  �  �  u   T `  av `    
x  �  a  =q  g  $�  `  .�  ,  	  -  3  �   .�  �  	  K  Q  �   T `  av `   
�  2  ��  =q  �g  T 5   L�  M=2    �  ��  =q  �g  T 5   L�  MC2    ��  `�  $�U  a5   T U2   ��  �  =q  �g  T 5   L�  M72    � �;  =q  �g  T 5   L�  MU2    ��  `\  $�U  a`  T Ik   N6  ��  g  N6  �?  g  N6  �� g  N6  ���  g  m�  
��  �  T `  Ik  Ik   $-�  j>H  '5�  
!x�  �  �  T Ik  Ik   ?�  
L�    T 5   U2  U2   'U�  
�  U2  6  T U2  �   $-�  j>�  Wd�  
!g�  6  T U2  U2    +l  
`  B  �  �  BF  �  a  {frg �0  XE3  	
�  |��  �   Yd^  	�  Z�  b4j  g    [�  OG  5   �  %�   cred %h^   �o  0�  �o  �F    %  �0   ?�o  �D  9  D  �0  �0   @�  �z  �0  \  g  �0  �0   tl  �    �  �   pU  �   �I   �   �D  !�    [r  "�  ( 
�  q  %  '�  '1Q  `  �  T &  [:   W�Q  '!=  `  T �  r:    dV  5�
  dh 8<  �0  -  [:   'pl  =�n  [:  G  [:   '�p  B�^  [:  a  [:   'lU  Ef|  [:  {  [:   '�I  I�  [:  �  [:   '�D  LE  [:  �  [:   .<3  Pfm  [:  �  �  �:   P�E  U�L  `  �  [:   P�_  Z�M  `    [:    c  djw      �:   ? c  gar  1  <  �:  �:   @�  i
J  �:  T  _  �:  �:   .��  op  [:  w  }  �:   �D  |+G  �  �  �:  [:   ��  ��z  �  �  �:  [:  [:   5>  ��@  �  �  �:  [:  [:   �F  �4\  �  	  �:  [:   2�  Dj  	  '	  �:  [:   ,O  $d  =	  M	  �:  [:  [:   ,�U  D�6  c	  s	  �:  [:  [:   ,�  x�E  �	  �	  �:  [:   , q  �nq  �	  �	  �:  [:   ,�9  1y  �	  �	  �:  [:   2�=  Ӏ  �	  �	  �:  [:   2�z  #�8  
  
  �:  [:   CL  0Nx  `  0
  6
  �:   CL  9�/  `  P
  j
  �:  [:  U2  �:  �:   A?3  ��    D �
  T &  Q�P  ��  A �   
  <�5  �W  5�}  5��  5��  5�G  5�a  5��  \   2Z|  �@  �
    �:  /   2�F  �V�    (  �:  [:   A�R  �/  T &  Q�P  ��  L /  A �   .H  5�  dh 8�4  �0  }  r:   'pl  =&i  r:  �  r:   '�p  B�Z  r:  �  r:   'lU  EP  r:  �  r:   '�I  I�f  r:  �  r:   '�D  L}S  r:  �  r:   .<3  PO]  r:      �:   P�E  U�g  `  8  r:   P�_  Z)?  `  S  r:    c  d8  g  m  �:   ? c  g~u  �  �  �:  �:   @�  i'O  �:  �  �  �:  �:   .��  oAs  r:  �  �  �:   �D  |�k  �  �  �:  r:   ��  ��0      �:  r:  r:   5>  ��A  '  7  �:  r:  r:   �F  �X  L  W  �:  r:   2�  �1  l  w  �:  r:   ,O  
e  �  �  �:  r:  r:   ,�U  DxT  �  �  �:  r:  r:   ,�  xfC  �  �  �:  r:   , q  �{l  �    �:  r:   ,�9  E}    &  �:  r:   2�=  �9  ;  F  �:  r:   2�z  #�`  [  f  �:  r:   CL  0�_  `  �  �  �:   CL  9�a  `  �  �  �:  r:  U2  �:  �:   A?3  ��    D �  T �  Q�P   �  XA �   
W  I�~  �5��  5��  5�  5��  5��  5��  \W   2Z|  �<R  I  T  �:  /   2�F  �/L  i  t  �:  r:   A�R  �/  T �  Q�P   �  XL /  A �    Z�  b4j  g    [�  /�  �  }clz �3  5   �  �    T �    ~��  �$�  O Q  5   �!  %�   %ʃ  %QS   
�  �U  H�	�  �U  ���  G  \  [:  �  0  �    ?�U  ���  p  {  [:  f:   @�  �
`D  l:  �  �  [:  f:   .��  ��b  `  �  �  [:  �    �U  �!   WS  �<  p �  �=  �%*   
&  �U  ��	�  \&   �U  �Pc  "  7  r:  0  �   5    ?�U  �z  K  V  r:  }:   @�  �4  �:  n  y  r:  }:   �  �<   H�D  ��   L$H  ��:  P�B  �%*  X 
�  %\  �	*  %\  �/  �  �  �:   ?%\  �l5  �  �  �:  �;   @�  ��h  �;      �:  �;   �E  ��:    
�  �R  �	a  e�  ��v  `  P  �:  f:  f:    �.   �	�  �.  �R�  �  �  �:   �E  �	�0   �o  �r:  �e  ��   $1|  �2*  u  ��=  �  �  p9  �:   fu  (�t  �  �  p9  �:   �  *�K  ;       p9  �:    �  ��o  �   9  D  p9  �    C�  L�g  �   ^  n  p9  �   �    ,�  ~��  �  �  p9  �    ,�I  �Ճ  �  �  p9  �   �     WV  1	e;  �   �  �  p9   �C  >;                         @       ]�v  @ �   ]�`  A �    '�~  H�U  �   9  �    '�.  W�N  �   S  �    ]QC  j<   =zz  l  '|  oK>  `  �  �    =́  |  =]C    ��D  �   ^�~  ��<  [:  �  �  p9  0   ^��  &q  r:  �  �  p9  5    ^FS  %n^  [:      p9  �    24  7:k  3  9  p9   2]  >�J  N  Y  p9  [:   �[  �
�:   �1  ��0  $�U  �?*  L  �s  �=  �	�    eu  �m;  (sz  �1  tZ  �0   
�  �4^  V�  ,�B  X�;  �  �  e9  p9   C�  [kt  �       e9  �    ,�I  _p3  )  9  e9  �   �    ,�  c"u  O  Z  e9  �    CV  g�c  �   t  �  e9  �   �    !ZD  lp9   sz  �1  tZ  �0   X�  
�  go   �  ��   �  �.  72   O%  5   ,  %�   %�  chex  R�  {  ��  {_  ��  |5   �  ~;  =  C  2   _�    S  2  5     )    t  z  &2   )  a  �  �  &2  �   )  �  �  �  &2  12   )  �  �  �  &2  72   )  *�  �  �  &2  =2   )  0x      &2  C2   (  8  /  :  &2  5     �  =O  I2  S  ^  &2      c  Q�  `  w  }  O2    c  T�  `  �  �  &2    m  X�  `  �  �  O2    R  \+  12  �  �  O2    R  `[  U2  �  �  &2    !  d�  [2      &2   f  �  ,  2  &2   �  �   �  �`  ��  %z�  h  s  U U2  &2  U2   T 5    
  �*  2h  �*  3Z(  �  �  a2   .	   6C  �  �  �  a2  �      <�   �  =5   �)  >  �   ?`  �'  @`  �#  A`  <  B`  �  C`  �*  E&  C  N  a2  5    ��*  >  \  a2  �    
�  Yp  J�#  ��  Nc�  �  P (  T 5   �3  5   `  5   5   5   X    �-  N�!  �  P (  T �   �3  �   `  5   5   5   X    �'  x<+  :  P (  T �   �3  �   5   5   5   X    ۮ  x��  w  P (  T 5   �3  5   5   5   5   X    �  ��+  �  T �   F (  �   �  �3   ��  ��  �  T 5   F (  5   �  �3   ��  NH�    P �5  T �2  �B  �2  `  5   5   5   X    ]�  N��  W  P �5  T �   �B  �   `  5   5   5   X    ��  N��  �  P �5  T   �B    `  5   5   5   X    ��  N5�  �  P �5  T �   �B  �   `  5   5   5   X    �  NG�    P a4  T �2  �K  �2  `  5   5   5   X    E�  Na�  _  P a4  T �   �K  �   `  5   5   5   X    ��  N��  �  P a4  T   �K    `  5   5   5   X    ��  N��  �  P a4  T �   �K  �   `  5   5   5   X    I�  N�  %  P 5  T �2  fP  �2  `  5   5   5   X    	 N�  g  P 5  T �   fP  �   `  5   5   5   X    �  Nm�  �  P 5  T   fP    `  5   5   5   X    ^�  N��  �  P 5  T �   fP  �   `  5   5   5   X    :�  N6�  -  P �3  T �2  mU  �2  `  5   5   5   X    {�  N��  o  P �3  T �   mU  �   `  5   5   5   X    N�  NI�  �  P �3  T   mU    `  5   5   5   X    ��  N��  �  P �3  T �   mU  �   `  5   5   5   X    ��  x�  0   P �5  T �2  �B  �2  5   5   5   X    @�  xo�  m   P �5  T �   �B  �   5   5   5   X    ��  x� �   P �5  T   �B    5   5   5   X    ��  xA�  �   P �5  T �   �B  �   5   5   5   X    /�  x' $!  P a4  T �2  �K  �2  5   5   5   X    N�  x��  a!  P a4  T �   �K  �   5   5   5   X    <�  xO�  �!  P a4  T   �K    5   5   5   X    ~�  xJ�  �!  P a4  T �   �K  �   5   5   5   X    ��  x`�  "  P 5  T �2  fP  �2  5   5   5   X    �  x�  U"  P 5  T �   fP  �   5   5   5   X    ��  x,�  �"  P 5  T   fP    5   5   5   X    �  x	�  �"  P 5  T �   fP  �   5   5   5   X    ��  x��  #  P �3  T �2  mU  �2  5   5   5   X    ^�  x��  I#  P �3  T �   mU  �   5   5   5   X    D�  x��  �#  P �3  T   mU    5   5   5   X    ���  x!�  P �3  T �   mU  �   5   5   5   X     x�  ��#  ��  �
�     O:�  5   �$  %u�   %e�  %a�  %��   R�  �%  o�  ׈  )$  /$  �2   o�  ��  D$  O$  �2  �1   o�  �  d$  t$  �2  �1  �     �  �  �1  �$  �$  �2    �  #��  �2  �$  �$  �2  �     @  '	7�  �   �$  �$  �2    
�  +p�  `  �$  �$  �2  $    �  3�  `  %  %  �2  $    ��  7	
�  �   7%  G%  �2  X   �     Ĉ  ?	ȉ  �   `%  k%  �2  X     R�  G�  $  �%  �%  �2  �   �    з  X�1   o Y	�   �  X    
$  R�  n'  o�  ��  �%  �%  �2   o�  �  �%  &  �2  �2   o�  ��  &  *&  �2  �2  �     �  �  �2  C&  I&  �2    �  #��  �2  b&  m&  �2  �     @  '	I�  �   �&  �&  �2    
�  +�  `  �&  �&  �2  �%    �  3k�  `  �&  �&  �2  �%    ��  7	!�  �   �&  �&  �2  �2  �     Ĉ  ?	g�  �   '  !'  �2  �2    R�  G��  �%  :'  J'  �2  �   �    з  X�2   o Y	�   �  �2   
�%  <j�  �'  2j�  "��  �'  �'  �2  �2  �    Aܨ  &�2   A@  '	�    
s'  X�  	

�'  g�  	�'  �  	*  �)  	E#  (  (  �3  3   q,  �		�)  q,  	�#  1(  <(  �3  �3   ?q,  	_   P(  [(  �3  �3   @�  		~-  �3  s(  ~(  �3  �3   p,  	�*  �(  �(  �3  5    .)  	"	�  �3  �(  �(  �3  �'   �$  	'a&  �(  �(  �3  X    �$  	1�  �(  �(  �3  �1   /�)  	>�3   /ܨ  	?{3  /7&  	@
�   �/)  	A`  �./�  		`�  �3  U)  `)  T X   �3  X    .d�  		u�  �3  )  �)  T s'  �3  s'   ec.  		�*  �3  �)  T �1  �3  �1    
(  .�  	H`*  (  �)  �)  �3   �#  	M�"  �)  �)  �3  �1   /.  	Q3   U(  3  �].  �   � h�  �;�  K�v  �+�  K�D  �7�  K�D  �7�
  Rmv  �+  �~  �  n*  t*  };   �~  e/  �*  �*  };  �  �1   �~  GZ  �*  �*  };  �1   f�~  !�b  �*  �*  };  �;   �~  #�.  �*  �*  };  �;   �~  (�Y  +  +  };  5     �  - R  �;  2+  =+  };  L*   �~  2J�  R+  X+  };   |  8�Y  m+  s+  };    f3  >C  `  �+  �+  };    Gc  B=K  `  �+  �+  };  ~1   �1  G	~1   e3  H`  tZ  �0   
L*  '�  
i  12  ,  T 5   12  12   `)  �@%  ,,  F (  �   �  �3   `)  ���  S,  F (  5   �  �3   (N#  8��  �,  T �   F (  ~\  �  �3   (�  3w�  �,  T X   F (  �2  �3   ( ���  �,  F �5  �B  X   �  �#  �7   (��  q��  -  F �5  �B  X   �  �#  �7   ($ '��  B-  F �5  �B  X   �  �#  �7   (`)  ��  j-  F (  s'  �  �3   `)  �O'  �-  F (  �1  �  �3   (� ���  �-  F a4  �K  X   �  �#  �7   (+�  qF�  �-  F a4  �K  X   �  �#  �7   (��  'Q�  '.  F a4  �K  X   �  �#  �7   (�  ��  Y.  F 5  fP  X   �  �#  �7   (��  q	�  �.  F 5  fP  X   �  �#  �7   (a�  '�  �.  F 5  fP  X   �  �#  �7   (�  �}�  �.  F �3  mU  X   �  �#  �7   (��  q�  !/  F �3  mU  X   �  �#  �7   (?�  '��  S/  F �3  mU  X   �  �#  �7   '�  iI�  n/  I2  I2   (e�  3ˑ  �/  T s'  F (  ��  �3   (�  3�%  �/  T �1  F (  K�  �3   ` ���  �/  A {9  {9  �1  �7   Q�  ���  0  A �8  �8  �1  �7   'ʳ  	
��  #�  60  T �   #�  #�   C ���  ]0  A �7  �7  �1  �7   ��  ���  �0  A �6  �6  �1  �7   Wvo  
j  #�  T �   #�  #�    D�  D�  �  
�0  �  �  D�  #Q  y1  #Q  C|  �0  �0  ~1   ?#Q  �B  1  1  ~1  �1   @�   k  �1  +1  61  ~1  �1   �~  �A  J1  P1  ~1   |  �  d1  j1  ~1   /̀  5     
�0  �0  
~1  y1  �0  H  �1  �map vU  0  �1  �1  �1  �    _]   �f  �1  �1  0  �     �1  `�  	eIB     _   
�1  F�1  `�  	��B       
2    
&2  <   )5   {  )    {  5   5   �  
a2  S:  s  S�  �  +�  $  
�2  �%  
�2  _   �%  
�2  �2  F�2  +|  
�2  n'  
�2  �2  s'  
�2  �2  �`�'  	wIB     Yr  o3  <&  I3  �<&  
9(  '3  -3  o3   _�  '%  =3  o3  �1    iD  +�  �'  i�  ,�  *  h}�   3  i3  -X   �3  1�    �'  
�3  (  
�3  �)  (  |�  DV4  |�  EW �3  �3  V4  �   �$  H6�  �3  �3  V4  X    �$  M��  4  4  V4  �1   �$  R��  +4  ;4  V4  �1  �    �  W�   ��  X	�    �3  
V4  '�  [
5  '�  \��  �4  �4  
5  M    �$  _1�  �4  �4  
5  X    �$  d��  �4  �4  
5  �1   �$  l��  �4  �4  
5  �1  �    ݨ  tM    ��  u	�    a4  

5  h�  x�5  h�  yo�  65  F5  �5  M   �    �$  |��  Z5  e5  �5  X    �$  �B�  y5  �5  �5  �1   �$  ���  �5  �5  �5  �1  �    ݨ  �M    �p  �	�   ��  �	�    5  
�5  I ��6  I ���  �5  6  �6   w�  ��  6  6  �6   �$  �3�  06  ;6  �6  X    �$  �'�  O6  Z6  �6  �1   �$  �v�  n6  ~6  �6  �1  �    ݨ  �M    �p  �	�   ��  �	�    �5  
�6  Z�6  ��   �
%��   %��  %E�  %��  %	�  %��  %S�  %��    [��6  ��  �7  ��  ��  7  ,7  �7  V4  �7   �  h�  @7  K7  �7  X    �  ��  _7  o7  �7  �1  �    �  ~�  �7  �7  �7  X   �  �#   /��  @V4   /��  A�7  F �3   �6  
�7  �#  ��  �8  ��  R�  �7  �7  �8  �5  �7   �  �  8  8  �8  X    �  ��  18  A8  �8  �1  �    �  ��  U8  j8  �8  X   �  �#   /��  @�5   /��  A�7  F 5   �7  
�8   Z9  ��  S�  �8  �8  Z9  
5  �7   �  �  �8  �8  Z9  X    �  4�  �8  9  Z9  �1  �    �  ��  !9  69  Z9  X   �  �#   /��  @
5   /��  A�7  F a4   �8  
Z9  �  
e9  �  
p9  `�  <:  ��  ��  �9  �9  <:  �6  �7   �  �  �9  �9  <:  X    �  ��  �9  �9  <:  �1  �    �  �  :  :  <:  X   �  �#   /��  @�6   /��  A�7  F �5   {9  
<:  S��  �  S	�    &  
[:  �  &  �  
r:  �  �  �  
�:    
�:  �
    [:  /  
�:  �
  
�:  W  
�:  �  W  r:  �  
�:  a  �1  �  �  -  ;  1�    
;  B�{  �  B�7    Bf    B]f  S  j=Y  a   �j�N  �   �Vn  �     B�7  �  -a  };  1�    L*  
};  �+  )L*  L*  *  �  D\  Dn  D�  D�  y  ��@     �      ��<  P (  T 5   ��  N�3  ���   N$5   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ��e�@     E       �<  i a5   �l ��@     -       �<  i d5   �h ��@     0       i f5   �d  -X   �<  1�    �  �3@     �      �">  P (  T �   ��  N�3  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ���4@     E       �=  i a5   �l �4@     -       >  i d5   �h 5@     0       i f5   �d  �  �1@     U       ��>  P (  T �   ��  x�3  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �T34i$  {	�     :  ��@     �       �Y?  P (  T 5   ��  x�3  �X�   x!5   �T3(  x-5   �Ph  x85   �L�)  y5   �H�D  yX   �D�@     ;       i$  {	�   �l  w  �0@     �       ��?  T �   F (  �  ��   �lfo �/�  �`��  �6�3  �X �	  �?  j�@     �      �@  	�  �:  ��n [:  ��u [:  �Xv [:  �Pw [:  �H �	  5@  ʑ@     �      �|@  	�  �:  ��n �[:  ��u �[:  �Xv �[:  �Pw �[:  �H �  |@     1       ��@  "O  U[:  �h -  �@            ��@  q,  =[:  �h 6�  
�@            �A  T &  "O  '[:  �h 6�  �@            �6A  T �  "O  'r:  �h   UA  Ȗ@     �      ��A  	�  �:  ��n r:  ��u r:  �Xv r:  �Pw r:  �H �  �A  (�@     �      �B  	�  �:  ��n �r:  ��u �r:  �Xv �r:  �Pw �r:  �H 8  h�@     1       �-B  "O  Zr:  �h �  L�@     �       ��B  T 5   F (  �  �5   �lfo �/�  �`��  �6�3  �X 6�+  95@     (       ��B  T 5   a 12  �hb #12  �` �5  �  �A     �      ��C  P �5  T �2  ��  N�B  ���   N$�2  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ���A     E       �C  i a5   �l a�A     -       �C  i d5   �h ��A     0       i f5   �d    z�A     �      �E  P �5  T �   ��  N�B  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ��j�A     E       �D  i a5   �l ��A     -       �D  i d5   �h ��A     0       i f5   �d  W  ��A     �      �KF  P �5  T   ��  N�B  ���   N$  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ����A     E       F  i a5   �l �A     -       +F  i d5   �h G�A     0       i f5   �d  �  *�A     �      �wG  P �5  T �   ��  N�B  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ��#�A     E       4G  i a5   �l r�A     -       WG  i d5   �h ��A     0       i f5   �d  ,  ,.@     J       ��G  F (  �  �!�   �Lfo �8�  �@��  �?�3  �� 7  �G  ��@     V      �H  	�  �:  �Xn �r:  �Ptl  �r:  �h�R  �r:  �` �  �{@            �JH  q,  L[:  �h �	  iH  .�@     H       ��H  	�  �:  �X"O  #[:  �P_�  $[:  �h {  m@            ��H  q,  I[:  �h 6  �{@            ��H  q,  8[:  �h �  I  ��@     V      �CI  	�  �:  �Xn �[:  �Ptl  �[:  �h�R  �[:  �` �	  bI  v�@            �I  	�  �:  �h"O  [:  �` &  �I  ��@            ��I  	�  �:  �h"O  r:  �` F  �I  "�@     H       �J  	�  �:  �X"O  #r:  �P_�  $r:  �h }  }�@            �2J  q,  =r:  �h �  QJ  ��@     �      �/K  	�  �:  ��n xr:  ��tl  {r:  �Ps �r:  �XTr  ��  ����@     �       �J  x �r:  �H ��@     z       �J  x �r:  �@ K�@     Q       K  .\  �r:  �� ��@     Q       .\  �r:  ��    ��@     1       �ZK  "O  Ur:  �h �  j�@            ��K  q,  Lr:  �h 6d  �@            ��K  q,  8r:  �h a4  �  ��A     �      ��L  P a4  T �2  ��  N�K  ���   N$�2  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ��{�A     E       �L  i a5   �l ��A     -       �L  i d5   �h ��A     0       i f5   �d    �A     �      �N  P a4  T �   ��  N�K  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ��ӿA     E       �M  i a5   �l "�A     -       �M  i d5   �h O�A     0       i f5   �d  _  ;�A     �      �:O  P a4  T   ��  N�K  ���   N$  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ��4�A     E       �N  i a5   �l ��A     -       O  i d5   �h ��A     0       i f5   �d  �  ��A     �      �fP  P a4  T �   ��  N�K  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ����A     E       #P  i a5   �l ۼA     -       FP  i d5   �h �A     0       i f5   �d  5  �  �A     �      ��Q  P 5  T �2  ��  NfP  ���   N$�2  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ���A     E       UQ  i a5   �l 3�A     -       xQ  i d5   �h `�A     0       i f5   �d  %  L�A     �      ��R  P 5  T �   ��  NfP  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ��<�A     E       �R  i a5   �l ��A     -       �R  i d5   �h ��A     0       i f5   �d  g  ��A     �      ��S  P 5  T   ��  NfP  ���   N$  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ����A     E       �S  i a5   �l �A     -       �S  i d5   �h �A     0       i f5   �d  �  ��A     �      �U  P 5  T �   ��  NfP  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ����A     E       �T  i a5   �l D�A     -       �T  i d5   �h q�A     0       i f5   �d  ,,  ��@     J       �mU  F (  �  �5   �Lfo �/�  �@��  �6�3  �� �3  �  T�A     �      ��V  P �3  T �2  ��  NmU  ���   N$�2  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ��M�A     E       \V  i a5   �l ��A     -       V  i d5   �h ɴA     0       i f5   �d  -  ��A     �      ��W  P �3  T �   ��  NmU  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��4  P�1  �Xݨ  S�<  ��k T5   ����A     E       �W  i a5   �l ��A     -       �W  i d5   �h !�A     0       i f5   �d  o  �A     �      ��X  P �3  T   ��  NmU  ���   N$  ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ���A     E       �X  i a5   �l U�A     -       �X  i d5   �h ��A     0       i f5   �d  �  e�A     �      �#Z  P �3  T �   ��  NmU  ���   N$�   ���'  N1`  ��3(  N?5   ��h  O5   ���)  O5   ���D  O#X   ��~4  P�1  �Xݨ  S�<  ��k T5   ��^�A     E       �Y  i a5   �l ��A     -       Z  i d5   �h گA     0       i f5   �d  �  �A     W       ��Z  P �5  T �2  ��  x�B  �h�   x!�2  �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�2    0   ��A     U       �G[  P �5  T �   ��  x�B  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �T34i$  {	�     m   �A     �       ��[  P �5  T   ��  x�B  �X�   x!  �P3(  x-5   �Lh  x85   �H�)  y5   �D�D  yX   �@A�A     ?       i$  {	�   �h  �   ìA     W       �~\  P �5  T �   ��  x�B  �h�   x!�   �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�     �   S,  ��@     N       ��\  T �   F (  �  8~\  �Hfo 8-�  �@��  84�3  �� �(  �\  6@     �       �]  	�  �3  �hs 	'X   �d �(  7]  �/@     �       �S]  	�  �3  �hstr 	1�1  �` "3  a]  �]  �  a:  &�B  ��  &�=  �%0  &�U  �6�    7S]  �[  �]  F{@     K       ��]  a]  �hj]  �dv]  �X�]  �P   �]  �q@     7      �-^  	�  �:  �Htl  �r:  �@"O  �"r:  ��*L  �r:  �X �  L^  np@     7      ��^  	�  �:  �Htl  �r:  �@"O  �!r:  ��M�  �r:  �X �  �^  �o@     j       ��^  	�  �:  �h"O  |r:  �` �  �^  z@     7      �_  	�  �:  �Htl  �[:  �@"O  �"[:  ��*L  �[:  �X a  �j@            �G_  q,  E[:  �h �  f_  �x@     7      ��_  	�  �:  �Htl  �[:  �@"O  �![:  ��M�  �[:  �X G  cj@            ��_  q,  B[:  �h 8<  �_  (p@     (       �`  	�  �:  �ha �!f:  �`b �1f:  �X }  1`  lx@     j       �M`  	�  �:  �h"O  |[:  �` "�  [`  e`  �  �:   *M`  �c  �`  *d@            ��`  [`  �h "  �`  �`  �  x:  &�=  �0  &�U  �)�   &$w  �65    7�`  �X  �`  x@     d       �a  �`  �h�`  �`�`  �X�`  �T 8�  0a  �o@            �=a  	�  �:  �h w  \a  |u@     �      ��a  	�  �:  ��"O  r:  ���/   r:  ��tl  r:  �X�  r:  �PpU  r:  �H �  ]u@            ��a  q,  Ir:  �h �  b  �r@     a      �fb  	�  �:  ��"O  Dr:  ��.\  D$r:  ��M�  Er:  �X*L  Fr:  �Ptl  Zr:  �H �  �q@            ��b  q,  Er:  �h �  Pp@            ��b  q,  Br:  �h 8�  �b  Rj@            ��b  	�  �:  �h �   l�A     W       �zc  P a4  T �2  ��  x�K  �h�   x!�2  �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�2    $!  �A     U       �d  P a4  T �   ��  x�K  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �T34i$  {	�     a!  x�A     �       ��d  P a4  T   ��  x�K  �X�   x!  �P3(  x-5   �Lh  x85   �H�)  y5   �D�D  yX   �@��A     ?       i$  {	�   �h  �!  !�A     W       �Ce  P a4  T �   ��  x�K  �h�   x!�   �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�     �!  ʪA     W       ��e  P 5  T �2  ��  xfP  �h�   x!�2  �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�2    "  u�A     U       �gf  P 5  T �   ��  xfP  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �T34i$  {	�     U"  ֩A     �       �g  P 5  T   ��  xfP  �X�   x!  �P3(  x-5   �Lh  x85   �H�)  y5   �D�D  yX   �@��A     ?       i$  {	�   �h  �"  �A     W       ��g  P 5  T �   ��  xfP  �h�   x!�   �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�     �,  
�@     G       ��g  T X   F (  �  3�2  �H��  3!�3  �@ �"  (�A     W       �zh  P �3  T �2  ��  xmU  �h�   x!�2  �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�2    #  ӨA     U       �i  P �3  T �   ��  xmU  �h�   x!�   �d3(  x-5   �`h  x85   �\�)  y5   �X�D  yX   �T34i$  {	�     I#  4�A     �       ��i  P �3  T   ��  xmU  �X�   x!  �P3(  x-5   �Lh  x85   �H�)  y5   �D�D  yX   �@[�A     ?       i$  {	�   �h  8m&  �i  "�A            ��i  	�  �2  �h "�%  �i   j  �  �2  Gcs  �2   *�i  ^�  #j  ȧA     Y       �4j  �i  �h�i  �` 8�$  Sj  v�@            �`j  	�  �2  �h "/$  nj  �j  �  �2  Gcs  �1   *`j  ~�  �j  �@     R       ��j  nj  �hwj  �` �#  p�A     W       �Ik  P �3  T �   ��  xmU  �h�   x!�   �`3(  x-5   �\h  x85   �X�)  y5   �T�D  yX   �P34i$  {	�     `  �  &�A     J       ��k  T `  x 
Ik  �Xy 
Ik  �Pyu  
`  �o 6�  �A            ��k  T Ik  x 
*Ik  �h �  ˦A     J       �l  T 5   x 
U2  �Xy 
U2  �Pyu  
5   �l �,  g�A     d       ��l  F �5  ��  ��B  �ht �*X   �d��  �<�  �X��  ��#  �`vsp �%�7  �P �,  ��A     �      �r  F �5  ��  q�B  ��t q(X   ����  q:�  ����  r�#  ��vsp r%�7  ���A           %m  �   x  �X #�!  ?m  �$ �?m  �@ <�  ��n  8�  ��  ^m  um  cm  ?m  nm  )?m   8�  ��  �m  �m  cm  �m  �m  
?m   98�  ��  �m  �m  cm   7�  �  �m  �m  cm  5    !~�  �r   !��  ��B  : {�   n  |�A     �       �^n  8�  �   8�  �   	�  ,n  �X
"r  �   ��   �T��  r  �X��  �B  �X# ;�  ��  �n  ��A     �       �8�  �   8�  �   	�  ,n  �X�   ��   �P��  r  �X��  �B  �X#  #�!  �n  �$ ��n  �� <�  �np  8�  7�  o  o  o  �n  o  )�n   8�  ��  +o  Ao  o  5o  ;o  
�n   98�  ��  Ro  Xo  o   7�  �  io  to  o  5    !~�  �r   !��  ��B  : � �o  ,�A     �       �p  ��  �   ��  �   	�  �o  �X
r  �   ��   �T��  r  �X��  �B  �X# ;�  ��  4p  R�A     �       ���  �   ��  �   	�  �o  �X�   ��   �P��  r  �X��  �B  �X#  # "  �p  �$ ��p  �� I��  �8�  ��  �p  �p  �p  �p  �p  )�p   8�  ��  �p  �p  �p  �p  �p  
�p   98�  ��  �p  �p  �p   7�  ��  
q  q  �p  5    !~�  �r   !��  ��B  : j�  fq  ܝA     �       ��q  ��  �   ��  �   	�  rq  �X
r  �   ��   �T��  r  �X��  �B  �X# ;�  ��  �q  �A     �       ���  �   ��  �   	�  rq  �X�   ��   �P��  r  �X��  �B  �X#   �  �p  ;o  �m  -  ǒA     �      �Dt  F �5  ��  '�B  ��~t ')X   ��~��  ';�  ��~��  (�#  ��~vsp (%�7  ��~�A     0       �r  i 85   �l ��A     �      �s  s A	�1  �`p E5   �\��A     J       s  i J5   �X ֖A     0       =s  i L5   �T �A     ,       as  i O5   �P 2�A     R       i Q5   �L  ��A     �      s V	�2  �@p Z5   ��y�A     V       �s  i _5   �� ϘA     0       �s  i a5   �� ��A     ,       !t  i d5   �� +�A     V       i f5   ��   B-  ��@           ��t  F (  ��  's'  ��fo <�  ����  C�3  ��p �t  �`��@     �      i �   �hҶ@     �      c 	�  �_   �  j-  .@     *       �>u  F (  �  � �1  �hfo �7�  �`��  �>�3  �X �  ]u  i@     �       ��u  	�  v9  �H@  %8�   �@WS  +0  �Xfra -[:  �P T  �u  �d@     �       ��u  	�  �:  �X"O  �r:  �P_�  �r:  �h =+  v  �h@     L       �v  	�  �;  �h   1v  �g@     �       �^v  	�  �:  �X"O  �[:  �P_�  �[:  �h �  }v  �f@     D      �3w  	�  v9  ���  45   ��WS  
0  �@�1  �   ���f  	�   �Xslb r:  ����  �:  �Pag@     ^       off �   �Hwg@     >       �  �:  ��   X+  Rw  �c@     O       �_w  	�  �;  �h �  ~w  :f@     X       ��w  	�  �:  �X_�  pr:  �h W  �w  ~e@     �       �x  	�  �:  �H"O  r:  �@B>  r:  �h`w  r:  �`�e@     I       M�  r:  �X  8�  7x  @d@     I       �`x  	�  a:  �Xp ��   �Padr �	�   �h "�*  nx  �x  �  �;    <    7`x  a4  �x  .b@     '       ��x  nx  �h "�*  �x  �x  �  �;  &�1  �1   7�x  S�  �x  �a@     2       �y  �x  �h�x  �` �-  c�A     d       �wy  F a4  ��  ��K  �ht �*X   �d��  �<�  �X��  ��#  �`vsp �%�7  �P �-  ��A     �      ��~  F a4  ��  q�K  ��t q(X   ����  q:�  ����  r�#  ��vsp r%�7  ����A           z  �   x  �X #!  -z  �$ �-z  �@ <�  ��{  8�  ��  Lz  cz  Qz  -z  \z  )-z   8�  � tz  �z  Qz  ~z  �z  
-z   98�  8�  �z  �z  Qz   7�  5 �z  �z  Qz  5    !~�  �r   !��  ��K  : �  {  x�A     �       �L{  8�  �   8�  �   	�  {  �X

  �   ��   �T��  r  �X��  �K  �X# ;�  ��  }{  ��A     �       �8�  �   8�  �   	�  {  �X�   ��   �P��  r  �X��  �K  �X#  #@!  �{  �$ ��{  �� <�  �\}  8�  � �{  |  �{  �{  |  )�{   8�  ��  |  /|  �{  #|  )|  
�{   98�  �  @|  F|  �{   7�  � W|  b|  �{  5    !~�  �r   !��  ��K  : ��  �|  (�A     �       ��|  ��  �   ��  �   	�  �|  �X
  �   ��   �T��  r  �X��  �K  �X# ;�  ��  "}  N�A     �       ���  �   ��  �   	�  �|  �X�   ��   �P��  r  �X��  �K  �X#  #p!  w}  �$ �w}  �� I��  �8�  q�  �}  �}  �}  w}  �}  )w}   8�  ��  �}  �}  �}  �}  �}  
w}   98�  E�  �}  �}  �}   7�  ��  �}  ~  �}  5    !~�  �r   !��  ��K  : �  T~  ؉A     �       ��~  ��  �   ��  �   	�  `~  �X
�~  �   ��   �T��  r  �X��  �K  �X# ;�  w�  �~  ��A     �       ���  �   ��  �   	�  `~  �X�   ��   �P��  r  �X��  �K  �X#   �}  )|  �z  �-  �~A     �      �,�  F a4  ��  '�K  ��~t ')X   ��~��  ';�  ��~��  (�#  ��~vsp (%�7  ��~�A     0       �  i 85   �l ��A     �      j�  s A	�1  �`p E5   �\��A     J       �  i J5   �X ҂A     0       %�  i L5   �T �A     ,       I�  i O5   �P .�A     R       i Q5   �L  ��A     �      s V	�2  �@p Z5   ��u�A     V       ��  i _5   �� ˄A     0       �  i a5   �� ��A     ,       	�  i d5   �� '�A     V       i f5   ��   '.  _~A     d       ���  F 5  ��  �fP  �ht �*X   �d��  �<�  �X��  ��#  �`vsp �%�7  �P Y.  �vA     �      �%�  F 5  ��  qfP  ��t q(X   ����  q:�  ����  r�#  ��vsp r%�7  ���vA           :�  �   x  �X #�   T�  �$ �T�  �@ <�  �ރ  8�  {�  s�  ��  x�  T�  ��  )T�   8�  #�  ��  ��  x�  ��  ��  
T�   98�  ��    Ȃ  x�   7�  ��  ق  �  x�  5    !~�  �r   !��  �fP  : ��  5�  trA     �       �s�  8�  �   8�  �   	�  A�  �X
1�  �   ��   �T��  r  �X��  fP  �X# ;�  n�  ��  �qA     �       �8�  �   8�  �   	�  A�  �X�   ��   �P��  r  �X��  fP  �X#  #�   ��  �$ ���  �� <�  ���  8�  $�  �  /�  �  ��  (�  )��   8�  �  @�  V�  �  J�  P�  
��   98�  	�  g�  m�  �   7�  �  ~�  ��  �  5    !~�  �r   !��  �fP  : ��  ڄ  $tA     �       ��  ��  �   ��  �   	�  �  �X
+�  �   ��   �T��  r  �X��  fP  �X# ;�  7�  I�  JsA     �       ���  �   ��  �   	�  �  �X�   ��   �P��  r  �X��  fP  �X#  #�   ��  �$ ���  �� I��  �8�  ��  ��  Ѕ  ��  ��  Ʌ  )��   8�  �  �  ��  ��  �  �  
��   98�  �  �  �  ��   7�  n �  *�  ��  5    !~�  �r   !��  �fP  : o {�  �uA     �       ���  ��  �   ��  �   	�  ��  �X
%�  �   ��   �T��  r  �X��  fP  �X# ;�  ��  �  �tA     �       ���  �   ��  �   	�  ��  �X�   ��   �P��  r  �X��  fP  �X#   �  P�  ��  �.  �jA     �      �S�  F 5  ��  'fP  ��~t ')X   ��~��  ';�  ��~��  (�#  ��~vsp (%�7  ��~�lA     0       ч  i 85   �l �mA     �      ��  s A	�1  �`p E5   �\�nA     J       (�  i J5   �X �nA     0       L�  i L5   �T �nA     ,       p�  i O5   �P *oA     R       i Q5   �L  |oA     �      s V	�2  �@p Z5   ��qpA     V       �  i _5   �� �pA     0       �  i a5   �� �pA     ,       0�  i d5   �� #qA     V       i f5   ��   6)  y�  ��@     *       ���  T X   	�  �3  �h�  	X   �d �.  [jA     d       ��  F �3  ��  �mU  �ht �*X   �d��  �<�  �X��  ��#  �`vsp �%�7  �P �.  �bA     �      ���  F �3  ��  qmU  ��t q(X   ����  q:�  ����  r�#  ��vsp r%�7  ���bA           ��  �   x  �X #�  ��  �$ ���  �@ <�  �G�  8�  ��  ܊  �  �  ��  �  )��   8�  `�  �  �  �  �  �  
��   98�  ��  +�  1�  �   7�  6�  B�  M�  �  5    !~�  �r   !��  �mU  : ��  ��  p^A     �       �܋  8�  �   8�  �   	�  ��  �X
��  �   ��   �T��  r  �X��  mU  �X# ;�  ��  �  �]A     �       �8�  �   8�  �   	�  ��  �X�   ��   �P��  r  �X��  mU  �X#  #    b�  �$ �b�  �� <�  ��  8�  ��  ��  ��  ��  b�  ��  )b�   8�  ��  ��  ��  ��  ��  ��  
b�   98�  � Ќ  ֌  ��   7�  ��  �  �  ��  5    !~�  �r   !��  �mU  : ��  C�   `A     �       ���  ��  �   ��  �   	�  O�  �X
��  �   ��   �T��  r  �X��  mU  �X# ;�  d ��  F_A     �       ���  �   ��  �   	�  O�  �X�   ��   �P��  r  �X��  mU  �X#  #P   �  �$ ��  �� I��  �8�  d "�  9�  '�  �  2�  )�   8�  �  J�  `�  '�  T�  Z�  
�   98�  <  q�  w�  '�   7�  ��  ��  ��  '�  5    !~�  �r   !��  �mU  : ��  �  �aA     �       �"�  ��  �   ��  �   	�  ��  �X
��  �   ��   �T��  r  �X��  mU  �X# ;�   S�  �`A     �       ���  �   ��  �   	�  ��  �X�   ��   �P��  r  �X��  mU  �X#   Z�  ��  �  !/  �VA     �      ���  F �3  ��  'mU  ��~t ')X   ��~��  ';�  ��~��  (�#  ��~vsp (%�7  ��~�XA     0       :�  i 85   �l �YA     �      ��  s A	�1  �`p E5   �\�ZA     J       ��  i J5   �X �ZA     0       ��  i L5   �T �ZA     ,       ِ  i O5   �P &[A     R       i Q5   �L  x[A     �      s V	�2  �@p Z5   ��m\A     V       O�  i _5   �� �\A     0       t�  i a5   �� �\A     ,       ��  i d5   �� ]A     V       i f5   ��   �  ۑ  �VA     ;       ��  	�  ,2  �h 6  6  ��@            ��  T U2  x 
.�  �h S/  �UA     �       ���  ��  iI2  �HJ�  i.I2  �@�UA     0       |�  tmp o5   �\ -VA     0       tmp s5   �X  �9  ��  �QA     �      �,�  	�  B:  ��}t X   ��}��  /�  ��}��  J�#  ��}  <�  	0rB     uTA     |       p 4	[2  �X  -_   <�  1�   
 
,�  �9  `�  �QA     )       �z�  	�  B:  �hc X   �d �9  ��  ZQA     1       ���  	�  B:  �hc �1  �`n )�   �X �)  ߓ  h-@     &       ���  	�  �3  �h/&  	M�1  �` �'  n/  �@     I       �K�  T s'  F (  �  3��  �H��  3!�3  �@ 2  �/  �,@     E       ���  T �1  F (  �  3K�  �H��  3!�3  �@ "(  ��  ��  �  �3  &�)  	�3   *��  �  �  �,@     4       ��  ��  �h��  �`    �  �Z@     �      �%�  	�  v9  ��~p �1�   ��~�Z@     �      ߕ  �  �5   �\bkt �:  �P`v  L*  ���  �:  ��d[@     *      ��  slb 	r:  �H �\@     �      slb 	r:  �@Cx  #L*  ��  �^@     �       @  :�   ��fra ;[:  ��Cx  =L*  ��~  9  D�  �MA     �      ���  	�  `9  ��}t X   ��}��  /�  ��}��  J�#  ��}  <�  	 qB     KPA     |       p 4	[2  �X  �8  Җ  bMA     )       ��  	�  `9  �hc X   �d �8  �  0MA     1       �2�  	�  `9  �hc �1  �`n )�   �X A8  Q�  bIA     �      ���  	�  �8  ��}t X   ��}��  /�  ��}��  J�#  ��}  <�  	�pB     !LA     |       p 4	[2  �X  �7  ߗ  8IA     )       ���  	�  �8  �hc X   �d 8  �  IA     1       �?�  	�  �8  �hc �1  �`n )�   �X o7  ^�  8EA     �      �͘  	�  �7  ��}t X   ��}��  /�  ��}��  J�#  ��}  <�  	�pB     �GA     |       p 4	[2  �X  "L  �  ��  U U2  �  ,2  &q  %U2   7͘  N�  "�  �DA     N       �3�  U U2  �  �X�  �P :  R�  �DA     )       �o�  	�  ,2  �h�  =   �` "�  }�  ��  �  ,2  &�  72   7o�  ��  ��  rDA     N       �Ǚ  }�  �X��  �P ,7  �  HDA     )       � �  	�  �7  �hc X   �d K7  �  DA     1       �F�  	�  �7  �hc �1  �`n )�   �X 6B  DA            �v�  T U2  x 
*U2  �h "C  ��  ��  �  !2    <    *v�  6.  ��  �+@            �Ú  ��  �h ")  њ  ۚ  �  !2   *Ú  9*  ��  �+@            ��  њ  �h �/  :=A     �      ��  A {9  ��  �{9  ��~s �)�1  ��~vsp �7�7  ��~|=A     �      ��  ��  ����  �#  �`�=A     c       ��  n ��   �h y@A     ~       Λ  w �5   �d �AA     �       q  	5   ��   "�9  �  #�  �  B:  &��  �6  Gvsp ,�7   *�  ��  F�  =A     *       �_�  �  �h
�  �`�  �X �(  ~�  �+@     ,       ���  	�  �3  �h�'  �  `)  ��  ��@     6       �՜  T s'  	�  �3  �h�  	s'  �P �)  ��  4+@     )       ��  T �1  	�  �3  �h�  	�1  �` "~(  %�  8�  �  �3    <    *�  *$  [�  (+@            �d�  %�  �h �)  ��  �*@     )       ���  	�  �3  �` �  ��  |V@     (       �̝  	�  k9  �h@  [�   �` 9  TU@     �       �[�  @  W0�   ��tc Y�   �`e b�   �Xf c�   �Pip d�   �His e�   �@�U@     :       i [�   �l  6  �T@            �˞  idx H6�   ��tc J�   �hs O5   �dip P�   �Xis Q�   �Pf R�   �H �/  D6A     �      ���  A �8  ��  ��8  ��~s �)�1  ��~vsp �7�7  ��~�6A     �      ��  ��  ����  �#  �`�6A     c       o�  n ��   �h �9A     ~       ��  w �5   �d �:A     �       q  	5   ��   "�8  ş  �  �  `9  &��  
5  Gvsp ,�7   *��  E�  
�  6A     *       �#�  ş  �hΟ  �`ڟ  �X �   60  s�@     +       �f�  T �   a 	#�  �hb 	##�  �` 60  N/A     �      �R�  A �7  ��  ��7  ��~s �)�1  ��~vsp �7�7  ��~�/A     �      ��  ��  ����  �#  �`�/A     c       
�  n ��   �h �2A     ~       -�  w �5   �d �3A     �       q  	5   ��   "�7  `�  ��  �  �8  &��  �5  Gvsp ,�7   *R�  |�  ��  $/A     *       ���  `�  �hi�  �`u�  �X kO�  %5   �A     �      �k�  H V�  A�  %��  ��yV�  fmt %-�1  ��y��  %Ak�  ��y��  &	5   �l�A     t      � 8�   �`h  B5   �\�U  [�   �XV \�   �T#p  ��  c 3X   ��~ #�  â  res �$�2  �Hc �X   �G #�  �  res �$�2  ��c �X   �� #   �  res �$�2  ��c �X   �� #0  R�  � �M   ��~c �X   ����  �5   �� #`  ��  � 	M   ��~c 
X   ����  5   �� #�  �  /�  5   ��W�  q�  ��z� 5M   ��~��  65   ��c 7X   ���A     F       c /#X   ��  � A     @      R�  res F$�2  ��c GX   ��~� _��  ��~ H�  � d[2  ��~   �   -X   ��  ��     �   ]0  X(A     �      �u�  A �6  ��  ��6  ��~s �)�1  ��~vsp �7�7  ��~�(A     �      ��  ��  ����  �#  �`�(A     c       -�  n ��   �h �+A     ~       P�  w �5   �d -A     �       q  	5   ��   "7  ��  ��  �  �7  &��  V4  Gvsp ,�7   *u�  ~�  ȥ  .(A     *       ��  ��  �h��  �`��  �X k��  %5   �A     �      ���  H e�  A�  %�  ��ye�  fmt %-�1  ��y��  %Ak�  ��y��  &	5   �l2A     t      � 8�   �`h  B5   �\�U  [�   �XV \�   �T#�  ��  c 3X   ��~ #   �  res �$�2  �Hc �X   �G #P  �  res �$�2  ��c �X   �� #�  :�  res �$�2  ��c �X   �� #�  u�  � �M   ��~c �X   ����  �5   �� #�  ��  � 	M   ��~c 
X   ����  5   �� #  .�  /�  5   ��W�  q�  ��z� 5M   ��~��  65   ��c 7X   ���A     F       c /#X   ��  A     @      u�  res F$�2  ��c GX   ��~� _��  ��~ H@  � d[2  ��~   6�0  �V@     +       �˨  T �   a #�  �hb ##�  �` "�  ٨  �  �  ,2  &�  *=2   7˨  %'  �  �)@     V       �#�  ٨  �h�  �` 8}  B�  (A            �O�  	�  ,2  �h "  ]�  p�  �  ,2    <    7O�  g  ��  �)@            ���  ]�  �h "_  ��  ��  �  ,2   7��    ש  �)@     #       ��  ��  �h 5�  aM   �A     2       �/�  M   �h5   �d�  �X  ?�  	HrB      -_   ?�  1�    
/�  ��  ,�   �A     ;      �R�  ݨ  ,$�2  ��|@  ,3�   ��|��  ,@�   ��|Q ,M�  ��|z�  -u3  �P�A     �       ��  �z  4
�   �hH�  ��  6�   ��}  �A     �       i G�   �`�A     �       �z  H�   �XH�  ��  J�   ��}    ��  ��   QA     ;      �`�  ݨ  ��   ��|@  �,�   ��|��  �9�   ��|Q �F�  ��|z�  �u3  �P�A     �       �  �z  �
�   �hH0  ��  �   ��}  �A     �       i �   �`�A     �       �z  �   �XH`  ��  �   ��}    ��  �5   A     D       ���  �  ��  �Xd ��  �o TM�  �5   �A            �֬  Q ��  �h T@�  �5   �A            �
�  Q ��  �h lo�  ��A            �:�  Q ��  �h F�  �5   tA     [       �g�  �  ��~ m��  �A     [       ���  �  ��~ m� �� A     [       ���  �  ��~ ��  �5   # A     �       �.�  out �.�  ���  �'�1  ����  �>k�  ��vs ��#  �@p ��5  �� M   ��  �5   o�@     �       ���  out �.�  ��~�  �&�1  ��~0��  �
�   ��~JC  �5   ��~ �  �		  9�@     6       ��  ػ  �.�  �hn �'�  �`�  �.5   �\Q �;�  �P  (�  	 rB      �   -_   (�  1�    
�  �  �		  ��@     �      ���  ػ  �.�  ��~n �&�  ��~Q �/�  ��}ݨ  �M   �X\�  �	�   �Pk �	�   �H ]�  �5   	�@     z       ���  �^  ��1  �Xez  �5   �l T��  �5   ��@            �(�  Q ��  �h T�  �5   ��@            �\�  Q ��  �h l�  ���@            ���  Q ��  �h :�  ~5   ��@     /       ��  �  ~�  �h�  ~)�  �`  ��  	rB      �  -_   ��  1�    
�  ��  y5   m�@     /       �U�  �  y�  �h�  y9[�  �`  ��  	rB      �  FU�  	 u�   ;�@     2       �ı  ݨ  u�2  �h@  u*�   �`��  u8�   �XQ uE�  �P ��  q�   	�@     2       �(�  ݨ  q�   �h@  q#�   �`��  q0�   �XQ q=�  �P ��  oH  ��@     .       �o�  H  �l�  �`  ��  	 rB      7�  nH  ��@     *       ���  �2  �l  (�  	�qB      �  mH  ��@     .       ���  �2  �l�  �`  �  	�qB      -_   �  1�    
��  .�  lH  `�@     #       �A�    (�  	�qB      (�  kH  5�@     +       ���  �  �h  �  	�qB      D�  j5   �@     .       �ǳ  �  �h5   �d  �  	�qB      >�  i5   ��@     /       ��  �2  �h�  �`  �  	�qB      -_   �  1�    
�  �  hH  ��@     .       �j�  �2  �l�  �`  �  	�qB      ��  g
��  x�@     2       ���  ��  �h5   �d�  �X  �  	�qB      �2  F��  '�  fH  M�@     +       ��  �  �h  �  	�qB      ~�  M5   p�@     �       ���  �^  M�1  ��z�  Nu3  �`�z  P	�   �hlen Q	�   �X��  ^	�   �P��@     O       ��  S
�   �H  ��  I5   Y�@            �̵  c I5   �l �  F5   5�@     $       ���  c F5   �l 3�  B5   �@     "       �@�  c B5   �l�  B�  �` x�  <5   ��@     I       ���  c <5   �\�  < �  �Pd =X   �o n3	 85   ��@            �n�  45   ��@            ���  05   ��@            ��  �  0�  �h ��  ,5   f�@            �6�  �  ,�  �h }�  (5   A�@     %       �z�  �^  ("2  �h�  (;�  �` ��  #5   ��@     P       ���  �^  #+2  �h�  #D�  �` 2�  5   ��@     "       � �  c 5   �l�  �  �` w�  5   ��@     K       �P�  c 5   �\�  !�  �Pd X   �o �  �M   ��@     �       ���  ݨ  �S   �X�1  �-�   �P�  �H�  �H  �  	�qB     ��@     �       i ��   �h��@     �       c �5   �d   ��  �5   k�@     D       �I�  �  ��  �Xc �X   �g5�  ��   �h ��  �5   <�@     /       ���  �2  �hk�  �`  ��  	�qB      ��  �5   �@     /       �׹  �2  �hk�  �`  (�  	�qB      ] �5   ��@     x       ��  �2  ��~0  �  	�qB      ��  �5   �@     x       �Y�  �2  ��~0  ��  	�qB      ��  �5   ��@     7       ���  ��  �h�   �`�2  �Xk�  �P  (�  	xqB      ��  �5   ��@     7       ��  ��  �h�   �`�2  �Xk�  �P  �  	hqB      -_   �  1�   	 
�  ��  �5   7�@     x       �o�  ��  ��~�   ��~�2  ��~0  ��  	`qB      ��  �5   ��@     x       �»  ��  ��~�   ��~�2  ��~0  (�  	PqB      [ �5   ��@     3       ��  �  �h�2  �`k�  �X  (�  	@qB      ��  �5   Y�@     3       �`�  �  �h�2  �`k�  �X  �  	0qB      \ �5   ��@     x       ���  �  ��~�2  ��~0  ��  	(qB      ��  �5   i�@     x       ���  �  ��~�2  ��~0  (�  	qB      ��  �5   6�@     3       �[�  ݨ  �$2  �h�  �C2  �`��  �Zk�  �X  ��  	qB      � �5   ��@     �       �н  ݨ  �S   ���  �>2  ����  �Uk�  ��vs ��#  �@p �a4  �� �  �5   ��@     �       �W�  ݨ  � S   ��~�1  �/�   ��~�  �2  ��~��  �1k�  ��~vs ��#  ��p �5  �� ��  �5   ��@     /       ���  �  �#2  �h��  �:k�  �`  �  	�pB      ��  �5   k�@     /       ��  �  �$2  �h��  �;k�  �` e�  �5   �@     `       ���  �  ��  �H�  �=2  �@��  �Tk�  ��z�  �u3  �h��	��  U��  n�  �  s�  V�  5    U��  ��  ��  s�  ��  )V�   U��  ��  ��  s�  ��  ��  
V�   U��  Ϳ  ӿ  s�   oh�  �X   ��  N�@     b       �%�  	�  X�  �Xc �	X   �oִ  ��   �` oo�  �X   L�  ��@     [       �|�  	�  X�  �X
s�  c �	X   �oִ  ��   �` !z�  �u3   !D�  �5    A�  �V�  �P ��  �5   ��@     }       ��  �  ��  ���  �>2  ����  �Uk�  ��vs ��#  �@p ��3  �� ��  �5   ��@     �       ���  ݨ  �#2  ��}�  �B2  ��}0��t�  V��  ~�  ��  ��  e�  5    V��  ��  ��  ��  ��  )e�   V��  ��  ��  ��  ��  ��  
e�   V��  ��  ��  ��   ph�  �X   �  ��@            ��  	�  O�  �h po�  �X   C�  ��@     0       �U�  	�  O�  �h
��   Aݨ  ��1   AD�  �5    A�  �e�  ��~��  ��   ��~JC  �	5   ��~ ��  z5   ��@     �       ��  ݨ  zS   ��~�  z=2  ��~0��  {
�   ��~JC  }5   ��~ �  s5   G�@     �       ���  ݨ  sS   ��~�1  s.�   ��~�  sO2  ��~0��  t
�   ��~JC  v5   ��~ g�  o5   ��@     x       ���  �  o"2  ��~0  �  	�pB      �� %�@     �       �#�  � �   �h@  0�   �di I�2  �X >�  �5   n�@     �       �w�  �  �#2  ��~0��  �
�   ��~JC  �5   ��~ >f�  �5   ��@     �       ���  �  ��  ��~�  �<2  ��~0��  �
�   ��~JC  �5   ��~ > �  �5   �@     �       �?�  �  ��  ��~�  �=2  ��~0��  �
�   ��~JC  �5   ��~ ��  ���@     2       ���  �  ��  �hݨ  �7S   �`  �  	�pB      >2�  ��  ��@     3       ���  �  �&2  �h)  �G2  �`�  �^�  �X  ��  	�pB      > �  �M   v�@     +       �8�  ݨ  �M   �h  �  	�pB      >s�  ��  S�@     #       �n�    ��  	�pB      >5�  �5   �@     5       ���  ��  �5   �l<�  �(�1  �`_�  �65   �hC�  �L�1  �X  (�  	�pB      >t�  �5   ��@     �       �S�  @�  ��1  �XC�  �*�1  �P  �  	�pB     ��@     /       e �	5   �l  >�  �5   n�@     +       ���  �  ��1  �h  �  	�pB      Z6  ��  �'A     O       ���  	�  �6  �Xstr ��1  �Pn �&�   �H�'A     8       i ��   �h  ;6  �  x'A     S       �Y�  	�  �6  �Xstr ��1  �P�'A     @       i ��   �h  6  x�  ,'A     L       ���  	�  �6  �hc �X   �d 6  ��  "&A     	      ��  	�  �6  �H  �  	;rB     G&A     �       �  �	�   �h��  �	M   �P  "�5  �  �  �  �6   *�  ;	 <�  �%A     .       �E�  �  �h �5  d�  �%A     O       ���  	�  �5  �Xstr ��1  �Pn �&�   �H�%A     8       i ��   �h  e5  ��  P%A     S       ��  	�  �5  �Xstr ��1  �P`%A     @       i ��   �h  8F5  %�  �$A     Q       �?�  	�  �5  �hc |X   �d ""5  M�  o�  �  �5  &ݨ  yM   &�p  y&�    *?�  ��  ��  �$A     6       ���  M�  �hV�  �`b�  �X 8�4  ��  d$A     c       ��  	�  5  �Xstr l�1  �Pn l&�   �Ht$A     P       i n�   �h  8�4  1�  �#A     g       �l�  	�  5  �Xstr d�1  �P$A     X       i f�   �h  8�4  ��  �#A     <       ���  	�  5  �hc _X   �d "n4  ��  ��  �  5  &ݨ  \M    *��  �  ��  �#A     &       ���  ��  �h��  �` 4  �  L#A     M       �E�  	�  \4  �hstr R�1  �`n R&�   �X �3  d�  �"A     e       ���  	�  \4  �Xstr M�1  �P �3  ��  �"A     H       ���  	�  \4  �hc HX   �d "�3  ��  ��  �  \4  &�  E�   *��  1  �  x"A     &       ��  ��  �h��  �` "�'  �  C�  �  �2  qݨ  "�2  q@  "(�    *�  ��  f�  �@     *       ��  �  �h(�  �`5�  �X �  ��  M@     6       ���  	�  g2  �`c 63�  �\�>  7�  �h r2  2��  ��  �  g2    <    7��  .  �  �)@            ��  ��  �h h  rN  2/�  >�  �  g2  �   7�  �  a�   )@     �       �r�  /�  �h8�  �` "�  ��  ��  �  g2   7r�  K  ��  �(@     \       ���  ��  �h �.  ^  �   �(@            ���  @  #�   �hp /�   �` 8P1  �  �M@            �&�  	�  �1  �h 61  E�  �M@     B       �e�  	�  �1  �h  u�  	rB      -_   u�  1�    
e�  6�  �M@            ���  x )�   �h "  ��  ��  �  �0   *��  1~  ��  :M@     Q       ���  ��  �h +i	  +J  s&  %*  "s�  %*  " ~   M;  �  �	 �  ��A     �      4 �  �9   �  �>  L   int Q  _   j   _   �  j   �o  _   �  	�  
�	 4_   R�A     H       ��   � 4e   �Xsrc 4<�   �Pn 59   �h q   �   
7
 0�   �A     7       �C  � 0�   �hsrc 0'C  �`len 03-   �X I  
�
 'L   ��A     ]       ��  e 'L   �\ݨ  '_   �P�	 ',-   �Hs (_   �h �	 
_   ~�A     @      ��  e 
L   �\s �   �h 
�	 
9  L�A     2       �9  9  �hD  �d-   �X  `  	 |B      D  9  |  D  q   `  9    P  
k
 -   !�A     +       ��  �  �h  �  	|B      K  �  q   �  9    �  �
 �
9  ��A     f       �@  s �!�  �Xc �,D  �T@  �6-   �Hr
  �  �`��A     H       i -   �h  �	 �
9  ��A     3       ��  ?  �h�  �`�  �X  �  	|B      9  �  G
 �
9  Y�A     /       ��  �  �h�  �`  �  	|B      �
 �-   *�A     /       �%  �  �h�  �`  �  	 |B      R	 �
9  ��A     .       �k  �  �hD  �d  `  	�{B      (
 �
9  ��A     /       ��  �  �h�  �`  `  	�{B      \
 �-   ��A     /       ��  �  �h�  �`  `  	�{B      0
 �
9  p�A     .       �=  �  �hD  �d  �  	�{B      u	 �L   =�A     3       ��  �  �h�  �`-   �X  `  	�{B       �L   
�A     3       ��  ?  �h�  �`-   �X  `  	�{B      ?
 �L   ��A     3       �'  �  �h�  �`-   �X  `  	�{B      �
 �L   ��A     /       �m  �  �h�  �`  `  	�{B      �
 �L   y�A     /       ��  �  �h�  �`  �  	�{B      }	 �
9  F�A     3       �  ?  �h�  �`-   �X  `  	�{B      d
 �
9  �A     /       �G  ?  �h�  �`  �  	�{B      l	 �
9  ��A     3       ��  9  �h�  �`-   �X  �  	�{B      q   �  9    �    �
9  ��A     3       ��  ?  �h�  �`-   �X  `  	�{B      �	 �
9  ~�A     3       �F  ?  �h�  �`-   �X  `  	�{B      �	 �
9  O�A     /       ��  ?  �h�  �`  �  	�{B      �	 ��  �A     2       ��  �  �h�  �`L   �\  �  	�{B      �  �
 �9   ��A     2       �/	  �  �h�  �`L   �\  `  	x{B      �	 �}	  ��A     2       �}	  �  �h�  �`L   �\  `  	p{B      �  �	 ��	  ��A     2       ��	  �  �h�  �`L   �\  �  	h{B      �  �	 �
  X�A     /       �
  �  �h�  �`  `  	`{B      E  �	 �l
  )�A     /       �l
  �  �h�  �`  �  	X{B      i	  �	 ��
  ��A     /       ��
  �  �h�  �`  �  	Q{B      J  Z	 �_   ��A     \       �
  s ��   �Xc �$L   �Ti �	-   �h U
 �_   r�A     ,       �_  s �e   �h
 �9�   �` �_   	�C      
 �_   H�A     *      ��  s �!e   �Xdel �;�   �Pm �R�  �H  �  	H{B     tok �_   �hp �_   �` _   �  	 �_   ��A     �       ��  s ��   �Hd	 �)�   �@��A     �       i �-   �h��A     x       �
 ��  �g��A     a       j �-   �X    l  �
 �-   (�A     m       ��  s ��   �X�	 �*�   �Pn �	-   �h  �_   ��A     p       �A  s ��   �Xc �"L   �Tp �	-   �`��A     J       i �-   �h  0 �_   J�A     n       ��  s ��   �X�	 �*�   �Pn �	-   �h �
 }-   ��A     m       ��  s }�   �X�	 }+�   �Pn ~	-   �h z
 r_   t�A     i       �#  s r�   �Xc r!L   �Ti s	-   �h �
 k�   �A     Y       ��  s kC  �Xc k!L   �T@  k+-   �Hr
 l�  �`2�A     ;       i m-   �h  �  �  �  �
 f-   ��A     3       �  � f!e   �hsrc f>�   �`�1  fJ-   �X  `  	@{B      ( UL   a�A     �       ��  a U�   �Xb U(�   �P�1  U2-   �Hi V	-   �hy�A     k       �
 Z�  �gN
 [�  �f  �
 PL   <�A     %       ��  a P�   �hb P(�   �` �
 @L   ��A     r       �R  a @�   �Xb @'�   �Pi A	-   �h��A     Z       �
 C�  �gN
 D�  �f  v	 5L   X�A     r       ��  a 5C  �Xb 5'C  �P@  51-   �Hh�A     [       i 6-   �hz�A     B       �
 7�  �gN
 8�  �f   �
 (_   ��A     �       �i  � ( e   �Hsrc (=�   �@�1  (I-   ���.  )_   �h�.  *�   �`i ,	-   �X �
 $_   ��A     ;       ��  � $e   �hsrc $<�   �` �
 _   �A     �       �&  �  e   �Hsrc 2�   �@�1  >-   ���.  _   �h�.  �   �`i 	-   �X �
 _   ��A     S       �� e   �Xsrc 1�   �P�.  _   �h�.  _   �`  �   �<  �  � �  ��A           : �  �  �  �  N   �  �  �  int �  �  �N   �  B     4q   �  �N   �  j   �  j   r  �  8 @x c   �   �  c    C ; c   �   c    � 0^ c   "  �  c      # � c   K  c   �   c   |   U , c   t  c     �      � � c   c   }  �       	�  �  
�  �   Y�A     C       ��  �  @�  �X)  @+c   �Tret Ac   �l �   �A     :       �  fd ;c   �l 	c   �   ��A     W       �|  �  0�  �X   0)c   �Tfd 05  �H_fd 1c   �l 	�   "  a�A     g       �  fd c   �\�  �   �Ps�  )c   �Xͨ  8|  �Hoff  	�   �h� !c   ret #}   �` 	�   K   �A     a       �}  fd c   �\buf   �P��  )�   �H5�  9  �@ret c   �l� c    	�  t  ��A     f       �fd c   �\ݨ  $}  �P��  3�   �HM C  �@ret c   �l  �   �=  �  � �   0          �; �  �:   )   �  �  �  E  6  std  ?  �  	�   q  	F  �  	?  	�  	�  �   �   �   
T   	�  	q  �   �   �   
T   T ?  v ?    f   �  	O  q  	F  �  	?  	�  	,  �     !  
c   	�  	�  �   9  ?  
c   T ?  v ?   �   � 	`u  �U  	a   T �   � 	[�  �U  	\Y  T Y   � 	`�  �U  	av  T    -�  	j>�  O !� �  �  T      � � �    T Y      -�  	j>�   � �  2  T �     -�  	j>a   l  ?    s   �   F  �   O  �  �  �  w  �  �  int �  �  
�:     4�  �  frg 	5  E3  	�  ��  �   d^  	�    4j  F    �  G  �  .  �   red h^   �o  0�  �o  �F  O  U  
?   �o  �D  i  t  
?  E   �  �z  K  �  �  
?  E   tl  Q   �  Q  pU  Q  �I   Q  �D  !Q   [r  "	  ( .  q  %dV  5�   h 8<  ?    �   pl  =�n  �  4  �   �p  B�^  �  N  �   lU  Ef|  �  h  �   �I  I�  �  �  �   �D  LE  �  �  �   	<3  Pfm  �  �  �  
�   !�E  U�L  ?  �  �   !�_  Z�M  ?  �  �    c  djw    
  
�    c  gar    )  
�  �   �  i
J    A  L  
�  �   	��  op  �  d  j  
�   "�D  |+G    �  
�  �   "��  ��z  �  �  
�  �  �   "5>  ��@  �  �  
�  �  �   "�F  �4\  �  �  
�  �   #�  Dj  	    
�  �   $O  $d  *  :  
�  �  �   $�U  D�6  P  `  
�  �  �   $�  x�E  v  �  
�  �   $ q  �nq  �  �  
�  �   $�9  1y  �  �  
�  �   #�=  Ӏ  �  �  
�  �   #�z  #�8  �    
�  �   %L  0Nx  ?    #  
�   %L  9�/  ?  =  W  
�  �  	       &?3  �Q   D �  T �  '�P  �  A �   �  (�5  �D  )�j  )��  )��  )�4  )�N  )��  *�   #Z|  �@  �  �  
  v   #�F  �V�  
    
  �   &�R  �v  T �  '�P  �  L v  A �   .H  5�   h 8�4  ?  j  �   pl  =&i  �  �  �   �p  B�Z  �  �  �   lU  EP  �  �  �   �I  I�f  �  �  �   �D  L}S  �  �  �   	<3  PO]  �  	  
	  
&   !�E  U�g  ?  %	  �   !�_  Z)?  ?  @	  �    c  d8  T	  Z	  
&    c  g~u  n	  y	  
&  1   �  i'O  7  �	  �	  
&  1   	��  oAs  �  �	  �	  
&   "�D  |�k  �	  �	  
&  �   "��  ��0  �	  �	  
&  �  �   "5>  ��A  
  $
  
&  �  �   "�F  �X  9
  D
  
&  �   #�  �1  Y
  d
  
&  �   $O  
e  z
  �
  
&  �  �   $�U  DxT  �
  �
  
&  �  �   $�  xfC  �
  �
  
&  �   $ q  �{l  �
  �
  
&  �   $�9  E}      
&  �   #�=  �9  (  3  
&  �   #�z  #�`  H  S  
&  �   %L  0�_  ?  m  s  
&   %L  9�a  ?  �  �  
&  �  	  =  =   &?3  �Q   D �  T �  '�P  �  XA �   D  +�~  �)��	  )��	  )��	  )��  )��  )��  *D   #Z|  �<R  6  A  
C  v   #�F  �/L  V  a  
C  �   &�R  �v  T �  '�P  �  XL v  A �    �  4j  F    �  ,��  �$�   Q  �  ��  �   ʃ  QS   �  �U  H�	�  �U  ���      
�  �  �  )    �U  ���  .  9  
�  �   �  �
`D  �  Q  \  
�  �   	��  ��b  ?  t    
�  Q   �U  ��   WS  ��  p �5   �=  ��   �  �U  ��	l  *�   �U  �Pc  �  �  
�  �  )   �   �U  �z  	    
�  �   �  �4  �  ,  7  
�  �   �  ��  H�D  �w  L$H  ��  P�B  ��  X �  -%\  �R  �	�  .�  ��v  ?  �  
  �  �    �.   �	�  �.  �R�  �  �  
N   �E  �	X   �o  ��  �e  ��   1|  ��  "u  ��=    #  
Y  �   /u  (�t  8  C  
Y  d   0�  *�K  j  \  g  
Y  d   1�  ��o  Q  �  �  
Y  )    %�  L�g  Q  �  �  
Y  Q  )    $�  ~��  �  �  
Y  Q   $�I  �Ճ  �  �  
Y  Q  )    1WV  1	e;  )       
Y   2C  >�                         @       3�v  @ ~  3�`  A ~   �~  H�U  )     w   �.  W�N  )   �  )    3QC  j�  zz  l5   |  oK>  ?  �  w   ́  |5   ]C  5   4�D  �5    5�~  ��<  �      
Y  �   5��  &q  �  4  ?  
Y  �   5FS  %n^  �  X  c  
Y  )    #4  7:k  x  ~  
Y   #]  >�J  �  �  
Y  �   �[  �
�   �1  �X  �U  ��  L  ��  �=  �	)    eu  ��  (6sz     6tZ  X   �  74^  V�  $�B  X�;  '  2  
  Y   %�  [kt  Q  L  W  
  )    $�I  _p3  m  }  
  Q  )    $�  c"u  �  �  
  Q   %V  g�c  Q  �  �  
  Q  )    8ZD  lY   6sz     6tZ  X   9 3  � D     
�   ݨ  �   '�  :   '� :    :� �  ;get  � �  Z  `  
�   <� %)�   "� P �  �  =�  
�   T     >�v  �+.  >�D  �7�  >�D  �7�  ?8 �	  � 0 �  �  
�   ݨ  �   @�  :   �'� :    A� �|  ;get   j  1  7  
�   <� %)�   "E � i  t  B�  i  C�   
�  �   T �   9� �  � � �  �  
   ݨ     '�  :   '� :    D+ ;get  t *  �  �  
0   <� %)|   "� � !  ,  B�  !  CY   
0  �   T     E�  E�  .  F�  F.  GE�  #Q    #Q  C|  y    
	   #Q  �B  �  �  
	     �   k    �  �  
	     �~  �A  �  �  
	   |  �  �  �  
	   H̀  �    X  X  	  F  FX  H  q  Imap vU  �  E  P  
q  )    J]   �f  `  
q  �  )        q  j %>  �  �  Kr  -�  �  L�  �  M:     F   3  �  �  F�  F�  �  Fl  F�  q  �  �  F�  F�  F�  F�  v  �    D  &  F�  FD  F�  �  C  �  N  �  Y  F�  F�  L5   �  M:    p  �{    �7  I  f  W  ]f  �  =Y  �  �N  �  Vn  �  �7  �  L�  �  M:    �  �  L�  �  N:   � 	  �      |    L�  *  M:    F  �  0  O@	  I  S  P�  ,   Q;  k v  ��A            �  RI  �h O!  �  �  P�  I  S�R  �v   T  ` �  ��A     $       ��  R�  �hR�  �  O�  �  �  P�  �   Q�  Y   ��A            �  R�  �h Fv  U�  ��A     
       �R  T   Vx *  �h O�  `  j  P�  T   TR  I �  d�A     7       ��  R`  �h O�  �  �  P�  !  S�R  �v   T�  6 �  @�A     $       ��  R�  �hR�  �  O  �    P�  
  Su  X+Y   Q�   7  &�A            �H  R�  �hR  �` O�  V  `  P�     QH   �  �A            ��  RV  �h O  �   �  P�  _  W�[  �-�   T�  o �  ��A     {       ��  R�  �XR�  �P O�  �  �  P�  �   Q�  F   n�A     %       �(  R�  �h O�  6  @  P�  �   Q(  f c  \�A            �l  R6  �h X�  �  N�A            ��  Y�  6  �h ZY  O�  �  �  B�  �  CY   P�  6  [�    T�  �   ��A     P       �   B�    CY   R�  �X\  ]�   R�  �P F  U�  ��A            �V  T Y  Vx .   �h X  u  ��A            ��  Y�  �  �h OE  �  �  B�  �  C�   P�  �  [�    T�  < �  ��A     P       �  B�  �  C�   R�  �X\�  ]�   R�  �P F2  U  ��A            �:  T �  Vx .  �h XA  Y  v�A            �f  Y�  �  �h On  y  �  =�  P�  �  ^ Tf  � �  J�A     ,       ��  =�  Ry  �h^ _P  �  ��A     R       �  Y�  w  �h`WS   (�  �``p  8)   �Xa  +  	�|B      L�  +  M:      b-  R  ��A     Q       ��  Y�  w  �X`p ()   �Pcptr Q  �ha  �  	�|B      L�  �  M:    �  dz �   ��A     �       �  e� (3  	�C     e� "	  	�C     e� '�  	�C      F|  Oe  "  ,  P�     Q  - O  4�A            �X  R"  �h f.  ^  Q  �(@            ��  `@  #)   �hVp /Q  �` �  i	  J  g�  �  "g�  �  " �   �D  �  � �  �1          �@ �  �5   �  �  �  �  V   �  V   �  �  int p   �  3  J   frg S  �  �   o   �   	�   �   
.  7Y   �  !  �  {,  �  |p   �  ~;  
    t   �       t  p     )    A  G  z   )  a  \  g  z  �    )  �  |  �  z  �   )  �  �  �  z  �   )  *�  �  �  z  �   )  0x  �  �  z  �   (  8  �    z  p    �  =O  �     +  z  �    c  Q�  �  D  J  �   c  T�  �  c  i  z   m  X�  �  �  �  �   R  \+  �  �  �  �   R  `[  �  �  �  z   !  d�  �  �  �  z   f  �  �  �  z   �  ��    �  ��  T p    �   p  J�  
.  �  7  �  �   e  S  �  ^  �  E  6  std  �  �  	�  q  	�  �  	�  �  	�  �  �  �  
   �  	q  �  �  �  
   T �  v �    �  �  	q  q  	�  �  	�  �  	,    =  C     �  	�    [  a     T �  v �   �  2  	��  q  	��  T p   �   �    �  	��  q  	��  T p   �   �    !6  	��  �  !6  	�?  �   l  �  "  �  �  "F    q  #�   	�|B     #�   	��B      
r  �z  
i    F�  
i   �:  
V    $�   �   %w   &p   %!  &�   %�   !  %p   p   ':  �  '�  �  �  �  |  �  #<  	�|B     (r  �  )D  +�  H  )�  ,�  M  *\z  p   I  +�   +σ  +�=  +�^  +mS   �1  �  ,it S   ,end S  -c  7�  �  �  �  �   C e   �  �  ,it �   ,end �  -c  օ  �  �  �  �   C V    fT  -  ,it �   ,end �  -c  �3  �    %  �   C �   � q_  .w�  r��    N  �  �  �    f�  #�   � 	j  l" 	  l" � �  �  �   �z  �  �  �  �  �   �:  F  �  �  �  �   �  �   �  �  �  �   /�z  5p    /�:  6_   '" 9	M  .�  <�   <  �    	    0� 
�  0w �    � �  ,it '   ,end S  -c  � �  �  �  -   C ^   � 	  ,it �   ,end �  -c  ! �  �  �  !   C ]    � N	  ,it �   ,end �  -c  1 �  @	  F	  8   C �   1^ Q�
  �
  2�
   3�  ~! v	  �	  L  W   3�  - �	  �	  L  ]   �  R �	  �	  L   4W UM   N	  �	  �	  L  �  c  i   4� q�   N	  
  !
  L  �  o  i   4^ ��   N	  A
  V
  L  �  u  i   4v  �   N	  v
  �
  L    {  i   5�  D N	  �
  �
  L  p    G k   N	  1� ,�
  x  3� � �
  �
  �  �   6� �   7� ,  �
  
    �  p    w�  0K�    -  =  �  ^  �   � D4"   U  e  �  ^  �   � WY! y  �  �  �  �   4W Z�   �
  �  �  �  �  c  i   4� ]w   �
  �  �  �  �  o  i   4^ `�   �
    (  �  �  u  i   4v  cQ   �
  H  ]  �    {  i   � g�  w j�  	 �
  8	 �5! �  8� � �   I  �  V   ]   �  �  �  �  �  -  �  %_  x  �  r %I    �  %j  %�  "� M  "� [  �  ^  j  -  	  8  9&  r  N	  L  &N	  %�
  %�  %=  %�  )   %	  �
  �  %x  :p   �  ; �  <Y�  �  %�  =�  =�  >(	  �  j�A            ��  ?�  >  �h >�    J�A            �  ?�  3  �h >  4  *�A            �A  ?�  �  �h >�  `  
�A            �m  ?�  �  �h >o  �  ��A            ��  ?�  �  �h @V
  �  ��A     X      �h  ?�  R  ��A  �3  ��A�1  �R{  ��Bst �i  ��C  x  	�}B     D� �j  �PEes �  �OF�A     �       Ecp �_  �HEcps ��  ��Gp1  Ee �  �l   He  x  I5    h  @!
  �  ~�A           �&  ?�  R  ��A  �@�  ��Bn �Nu  ��Bst �i  ��C  6  	 ~B     D� �I  �PEds �x  �HF��A     !       Ee �  �l  He  6  I5    &  @�	  Z  6�A     G      ��  ?�  R  ��A  q9�  ��A�1  qRo  ��Bst ri  ��C  x  	P~B     D� uI  �PEds vx  �HF��A     $       Ee z  �l  @�	    ��A     K      ��  ?�  R  ��A  U.�  ��A�1  UIc  ��Bst Vi  ��C  �  	b~B     D� YI  �@Eds Zx  ��F��A     $       Ee ^  �\  He  �  I5    �  J�
  Q�  �  K�  R  K  w    L�  �! �  ��A     +       ��  M�  �h L�  S   ��A     -       �#  M�  �h N�	  1  ;  K�  R   L#  � ^  X�A     7       �g  M1  �h O}  ��A            ��  D� �-  	�C      P:  ��  ��A            ��  ?�  �  �hBnc �/�  �dBwc �>�  �X Q�  ?�A     g       �  D �5N	  	�C      N�
  $   7  K�  �  K  w    L  �! Z  �A     +       �c  M$  �h R  / �  ��A            ��  M$  �h @(  �  ��A     |       ��  ?�  �  �XA  <.  �PA�1  <O	  �HEwc =	V   �lC  
  	~B      He  
  I5   
 �  @�  .  R�A     �      �k  ?�  �  �XBseq 4�  �PEuc 	<   �oC  
  	@~B      S�  V   �  @�A            ��  ?�  �  �h S�  p   �  0�A            ��  ?�  �  �h N�  �  �  K�  �   R�  �    �A             �  M�  �h Ne    ?  K�  �  T�  W�  T� W8�   R  � b  ��A     =       �{  M  �hM&  �dM2  �` i	  J   (   �I  �  �# �  �2          }G �  �  �<   �  �  E  6  �  �  �  p   �  p   �  �  int �   3  	d   std    �  
  	q  
!  �  
  
�  
�  �   �   �   /   
�  
q  �   	    /   T   v     �   �  
�  	q  
!  �  
  
�  
,  >  b  h  >   
�  
�  >  �  �  >   T   v    $  2  
��  	q  
�!  T �   �  �	    �  
��  	q  
�!  T �   �  �	    6  
��  !  6  
�?  !   l      �     F  1  �  frg 	�	  �  R  o   [  �   �  .  7�	   %  �   ,�  �   �  hex  �  �  �  {  �  |�   �  ~;  �  �  �	    �    �  �	  �     !)      #  �	   !)  a  8  C  �	  "R   !)  �  X  c  �	  "�	   !)  �  x  �  �	  "�	   !)  *�  �  �  �	  "�	   !)  0x  �  �  �	  "�	   !(  8  �  �  �	  �    #�  =O  �	  �    �	  "�   #c  Q�       &  �	   #c  T�    ?  E  �	   #m  X�    ^  d  �	   #R  \+  �	  }  �  �	   #R  `[  �	  �  �  �	   #!  d�  
  �  �  �	   f  �  �  �  �	   $�  ��   $�  �  T �    �  �*  2�  �*  3Z(  #  )  
   
	   6C    A  L  
  "�   $   <�   $�  =�   $�)  >�  $�   ?  $�'  @  $�#  A  $<  B  $�  C  %�*  E&  �  �  
  �    &�*  >  �  
  "<      'p  J�  (�-  N�!  <  P �  T p   "�  "p   "  "�   "�   "�   "�	   (�'  x<+  y  P �  T p   "�  "p   "�   "�   "�   "�	   )�  ��+  T p   F �  "p   "  "�    �  
�  �  �  �  �  �)  E#  �  �  �  "S
   q,  �	a  q,  �#      �  "�   *q,  _   *  5  �  "�   +�  	~-  �  M  X  �  "�   p,  �*  l  w  �  �    
)  "	�  �  �  �  �  "�   �$  'a&  �  �  �  "�	   �$  1�  �  �  �  "�	   ,�)  >�   ,ܨ  ?�  ,7&  @
0   �,)  A  �
�   	  �  /  :  T p   �  "p    -c.  	�*  �  U  T �	  �  "�	    �  
�  H`*  �  ~  �  �   !�#  M�"  �  �  �  "�	   ,.  QS
   .U(  S
  /].  <   � 0�  1�  
i  �	  �  T �   "�	  "�	   (`)  �@%  	  F �  "p   "  "�   (`)  �O'  ?	  F �  "�	  "  "�   2N#  3�  i	  T p   F �  "�  "�   3�  3�%  T �	  F �  "  "�    4`  	p~B     �	  �	  �  �	  4y  	��B     �  �	  �  �	  5�   6�   5�  6�  5�  �  5�   �     
  7:  �  7�  �  �  |  4�  	�~B     'r  �  <&  �
  8<&  
9(  u
  {
  �    �  '%  �
  �  "�	    9D  +�  �  9�  ,�  �  f�  #�   �$ �  
�$ =$   �
  �
  �   
�" �"       �  "�
   
d$ m$   )  4  �  "�
   
�$ �#   L  W  �  "�
   
�" �#   o  z  �  "�
   
�$ �$   �  �  �  "�
   
�" q#   �  �  �  "�
   
�" y"   �  �  �  "�
   
�$ �"   �    �  "�
   
�$ �"     )  �  "�
   
�# #   A  L  �  "�
   
# 7#   d  o  �  "�
   
$ �# �
  �  �  �  "�
   -�$  $ �
  �  �  "�
    :�$ �
T# �   S
  �
  �  �  �  �  �  5a  5�  ;�	    <<    =�  =  >�  /  6@     �       �I  ?�  �  �h@s '�	  �d A�  95@     (       ��  T �   @a �	  �h@b #�	  �` B�  �3@     �      ��  P �  T p   C��  N�  ��C�   N$p   ��C�'  N1  ��C3(  N?�   ��Ch  O�   ��C�)  O�   ��C�D  O#�	  ��D4  P�	  �XDݨ  S�  ��Ek T�   ��F�4@     E       o  Ei a�   �l F�4@     -       �  Ei d�   �h G5@     0       Ei f�   �d  ;�	  �  <<    B<  �1@     U       �T  P �  T p   C��  x�  �hC�   x!p   �dC3(  x-�   �`Ch  x8�   �\C�)  y�   �XC�D  y�	  �THIi$  {	p     By  �0@     �       ��  T p   F �  C�  �p   �l@fo �/  �`C��  �6�  �X >�  �  �/@     �       ��  ?�  �  �h@str 1�	  �` B�  ,.@     J       �7  F �  C�  �!p   �L@fo �8  �@C��  �?�  �� B	  .@     *       ��  F �  C�  � �	  �h@fo �7  �`C��  �>�  �X 5w   B?	  %-@     C       ��  T p   F �  J�  3�  �HJ��  3!�  �@ >�  �  h-@     &       �  ?�  �  �hC/&  M�	  �` 5�	  Bi	  �,@     E       �b  T �	  F �  J�  3  �HJ��  3!�  �@ K�  p  �  L�  �  M�)  �   Nb  �  �  �,@     4       ��  Op  �hOy  �` K�  �  �  L�  �	  L  �    N�  6.  �  �+@            �  O�  �h K�      L�  �	   N  9*  B  �+@            �K  O  �h >  q  ^+@     (       ��  T p   ?�  �  �hC�  p   �d >w  �  �+@     ,       ��  ?�  �  �hP�  �  >:  �  4+@     )       �  T �	  ?�  �  �hC�  �	  �` KX    $  L�  �  L  �    N  *$  G  (+@            �P  O  �h >f  o  �*@     )       �|  ?�  �  �` K�  �  �  L�  �	  M�  *�	   Q|  %'  �  �)@     V       ��  O�  �hO�  �` K�  �  �  L�  �	  L  �    Q�  g    �)@            �!  O�  �h K  /  9  L�  �	   Q!    \  �)@     #       �e  O/  �h A�  ��A            ��  D�$ ��
  	�C      R�  ��  8�A     �       ��  ?�  �  ��~@c �'�
  ��~ Ro  v�  ��A     �       �  ?�  �  ��~@c v'�
  ��~ RL  m5  ��A     �       �Q  ?�  �  ��~@c m"�
  ��~ R)  ds  �A     �       ��  ?�  �  ��~@c d"�
  ��~ R  [�  R�A     �       ��  ?�  �  ��~@c ["�
  ��~ R�  R�  t�A     �       �  ?�  �  ��~@c R"�
  ��~ R�  I-  ��A     �       �I  ?�  �  ��~@c I"�
  ��~ R�  @k  ��A     �       ��  ?�  �  ��~@c @"�
  ��~ Rz  1�  ��A           ��  ?�  �  ��~@c 1"�
  ��~ RW  (�  ��A     �       �  ?�  �  ��~@c ("�
  ��~ R4  %   �A     �       �A  ?�  �  ��~@c #�
  ��~ R  c  f�A     �       �  ?�  �  ��~@c "�
  ��~ R�
  �  ��A     �       ��  ?�  �  ��~@c "�
  ��~ S�
  �  ��A            ��  ?�  �  �h T�  2�    L�  
  L  �    Q�  .  3  �)@            �<  O�  �h 5�  T�  2S  b  L�  
  "<   QB  �  �   )@     �       ��  OS  �hO\  �` K  �  �  L�  
   Q�  K  �  �(@     \       ��  O�  �h U.  ^  D  �(@            �  C@  #0   �h@p /D  �` i	  J   %   O  �  % �  ��A     A       .T �  �  �  E  6  std  �  �  �   q  �  �  �  �  �  s   �   �   	�   �  q  s   �   �   	�   
T �  v �    Y   �  B  q  �  �  �  �  ,  �       	�   �  �  �   ,  2  	�   
T �  v �   �   2  �t  q  ��  
T   �  D    �  ��  q  ��  
T   �  J    6  ��  �  6  �?  �   l  �    f   �   F  �   B  �  �  �  �  �  int   frg 	�  �  +  o   4  �   `  .  7   �  �  �  {�  �  |  �  ~;  �  �  	,   �    �  	,  	    )    �  �  	2   )  a  �  �  	2  +   )  �      	2  8   )  �  ,  7  	2  >   )  *�  L  W  	2  D   )  0x  l  w  	2  J   (  8  �  �  	2  	   �  =O  P  �  �  	2  `   c  Q�  �  �  �  	V   c  T�  �  �  �  	2   m  X�  �      	V   R  \+  8  1  7  	V   R  `[  \  P  V  	2   !  d�  b  o  u  	2   f  �  �  �  	2    �  �m    �  ��  
T    `  !p  J�  
�  �  �  �  i  �)  E#  �    	d  �   "q,  �  H`*    !  '  	d   �#  M�"  <  G  	d     #.  Q�   $U(  �  %].  4   � &�  �)  E�&  �  �  	|  �   "q,  �  H�#  �  �  �  	|   �#  M�  �  �  	|     #.  Q�   $U(  �  %].  4   �  '9  	�B         �    'R  	��B     m  `  (  )  (�  )`  (`  �  (    *:  T  *�  �  �  |  '�  	��B     +r  N  <&  �  ,<&  
9(  �  �  	N   �  '%  �  	N      P(  -  ,P(  6"      	Y   �  �'  !  	Y      -D  +�  �  -�  ,�  i   �  N  �  Y  �  .-  $	�C     i  .=  	%	�C     /�  /�  0  �  �A     !       ��  1�  _  �h2/&  )  �` 0�  �  ��A            �  1�  T  �h2/&  (  �` i	  J   �   R  �  �% �  �4          jU �  �  �<   �  �  E  6  �  b   �  �  �  |   �  �  �  J  �   int �   �% )   �  �<   4  	�   �   �  	�   ,  	V   3  	p     	4�   std  z  �  
  	q  
�  �  
z  
�  
�  '  K  Q  �   
�  
q  '  i  o  �   T z  v z      �  
�  	q  
�  �  
z  
�  
,  �  �  �  �   
�  
�  �  �  �  �   T z  v z   �  2  
�(  	q  
��  T �   �  L
    �  
�U  	q  
��  T �   �  R
    6  
��  �  6  
�?  �   l  z        F  �  �  �  frg 	�	  �  �  o   �  �   �  .  7

   %  �   ,  �   �  hex  �  b  �  {m  �  |�   �  ~;  K  Q  *
    �    a  *
  �     !)    �  �  5
   !)  a  �  �  5
  "�   !)  �  �  �  5
  "@
   !)  �  �  �  5
  "F
   !)  *�  �    5
  "L
   !)  0x    (  5
  "R
   !(  8  =  H  5
  �    #�  =O  X
  a  l  5
  "   #c  Q�  z  �  �  ^
   #c  T�  z  �  �  5
   #m  X�  z  �  �  ^
   #R  \+  @
  �  �  ^
   #R  `[  d
      5
   #!  d�  j
     &  5
   f  �  :  @  5
   $�  �   $�  �z  T �      �*  2N  �*  3Z(  �  �  p
   
	   6C  g  �  �  p
  "�   $   <�   $�  =�   $�)  >  $�   ?z  $�'  @z  $�#  Az  $<  Bz  $�  Cz  %�*  E&  *  5  p
  �    &�*  >  B  p
  "�    g  'p  J	  (' Nw( �  P T  T <   "�  "<   "z  "�   "�   "�   "
   (�& x2% �  P T  T <   "�  "<   "�   "�   "�   "
   )( ��% T <   F T  "<   "g  "�    �  
	  �    *�  �  0	  �)  E�&  I  T  �  "�
   q,  �	�  q,  �&  u  �  �  "�   +q,  N"  �  �  �  "�   ,�  	�   �  �  �  �  "�   p,  �"  �  �  �  �    
)  "	�(  �  �    �  "	   �$  'r    #  �  "
   �$  1�,  7  B  �  "
   -�)  >�   -ܨ  ?*  -7&  @
0   �-)  Az  �
�3  	_' �  �  �  T �  �  "�   .c.  	�$  �  �  T 
  �  "
    T  
�  H�#  T  �  �  �   !�#  M�  	  	  �  "
   -.  Q�
   /U(  �
  0].  <   � 1�  
i  @
  V	  T �   "@
  "@
   (f  �Q& }	  F T  "�
  "g  "�   (f  ��  �	  F T  "
  "g  "�   2�' 3�( �	  T �  F T  "�  "�   3   3n$  T 
  F T  "�  "�    4�  	 �B     
  
  �  
  4�  	��B       *
    5
  5�   6�   5b  6  5  b  5�   �   g  p
  7:    7�  5  �  |  �
  84  	�B     'r  $  P(    9P(  6"  �
  �
  $    �  �'  �
  $  "
    :D  +�  #  :�  ,�  (   �
  ;
  :  <<    =�  >,% ?i3  �   @�~  f  l  �   @|  |  �  �   $H& !
�    $�1  $�     A	:  BH  ?  �  (  �  T  �  5�  5T  BU  Bg  C    b5@     �       �  D�  �  �hEs '
  �d F0	  95@     (       �X  T �   Ea @
  �hEb #@
  �` G_  c�A     �      ��  P T  T <   H��  N�  ��H�   N$<   ��H�'  N1z  ��H3(  N?�   ��Hh  O�   ��H�)  O�   ��H�D  O#
  ��~I4  P
  �XIݨ  S�  ��Jk T�   ��K\�A     E       A  Ji a�   �l K��A     -       d  Ji d�   �h L��A     0       Ji f�   �d  ;
  �  <<    G�  �A     W       �&  P T  T <   H��  x�  �hH�   x!<   �`H3(  x-�   �\Hh  x8�   �XH�)  y�   �TH�D  y
  �PMNi$  {	<     G�  m�A     �       �}  T <   F T  H�  �<   �hEfo �/g  �`H��  �6�  �X C#  �  v.@     �       ��  D�  �  �hEstr 1
  �` GV	  ��A     }       �  F T  H�  � �
  ��Efo �7g  ��H��  �>�  �� G}	  �-@     *       �[  F T  H�  � 
  �hEfo �7g  �`H��  �>�  �X C�  z  �,@     &       ��  D�  �  �hH/&  M
  �` 5�  G�	  ��A     E       ��  T �  F T  O�  3�  �HO��  3!�  �@ 5

  G�	  �+@     E       �6  T 
  F T  O�  3�  �HO��  3!�  �@ Pa  D  Z  Q�  �  R�)  �   S6  �  }  �+@     4       ��  TD  �hTM  �` PQ  �  �  Q�  0
  Q  �    S�  6.  �  �+@            ��  T�  �h P7  �  �  Q�  0
   S�  9*    �+@            �  T�  �h C�  >  �*@     ,       �S  D�  �  �hU	  �  Cz  y  ��A     )       ��  T �  D�  �  �hH�  �  �` C�  �  �*@     )       ��  T 
  D�  �  �hH�  
  �` P�  �  �  Q�  �  Q  �    S�  v(    t*@            �$  T�  �h C�  C  J*@     )       �P  D�  �  �` P�  ^  t  Q�  ;
  R�  *L
   VP  %'  �  �)@     V       ��  T^  �hTg  �` P(  �  �  Q�  ;
  Q  �    V�  g  �  �)@            ��  T�  �h Pm      Q�  ;
   V�    0  �)@     #       �9  T  �h W�' <1T�A     .       �v  Eptr <Nv  �XIHx  =�  �h �   X�' 00�   
�A     J       ��  Eptr 0Mv  �XIHx  1�  �h Yd( +1��A     f       �Zl  �  ��A            �  D�  �  �h CV  "  @�A     J       �<  D�  �  �XJv �   �l C�  [  M@     6       ��  D�  v
  �`Ec 63�  �\I�>  7g  �h [  2�  �  Q�  v
  Q  �    V�  .  �  �)@            ��  T�  �h 5N  [5  2�  �  Q�  v
  "�   V�  �     )@     �       �/  T�  �hT�  �` Pt  =  G  Q�  v
   V/  K  j  �(@     \       �s  T=  �h \.  ^  �  �(@            ��  H@  #0   �hEp /�  �` i	  J   %U   :;9I  $ >  $ >  & I  :;9   :;9I8   :;9I8  	   
 I  :;9n  I  ! I/  ;   .?n4<d   I4  4 :;9I?<   :;9I  I   I    :;9   :;9I8   :;9I8  :;9   :;9I  >I:;9  (   (    <  :;9    :;9I8  !4 :;9I?  "4 :;9I?  #:;9  $.?:;9n2<d  %.?:;9nI2<d  & :;9I82  ' :;9I82  (/ I  ).?n42<d  *4 I?4<  +. 4@�B  ,.Gd   - I4  ..1nd@�B  / 1  0.4@�B  1 :;9I  2.Gd@�B  3 I4  4 :;9I  54 :;9I  6  74 :;9I  8.Gd@�B  9.G:;9d   :.1nd@�B  ;  <.?:;9I@�B  =4 :;9I  >4 :;9I  ?.?:;9n@�B  @.?:;9nI@�B  A I   %  . @   %  $ >   :;9I  $ >  .?:;9'@�B   :;9I   %  $ >   :;9I  ;   $ >  & I     9:;9  	4 :;9nI?<  
.?:;9nI<   I  . ?:;9nI<  . ?:;9n�<  .?:;9n<  .?:;9n�<  9:;  :;9   :;9I?<l   .?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I  9:;9   :;9  4 :;9I<l  9:;9   4 :;9I<l  !:;9  ":;9  # :;9I  $.?:;9n<d  %.?:;9n<d  &.?:;9n2<d  '.?:;9nI2<d  ( :;9I8  )9 :;9  * <  +4 G  , I  -B I  .4 nG  /4 G  0. ?:;9n@�B  1. ?:;9I@�B  2.G@�B  3 :;9I  4.G@�B  54 :;9I  64 :;9I  7. G@�B  8 :;9I  94 I4  :I  ;! I/   %U  $ >   :;9I  ;   9:;  :;9   :;9I?<l   .?:;9nI<d  	 I4  
/ I  0 I  & I  ��  / I  4 :;9nI?<l   4 nG   I     $ >  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  *.?:;9n<�d  +.?:;9nI<�d  , :;9I82  -.?:;9nI<d  ./ I  /0 I  0.?:;9nI<  1.?:;9n<  2.?:;9n<  34 G  4 I  5B I  64 nG  7.?:;9n<�d  84 :;9nI?<  9I  :! I/  ;4 G  <.Gd@�B  = I4  > :;9I  ?.G@�B  @.G@�B  A :;9I  B4 :;9I  C4 :;9I  D  E  F  G4 :;9I  H :;9I  I.Gd   J I4  K :;9I  L.1nd@�B  M 1  N I  O.1nd@�B  P.?:;9@�B  Q.G:;9d   R.?:;9nI@�B   %   :;9I  $ >  .?:;9I@�B   :;9I  4 :;9I     I  	& I  
 :;9I  4 :;9I       7 I  &   $ >    I   I4   :;9I  4 :;9I  / I  & I   :;9I   I4  	.Gd@�B  
4 :;9I  4 :;9I   :;9I8   I   I   :;9I  4 :;9I   1    .G@�B  .?:;9n2<d  4 I4  :;9   I4  .?:;9n<d  .?:;9I@�B  .?:;9nI<   :;9I  $ >  .?:;9n2<d  I  .Gd    .?:;9nI<d  !! I/  " :;9I  #  $.?:;9I@�B  %(   &.?:;9nI2<d  '.?:;9n<d  ( :;9  )4 nG  *.1nd@�B  + :;9I  ,.?:;9n<�d  -.?:;9nI<�d  ..G@�B  / :;9I8  0.?:;9nI2<d  1 :;9I?<l   2.Gd@�B  3 :;9I82  4/ I  5.1nd@�B  64 G  7m>I:;9  8.?:;9n<  9.?:;9nI2<  : :;9I82  ;0 I  <4 G  =7 I  > I  ?.?:;9�@�B  @4 :;9I?<  A:;9n  B :;9  C.?:;9n<d  D9:;9  E9  F: :;9  G I8  H :;9I?<l   I.?:;9nI<d  J :;9I  KB I  L
 :;9  MU  N.?:;9@�B  O :;9I?<l   P :;9I?<l   Q4 :;9I<l  R(   S:;9  T.?:;9nI<d  U <  V4 :;9I<l  W.?:;9nI<  X.?:;9nI2<  Y.?:;9n2<�d  Z.?:;9n<  [0 I  \��  ]/ I  ^4 :;9nI?<l   _4 nG  `4 :;9nI?<  a.?:;9nI<cd  b4 nG  c.G:;9d   d IJ  e%U  f$ >  g   h9:;9  i:;9  j :;9I?<l   k :;9I82  l :;9I82  m9:;9  n4 :;9I<l  o:;9  p :;9I  q.?n4<d  r.?n4<d  s.?:;9n<  t0 I  u4 :;9I<
l  v:;9  w:;9  x.?:;9nI<  y:;9  z.?:;9nI2<�d  { :;9I?<
l   | :;9I?<l   }:;9  ~ :;9I8  4 Gn  �! I/  �;   �9:;  �&   �.?:;9n<�d  �.?:;9nI<d  �4 :;9I<  �4 :;9I?  �4 nG  �. 4@�B  �.4@�B  �  �4 :;9I  �.?:;9@�B  �.?:;9I@�B  �.?:;9I@�B  �I  �   �. ?:;9I@�B  �.?:;9nI@�B  �4 :;9Il   %U   :;9I  $ >  & I   :;9I  ;   $ >  :;9  	 :;9I8  
9:;   :;9I?<l   .?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I   .?:;9n<d  !.?:;9n<d  ".?:;9n2<d  # I  $.?:;9nI2<d  %.?n4<d  &9 :;9  '/ I  (.?:;9n<�d  ).?:;9nI<�d  * :;9I82  +.?:;9nI<d  ,0 I  - <  ..?:;9n<  /.?:;9n<  04 G  1 I  2B I  34 nG  49:;9  5.?:;9n<�d  64 :;9nI?<  7 :;9I8  8.?:;9nI<cd  9<  :.?:;9nI<  ;9  <>I:;9  =: :;9  >I  ?! I/  @4 G  A.Gd@�B  B I4  C :;9I  D.G@�B  E :;9I  F :;9I  G.Gd   H I4  I :;9I  J.1nd@�B  K 1  L I  M.Gd@�B  N  O4 :;9I  P :;9I  Q.1nd@�B  R.?:;9I@�B  S4 I4  T :;9I  U4 :;9I  V.?:;9I@�B  W.G@�B  X4 :;9I  Y.G:;9d     I   I4   :;9I  / I   I4  & I   :;9I8  .Gd@�B  	4 :;9I  
 I  .?:;9nI2<d   I   1  .?:;9n2<d  4 :;9I  .G@�B  4 :;9I   :;9I  4 :;9I   I4  :;9   :;9I  .?:;9n<d    .Gd   .?:;9nI<  $ >  .?:;9n2<d  .Gd@�B   :;9I  .?:;9nI<d   .?:;9n<d  ! :;9  ".1nd@�B  #  $ :;9I  %I  &! I/  '.G@�B  (.1nd@�B  ).?:;9n<�d  *.?:;9nI<�d  +/ I  , :;9I  - :;9I?<l   .4 nG  /(   0.?:;9nI2<d  14 :;9I?<  2 :;9I82  3 :;9I82  44 I4  5.?:;9n<  64 G  7B I  8.?:;9nI2<  90 I  ::;9  ;.?:;9n<  <4 G  =.?:;9I@�B  > :;9  ?9:;9  @9  A: :;9  Bm>I:;9  C I8  D :;9I?<l   E.?:;9nI<d  F.?:;9n<d  G.?:;9nI2<d  H :;9I  I0 I  J��  K/ I  L4 :;9nI?<l   M.?:;9nI<  N4 :;9I<l  O(   P.?:;9nI2<  Q:;9  R.?:;9nI<d  S.?:;9n2<�d  T4 :;9I<l  U4 nG  V4 :;9nI?<  W.:;9<  X4 nG  Y  Z :;9I  [ :;9I  \.G:;9d   ] IJ  ^%U  _$ >  `   a;   b9:;  c9:;9  d4 :;9I<
l  e:;9  f.?:;9nI<  g:;9  h.?:;9nI2<�d  i :;9I?<
l   j :;9I?<l   k:;9  l :;9I8  m9:;9  n4 :;9I<l  o:;9  p :;9I  q.?n4<d  r.?n4<d  s.?:;9n<  t0 I  u <  v.?:;9nI<d  w&   x.?:;9n<�d  y4 :;9I<  z. :;9<  {. :;9I<  |.:;9I<  }4 :;9I?  ~4 I?4<  4 nG  �4 :;9I  �4 :;9I  �1  �4 1  �1  �4 1  � I  �.?:;9nI@�B   %  4 :;9I?  $ >   I  $ >    I   I4  / I   I4   :;9I  .Gd@�B  & I  4 :;9I  	 :;9I  
4 :;9I   I   :;9I8   I   1  .?:;9nI<d     I4  :;9   :;9I  .?:;9n<d  4 :;9I  .G@�B  4 :;9I    .?:;9n2<d   :;9I  .Gd   .?:;9nI<  / I   :;9I82  .?:;9n2<d   .1nd@�B  !$ >  ".G@�B  #(   $.?:;9n<d  %I  &! I/  '.?:;9nI2<d  (.?:;9nI2<d  ) :;9  * :;9I  +4 I4  ,.1nd@�B  -.?:;9I@�B  ./ I  /.?:;9n<�d  0.?:;9nI<�d  1.Gd@�B  24 G  3 :;9I  4 :;9I?<l   54 nG  6.?:;9n<  74 :;9I?<  8B I  94 G  :4 1  ;4 1  <m>I:;9  =0 I  > I8  ?.?:;9nILM2<d  @.?:;9nILM2<d  A.:;9I<  B :;9  C.?:;9n<d  D9:;9  E9  F.?:;9nI2<  G :;9I82  H.?:;9nI<d  I.?:;9n<  J��  K4 :;9I<  L I  M.?:;9nI<d  N4 :;9I<l  O: :;9  P:;9  Q :;9I?<l   R I82  S :;9I2  T :;9I  U4 G:;9  V.G:;9d   W  X4 I4  Y1  Z IJ  [0 I  \��  ]9 :;9  ^4 :;9nI?<l   _4 :;9I<l  `(   a:;9  b0 I  c.?:;9nI<  d.?:;9nI2<  e:;9  f.?:;9nI<  g.?:;9n2<�d  h.?:;9nI2<d  i.?:;9nI<d  j4 nG  k.?:;9n<�d  l4 :;9nI?<  m:;9  n.?n4<�d  o4 nG  p��:;9  q.?:;9@�B  r.4<d  s.4d@�B  t.I4d@�B  u.4@�B  v4 :;9I  w1  x%U  y$ >  z   {;   |9:;  }9:;9  ~9:;9  4 :;9I<l  �:;9  � :;9I  �.?n4<d  �.?n4<d  �.?:;9n<  �4 :;9I<
l  �:;9  �.?:;9nI2<�d  � :;9I?<
l   � :;9I?<l   �:;9  � :;9I8  �:;9  � I84  �.?:;9nL<d  �.?:;9nILM<d  �4 :;9I<  �.?:;9nI<d  �.?:;9nILM<d  � :;9I82  �.?nL4<d  �.:;9<d  �.:;9<d  �: :;9  �4 nG  �  �I  �   � I  �4 I?4<  �. 4@�B  �.4@�B  �.1d@�B  �1  �.1d@�B  � :;9I  � :;9I  �4 :;9I  �.?:;9nI@�B    I   :;9I   I4  / I   :;9I  4 :;9I  4 :;9I  4 :;9I  	 I4  
& I  4 I4     I  .G@�B     :;9I  4 :;9I  .Gd@�B  .?:;9I@�B   :;9I8   I   1  / I   I  .?:;9n<d  .?:;9n<   :;9I  .?n4<d  :;9   I4  .?:;9n2<d   .?:;9nI2<d  ! :;9I8  ".Gd   #U  $ :;9I  %(   & :;9I  '.?:;9nI<  (.?:;9n<  )B I  *.1nd@�B  +$ >  ,.?:;9n2<d  -I  ..?:;9nI<d  / :;9I82  0   1! I/  2.?:;9n<d  3  44 :;9I  5 :;9  6.G@�B  7.1nd@�B  8.Gd@�B  9.?n4<�d  :.?n4d@�B  ;.?n4d@�B  <:;9  = :;9I?<l   >.?:;9I@�B  ?.?:;9n<�d  @.?:;9nI<�d  A :;9I82  B4 nG  C.?:;9nI2<d  D4 G  E4 :;9I?<  F7 I  G :;9I  HU  I:;9  J :;I8  K :;9I  L��  M/ I  N4 :;9nI?<l   Om>I:;9  P.?:;9nI2<  Q0 I  R:;9  S4 nG  T.?:;9I@�B  U.4<d  V.42<d  W.?:;9nI<  X :;9  Y9:;9  Z9  [: :;9  \ I8  ] :;9I?<l   ^.?:;9nI<d  _.?:;9n<d  `4 G  a0 I  b4 :;9I<l  c(   d.?:;9nI2<  e.?:;9nI<d  f.?:;9n2<�d  g4 :;9I<l  h <  i4 :;9nI?<  j4 nG  k.:;9I@�B  l.?:;9@�B  m.?:;9@�B  n. ?:;9I@�B  o.:;9Id@�B  p.:;9I2d@�B  q :;9I  r.G:;9d   s IJ  t%U  u$ >  v I  w:;  x   y;   z9:;  {9:;9  |4 :;9I<
l  }.?:;9nI<  ~:;9  .?:;9nI2<�d  � :;9I?<
l   � :;9I?<l   �:;9  �9:;9  �4 :;9I<l  �:;9  � :;9I  �.?n4<d  �.?:;9n<  �0 I  �9 :;9  �.?:;9nI<d  �&   �.?:;9n<�d  �>I:;9  �4 nG  �! I/  �:;9  �:;9  �.:;9@�B  �.?:;9@�B  �.?:;9nI@�B   %   :;9I  $ >  4 :;9I?<  $ >   I  7 I  & I  	   
.?:;9I@�B   :;9I   :;9I  4 :;9I  &   .?:;9I@�B   I  4 I4  I  ! I/  .?:;9I@�B   :;9I   :;9I  4 :;9I    .?:;9I@�B  4 :;9I  4 :;9I  .?:;9I@�B   %  $ >   :;9I  $ >  9:;9  .?:;9nI<   I  .?:;9nI<  	 I  
& I  .G@�B   :;9I  4 :;9I   :;9I  4 :;9I     &   .G@�B   %U   :;9I  & I  $ >  ;   9:;  :;9   :;9I?<l   	.?:;9nI<d  
 I4  / I  0 I  .?:;9nI<   I  4 nG   I  $ >  9:;9   :;9  4 :;9I<
l  9:;9  9  4 :;9I<l  : :;9  m>I:;9  (   (   .?:;9n<d  .?:;9n<�d  .?:;9nI<�d   :;9I8   .?:;9nI2<  !.?:;9nI2<  ".?:;9n2<d  #.?:;9n<d  $.?:;9n2<d  %.?:;9nI2<d  & :;9I82  '0 I  (:;9  ) :;9  * I8  +:;9  ,:;9  - <  ..?:;9nI<d  /.?:;9n2<�d  0.?:;9nI2<�d  1.?:;9nI2<d  2 :;9I?<
l   3 :;9I?<l   4 :;9I?<l   5.?:;9nI<d  6/ I  7:;9  8 :;9I8  9�:;9  :�:;9  ;.?:;9nI2<d  < :;9I�8  =��   > :;9I  ?�:;9  @0 I  A�:;9  B��  C/ I  D�:;9  E4 G  F I  G   H :;9I82  I.?:;9nI<d  J.?:;9n<d  K9 :;9  LI  M! I/  N! I/  O.Gd   P I4  Q.1nd@�B  R 1  S :;9I  T.1nd@�B  U.G@�B  V :;9I  W :;9I  X.Gd@�B  Y I4  ZB I  [��:;9  \��:;9  ] 1  ^�� :;9  _.G:9d@�B  ` :;9I  a4 I4  b.G:;9d@�B  c4 :;9I  d.?:;9nI@�B  e4 :;9I  f.?:;9nI@�B  g IJ   %U   :;9I  $ >  & I  $ >  9:;9   :;9  4 :;9I<l  	9:;9  
4 :;9I<l  :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  9 :;9   <   I  ;   9:;  :;9   :;9I?<l   .?:;9nI<d  0 I  ��   / I  !4 :;9nI?<l   "4 nG  #4 G  $   % I  &B I  '4 nG  (9:;9  )4 :;9nI?<  *m>I:;9  +(   , :;9I8  -.?:;9nI<cd  ..?:;9nI<d  / :;9I82  0 :;9I?<l   1:;9  2 I8  3.?n4<d  4.?:;9nILM<d  5.?nL4<d  6 I84  7.?:;9nL<�d  8. ?:;9nI<  94 I?4<  :I  ;   < I  =4 G  >.Gd@�B  ? I4  @.Gd@�B  A :;9I  B :;9I  C4 I4  D4 :;9I  E4 :;9I  F  GU  HI  I! I/  J.G:;9d   K I4  L.1nd@�B  M 1  N.Gd   O.G@�B  P.G:;9d@�B  Q.G@�B  R.1nd@�B  S.GId@�B  T :;9I   %U  $ >   :;9I  ;   & I  $ >  9:;  :;9  	 :;9I?<l   
.?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I     9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  *.?:;9n<�d  +.?:;9nI<�d  , :;9I82  -.?:;9nI<d  ./ I  /0 I  0 <  1.?:;9nI<  2.?:;9n<  3.?:;9n<  44 G  5 I  6B I  74 nG  8.?:;9n<�d  94 :;9nI?<  :. ?:;9nI<  ;I  <! I/  =4 G  >.Gd@�B  ? I4  @ :;9I  A.G@�B  B.G@�B  C :;9I  D4 :;9I  E4 :;9I  F  G  H  I4 :;9I  J :;9I  K.Gd   L I4  M :;9I  N.1nd@�B  O 1  P I  Q.1nd@�B  R.G:;9d@�B  S.G:;9d@�B  T.G:;9d   U.?:;9nI@�B   %  $ >  ;   9:;  :;9   :;9I?<l    :;9I  .?:;9nI<d  	 I4  
/ I  0 I  & I  ��  / I  4 :;9nI?<l   4 nG   I  $ >  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  :;9  :;9   :;9I  .?:;9n<d  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d    :;9I8  !9 :;9  " <  # :;9I82  $/ I  %0 I  &:;9  '4 G  ( I  )B I  *4 nG  +9:;9  ,.?:;9n<�d  -4 :;9nI?<  .4 G:;9  /4 G  0.G:;9d@�B  1 I4  2 :;9I   %U  $ >   :;9I  ;   $ >  & I  9:;  :;9  	 :;9I?<l   
.?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I     9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  * <  +.?:;9n<�d  ,.?:;9nI<�d  - :;9I82  ..?:;9nI<d  // I  00 I  1.?:;9nI<  2.?:;9n<  3.?:;9n<  44 G  5 I  6B I  74 nG  8&   9.?:;9n<�d  :4 :;9nI?<  ;I  <! I/  =9  >:;9  ? :;9I<l   @.:;9<d  A: :;9  B4 G  C.Gd@�B  D I4  E :;9I  F.G@�B  G.G@�B  H :;9I  I4 :;9I  J4 :;9I  K  L  M  N4 :;9I  O :;9I  P.Gd   Q I4  R :;9I  S.1nd@�B  T 1  U I  V.1nd@�B  W.?:;9@�B  X.?:;9I@�B  Y. ?:;9@�B  Z.Gd@�B  [.G:;9d   \.?:;9nI@�B   �   �  �      /home/computerfido/.local/share/lemon/sysroot/usr/include/gfx /home/computerfido/.local/share/lemon/sysroot/usr/include/gfx/window /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/sysroot/usr/include/bits /home/computerfido/.local/share/lemon/sysroot/usr/include/lemon /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include/freetype/config /home/computerfido/.local/share/lemon/sysroot/usr/include/freetype  graphics.h   window.h   main.cpp    list.h   types.h   stdint.h   fb.h   stddef.h   surface.h   types.h   stdio.h   ipc.h   unistd.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h    G 	L@     
�ff!.  tt!.�  	�@     �*  	]@     � 	�'
�' t �	�K t��+��<tKxfftK� ot�>	�'
� t�K
�+�( t ���<tKK +mt%����'��= jt�>Zt<ZK
�H<
t&$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�.K�k�<60B�4�B �8R:�<(.*�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9%$/AtK/Z/��T���.��u	,(!
 <,�, t � / �kv>f�.�f�.��u,fftJg,fftJg�& J( t��& J( t�tf � ��"u%�* f�/f�, �9 fG �; �  .Y �f fM �t �� f� �� �h .���u�<f5 J; t& <K+f �7.Df9�J�trX�t<K'f�J='f�JZ'f�)J<='f�)J<">4<;tf6K�K- g.�� J	�w  �" t f�	u*ut �* f �8 �H fY �J �, .k �{ f_ �� �� f� �� �} .�!u�<f: J@ �( <�t���<K)f�J=)f�JZ)f�+J<=)f�+J<! >3 <: t f8 K � K0���t � t�tJ" X' t <Y$�)t/<�h$�(t�.L�K00tg\+tgZy.mh $X4 tg t f eClRfIfY<<4.t��*[� f�}���<J  	�@     ����  	�@     � 
�u  	@     � �  	*@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K  	X@     �  	z@     )�#���tY��Y����  	H@     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	�@     	 � t J / �    '   �       src/gfx/sse2.asm      	@"@     !>==ALLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""�� �    �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include  syscall.c   types.h   stdint.h    g 	N$@     �� �   !  �      ../sysdeps/lemon/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../options/ansi/include/bits/ansi ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg  lemon.cpp   stddef.h   pid_t.h   time_t.h   types.h   stdint.h   debug.hpp   type_traits   sysdeps.hpp   string.hpp 	  optional.hpp 	  logging.hpp 	  <built-in>    formatting.hpp 	    	�$@     

�(5>� �
�J
�	%tY
vY00
�Y$0
�'>K�2
�	'
u=:0
0	&�
�uY00�Y%0�Y2	KY1L �	   {  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/mlibc  new   formatting.hpp   ensure.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   type_traits   string.hpp   debug.hpp   <built-in>     2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	y&@     &�,�!  # +�� # 6���?&�+�!  # +�� # 6���  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/  	J*@     � �/  	t*@     � 	 	�*@     
�/K 	 	�*@     
�/K 	 	�*@     !�t��K  	�*@     � �/  	(+@     � 	 	4+@     
�/K 	 	^+@     
�/K 	 	�+@     !�t��K  	�+@     � �  	�+@     � �  	�+@     -�1%  	�+@     ��2  	C,@     ��0  	�,@     � �/  	�,@     -�1%  	�,@     ��2  	%-@     ��0  	h-@     � �/  	�-@     �=/  	�-@     �/4  	.@     �=/  	,.@     �/4  	v.@     0��  � .��gt��������y�	X  	G/@     �	/fY%* � � � .�%  	�/@     0��  � .��gt��������y�	X  	�0@     �	/fY%* � � � .�%  	Q1@     � �3  	�1@     � �3  	�1@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�3@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	95@     �� J J . K  	b5@     &  � .��gt���J�����  	6@     &  � .��gt���J����� �   �   �      ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  essential.cpp   stddef.h    . 	�6@     �� � � � W	vKN0�� � � � � < -	vK90��� � � � � < -w �. �5 � � �5 � < -	wK0	�� � ! W	vK �/   �  �      ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  random.hpp   new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   stdlib-stubs.cpp   optional.hpp   strtofp.hpp   logging.hpp   utility.hpp   mutex.hpp   errno.h   types.h   stdint.h   stddef.h   locale_t.h 	  stdlib.h   string.hpp   type_traits   debug.hpp   charcode.hpp   mbstate.h   <built-in>      	fJ@     �  	�J@     
�� � �# u( �+ <4 �9 �< <> �- < .H f �F � . � �"  	4K@     ���� t � �, t/ f1 � X Y �  � X0 .3 f& f J �k t � �, t/ f1 � X Y �& �! X6 .9 f, f J �k�,t.fXY!�X1.4f'f.	�����f=fX=fX=f
>= 2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	M@     5//
�!  	:M@     �F  	�M@     ��  	�M@     �6J7tXK�  	�M@     �Ju ! 	N8@     �X�/�Y/�Y%/�YE/�+t�D/�/K/$�0��M/2	tKt�X	LU0$ ��KtK	K[g f�#X\�	tKt J tK<$�X	xzX	.u� f t .J!S/0YX00��	w�<g��1g	u�<	�g�<g f  fgt  J t
K�gYvg f t X&=	f&/$f	 =�u�XKg�X�� J t X?�# f J4 f, J> f��u! r�<g]>	 g	�gtKu f � JuK]/0Y2-L<�Y0���=>�?X��4>��	g
�	v L)/�K
uu	�K3K ��	YY'/���Y���� ����/�	��
��
�<uA���gg	
g�%�i �	�Y/0v �*�&�	tK �+�'�
tK<X
N�� � �
 � g � � < / � co  ��>���#��"��	t=�	=K&/�2��-�#6�,�6�,K)�,�L�A;�#�&g�J KQu��AX�� �� �� �� ���t<	/Y&/�A�#=�//�3�)�3.L;v+�Jg
�2i#�Jg�J
�K	�.
g LX0=�"!�f��� ���Y5�?����!>!%�Z!�fK����	�K'0�'��!�fK��  +��	�K;0KJ
g��t
Yu7�".!
uw <�	�Y[v=�� f�}���<J  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/ 	 	�M@     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	ZY 	 	CP@     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	LY 	 	�R@     	�t�t J tKZt J! � <1 J6 �( <K�Z K&�J� t � J K��X�!�
�f�S6����<# J( � <8 J= �/ <K��YX"L)����	s.<
z<'u�g	�= 
 	�*@     � �/ 
 	(+@     � 
	 	4+@     
�/K 
	 	�+@     !�t��K 
	 	�T@     
�/K  	�T@     � v
�<g�ut�t!J�u �&�)J�  	TU@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	RV@     ��Y  	|V@     �
�t�  	�V@     �
=*t/ 
 	�V@     �� X J . K  	�+@     � �  	�+@     � � 
 	�,@     -�1%  	�,@     ��2 
 	h-@     � �/  	�V@     ��2  	DW@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	�Z@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	\_@     �Nu�u
/� ���g�u � .
�f�*�$t��	�gu	�g
0� � � .� � � .��g	hgu%u	�/
0_J #�  	.@     �=/  	a@     �=/S  	�a@     $�/�  	.b@     '��K�  	Vb@     ��=��'g !3�(�	<(g" � � � .�	jY  	c@     ����uf	u.u
fy.�"k  	�c@     7� � � .���  	*d@     ���  	@d@     �	���# f- �+ � < f t Y  	�d@     ���fK/[���fKg0#�fKg0t�X  	~e@     ����uf	u.u
fy.�"k  	:f@     � ��uu���
0K  	�f@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�g@     ���fK/[���fKg0#�fKg0t�X  	�h@     1� � � .���  	i@     � � � .�t�J/	PK 
 	�/@     0��  � .��gt��������y�	X  	�i@     �	=fY&* � � � .�&  	Rj@     �  �u  	cj@     � �(�K  	�j@     � �)�K  	�j@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	m@     � �/�K  	 m@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�o@     �  �u  	�o@     � � � � .��/1  	(p@     ����  	Pp@     � �(�K  	np@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�q@     � �)�K  	�q@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	�r@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	]u@     � �/�K  	|u@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	x@     �6h:J  	lx@     � � � � .��/1  	�x@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	z@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	F{@     �3g71  	�{@     � �4  	�{@     7��  	�{@     � �-�K  	|@     � �uu�(<g  	N|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	�@     <�*�=  	.�@     ���u�<L�0#  	v�@     ���  	��@     ���  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�@     7��  	"�@     ���u�<L�0#  	j�@     � �-�K  	��@     � �uu�(<g  	��@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	}�@     <�*�=  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	��@     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��@     � �uu�(<g  	ʑ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	j�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	
�@     &
�Y  	�@     &
�Y  	(�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	Ȗ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	h�@     � �uu�(<g 
 	95@     �� J J . K 
 	6@     &  � .��gt���J����� g	   
  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/ansi/include ../options/internal/include/bits ../options/internal/include ../subprojects/cxxshim/stage2/include  formatting.hpp   charcode.hpp   charset.hpp   ctype-stubs.cpp   optional.hpp   string.hpp   logging.hpp   stddef.h   wctype.h   types.h   stdint.h   mbstate.h   type_traits   debug.hpp   <built-in>      	�(@     2&�*M  	�)@     1�  	��@     /KJ	=J J �K�)�&�)�(K%�(�K$0�JgZ �� �� Y - 	��@     !1u" f1 f? f1 � t 
Y  	��@     #���
g+u.J =0#���
g+u.J =0#���
g,u/J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g"u%� =0#���
gu� =4)��t
g+u.J =0)��t
g+u.J =0)��t
g,u/J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g"u%� =!.!�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 Ju�/�5 T��	� Y 0��#���
g+Y K0#���
g+Y K4���  	�)@     �<  	�)@     7�  	�@     �h��K;0  	4�@     *��JYu � �gt�$J�K r
wY  	�*@     � �/  	(+@     � 	 	4+@     
�/K 	 	�+@     !�t��K  	�+@     � �  	�+@     � �  	�,@     -�1%  	�,@     ��2  	h-@     � �/  	.@     �=/  	�/@     0��  � .��gt��������y�	X �)   O  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   environment.cpp   optional.hpp   string.hpp   logging.hpp   vector.hpp   utility   mutex.hpp   utility.hpp   errno.h   stdio.h   stddef.h   types.h   stdint.h   type_traits   debug.hpp   <built-in>      	:M@     �F  	�M@     ��  	�M@     �6J7tXK�  	�M@     �Ju 2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	M@     5//
�!  	�@     ��#f 2 	��@     % �"�#JK� � �" �1  	 7: � ���K vf
�u4�CK �B JC X	8u0������ � � � � �v�
�w�
 Q0)� #�gu�J.[ ��J�=�
��/��� #�g t � .�   < t X J)��4��w
�� ��*
u!�"J!� t%�,�/� = 0�/�u�Y	5Y@v"����!�0 57��	��� 2� ��Y	D Y ��Y	&Y  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/  	�@     �h��K;0 	 	�@     6" �  �gt�Y dxu 	 	�*@     � �/ 	 	(+@     � 		 	4+@     
�/K  	d�@     
�u 	 	v�@     &
�� 		 	��@     
�/K 		 	�+@     !�t��K  	��@     � = t � .�1t#  	4�@     *��JYu � �gt�$J�K r
wY 
 	0�@     �N.R$ 
 	��@     �� � � fvJ�� 
 	Ĳ@     � 
�� 
 	ֲ@     � � � � fv� 
 	
�@     ���/��J<��
=K 
 	��@     ��2/���J<�u
=K 
 	�@     � 
���= 
 	*�@     � 
����= 
	 	P�@     � 
�� ! 	b�@     0�u  	s�@     ��
K�
u�u 
 	´@     ��="�!�t	�K  	�+@     � �  	�+@     � � 	 	�,@     -�1%  	�,@     ��2  	�@     ��6 	 	h-@     � �/  	T�@     �#f ! 	~�@     0�u  	�T@     � v
�<g�ut�t!J�u �&�)J�  	TU@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	RV@     ��Y 
 	��@     ��	��� � �# g, �" � � � ew � � fvJ���t�   	.@     �=/  	��@     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	DW@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	|V@     �
�t� 	 	�/@     0��  � .��gt��������y�	X 	 	6@     &  � .��gt���J�����  	��@     �=7  	�a@     $�/�  	.b@     '��K�  	Vb@     ��=��'g !3�(�	<(g" � � � .�	jY  	c@     ����uf	u.u
fy.�"k  	�c@     7� � � .���  	*d@     ���  	@d@     �	���# f- �+ � < f t Y  	�d@     ���fK/[���fKg0#�fKg0t�X  	�Z@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	,.@     �/4  	Rj@     �  �u  	�h@     1� � � .���  	cj@     � �(�K  	�j@     � �)�K  	�j@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	m@     � �/�K  	 m@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�o@     �  �u  	�o@     � � � � .��/1  	(p@     ����  	Pp@     � �(�K  	np@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�q@     � �)�K  	�q@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	~e@     ����uf	u.u
fy.�"k  	:f@     � ��uu���
0K  	�f@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�g@     ���fK/[���fKg0#�fKg0t�X  	i@     � � � .�t�J/	PK  	�0@     �	/fY%* � � � .�%  	�{@     7��  	�{@     � �-�K  	|@     � �uu�(<g  	N|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	�@     <�*�=  	.�@     ���u�<L�0#  	v�@     ���  	��@     ���  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�@     7��  	]u@     � �/�K  	"�@     ���u�<L�0#  	j�@     � �-�K  	�r@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	|u@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	x@     �6h:J  	lx@     � � � � .��/1  	�x@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	z@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	F{@     �3g71  	�1@     � �3  	��@     � �uu�(<g  	ʑ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	j�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	
�@     &
�Y  	�@     &
�Y  	}�@     <�*�=  	��@     � �uu�(<g  	(�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	Ȗ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�3@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	h�@     � �uu�(<g 
 	95@     �� J J . K D    >   �      ../options/ansi/generic  errno-stubs.cpp    �5   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include/mlibc ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/posix/include/bits/posix  new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   file-io.cpp   optional.hpp   list.hpp   logging.hpp   utility.hpp   allocation.hpp   utility   intrusive.hpp   mutex.hpp   file-io.hpp   errno.h   stddef.h   types.h   stdint.h 	  ssize_t.h 
  stdio.h   off_t.h 
  type_traits   string.hpp   debug.hpp   <built-in>     2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	:M@     �F  	�M@     ��  	�M@     �6J7tXK�  	�M@     �Ju  	�@     /V�D��������!�/> K��Y�Y���Y��-��Yv<
����Z��"MB' ���XK!��0��g��tY�
�� J �Y�Y������ g� g�;�)g��tY���!$ ��/�-�fBJ� ��JY�	� YT>' ���XK!��� �1��g�� ��
���Y g� g�� J �Y�Y��� ��(�&�:�X:<wK�,Y�u�
tuM ���	t��<"��+Y�3��<'�0��7��<�����-��$�:��<��g�XKw	 Y#> ��
����<g5L� J�	�Y0������L���Y�g[�
gY	�Y00.���
g)Z#�;<3� <t	u Y30/�
g�&g �8<0�<6��<�/[ f f1��<g/^	� Y!>�t
K"v�f
gY �	�Y$>�t
K v�!<XKu �	�Y">��
g���
Y�tVZ��3<��g��� �� J���V�3�A��f&�$�J.g/Z ��gxf	XY >! 
g����/<�9��g��5�?���
Z	v Y0��
g�tY J� J���	�Y*0� ���[$�g�$B$/(/L	�u>!��Y�Y��<
g	YY0>�"	g
�u	�
�v >30��	�
��<	g
�u	�
�v�&X��ZJ>v�
gY	� YQ>v�
gY	� YC>g�
g	YY
<�L" 1 � / �g�Y� � �]&D� t � X K �0��&-<E�7�S�&<S�&<S�1U��"<��K
g���K
g�	v��6�7�?�K����	���K�	�K�	�
Ku��7�? K���v�X�	g
�5v'�TY X f Y&6E�7�S�&<S�&<S�(z�u�Y��5�'�TY X fY0� t � X K u � XKu��XKu	�=50/ t � X K �	g�	vY0� t � X L X	g�	� K&0� t � X K � X
K	uY/��C0h t � X K"g<
��v"g<
g�v"g<
g�	w�	wY0� t � X K Y /$>� t � X K	 = = 0� t � X K ��{<�Kv.�*K3�*<	�3�	J3�=��Kv.�*K3�*<	�3�	J3�=��� ��{���X�X�X��&<J  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/  	J�@     � "�&f  	l�@     3�7�  	��@     �  � � .(�� � � .� � � .� � � .��Y���.K�f>�.Kg 	 	�*@     � �/ 	 	(+@     � 		 	4+@     
�/K 		 	�+@     !�t��K  	�T@     � v
�<g�ut�t!J�u �&�)J�  	TU@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	RV@     ��Y  	2�@     � � � � .�g  	��@     � � � .� � � .1�!.�,K.�JY  � .�� 0 � .�J�Nu � � .�J�� / � .#�. ��.? � � .�.u.�.
LK 	 	J*@     � �/ 	 	t*@     � 		 	�*@     
�/K 		 	�*@     !�t��K 

 	s�@     �� X J . K 

 	�V@     �� X J . K 		 	��@     
�/K  	|V@     �
�t�  	��@     �(�%  	��@     ��K  	�@     ;�.=  	F�@     ?��uK  	x�@     4�u 		 	��@     
/K  	��@     �v/�#  	��@     �K  	�+@     � �  	�+@     � �  		�@     
�K  	�@     $��� ! 	H�@     0�u  	Z�@     1�� 	 	�,@     -�1%  	�,@     ��2 	 	h-@     � �/  	DW@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�   	 	�+@     -�1%  	�+@     ��2 	 	�,@     � �/  	t�@     ��0  	�Z@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	��@     8�t� 	 	��@     ,� ��  	
�@     ��4  	R�@     �=� 
 	��@     !��  	��@     ��  	.@     �=/  	�a@     $�/�  	.b@     '��K�  	Vb@     ��=��'g !3�(�	<(g" � � � .�	jY  	c@     ����uf	u.u
fy.�"k  	�c@     7� � � .���  	*d@     ���  	@d@     �	���# f- �+ � < f t Y  	�d@     ���fK/[���fKg0#�fKg0t�X  	�-@     �=/  	��@     �/4  	~e@     ����uf	u.u
fy.�"k  	:f@     � ��uu���
0K  	�f@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�g@     ���fK/[���fKg0#�fKg0t�X  	�h@     1� � � .���  	i@     � � � .�t�J/	PK  	�@     �K��/[4��K � � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY s�k�$  
 	>�@     �K 	 	�/@     0��  � .��gt��������y�	X  	Rj@     �  �u  	cj@     � �(�K  	�j@     � �)�K  	�j@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	m@     � �/�K  	 m@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�o@     �  �u  	�o@     � � � � .��/1  	(p@     ����  	Pp@     � �(�K  	np@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�q@     � �)�K  	�q@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1 	 	v.@     0��  � .��gt��������y�	X  	L�@     �	/fY%* � � � .�%  	�r@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	]u@     � �/�K  	|u@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	x@     �6h:J  	lx@     � � � � .��/1  	�x@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	z@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	F{@     �3g71  	�{@     7��  	�{@     � �-�K  	|@     � �uu�(<g  	N|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	�@     <�*�=  	.�@     ���u�<L�0#  	v�@     ���  	��@     ���  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�@     7��  	"�@     ���u�<L�0#  	j�@     � �-�K  	��@     � �Fg	<Y3,3  	��@     � �uu�(<g  	��@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	}�@     <�*�=  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	��@     � �uu�(<g  	ʑ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	j�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	
�@     &
�Y  	�@     &
�Y  	(�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	Ȗ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�3@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��@     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	h�@     � �uu�(<g 

 	95@     �� J J . K 	 	6@     &  � .��gt���J�����  	�@     � �!  	B�@     � � �~   �  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   stdio-stubs.cpp   optional.hpp   utility.hpp   logging.hpp   utility   mutex.hpp   string.hpp   errno.h   <built-in>    stdarg.h   stddef.h   ssize_t.h   stdio.h   types.h   stdint.h 	  type_traits   debug.hpp   list.hpp     	:M@     �F  	�M@     ��  	�M@     �6J7tXK�  	�M@     �Ju 2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	M@     5//
�!  	�@     ��#f  	x"A     � �f  	�"A     � 	���  	�"A     � 	*	�/  	L#A     � 	=�g  	�#A     � �f  	�#A     � �
t�<g��  	�#A     � � � ! � t � < < /	 � �x  	d$A     � � � � � t � < < /	 � �x  	�$A     � )�-#  	�$A     � ���Yt�<g��  	P%A     �� � !
 � �v  	�%A     �> � �
 � �v  	�%A     �&�*#  	"&A     ����)�"� �3t5�@�K �
��
t	�t�
�� J�  	,'A     �	�
t�<g��  	x'A     �� � !
 � �v  	�'A     �= � �
 � �v " 	n�@     ��4���	��vX	g�	vYV/Y�K��f�=?���J?Y-	&gI/Y-	&g00Y-	)gL.�-�0�0�0� 0� 0�0�2�"/�<Y\�Y-	*gJ/Y-	&g@�	�0�t�t	�Ov.YX�-&g[/>�02KA�tuJYt � fY0�tuJYt� � fYZl.= t � X J � �' f !@/��@/�7�"
u�'��5J)�f*<,<= K[�>�02JJ<=K`/=@�Y?�YL�<K�<�YJ�YW�tV�t-�Y,�Y9��8��ؼ�
u	u uP0= t���g�=i�
fu�=iw�[g�=`f"XY)0�g�t
K	u Y /�L0�/'t
K	uYC/�/!0��0��0K!0K!(0�g�t
K	u =/�0�g/��08�� X � X	 L ��'WLu	JYww�.�X
K	w Y0�=�. ��9����׺�J��׬ ��H�uuP0uuC0�3�� ���>�$t=0�$t= 0�� t t
K	"+:B� �	���	���
Y��2u<X��fK�
��=�=�E�O1�����F�g3�Y-	&gD0>��
2�JJ<=JuK2!�NX��>!�PX��>!�QX��)>��$>�$t=&0�$t="0
��t
K	uJ =Q0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��&�-�t�WM�Y��/t]s�
X&� mf
�vX0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��-�4�t�WM�Y��/t]s�
X&� mf
�v+0/�y�	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=�}.	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=  	�)@     �<  	�)@     7�  	(A     � 
��  	�)@     )���u�K&<f/ 
 	�V@     �� X J . K  	.(A     #�'f  	X(A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	$/A     #�'f  	N/A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X 
 	s�@     �� X J . K  	6A     #�'f  	D6A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	�T@     � v
�<g�ut�t!J�u �&�)J�  	TU@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	|V@     �
�t� 	 	�*@     � �/ 	 	(+@     � 		 	4+@     
�/K 		 	��@     
�/K 		 	�+@     !�t��K  	=A     #�'f  	:=A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	�+@     � �  	�+@     � � 
! 	DA     0�g  	DA     =�  	HDA     K  	rDA     "=�/  	�DA     <�/K  	�DA     $(=�K  	8EA     (5+�'Z+�'Z+�'Z �� �� �� �� �� f�.t�Z ��	�.�J�[2���  	IA     =�  	8IA     K  	bIA     (5+�'Z+�'Z+�'Z �� �� �� �� �� f�.t�Z ��	�.�J�[2���  	0MA     =�  	bMA     K  	�MA     (5+�'Z+�'Z+�'Z �� �� �� �� �� f�.t�Z ��	�.�J�[2���  	�Z@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
 	 	�,@     -�1%  	�,@     ��2  	�@     ��6 	 	h-@     � �/  	ZQA     =�  	�QA     K  	�QA     (5+�'Z+�'Z+�'Z �� �� �� �� �� f�.t�Z ��	�.�J�[2���  	�UA     � �  J �*KJJ�	�' J � < KJ�*>�0./�	<' J �!KJ�)>� 1��� 
 	��@     �K  	�VA     � � � � .�K  	�VA     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	�]A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	p^A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	F_A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	 `A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�`A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�aA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	�bA     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	[jA     ��_/0 � .� 		 	��@     
/K  	�jA     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	�qA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	trA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	JsA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	$tA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�tA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�uA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	�vA     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	_~A     ��_/0 � .�  	�~A     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	��A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	x�A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	N�A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	(�A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	��A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	؉A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��A     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	c�A     ��_/0 � .�  	�a@     $�/�  	.b@     '��K�  	@d@     �	���# f- �+ � < f t Y  	~e@     ����uf	u.u
fy.�"k  	:f@     � ��uu���
0K  	�c@     7� � � .���  	�f@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�g@     ���fK/[���fKg0#�fKg0t�X  	�h@     1� � � .���  	�d@     ���fK/[���fKg0#�fKg0t�X  	i@     � � � .�t�J/	PK  	.@     �=/  	��@     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	ǒA     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	��A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	|�A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	R�A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	,�A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	ܝA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��A     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	g�A     ��_/0 � .� 
 	˦A     ��
=�
g�g 
! 	�A     0�u 
 	&�A     ��
=�
g�g  	p�A     � �4  	�@     �h��K;0 	 	v�@     &
��  	ȧA     �h�K;0 	 	"�A     &
��  	4�A     � �Fu	Ju4,4  	ӨA     � �3  	(�A     � �4  	
�@     ��4  	�A     � �4  	֩A     � �Fu	Ju4,4  	u�A     � �3  	ʪA     � �4  	!�A     � �4  	x�A     � �Fu	Ju4,4  	�A     � �3  	l�A     � �4  	Rj@     �  �u  	Pp@     � �(�K  	�q@     � �)�K  	�r@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	]u@     � �/�K  	|u@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�o@     �  �u  	x@     �6h:J  	*d@     ���  	lx@     � � � � .��/1  	(p@     ����  	cj@     � �(�K  	�x@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�j@     � �)�K  	z@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	�o@     � � � � .��/1  	np@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�q@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	F{@     �3g71 	 	�/@     0��  � .��gt��������y�	X 	 	6@     &  � .��gt���J�����  	��@     �=7  	ìA     � �4  	�A     � �Fu	Ju4,4  	��A     � �3  	�A     � �4  	e�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	T�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��@     �/4  	��A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	L�A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	;�A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�@     7��  	j�@     � �-�K  	��@     � �uu�(<g  	��@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	}�@     <�*�=  	"�@     ���u�<L�0#  	��@     ���  	v�@     ���  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�{@     7��  	m@     � �/�K  	.�@     ���u�<L�0#  	�{@     � �-�K  	��@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	,.@     �/4  	*�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	z�A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	95@     �� J J . K  	L�@     �	/fY%* � � � .�%  	h�@     � �uu�(<g  	(�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	Ȗ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	
�@     &
�Y  	�@     <�*�=  	|@     � �uu�(<g  	ʑ@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	j�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�0@     �	/fY%* � � � .�%  	��@     � �Fg	<Y3,3  	�1@     � �3  	�3@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��@     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h �   �   �      ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  string-stubs.cpp   errno.h   stddef.h    6 	��A     ���	t K�<�-0	uKH/�	��t J ��<�/V
2��=V	2KA0��	YKS/=���	K�t J ��<�/V2	uK70� �8��8g�g�u� zt	|Y*/	���=�= fgv�u�uY/+0�/<0	���u�=�= fgv�u�uY/T/=1��� ���<2K �	wY$/	��	!#Y�U3"g	�Y1/	�
�� J �  X t XKgV 20/	��!�f#K�U	3Y%/�� ����*Y.� �	xY0/	�
��  J �  X t XKgV 22/� �YK �!� J �+ � �
MK+|#g u�	�YU/= ��u�t	YJ
��t J t  X t XKW3�t J t  X t XKW1tKu
J�ZJ	vKD/��'1	��	!#Y�U!3�@0�?��F��C�.I�.M�.S�.A��J�<�<7�<A��J�<.��/��7�<E�<7�<+��2��4��,��1��3��W�<<��� ��J)Y,� �	wY 0�.�.�v35�Y.�Y2�Y3�Y0�Y4�Y0�Y&�Y5�/9�/-�/D�/9�/7�/*�/1�/7�0�K33/	�h�t
K	uY80=*�uA0���� �   $  �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  filesystem.cpp   types.h   stdint.h   stddef.h   ssize_t.h   off_t.h    K 	��A     
h'�tg
v YE0j'<Yv
� YD0])�uv
� Y81
0&<Kv
� Y0
�(Y00�	L<K�u Y �   �  �      ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/internal/generic ../subprojects/frigg/include/frg /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  new   allocator.hpp   allocator.cpp   eternal.hpp   utility   slab.hpp   rbtree.hpp   stddef.h   type_traits   types.h   stdint.h   mutex.hpp   <built-in>    sysdeps.hpp    2 	�(@     	�K  	4�A     �� ! 	��A     (� � J=u � J<' �; J1 �< J��0B� ��K@>= ��  	J�A     ��  	v�A     *�K  	��A     �K  	��A     '���  	��A     *�K  	��A     �K  	��A     '���  	N�A     *�K  	\�A     �t  	n�A     ��  	��A     �/ G X  
  	�A     ��  	&�A     ���  	@�A     ����  	d�A     ��( ! 	��A     �  	��A     � ��  	��A     ����  	��A     � �� �   �  �      ../options/internal/include/mlibc ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include  charcode.hpp   charcode.cpp   stddef.h   types.h   stdint.h   optional.hpp   string.hpp   logging.hpp   type_traits   mbstate.h   debug.hpp   hash.hpp   formatting.hpp   <built-in>      	��A     � S!W(  	�A     � J  	0�A     �'f  	@�A     �#t  	R�A     .�)t	<=f�JL��u�u��u�u��u�u� � ��x ��t$Xt.uf
�t�Y  	��A     ;=	tY f
�tYt�t�Y  	��A     +�X�*��5K � J
5uB0��Y)0
Lu  	X�A     � E�I(  	��A     � �!  	��A     � �  	��A     � � ��/� � � t X�Xg�LJuKut�/tt�XKu Y  	6�A     � v ��/� � � t X�Xg�KJvKu�t/tt�XKu Y  	~�A     �v ��/���XgZKJvKuv XKu Y  	��A     �v ��1 � � t X�tY<K�+��K�
hgZ ��t�Jx�y XJtYu Y  	��A     
�t�  	
�A     
�t�  	*�A     
�t�  	J�A     
�t�  	j�A     
�t� �   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   charset.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   string.hpp   debug.hpp   charcode.hpp   charset.hpp   <built-in>     2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1� # 	��A     	�Y%>u# � � J t X!K �! �. �! �9 X! .9 X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y&0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X)�z� �+ �7 �C �� � �* �6 �B �� � �� � �) �5 �A ��� � �* �6 �B � � � �) � �1 X) 	.1 	X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��)�3��	�Y%>u# � � J t XGK �  �- �: �G 
� �O XG .O X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y*0u# � � J t XK �����-X�	�g*0u# � � J t XK �����-X�	�g0
Lu  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/  	�*@     � �/  	(+@     � 	 	4+@     
�/K 	 	�+@     !�t��K 	 	^+@     
�/K  	�+@     � �  	�+@     � �  	�,@     -�1%  	�,@     ��2  	h-@     � �/  	%-@     ��0  	.@     �=/  	,.@     �/4  	�/@     0��  � .��gt��������y�	X  	�0@     �	/fY%* � � � .�%  	�1@     � �3  	�3@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	95@     �� J J . K  	6@     &  � .��gt���J����� 8     �      ../options/internal/generic ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/include/mlibc  debug.cpp   type_traits   optional.hpp   string.hpp   logging.hpp   debug.hpp   <built-in>    formatting.hpp    1 	��A     
��2L��    �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/gcc /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   guard-abi.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   string.hpp   debug.hpp   <built-in>     2 	�(@     	�K  	�(@     2&�*M  	 )@     1��  	�)@     1�  	M@     5//
�!  	@�A     �"u!��N�+$0��uF<��)�3���R>���J8<XK
�vZS/��Ju�  	�)@     �<  	�)@     7�  	�)@     )���u�K&<f/  	J*@     � �/  	t*@     � 	 	�*@     
�/K 	 	��A     
�/K 	 	�*@     !�t��K  	�+@     � �  	�+@     � �  	�+@     -�1%  	�+@     ��2  	��A     ��2  	�,@     � �/  	�-@     �=/  	��A     �=/S  	v.@     0��  � .��gt��������y�	X  	m�A     �	=fY&* � � � .�&  	�A     � �4  	c�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	95@     �� J J . K  	b5@     &  � .��gt���J�����      extensions FT_ENCODING_APPLE_ROMAN FT_Face_Internal FT_ENCODING_ADOBE_EXPERT xMin bbox tail user /home/computerfido/Desktop/Lemon/Applications/Init FT_StreamRec_ 20bitmap_info_header_t fbInfo FT_Face_InternalRec_ closeButtonBuffer num_faces FT_Size_InternalRec_ _ZN8ListNodeIP8Window_sEC4Ev FT_SubGlyph FT_DriverRec_ senderPID FT_Glyph_Format_ _ZN4ListIP8Window_sE10get_lengthEv FT_ENCODING_MS_BIG5 _ZN4ListIP8Window_sEixEj windows __mlibc_uintptr n_contours FT_ENCODING_NONE FT_UShort FT_ENCODING_MS_GB2312 FBInfo lsb_delta __buffer_size lastKey platform_id FT_Generic charmap 10win_info_t FT_ENCODING_UNICODE RemoveDestroyedWindows recieverPID renderPos horiBearingX horiBearingY FT_Bitmap descriptor FT_Vector_ main fb_info_t FT_Stream_IoFunc glyph_index mouseDown remove_at _ZN4ListIP8Window_sEC4Ev main.cpp uint8_t FT_Generic_Finalizer _ZN4ListIP8Window_sE8add_backES1_ FT_ENCODING_JOHAB compression FT_LibraryRec_ mouseX mouseY FT_ListRec_ library environ unsigned char FT_Stream ownerPID FT_Int realloc linePadding FT_ListNodeRec_ vertAdvance FT_ListNode add_front _ZN4ListIP8Window_sE10replace_atEjS1_ y_ppem yMax num_subglyphs FT_BBox_ mouseData underline_position __dirty_begin glyph __offset FT_SizeRec_ 20bitmap_file_header_t _ZN4ListIP8Window_sE6get_atEj windowInfo other hdrSize rows _ZN4ListIP8Window_sED2Ev vector2i_t decltype(nullptr) FT_ENCODING_ADOBE_STANDARD FT_Vector __mlibc_uint16 replace_at __static_initialization_and_destruction_0 FT_ENCODING_PRC operator+ stdin stream windowFound stdout vres __io_offset Vector2i FT_ENCODING_MS_SYMBOL descender _Z13AddNewWindowsv encoding outline keyMsg memory FT_StreamDesc_ ascender finalizer ListNode<Window_s*> __mlibc_int8 style_name FT_ListRec FT_CharMapRec_ clear AddNewWindows __mlibc_uint32 linearHoriAdvance __dirty_end RGBAColour FT_Encoding_ _ZN10win_info_tC2Ev family_name optind closeButtonLength _ZplRK8Vector2iS1_ FT_Generic_ __priority available_sizes format mouseDevice add_back FT_GLYPH_FORMAT_BITMAP FT_Size num_fixed_sizes operator[] rsb_delta FT_Size_Metrics this active uintptr_t FT_String FT_ENCODING_MS_WANSUNG FT_Library FT_ENCODING_SJIS _GLOBAL__sub_I_keymap_us colourNum closeButtonSurface pixel_mode List<Window_s*> __mlibc_uint64 __initialize_p FT_Face long long int __mlibc_uint8 internal FT_StreamDesc yMin depth num_glyphs mouseEventMessage underline_thickness FT_SubGlyphRec_ 13ipc_message_t FT_Fixed FT_FaceRec_ float rgba_colour_t x_scale renderBuffer FT_Glyph_Format FT_GLYPH_FORMAT_OUTLINE GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions FT_Bitmap_ palette FT_Size_Metrics_ __io_mode importantColours FT_ENCODING_ADOBE_CUSTOM FT_Encoding FT_ENCODING_MS_JOHAB FT_UInt32 FT_Glyph_Metrics autohint y_scale FT_UInt pathname FT_Bitmap_Size_ _ZN4ListIP8Window_sE9add_frontES1_ fbSurface FT_GLYPH_FORMAT_COMPOSITE __buffer_ptr FT_BBox __valid_limit FT_CharMap FT_Short x_ppem long double FILE data2 get_front _Z10DrawWindowP8Window_s FT_Size_Internal info FT_Glyph_Metrics_ FT_MemoryRec_ FT_Pos mainFont optopt _Z22RemoveDestroyedWindowsv style_flags FT_ENCODING_BIG5 surface_t n_points uint16_t palette_mode FT_Driver _ZN4ListIP8Window_sED4Ev DrawWindow FT_GLYPH_FORMAT_NONE FT_Outline_ opterr mousePos FT_ENCODING_GB2312 FT_GlyphSlot max_advance control_data FT_ENCODING_ADOBE_LATIN_1 FT_Stream_CloseFunc ~List num_grays xMax metrics get_back encoding_id FT_ENCODING_WANSUNG get_at FT_Alloc_Func num_charmaps max_advance_width _ZN4ListIP8Window_sE5clearEv horiAdvance FT_Bitmap_Size _ZN4ListIP8Window_sEC2Ev driver _ZN10win_info_tC4Ev stderr handle_t short int uint64_t bitmap generic drag colourPlanes linearVertAdvance redrawWindowDecorations FT_GLYPH_FORMAT_PLOTTER _ZN4ListIP8Window_sE9remove_atEj backgroundColor FT_Long get_length _ZN8ListNodeIP8Window_sEC2Ev FT_Slot_Internal FT_Free_Func windowHandle FT_Slot_InternalRec_ vertBearingX vertBearingY face_flags __dso_handle uint32_t dragOffset optarg _ZN4ListIP8Window_sE8get_backEv _windowCount title short unsigned int magic pitch closeInfoHeader control_len hres FT_ENCODING_OLD_LATIN_2 FT_Outline max_advance_height sizes_list __in_chrg units_per_EM _ZN4ListIP8Window_sE9get_frontEv bitmap_top tags __mlibc_int32 FT_ENCODING_MS_SJIS closeButtonFile FT_Memory __status_bits FT_GlyphSlotRec_ FT_Realloc_Func next face_index prev cursor bitmap_left /home/computerfido/Desktop/Lemon/LibC/build syscall arg0 arg1 arg2 arg4 ../sysdeps/lemon/generic/syscall.c GNU C17 8.2.0 -mtune=generic -march=x86-64 -g -fno-builtin -fPIC arg3 _ZNK3frg8optionalIiE9has_valueEv _millis sys_anon_allocate stack_buffer_logger<mlibc::InfoSink, 128> sys_exit _ZN5mlibc14sys_libc_panicEv _ZNSt17integral_constantIbLb0EE5valueE _ZSt18is_constructible_vIiJON3frg8optionalIiEEEE _fmt_basics wchar_t null_opt_type _ZNKSt17integral_constantIbLb0EEcvbEv Args _ZN3frg8optionalIiEptEv operator() endlog operator std::integral_constant<bool, true>::value_type _ZN3frg8optionalIiE13storage_unionD4Ev _ZNSt17integral_constantIbLb1EE5valueE has_value sys_anon_free _ZNSt16is_constructibleIiJON3frg8optionalIiEEEE5valueE ~storage_union long long unsigned int _ZN3frg8optionalIiEcvbEv _ZN5mlibc17sys_anon_allocateEmPPv __cxa_atexit _ZN5mlibc8sys_exitEi _ZN5mlibc12sys_libc_logEPKc _ZN3frg8optionalIiEdeEv _ZN5mlibc14sys_futex_waitEPii _ZNKSt17integral_constantIbLb1EEclEv operator std::integral_constant<bool, false>::value_type object _ZN5mlibc10sys_getpidEv clock _ZN3frg8optionalIiED4Ev sys_clock_get _ZNSt16is_constructibleIiJRKN3frg8optionalIiEEEE5valueE mlibc status time_t GNU C++17 8.2.0 -mtune=generic -march=x86-64 -g -std=c++17 -fno-builtin -fno-rtti -fno-exceptions -fPIC sys_getpid _ZN3frg8optionalIiEC4EOi pid_t expected operator-> _ZNKSt17integral_constantIbLb1EEcvbEv operator* _pid _ZN3frg8optionalIiEC4ENS_13null_opt_typeE operator= sys_libc_panic _ZN5mlibc11panicLoggerE endlog_t optional<int> _stor _ZN5mlibc13sys_anon_freeEPvm nanos _ZSt18is_constructible_vIiJRKN3frg8optionalIiEEEE small_digits _ZN3frg8optionalIiE13storage_unionC4Ev sys_libc_log null_opt _ZN3frg8optionalIiEC4EOS1_ _ZNK3frg8optionalIiEcvbEv panicLogger _non_null is_constructible<int, frg::optional<int>&&> _ZN3frg8optionalIiEC4ERKS1_ _ZN3frg8optionalIiE6_resetEv ~optional is_constructible<int, const frg::optional<int>&> operator bool _ZNKSt17integral_constantIbLb0EEclEv integral_constant<bool, false> stack_buffer_logger<mlibc::PanicSink, 128> _to_string_impl sys_futex_wait _Z19__mlibc_do_finalizev _ZN3frg8optionalIiEC4Ev _secs is_constructible_v _ZN5mlibc14sys_futex_wakeEPi _reset _ZN5mlibc13sys_clock_getEiPlS0_ _ZN5mlibc10infoLoggerE _ZN3frg8optionalIiEC4ERKi ../sysdeps/lemon/generic/lemon.cpp integral_constant<bool, true> sys_futex_wake __func__ __mlibc_do_finalize _ZNK3frg8optionalIiEdeEv infoLogger _ZN3frg8optionalIiEaSES1_ _ZN3frg3maxIiEERKT_S3_S3_ decimal _ZN3frg14format_optionsC2ERKS0_ format_integer<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> format<char const*, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg14format_optionsC4ERKS0_ _ZnwmPv format_object<frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ alt_conversion _ZN3frg14format_optionsC2Ev _ZN3frg8optionalIiED2Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg14format_options15with_conversionENS_17format_conversionE max<int> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ format<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg8optionalIiEC2Ev _sink format_integer<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> minimum_width _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ fill_zeros with_conversion format<char const*, frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4ERKS4_ left_justify number operator<< <unsigned int> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemaSERKS4_ print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic _ZN5mlibc9PanicSinkC4Ev _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4ERKS4_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD4Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEC4ES2_ format<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _emit plus_becomes_space _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev absv _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ append _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ format_conversion _ZN5mlibc8InfoSinkclEPKc _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ function _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ ../options/internal/generic/ensure.cpp message _off InfoSink _ZN3frg14format_optionsD4Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEC4ES2_ _ZN3frg8optionalIiEC2ERKS1_ __ensure_warn _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ _ZN5mlibc9PanicSinkclEPKc always_sign negative print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> radix _ZN5mlibc8InfoSinkC4Ev PanicSink _ZN3frg14format_optionsC4Ev _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE _emitted operator<< print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> format_object<frg::stack_buffer_logger<mlibc::InfoSink>::item> precision stack_buffer_logger _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg8optionalIiE13storage_unionC2Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv assertion ~format_options _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD4Ev _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ ~item _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ __ensure_fail _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemaSERKS4_ print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> operator new _ZN3frg14format_optionsD2Ev _ZN3frg8optionalIiE13storage_unionD2Ev Limit operator<< <char const*> strlen src_bytes ../options/internal/generic/essential.cpp dest_bytes mb_chr _ZN3frg11unique_lockI13AllocatorLockEC4EOS2_ size_to_bucket _ZN3frg7mt19937C2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC4Ev alignment _ZN3frg11unique_lockI13AllocatorLockEC4ENS_11dont_lock_tERS1_ replacement _ZN3frg7mt199371nE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ mag01 _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ item_size code_seq<char const> wseq mbstowcs max_size lldiv _tree_mutex strtold _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ nptr strtoll print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> lsbs get_root dont_lock_t __mlibc_rand_engine _is_locked _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg10bitop_implImE3clzEm _ZN5mlibc8code_seqIwEcvbEv operator<< <void*> _verify_integrity _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameaSERKS4_ _ZN3frg11unique_lockI13AllocatorLockED2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC4ERKS4_ tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE12huge_paddingE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14small_base_expE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ atof rotateRight _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ locale_t __cpoint _ZN5mlibc7strtofpIeEET_PKcPPc _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE12numUsedPagesEv endptr _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC4EPNS_9slab_poolIS1_S2_EE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11_find_frameEm _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ aggregate_node _usedPages atoi atol illegal_input address_ frame_hook _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC4ERS1_ wctomb _ZN3frg7mt199378matrix_aE insert_right left_ptr _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE23test_bucket_calculationEj __mlibc_errno copy _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ area_size seed _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ _ZN13AllocatorLock4lockEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ _ZN5mlibc7strtofpIfEET_PKcPPc type_ abort _ZN13AllocatorLockC4ERKS_ partial_hook slab_allocator tiny_sizes _ZN3frg11unique_lockI13AllocatorLockE9is_lockedEv result num_buckets slabsize _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ 7lldiv_t pool_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameaSERKS4_ num_reserved insert_root rbtree successor huge_padding _ZN3frg9_redblack11hook_structC4ERKS1_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ bucket_mutex isRed link _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ fix_insert _ZN3frg9_redblack11hook_structC4Ev llabs color_type mblen_state 5div_t _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ VirtualAllocator was_unavailable tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::_redblack::null_aggregator> deallocate predecessor mblen _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EaSERKSB_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE23_verify_frame_integrityEPNS3_5frameE _ZN3frg11unique_lockI13AllocatorLockE8protectsEPS1_ print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> compare _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEaSERKS3_ malloc check_invariant _frame_tree succ _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE9page_sizeE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14size_to_bucketEm replace_node _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EaSERKSB_ rand_r _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ Member frame_type program_invocation_name AllocatorLock _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ strtoul cutlim atoll aggregate<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame> dot_end _ZN3frg11unique_lockI13AllocatorLockEaSES2_ strtofp<double> _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ grand frame_less format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _construct_large address 6ldiv_t _Exit output_overflow _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ code_seq<wchar_t> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ get_right _ZN16VirtualAllocator3mapEm _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj frame_tree_type slab_frame length_ remove_half_leaf reallocate format<void*, frg::stack_buffer_logger<mlibc::InfoSink>::item> numUsedPages tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::_redblack::null_aggregator> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15max_bucket_sizeE _ZN3frg11unique_lockI13AllocatorLockE6unlockEv _ZN3frg11unique_lockI13AllocatorLockED4Ev _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg11unique_lockI13AllocatorLockEC4ERS1_ Mutex _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ _plcy _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm freelist child _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ unmap _verify_frame_integrity bsearch _ZN3frg7mt19937C4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv slab_allocator<VirtualAllocator, AllocatorLock> _redblack _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE16_construct_largeEm mb_string input_underflow _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ wcstombs isBlack _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEv system small_step_exp _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ _ZN3frg11unique_lockI13AllocatorLockEC4ERKS2_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frame8containsEPv tree_crtp_struct _ZN3frg7mt199374lsbsE protects _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC4Emmi _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC2Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10reallocateEPvm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ partial_tree calloc _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14small_step_expE strtoull _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11num_bucketsE _ZN16VirtualAllocator5unmapEmm qsort overhead _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE7reallocEPvm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistaSERKS4_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ new_size _ZN3frg3maxImEERKT_S3_S3_ enable_checking _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ _ZN13AllocatorLockaSERKS_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE17_verify_integrityEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ get_parent _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv _ZN3frg7mt199373msbE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8slabsizeE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ max<long unsigned int> program_invocation_short_name hook_struct head_slb _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8allocateEm strtofp<float> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5firstEv mb_limit mbtowc get_left rotateLeft new_length null_aggregator _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15_construct_slabEi _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ quot parent_color _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4ERKSB_ u_bytes _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm wc_limit ULONG_MAX _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC4ERKS3_ _ZN3frg7mt199374seedEj slab_pool _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv _bkts new_pointer mktemp _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4ERKSB_ bucket_guard unique_lock<AllocatorLock> matrix_a rbtree_hook at_quick_exit _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ small_base_exp aligned_alloc v_bytes index_ strtod strtof _GLOBAL__sub_I_stdlib_stubs.cpp strtol right_ptr _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4Ev func tree_guard _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC4ERKS4_ charcode_error element Policy max_bucket_size aggregate_path _ZN3frg9_redblack11hook_structaSERKS1_ __progress strtofp<long double> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10tiny_sizesE unlock _ctr test_bucket_calculation srand partial_tree_type _ZN13AllocatorLockC4Ev tree_struct _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ _ZN3frg9_redblack11hook_structC2Ev ../options/ansi/generic/stdlib-stubs.cpp cutoff strtod_l ~unique_lock _find_frame bucket_to_size tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> aggregate<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _futex _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ contains insert_left page_size _ZN5mlibc7strtofpIdEET_PKcPPc _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC4ENS3_10frame_typeEmm __shift mt19937 _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE4freeEPv _ZN5mlibc8code_seqIKcEcvbEv _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ slab_pool<VirtualAllocator, AllocatorLock> wc_string dont_lock _construct_slab dirty _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10deallocateEPvm denom posix_memalign bitop_impl<long unsigned int> pred _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC4Ev _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN13AllocatorLock6unlockEv fix_remove _ZN3frg11unique_lockI13AllocatorLockEC4Ev _ZN3frg7mt199371mE _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN3frg7mt19937clEv srandom _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC4ERKS4_ _ZN5mlibc8code_seqIjEcvbEv iswlower iscntrl isalnum _ZN3frg17basic_string_viewIcE10find_firstEcm _ZNK3frg17basic_string_viewIcE4sizeEv isprint isdigit isspace ct_digit _ZN3frg17basic_string_viewIcEC2EPKc ct_space iswspace ispunct _ZN5mlibc13wide_charcode7promoteEwRj _ZNK3frg17basic_string_viewIcEneES1_ isupper ct_punct iswcntrl toupper generic_is_control iswdigit iswpunct isgraph iswprint ct_graph isalpha basic_string_view towupper ct_alpha _ZN5mlibc18generic_is_controlEj _ZNK3frg17basic_string_viewIcEixEm iswxdigit _ZN3frg17basic_string_viewIcEC4EPKc basic_string_view<char> _ZN3frg17basic_string_viewIcEC4EPKcm ct_alnum isblank sub_string ct_blank codepoint _ZNK3frg17basic_string_viewIcEeqES1_ ct_cntrl iswblank find_first ct_upper iswalpha find_last iswctype _ZN3frg17basic_string_viewIcEC4Ev iswupper tolower operator== ct_print operator!= ct_xdigit wint_t towlower isascii _ZN5mlibc20polymorphic_charcode7promoteEcRj promote _ZNK3frg17basic_string_viewIcE4dataEv iswgraph ct_count isxdigit ct_null _ZN3frg17basic_string_viewIcE9find_lastEc iswalnum islower code_seq<unsigned int> Char _ZN3frg17basic_string_viewIcE10sub_stringEmm wctype_t ct_lower ../options/ansi/generic/ctype-stubs.cpp getenv unsetenv self _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ _ZN3frg10escape_fmtC4EPKvm update_vector _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED4Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEaSES6_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ES5_ push _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv new_capacity push_back get_vector _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm move<char*&> remove_reference<char*&> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4EOS6_ ../options/ansi/generic/environment.cpp _ZSt4swapIPcEvRT_S2_ unassign_variable operator<< <frg::escape_fmt> remove_reference<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv escape_fmt _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ remove_reference_t _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv ~vector _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backEOS1_ _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ empty_environment overwrite _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ES5_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backERKS1_ _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEENSt16remove_referenceIT_E4typeEOS7_ _ensure_capacity format<frg::escape_fmt, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERKS6_ move<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> vector<char*, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv putenv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv swap<char*> _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZN3frg10escape_fmtC2EPKvm new_array empty _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv start_from _ZN3frg17basic_string_viewIcEC2EPKcm find_environ_index _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5emptyEv _elements _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ ../options/ansi/generic/errno-stubs.cpp _ZN5mlibc13abstract_file5closeEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE4backEv default_list_hook _ZN5mlibc13abstract_file9_save_posEv chunk _ZN5mlibc13abstract_file7io_readEPcmPm _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ _vptr.abstract_file format_integer<int, frg::stack_buffer_logger<mlibc::InfoSink>::item> owner intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*> fclose _init_bufmode _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC4Ev _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ __vtbl_ptr_type _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> pipe_like whence erased remove_reference<int&> stdout_file forward<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > ssize_t rewind _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ ~fd_file fileno _write_back destruct<mlibc::abstract_file, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN5mlibc7fd_fileD2Ev _ZN3frg3minImEERKT_S3_S3_ _ZN5mlibc13abstract_file14determine_typeEPNS_11stream_typeE _ZN5mlibc13abstract_file6_resetEv composition<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > ~<lambda> _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8pop_backEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN5mlibc13abstract_file8io_writeEPKcmPm _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ _save_pos _init_type _ZN5mlibc13abstract_file10_init_typeEv _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ fileno_unlocked unknown _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN5mlibc13abstract_file13_init_bufmodeEv abstract _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5emptyEv OwnerPointer _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE _void_impl determine_bufmode intrusive_traits<mlibc::abstract_file, mlibc::abstract_file*, mlibc::abstract_file*> _ZN5mlibc13abstract_fileC4EPFvPS0_E __closure stream_type format<char, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN5mlibc13abstract_file7disposeEv fdopen _ZN3frg6formatIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc13abstract_fileD4Ev file_like update_bufmode iterator _ZN5mlibc7fd_fileC4EiPFvPNS_13abstract_fileEE _ZN5mlibc13abstract_file4seekEli _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ setvbuf io_read _GLOBAL__sub_I_file_io.cpp _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic new_offset line_buffer io_size operator<< <int> intrusive_list Locate _ZN5mlibc13abstract_fileaSERKS0_ _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE10push_frontES6_ unget _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ __for_range _ensure_allocation print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> has_plus _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN5mlibc13abstract_file5purgeEv _ZN5mlibc13abstract_file5ungetEc _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _current _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6spliceENS9_8iteratorERS9_ _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE _ZN5mlibc13abstract_file18_ensure_allocationEv io_write format<int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE _ZN5mlibc7fd_file2fdEv _ZN5mlibc13abstract_fileD0Ev _ZN5mlibc7fd_fileD4Ev print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> borrow_pointer _ZN5mlibc7fd_file5closeEv _ZN5mlibc13abstract_file7io_seekEliPl push_front BorrowPointer fseek ftell _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEi _ZN5mlibc13abstract_fileC4ERKS0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv forward<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > _ZN5mlibc7fd_fileC4ERKS0_ __for_begin _ZN5mlibc13abstract_file11_write_backEv off_t _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev previous __fpurge _ZN5mlibc13abstract_file4readEPcmPm current_offset ~abstract_file globallyDisableBuffering global_file_list _ZN5mlibc13abstract_file5flushEv _ZN5mlibc13abstract_fileC2EPFvPS0_E intrusive_list_hook _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ min<long unsigned int> stderr_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC4ES6_ io_seek _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIiEERS4_T_ actual_size __for_end _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE full_buffer _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv _ZN5mlibc7fd_fileD0Ev <lambda(mlibc::abstract_file*)> remove_reference<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6insertENS9_8iteratorES6_ operator void (*)(mlibc::abstract_file*) move<mlibc::abstract_file*&> args#1 fopen _result_of_impl splice owner_pointer determine_type locate_tag remove_reference<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > args#0 _ZN5mlibc13abstract_file5writeEPKcmPm decay _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5frontEv pop_front _ZN5mlibc7fd_file7io_seekEliPl operator<< <char> remove_reference<mlibc::abstract_file*&> operator++ borrow _ZN5mlibc7fd_fileC4EOS0_ buffer_mode _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ _do_dispose pop_back _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC4Ev remove_reference<frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>&> intrusive_list<mlibc::abstract_file, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > ungetc erase no_buffer flush_line get<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > seek_offset global_stdio_guard ../options/ansi/generic/file-io.cpp _ZN5mlibc7fd_file7io_readEPcmPm _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic in_list ~stdio_guard _ZN5mlibc13abstract_file4tellEPl stdin_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ _ZN5mlibc13abstract_fileD2Ev _ZN5mlibc13abstract_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc7fd_file8io_writeEPKcmPm iterator_to forward<int&> _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE fflush _FUN fflush_unlocked _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9pop_frontEv print_int<StreamPrinter, long int> _ZN3frg17basic_string_viewIwE9find_lastEw do_printf_ints<StreamPrinter> fgetc printf_format<PrintfAgent<StreamPrinter> > print_int<StreamPrinter, long unsigned int> fgets _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev vfprintf _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN11PrintfAgentI14LimitedPrinterEclEc _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_digits<BufferPrinter, long int> vswscanf fread_unlocked print_digits<ResizePrinter, long unsigned int> _ZN13ResizePrinter6expandEv BufferPrinter renameat fputws _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev vasprintf _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _vsp putchar __mlibc_intmax print_digits<BufferPrinter, long long unsigned int> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev is_constructible<int, int&&> print_int<ResizePrinter, long long unsigned int> fgetpos _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ clearerr _ZN13ResizePrinterC4Ev _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic SCANF_TYPE_INT print_int<ResizePrinter, long int> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ fputs_unlocked _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic ftrylockfile SCANF_TYPE_SIZE_T vfscanf _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN13StreamPrinter6appendEPKc print_digits<BufferPrinter, long unsigned int> do_scanf<sscanf(char const*, char const*, ...)::<unnamed class> > swap<int> _ZN3frg4swapERNS_8optionalIiEES2_ _ZNK3frg17basic_string_viewIwEneES1_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ print_digits<LimitedPrinter, long int> bytes_read feof_unlocked print_int<BufferPrinter, unsigned int> default_size print_int<ResizePrinter, long unsigned int> _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ vscanf _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN3frg17basic_string_viewIwEC2EPKw PrintfAgent _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ filename <lambda(auto:1)> fgetwc getwchar _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_int<LimitedPrinter, long int> fgetws vwprintf _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ do_printf_chars<LimitedPrinter> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE native_size _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ __builtin_va_list do_scanf<vfscanf(FILE*, char const*, __va_list_tag*)::<unnamed struct> > _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ do_printf_floats<LimitedPrinter> __gnuc_va_list handler _ZNK3frg17basic_string_viewIwE4sizeEv clearerr_unlocked _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZN11PrintfAgentI13StreamPrinterEC4EPS0_PN3frg9va_structE move<bool&> _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic print_int<BufferPrinter, long unsigned int> fwrite_unlocked _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE print_digits<StreamPrinter, long unsigned int> do_printf_chars<BufferPrinter> _ZN13BufferPrinterC2EPc _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic ungetwc fp_offset ptrdiff_t new_limit _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg8optionalIiEC4IRivEEOT_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ vsnprintf _ZN11PrintfAgentI13BufferPrinterEclEc new_path _ZSt4swapIiEvRT_S1_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ new_buffer vswprintf szmod _ZNK3frg17basic_string_viewIwEixEm print_int<LimitedPrinter, long unsigned int> fwide _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic _ZN14LimitedPrinter6appendEPKcm funlockfile _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _ZSt18is_constructible_vIiJRiEE putchar_unlocked _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic print_int<StreamPrinter, unsigned int> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE putwchar print_int<ResizePrinter, unsigned int> _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ SCANF_TYPE_PTRDIFF _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN3frg17basic_string_viewIwE10find_firstEwm print_digits<StreamPrinter, long int> rename _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ print_digits<ResizePrinter, long int> <lambda(auto:2)> do_printf_ints<BufferPrinter> print_digits<LimitedPrinter, long long unsigned int> _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ ferror vfwprintf _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic print_int<StreamPrinter, long long unsigned int> unused _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ args _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN13ResizePrinter6appendEc _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic _ZNSt16is_constructibleIiJOiEE5valueE _ZN3frg17basic_string_viewIwEC4Ev _ZN11PrintfAgentI13ResizePrinterEC4EPS0_PN3frg9va_structE _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE PrintfAgent<ResizePrinter> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic printf_size_mod second printf_format<PrintfAgent<BufferPrinter> > StreamPrinter _ZN3frg8optionalIiEC2EOi PrintfAgent<StreamPrinter> _ZN13StreamPrinter6appendEPKcm _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN11PrintfAgentI13BufferPrinterEC4EPS0_PN3frg9va_structE SCANF_TYPE_SHORT _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN11PrintfAgentI13ResizePrinterEclEc gp_offset _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE vprintf _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN11PrintfAgentI13BufferPrinterEclEPKcm perror move<int&> consume fputc_unlocked _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN14LimitedPrinter6appendEc _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN11PrintfAgentI13StreamPrinterEclEc _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE agent optional<int&> _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN13ResizePrinter6appendEPKcm overflow_arg_area _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev operator()<long unsigned int> fsetpos _ZN14LimitedPrinter6appendEPKc _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZN13BufferPrinterC4EPc <lambda(auto:3)> SCANF_TYPE_LL setbuf feof _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE print_int<BufferPrinter, long int> intmax_t LimitedPrinter expand __opts _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic olddirfd _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg8optionalIiEC2IRivEEOT_ swap<bool> va_struct _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE swap _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE fgets_unlocked num_consumed _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13ResizePrinterEclEPKcm _ZN3frg17basic_string_viewIwEC4EPKwm reg_save_area getdelim _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN14LimitedPrinterC2EPcm _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE invert _ZN13StreamPrinter6appendEc _ZN11PrintfAgentI14LimitedPrinterEC4EPS0_PN3frg9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev getchar_unlocked print_int<LimitedPrinter, unsigned int> old_path print_digits<BufferPrinter, unsigned int> _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic match_count ~<constructor> _ZNSt16is_constructibleIiJRiEE5valueE print_int<BufferPrinter, long long unsigned int> _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic __formatter _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev longlong_size _ZN14LimitedPrinterC4EPcm remove_reference<bool&> vsscanf do_printf_ints<ResizePrinter> ../options/ansi/generic/stdio-stubs.cpp SCANF_TYPE_CHAR _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ fputs vwscanf _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev getline _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN13BufferPrinter6appendEPKc _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZSt4swapIbEvRT_S1_ do_printf_ints<LimitedPrinter> _ZNK3frg17basic_string_viewIwEeqES1_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev _ZN3frg17basic_string_viewIwE10sub_stringEmm print_int<LimitedPrinter, long long unsigned int> _ZNK3frg17basic_string_viewIwE4dataEv freopen print_digits<StreamPrinter, long long unsigned int> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ print_digits<ResizePrinter, long long unsigned int> tmpnam _ZN13ResizePrinter6appendEPKc SCANF_TYPE_INTMAX scanset newdirfd look_ahead tmpfile print_digits<StreamPrinter, unsigned int> auto:2 auto:3 _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN13BufferPrinter6appendEc ferror_unlocked print_digits<ResizePrinter, unsigned int> SCANF_TYPE_L fread _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ do_printf_floats<StreamPrinter> fputc auto:1 do_printf_chars<StreamPrinter> print_digits<LimitedPrinter, long unsigned int> _ZN13BufferPrinter6appendEPKcm _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE fpos_t _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ PrintfAgent<LimitedPrinter> fgetc_unlocked _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev basic_string_view<wchar_t> _ZN3frg17basic_string_viewIwEC4EPKw fputwc _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev typed_dest store_int is_constructible<int, int&> PrintfAgent<BufferPrinter> _ZN13StreamPrinterC2EP17__mlibc_file_base vfwscanf _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ printf_format<PrintfAgent<ResizePrinter> > _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev vsprintf do_printf_floats<BufferPrinter> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev ResizePrinter _ZN13StreamPrinterC4EP17__mlibc_file_base _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ flockfile do_printf_floats<ResizePrinter> do_printf_chars<ResizePrinter> printf_format<PrintfAgent<LimitedPrinter> > _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZSt18is_constructible_vIiJOiEE operator()<unsigned int> _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ typedef __va_list_tag __va_list_tag fwrite print_digits<LimitedPrinter, unsigned int> getchar _ZN13ResizePrinterC2Ev wcsrchr strchrnul pattern wmemmove wmemcmp wcsncat bufsz wmemset wcstod wcscpy wcstof wcsncpy stpcpy wcstok wcstold wcstoull wcstol chrs wcstoll strerror ../options/ansi/generic/string-stubs.cpp delimiter strtok_r wcspbrk wcschr mempcpy wcsncmp wcsstr b_byte strtok wcscspn wcscat wcslen s_bytes strchr strncat strcspn wcstoul wcscmp strncpy strerror_r strcoll strcpy a_byte strxfrm wmemchr strspn wcscoll found wcsspn strcat strcmp saved strstr wcsxfrm strrchr wmemcpy strncmp strpbrk sys_access sys_close written sys_read _ZN5mlibc8sys_openEPKciPi _ZN5mlibc10sys_accessEPKci ../sysdeps/lemon/generic/filesystem.cpp sys_write sys_open _ZN5mlibc8sys_seekEiliPl sys_errno _ZN5mlibc9sys_writeEiPKvmPl _ZN5mlibc9sys_closeEi sys_seek _ZN5mlibc8sys_readEiPvmPl _ZN3frg15aligned_storageILm456ELm8EEC2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC2ERS1_ remove_reference<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less&> _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _ZN3frg15aligned_storageILm1ELm1EEC2Ev heap Align _ZN3frg7eternalI16VirtualAllocatorE3getEv aligned_storage<8, 8> aligned_storage eternal<> _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC4IJRS2_EEEDpOT_ eternal<VirtualAllocator&> _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEE3getEv move<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less&> remove_reference<frg::slab_pool<VirtualAllocator, AllocatorLock>*> _ZSt7forwardIPN3frg9slab_poolI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ eternal<frg::slab_allocator<VirtualAllocator, AllocatorLock> > MemoryAllocator getAllocator _ZSt4moveIRN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ _ZN3frg15aligned_storageILm8ELm8EEC4Ev forward<VirtualAllocator&> aligned_storage<456, 8> _ZN3frg7eternalI16VirtualAllocatorEC4IJEEEDpOT_ eternal<frg::slab_pool<VirtualAllocator, AllocatorLock>*> eternal<VirtualAllocator> virtualAllocator forward<frg::slab_pool<VirtualAllocator, AllocatorLock>*> _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2EPNS_9slab_poolIS1_S2_EE _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv _Z12getAllocatorv eternal<frg::slab_pool<VirtualAllocator, AllocatorLock> > _ZN3frg15aligned_storageILm8ELm8EEC2Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE aligned_storage<1, 1> _ZN3frg15aligned_storageILm456ELm8EEC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev _ZN13AllocatorLockC2Ev _ZN3frg15aligned_storageILm1ELm1EEC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC2Ev singleton ../options/internal/generic/allocator.cpp remove_reference<VirtualAllocator&> global_wide_charcode code_seq<unsigned int const> _ZN5mlibc16current_charcodeEv _ZN5mlibc8code_seqIKwEcvbEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate promote_wtranscode has_shift_states_ _ZN5mlibc20polymorphic_charcodeC2Ebb platform_wide_charcode _ZN5mlibc20polymorphic_charcodeD4Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED4Ev preserves_7bit_units _ZN5mlibc20polymorphic_charcodeC4ERKS0_ decode_wtranscode utf8_charcode code_seq<char> _ZN5mlibc13utf8_charcode16has_shift_statesE _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4Ev decode_wtranscode_length _ZN5mlibc20polymorphic_charcode17decode_wtranscodeERNS_8code_seqIKcEERNS1_IwEER15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode6decodeERNS_8code_seqIKcEERNS1_IjEER15__mlibc_mbstate _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4ERKS2_ auto has_shift_states _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE encode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate decode polymorphic_charcode_adapter<mlibc::utf8_charcode> _ZN5mlibc13utf8_charcode20preserves_7bit_unitsE code_seq<wchar_t const> _ZN5mlibc8code_seqIcEcvbEv _ZN5mlibc13utf8_charcode12decode_stateC4Ev global_charcode _ZN5mlibc20polymorphic_charcodeD2Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE ../options/internal/generic/charcode.cpp decode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _vptr.polymorphic_charcode current_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN5mlibc20polymorphic_charcode24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode17encode_wtranscodeERNS_8code_seqIcEERNS1_IKwEER15__mlibc_mbstate ~polymorphic_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13utf8_charcode12decode_state6cpointEv encode_wtranscode _ZN5mlibc13utf8_charcode12decode_stateC2Ev _ZN5mlibc13utf8_charcode12decode_state8progressEv preserves_7bit_units_ ~polymorphic_charcode_adapter _ZN5mlibc8code_seqIKjEcvbEv _ZN5mlibc22platform_wide_charcodeEv _ZN5mlibc20polymorphic_charcodeC4Ebb _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4EOS2_ _ZN5mlibc20polymorphic_charcodeD0Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev encode_state _ZN5mlibc20polymorphic_charcode18promote_wtranscodeEcRw decode_state _ZN5mlibc7charset8is_blankEj is_graph _ZN5mlibc7charset8is_alphaEj is_alpha _ZN5mlibc7charset8is_spaceEj is_alnum is_blank _ZN5mlibc7charset8is_printEj is_upper _ZN5mlibc7charset8is_lowerEj _ZN5mlibc7charset8is_upperEj _ZN5mlibc15current_charsetEv _ZN5mlibc7charset8is_graphEj _ZN5mlibc7charset9is_xdigitEj ../options/internal/generic/charset.cpp is_lower _ZN5mlibc7charset8to_lowerEj _ZN5mlibc7charset8is_alnumEj to_lower _ZN5mlibc7charset8to_upperEj _ZN5mlibc7charset17is_ascii_supersetEv is_digit _ZN5mlibc7charset8is_digitEj is_space global_charset is_ascii_superset is_punct _ZN5mlibc7charset8is_punctEj is_print is_xdigit current_charset to_upper ../options/internal/generic/debug.cpp Guard _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic __mlibc_int64 ../options/internal/gcc/guard-abi.cpp _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ complete _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ __cxa_guard_acquire __cxa_guard_release format<void*, frg::stack_buffer_logger<mlibc::PanicSink>::item> format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> __cxa_pure_virtual _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_                 ]@     L@     L@     �@     �@     �@     �@     �@     �@     @     @     *@     *@     W@     X@     z@     z@     H@     H@     �@     �@     �@                     y&@     �(@     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     �)@     �)@     �)@     �)@     �)@     J*@     J*@     s*@     t*@     *@     �*@     �*@     �*@     �*@     �*@     �*@     �*@     '+@     (+@     3+@     4+@     ]+@     ^+@     �+@     �+@     �+@     �+@     �+@     �+@     �+@     �+@     �+@     �+@     C,@     C,@     �,@     �,@     �,@     �,@     �,@     �,@     %-@     %-@     h-@     h-@     �-@     �-@     �-@     �-@     .@     .@     ,.@     ,.@     v.@     v.@     G/@     G/@     �/@     �/@     �0@     �0@     Q1@     Q1@     �1@     �1@     �1@     �1@     �3@     �3@     95@     95@     a5@     b5@     6@     6@     �6@                     AO@     P@     P@     P@                     �Q@     TR@     ZR@     [R@                     �S@     �T@     �T@     �T@                     N8@     eJ@     fJ@     �J@     �J@     3K@     4K@     M@     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     M@     :M@     :M@     �M@     �M@     �M@     �M@     �M@     �M@     �M@     �)@     �)@     �)@     �)@     �)@     J*@     �M@     CP@     CP@     �R@     �R@     �T@     �*@     '+@     (+@     3+@     4+@     ]+@     �+@     �+@     �T@     �T@     �T@     TU@     TU@     QV@     RV@     {V@     |V@     �V@     �V@     �V@     �V@     �V@     �+@     �+@     �+@     �+@     �,@     �,@     �,@     %-@     h-@     �-@     �V@     DW@     DW@     �Z@     �Z@     \_@     \_@     a@     .@     ,.@     a@     �a@     �a@     .b@     .b@     Ub@     Vb@     c@     c@     �c@     �c@     )d@     *d@     @d@     @d@     �d@     �d@     ~e@     ~e@     :f@     :f@     �f@     �f@     �g@     �g@     �h@     �h@     i@     i@     �i@     �/@     �0@     �i@     Qj@     Rj@     cj@     cj@     �j@     �j@     �j@     �j@     m@     m@     m@      m@     �o@     �o@     �o@     �o@     (p@     (p@     Pp@     Pp@     np@     np@     �q@     �q@     �q@     �q@     �r@     �r@     ]u@     ]u@     {u@     |u@     x@     x@     lx@     lx@     �x@     �x@     z@     z@     E{@     F{@     �{@     �{@     �{@     �{@     �{@     �{@     |@     |@     M|@     N|@     �@     �@     .�@     .�@     v�@     v�@     ��@     ��@     ��@     ��@     �@     �@     "�@     "�@     j�@     j�@     ��@     ��@     ��@     ��@     }�@     }�@     ��@     ��@     ��@     ��@     ��@     ��@     ɑ@     ʑ@     j�@     j�@     
�@     
�@     �@     �@     (�@     (�@     Ȗ@     Ȗ@     h�@     h�@     ��@     95@     a5@     6@     �6@                     ��@     ��@     �(@      )@     �)@     �)@     ��@     ��@     ��@     �@     �)@     �)@     �)@     �)@     �@     4�@     4�@     ��@     �*@     '+@     (+@     3+@     4+@     ]+@     �+@     �+@     �+@     �+@     �+@     �+@     �,@     �,@     �,@     %-@     h-@     �-@     .@     ,.@     �/@     �0@                     ��@     �@     :M@     �M@     �M@     �M@     �M@     �M@     �M@     �M@     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     M@     :M@     �@     �@     �)@     �)@     �)@     �)@     �)@     J*@     �@     4�@     �@     c�@     �*@     '+@     (+@     3+@     4+@     ]+@     d�@     u�@     v�@     ��@     ��@     ��@     �+@     �+@     ��@     0�@     4�@     ��@     0�@     ��@     ��@     ò@     Ĳ@     ֲ@     ֲ@     
�@     
�@     ��@     ��@     �@     �@     )�@     *�@     O�@     P�@     b�@     b�@     s�@     s�@     ´@     ´@     �@     �+@     �+@     �+@     �+@     �,@     �,@     �,@     %-@     �@     T�@     h-@     �-@     T�@     ~�@     ~�@     ��@     �T@     TU@     TU@     QV@     RV@     {V@     ��@     ��@     .@     ,.@     ��@     ��@     DW@     �Z@     |V@     �V@     �/@     �0@     6@     �6@     ��@     �@     �a@     .b@     .b@     Ub@     Vb@     c@     c@     �c@     �c@     )d@     *d@     @d@     @d@     �d@     �d@     ~e@     �Z@     \_@     ,.@     v.@     Rj@     cj@     �h@     i@     cj@     �j@     �j@     �j@     �j@     m@     m@     m@      m@     �o@     �o@     �o@     �o@     (p@     (p@     Pp@     Pp@     np@     np@     �q@     �q@     �q@     �q@     �r@     ~e@     :f@     :f@     �f@     �f@     �g@     �g@     �h@     i@     �i@     �0@     Q1@     �{@     �{@     �{@     |@     |@     M|@     N|@     �@     �@     .�@     .�@     v�@     v�@     ��@     ��@     ��@     ��@     �@     �@     "�@     ]u@     {u@     "�@     j�@     j�@     ��@     �r@     ]u@     |u@     x@     x@     lx@     lx@     �x@     �x@     z@     z@     E{@     F{@     �{@     �1@     �1@     ��@     ɑ@     ʑ@     j�@     j�@     
�@     
�@     �@     �@     (�@     }�@     ��@     ��@     ��@     (�@     Ȗ@     Ȗ@     h�@     ��@     }�@     ��@     ��@     �3@     95@     h�@     ��@     95@     a5@                     �@     I�@     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     :M@     �M@     �M@     �M@     �M@     �M@     �M@     �M@     �)@     �)@     �)@     �)@     �)@     J*@     J�@     l�@     l�@     ��@     ��@     2�@     �*@     '+@     (+@     3+@     4+@     ]+@     �+@     �+@     �T@     TU@     TU@     QV@     RV@     {V@     2�@     ��@     ��@     s�@     J*@     s*@     t*@     *@     �*@     �*@     �*@     �*@     s�@     ��@     �V@     �V@     ��@     ��@     |V@     �V@     ��@     ��@     ��@     �@     �@     F�@     F�@     x�@     x�@     ��@     ��@     ��@     ��@     ��@     ��@     	�@     �+@     �+@     �+@     �+@     	�@     �@     �@     H�@     H�@     Y�@     Z�@     t�@     �,@     �,@     �,@     %-@     h-@     �-@     DW@     �Z@     �+@     �+@     �+@     C,@     �,@     �,@     t�@     ��@     �Z@     \_@     ��@     ��@     ��@     
�@     
�@     Q�@     R�@     ��@     ��@     ��@     ��@     ��@     .@     ,.@     �a@     .b@     .b@     Ub@     Vb@     c@     c@     �c@     �c@     )d@     *d@     @d@     @d@     �d@     �d@     ~e@     �-@     �-@     ��@     �@     ~e@     :f@     :f@     �f@     �f@     �g@     �g@     �h@     �h@     i@     i@     �i@     �@     >�@     >�@     L�@     �/@     �0@     Rj@     cj@     cj@     �j@     �j@     �j@     �j@     m@     m@     m@      m@     �o@     �o@     �o@     �o@     (p@     (p@     Pp@     Pp@     np@     np@     �q@     �q@     �q@     �q@     �r@     v.@     G/@     L�@     ��@     �r@     ]u@     ]u@     {u@     |u@     x@     x@     lx@     lx@     �x@     �x@     z@     z@     E{@     F{@     �{@     �{@     �{@     �{@     |@     |@     M|@     N|@     �@     �@     .�@     .�@     v�@     v�@     ��@     ��@     ��@     ��@     �@     �@     "�@     "�@     j�@     j�@     ��@     ��@     ��@     ��@     ��@     ��@     }�@     }�@     ��@     ��@     ��@     ��@     ɑ@     ʑ@     j�@     j�@     
�@     
�@     �@     �@     (�@     (�@     Ȗ@     Ȗ@     h�@     �3@     95@     ��@     �@     h�@     ��@     95@     a5@     6@     �6@     �@     A�@     B�@     m�@                     �A     uA     zA     {A                     �A     `A     eA     fA                     A     �A     �A     �A                     �A     �A     �A     �A                     �A     A     �A     �A                     �A     �A     �A     �A                     �A     pA     �A     �A                     pA     �A     �A     �A                     �A     sA     �A     �A                     sA     A     �A     �A                     A     A     �A     �A                     XA     �A     �A     �A                     �A     �A     a"A     d"A                     {A     �A     A"A     D"A                     �A     /A     D"A     G"A                     /A     yA     G"A     J"A                     yA     2A     J"A     M"A                     2A     �A     M"A     P"A                     �A     � A     P"A     Q"A                     "A     A"A     d"A     e"A                     �dA     �eA     �eA     �eA                     �eA     �fA     �fA     �fA                     �fA     �gA     �gA     �gA                     �xA     �yA     �yA     �yA                     �yA     �zA     �zA     �zA                     �zA     �{A     �{A     �{A                     �A     ��A     ��A     ��A                     ��A     ��A     ��A     ��A                     �A     ��A     ��A     �A                     �A     ��A     ��A     ��A                     �A     ��A     ��A     �A                     �A     ��A     ��A     �A                     n�@     w"A     :M@     �M@     �M@     �M@     �M@     �M@     �M@     �M@     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     M@     :M@     �@     �@     x"A     �"A     �"A     �"A     �"A     K#A     L#A     �#A     �#A     �#A     �#A     �#A     �#A     c$A     d$A     �$A     �$A     �$A     �$A     O%A     P%A     �%A     �%A     �%A     �%A     "&A     "&A     +'A     ,'A     x'A     x'A     �'A     �'A     (A     �)@     �)@     �)@     �)@     (A     .(A     �)@     J*@     �V@     �V@     .(A     X(A     X(A     $/A     $/A     N/A     N/A     6A     s�@     ��@     6A     D6A     D6A     =A     �T@     TU@     TU@     QV@     |V@     �V@     �*@     '+@     (+@     3+@     4+@     ]+@     ��@     ��@     �+@     �+@     =A     :=A     :=A     DA     �+@     �+@     �+@     �+@     DA     DA     DA     GDA     HDA     qDA     rDA     �DA     �DA     �DA     �DA     8EA     8EA     IA     IA     7IA     8IA     aIA     bIA     0MA     0MA     aMA     bMA     �MA     �MA     ZQA     �Z@     \_@     �,@     �,@     �,@     %-@     �@     T�@     h-@     �-@     ZQA     �QA     �QA     �QA     �QA     �UA     �UA     �VA     ��@     	�@     �VA     �VA     �VA     �]A     �]A     o^A     p^A     F_A     F_A     `A      `A     �`A     �`A     �aA     �aA     �bA     �bA     [jA     [jA     �jA     ��@     ��@     �jA     �qA     �qA     srA     trA     JsA     JsA     #tA     $tA     �tA     �tA     �uA     �uA     �vA     �vA     _~A     _~A     �~A     �~A     ��A     ��A     w�A     x�A     N�A     N�A     '�A     (�A     ��A     ��A     ׉A     ؉A     ��A     ��A     c�A     c�A     ǒA     �a@     .b@     .b@     Ub@     @d@     �d@     ~e@     :f@     :f@     �f@     �c@     )d@     �f@     �g@     �g@     �h@     �h@     i@     �d@     ~e@     i@     �i@     .@     ,.@     ��@     ��@     ǒA     ��A     ��A     {�A     |�A     R�A     R�A     +�A     ,�A     �A     �A     ۝A     ܝA     ��A     ��A     g�A     g�A     ˦A     ˦A     �A     �A     &�A     &�A     p�A     p�A     ǧA     �@     4�@     v�@     ��@     ȧA     !�A     "�A     4�A     4�A     ӨA     ӨA     (�A     (�A     �A     
�@     Q�@     �A     ֩A     ֩A     u�A     u�A     ʪA     ʪA     !�A     !�A     x�A     x�A     �A     �A     l�A     l�A     ìA     Rj@     cj@     Pp@     np@     �q@     �q@     �r@     ]u@     ]u@     {u@     |u@     x@     �o@     �o@     x@     lx@     *d@     @d@     lx@     �x@     (p@     Pp@     cj@     �j@     �x@     z@     �j@     �j@     z@     E{@     �o@     (p@     np@     �q@     �q@     �r@     F{@     �{@     �/@     �0@     6@     �6@     ��@     �@     ìA     �A     �A     ��A     ��A     �A     �A     e�A     e�A     �A     �A     ��A     ��A     T�A     T�A     ��A     ��@     �@     ��A     ��A     ��A     L�A     L�A     �A     �A     ��A     ��A     ;�A     ;�A     �A     �A     ��A     ��A     *�A     �@     "�@     j�@     ��@     ��@     ��@     ��@     }�@     }�@     ��@     "�@     j�@     ��@     ��@     v�@     ��@     ��@     ��@     �{@     �{@     m@     m@     .�@     v�@     �{@     |@     ��@     �@     ,.@     v.@     *�A     ��A     ��A     z�A     z�A     �A     �A     ��A     95@     a5@     L�@     ��@     h�@     ��@     (�@     Ȗ@     Ȗ@     h�@     �@     (�@     
�@     �@     �@     .�@     |@     M|@     ʑ@     j�@     j�@     
�@     �0@     Q1@     ��@     ��@     �1@     �1@     �3@     95@     ��@     �@                     ��A     4�A     �(@     �(@     4�A     I�A     J�A     v�A     v�A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     N�A     N�A     \�A     \�A     n�A     n�A     ��A     ��A     �A     �A     &�A     &�A     @�A     @�A     d�A     d�A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     ��A                     M�A     x�A     ��A     ��A                     ��A     ��A     ��A     �A     �A     0�A     0�A     @�A     @�A     Q�A     R�A     ��A     ��A     X�A     X�A     ��A     ��A     ��A     ��A     ��A     ��A     5�A     6�A     }�A     ~�A     ��A     ��A     ��A     ��A     	�A     
�A     )�A     *�A     I�A     J�A     i�A     j�A     ��A                     ��A     ��A     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     �)@     �)@     �)@     �)@     �)@     J*@     �*@     '+@     (+@     3+@     4+@     ]+@     �+@     �+@     ^+@     �+@     �+@     �+@     �+@     �+@     �,@     �,@     �,@     %-@     h-@     �-@     %-@     h-@     .@     ,.@     ,.@     v.@     �/@     �0@     �0@     Q1@     �1@     �1@     �3@     95@     95@     a5@     6@     �6@                     @�A     ��A     �(@     �(@     �(@      )@      )@     �)@     �)@     �)@     M@     :M@     �)@     �)@     �)@     �)@     �)@     J*@     J*@     s*@     t*@     *@     �*@     �*@     ��A     ��A     �*@     �*@     �+@     �+@     �+@     �+@     �+@     �+@     �+@     C,@     ��A     ��A     �,@     �,@     �-@     �-@     ��A     m�A     v.@     G/@     m�A     �A     �A     c�A     c�A     �A     95@     a5@     b5@     6@                                                        � @                    @                   Q�A                   `�A                   `�B                   8�B                   8�B                   P�B                  	 `�B                  
 p�B                    �B                   ` C                                                                                                                                                                                                                                             ��                     P�B                 	 `�B             (     `�B             ;     0@             =     `@             P     �@             f     ` C            u     h C            �     0@             �     � C     0           ��                �     X�B             �     0�B             �     �A             �    ��                	     #@                ��                    �@     >       G    7@            `   ��                g   ��                v   ��                �   ��                �   ��                �   ��                �     M"@             �     q"@             �     �"@             �     �"@             �     #@                  #@                  #@            &   ��                /   ��                8   ��                B   ��                L    ��A            _   
 p�B            �    ��A            �    ��A            �   ��                L    �A            _   
 x�B            �    �A            �   ��                �   ��                L    @�A            _   
 ��B            �    R�A            �    S�A                T�A            7    U�A            `    1B            �                   �    �B            �    �B            �    �B            �    �B                 �B                �B            /    �B            D    �B            Z    �B            l    �B                �B            �    �B            �    �B            �    B            �    B            �    B            �    B     	           (B     	       &    8B            D    HB     	       [    �B            �    �B            �    �B                !J@     /       �    PJ@            �   ��                L    �B            _   
 ��B            �    �B                8B            =    @B     	       T    PB     	       k    `B     	       �   ��                �    pB                qB            7    rB            `    �*B            L    �B            _   
 ��B            �    �B            �    �C            �    ��@     �      �    �C             $    �C            O    Z�@     o       o    ɩ@     �       �    ��@     ?      �     +B            %    ի@     r      g    +B            �    "+B            �    )+B            �    0+B            �   ��                	   ��                L    @+B            _   
 ��B            �    R+B            �    S+B                T+B            7    U+B            `    jHB            	    �+B            C	    �C            n	    oHB            �	    tHB            �	    zHB            �	    �HB            @
    �HB            l
    �HB            �
    �HB            �
    �HB                �HB            3    �HB            m    �HB            �     C     x       �    �C     x       �     C     x           ��@            2    ��@            U    ��@     �       x    ��@     �       �    xC            �    ,�@     *       �    V�@            "    v�@            V    +�@     �       �    ��@     *           ��@            F    �@            {    ��@     �       
    �@            a    ��@                A�@     �       �    4�@            �   ��                �    IB                	IB            7    
IB            `    rB            L    eIB            _   
 ��B            �    wIB            �    ;rB                �pB                 �pB            5    �pB     	       L    �pB            b    �pB            w    �pB            �    �pB            �    %�@     �       �    �pB            �    ��@            �    ��@     0            �A     �      1    N�@     b       P    ��@     [       k    �A     �      �    �pB            �    qB            �    qB     	       �    (qB            �    0qB     
           @qB     	       $    PqB     	       ;    `qB            Q    hqB     
       i    xqB     	       �    �qB            �    �qB            �    �qB     	       �    �qB            �    �qB            �    �qB                �qB                �qB            +    �qB            @    �qB            T    �qB            h    �qB     	           �qB            �    �qB     	       �     rB            �    rB            �    rB            �     rB     	           HrB            !    �pB            ~    �pB            �     qB            9    0rB            �   ��                �    @{B            �    H{B     	       �    �C            �    Q{B            �    X{B                `{B            &    h{B            ;    p{B            Q    x{B            g    �{B     	       ~    �{B            �    �{B            �    �{B            �    �{B     	       �    �{B            �    �{B                �{B                �{B            ,    �{B            B    �{B            X    �{B            n    �{B            �    �{B            �    �{B            �    �{B            �     |B            �    |B            �    |B                |B                 |B            g   ��                /   ��                �    (|B                )|B            7    *|B            =    �C            c    �C            �    �C     �      �    �C            �    �C            �    �C            �    �|B            $    �|B            N   ��                L    �|B            _   
 ��B            �    �|B            [    @~B            �    ~B            �    �C            #    �C            V    �C            �    b~B                P~B            �     ~B            !    �}B            �   ��                L    p~B            _   
 ��B            �    �~B            �    �C            �   ��                L    �B            _   
 ��B            �    ��B            �   ��                L     �B            _   
 ��B            �    �B            �    �B                @�A     J       <    ��A            ]    `�@     #       f  "  ,.@     J       �  "  ��A     �       M  "  �@            �    R�A     H       �    Y�@            �  "  �jA     �      6  "  6A     *       p    8�A     �       �    ��A     S       �    �@     �      �  "  �(@     \       �  "  $tA     �       c     ��@     n       �     ��@     >       �   "  �)@     V       �   "  _~A     d       !    ��A     �       0!  "  F�@     2       �!  "  ��A     �      /"  "  v.@     �       v"  "  �+@     4       �"  "  �DA     N       �"  "  Q1@     U       >#  "  (+@            }#    S�@     #       �#     �B            �#    ��A     �       �#  "  �DA     )       �#    ��@     /       �#  "  �#A     &       �#  ! 
 ��B     @       $    H�A     *      $    ��A     3       $     @     (       M$    � C     (       ��    n�@     �       Z$    X C            a$    ��@     �       j$  "  �)@     #       �$    )�A     /       �$  "  �A     �       %  "  �@     R       +%    ��@     7       5%    ��@     �      Y%  "  b�@            �%  "  �+@     4       D�    ��@     I       �%  "  J�@     "       ]&  "  0MA     1       �&  "  *�A            �&  "  |V@     (       �&    ��@     B       �&  "  �q@     7      �'  "  �@     S       (    ~�A     @      (    Y�A     C       /(  "  .@     *       �(  "  DA     1       �(  "  �i@     �       ?)    �@     .       R)  "  �`A     �       �)  "  x"A     &       �)  "  JsA     �       �    i7@     �       y*    ��@     T       �*  "  �f@     D      �*  "  R�@     1       G+  "  ֩A     �       �E    G�@     �       �+  "  x@     d       �+    N$@     >       �+  "  ��A     =       �+  "  (�A     �       w,   ��A     W       �,  "  ��@           
-    ��@     4       -  "  �bA     �      �-  "  
�@     G       �-  "  �V@     +       �-    �A     2       �-  "  �@     -       .    �8@     $       .    ��A            /.  "  
�@     w       �.  "  F{@     K       �.  "  �*@     )       .�    f�@            /  "  P�@            a/    ��A            �/  "  �]A     �       0  "  �+@            *0    G�@     �       10  "  RV@     )       t0    !�A     +       {0    q�@     H       �0  "  �#A     <       �0    �@     :       �0    ,�@     S       �0  "  �!@            �0  "  }�@            �1    ?9@     9       �1    ��@     V       ݰ    B@     +       �1    ��A     2       �1    ��@     S       �1    Ҟ@     S       �1    �?@     �       �1    �@     �      2  "  ��@     V      �2  "  ��@     V      �3  "   )@     �       �3  "  l�A     W       :4  "  �T@     )       �4  "  u�A     U       �4    6�@     3       �4   �%@     c       �4  "  �*@     )       25  "  T�A     �      t5  "  �M@     M      �5    �@@           �5  "  �A             �5    ��A     .       �5  "  �V@     0       6  "  j�@     �      �6  "  ��A     )       G�    ��@     �       A7    ��@     �       G7  "  �-@     *       �7    �@     /       �7    e@     �      �7    ��@     S       �7  "  ��A     �       X8  "  �uA     �       �8  "  �qA     �       U9  "  �DA     N       t9    ��@     �       �9  "  *d@            �9  "  *�A     �      ��    ��@            ":    ��@     �       ?:  "  ��A     +       �:  "  ,�A     �       �:  "  ��A     U       ;;  "  X@     "       Q    7@     Z       X;    �A     !       r;  "  L@     I       �;  "  TU@     �       �;    k�@     �       �;   ` C             �;  ! 
 h�B     @        <  "  ��@     #       �<    �@     5       �<    	�@     z       �<  "  �M@            �<  "  	�@            "=  "  �x@     7      >  	 h�B             >    ��A            ;>  "  ìA     W       x>  "  �+@     ,       �>  "  h-@     &       ?  "  ��@     "       �    p�@     �       �?  "  ȧA     Y       �?  "  d�A     7       @    C            @   a�A     g       (@    ��@     V       0@    ��A            T@    ��@     5       ]@    ��@     Q       e@  "  |u@     �      UA    �A     +       yA  "  Z�@            B  "  bIA     �      fB  "  ��A     {       �B    ˟@     S       �B  "  �A     �       �B  "  ��A     P       TC    �?@     +       [C    ��@            `C  "  x�@            �C    x�@     2        D    ��A     /       D  "  CP@     L      &D    ��A     2       -D    ��@     �       JD  "  �A     �      �D  "  g�A     d       �D    �G@     �       �D    n�@     +       tz    e?@     *       E    %�@     S       E  "  :=A     �      YE  "  4�A            pE    (C            yE  "  �A     �      �E    ��@     �       �E    �:@     +       �E    2�@     u       �E  "  x�A     �       yF  "  l�@     *       �F  "  �'A     O       �F    ��@            �F    ��A     3       �F  "  ��@     *       BG    �:@     G      JG    �B             WG  "  (A            pG  "  ��A     -       �G    Y�A     /       �    ��@     x       �G  "  �@     (       UH  "  j�A            qH  "  �#A     &       �H  "  �VA     �      �H    �?@     +       �H    $�@     ?       I    �@     V       !I  "  IA     1       KI  "  l�@     *       �I    �C            �I  "  ��A     =       �I    E@     .       �I   `%@     6       �I  "  �"A     H       J    |F@     3       
J  "  X@     "       'J  "  @�A     $       �J  "  �)@     V       �J    7@     0       �J  "  t*@            4K  "  �3@     �      �K  "  z@     �       �K  "  ��@     �      `L    �!@     +       �L    �A            �L    �@     V       �L    <�@     /       �L    κ@     /       �L  "  �{@     W       *M    �A     7       2M    Q�@            9M  "  H�@            �M  "  �M@            �M  ! 
 ��B     P       �M  "  >�@            PN  "  t�@     C       �N  "  P%A     S       �N  "  N/A     �      O    f�A     �       -O  "  ��@     1       P  "  �c@     O       AP    �@     /       SP    ?E@     =      \P    ��A            �P  "  x�A     �       �P    �@     �       �P  "  ��@     C       Q    ��A     3       Q  "  �MA     �      lQ  "  "@            sQ  "  L#A     M       �Q  "  m�A     �       R    ��@     7       R  "  �j@     a      S    P?@            S  "  ��@     �      �S  "  m@            �T    b�@     m       �T  "  �Z@     �      �T    C            �T  "  Ĳ@            9U    )�B            IU    �>@     #       OU  "  @     "       hU  "  rDA     N       �U    � C            �U  "  �+@     E       �U    ��A     /       �U  "  @d@     I       )V  "  ��A     
       �V    tA     [       �V    E�@     V       �V    � @             �V  " �%@     ;       �V  "  Rj@            �W  "  ��A            �X    ��A     �       �X  "  �@            xY    x9@     J      Y  "  4�A     �       �Y  "  J�@     "       KZ    ��@     /       SZ    �C     �	      gZ    ��A     /       nZ    �B@           tZ    x�@     S       }Z  "  h�@     1       d[  "  �/@     �       �[    j�@     �       V     �B            �[  "  p^A     �       I\    C            Q\    �C            X\  "  6A     *       �\  "  [jA     d       �\  "  ��A            A]    ��@     �       H]  "  �@     2       \]    F@            w]  "  d�@            �]  "  L�A     �      �]    ]@           �]  "  X�A     7       =^  "  0�@     P       �^  "  ��A     �      �^    ��A     p       �^  "  N�A            &_    x!@     1       I_    O�A     /       P_    i>@     V       W_    d"@             m_  "  ��@            \`  "  :f@     X       >a    C            Ha  "  @�A     $       �a    �8@     3       �a  "  n�A     %       b  "  4K@     �      *b  "  &�A     J       >b  "  ZQA     1       gb  "  fJ@             {b    ��A     f       �b    N8@     -       �b    @ C            ��    �@     �       �b    ��@     P       �b    �@     S       �b  "  d$A     c       �b  "  T�@     *       �b  "  Pp@            �c    ��A     Q       �c    �@     �       
d  "  Z�@            �d  "  ʑ@     �      �e    ��A     ;       �e    �'@           �    ��@     .       �e  "  �%A     .       �e    R�A     �       �e  "  b5@     �       f    y=@     +       f  "  J*@     )       Uf    k�@     /       ]f    @C     (       pf  "  J�A            �f  "  np@     7      zg  "  R�A     �       �g   �%@            h  "  ��A     �      Vh  "  R�A     �      ,%    ��@     x       �h  "  ,'A     L       �h     �@     �       �h    �"@             �h  "  �QA     �      (i  "  $/A     *       ci    E�@     f       ii  "  rDA     N       �i  "  ��A     K      �i  "  ��@     C       Bj  "  J�A     ,       rj  "  ��@            �j  "  �+@            �j  "  ��A            �k    9�@     6       �k    ��@     U       �k    :�@           �k  ! 
 �B     P       l    X�A     /       |b    �A     Y       l    0#@     �       +l  "  ~e@     �       m  "  t*@            Qm   X&@            nm    P C            tm  "  �#A     g       �m  "  �@     2       �m    ��A            �m  "  ;�A     �      n    t�A     �       n  "  *d@            `n  "  
�A            �     @     &       {n    T�@            �n  "  v�A            �n    ��@            �n    ��A     �       �n  "  c�A     �      Eo  "  x@     d       "�    _=@            �o   ��A     f       �o  "  ��@     N       p  "  ��@     �       dp  "  .(A     *       �p  "  �A     W       �p  "  ��@     �      Fq  "  ��A            $r    ��@     .       -r  "  ��@     �      �r    <�A     %       �r    ��@     h       �r    ��@     V       �r  "  �A            s  "  =A     *       =s    a�A     �       Es  "  H@     �       cs  "  ��A     $       	t  "  �R@           't     C            /t    L�A     2       7t  "  "@            ?t    ]@     S       Zt    �A     �       �     ��@     �      bt  "  \�A            �t  "  ��A     $       /u    �C            Mu  "  (�A     W       �u    ��@     E       �u  "  �d@     �       Uv  "  p�A     W       �v  "  ȧA     Y       �v  "  ��A            �w    A     [       �w  "  x'A     S       �w   F&@            �w  "  =A     *       x    ��@     J       x  "  �UA     �       6x    OH@     �       >x  "  �a@     2       kx    hC            wx    |�@     *       �x  "  �@     -       �x  "  ӨA     U       �x    ��A     �       �x    g&@            �x  "  v�@            #y    ~@     "       Hy  "  �T@            �y  "  ��A     �       z  "  �"A     e       *z    r�A     ,       1z  "  d�A     7       qz    ?@     +       ��    X�A     r       z  "  �)@            �z    C            �z  "  �A     �      �z    '�@     �       �z  "  fJ@             �4    ��@     �       �z    �@     '      !{    �@     �       ={    ��@     V       E{  "  �A             p{    ��A     /       x{  "  j�@            a|    ��A     2       i|    ��A     �       q|  "  c@     �       M}  "  ��A            �}  "  ��@     0       0~    p�A     .       7~  "  ��@     3       �~  "  (�@     �      �  "  �@     *       �    �#@     p       �  "  �@     -       �  "  s�@     +       "�  "  �)@            :�    	�@     2       @�  "  X(A     �      ��  "  8EA     �      ߀  "  "�@     H       ΁    ��@     E       ��  "  lx@     j       �    ��@     x       ނ  "  ��A     �       �  "  ��A     E       u�    4=@     +       ~�  "  �-@     J       �  "  ��A     }       V�  "  �vA     �      ��  "  �$A     6       ؄    ��@     E      ބ    ` C             �    F�A     3       �    �@     &       �  "  �@     !       f�    ��@     *       0t    �6@     F       o�  "  ʪA     W       ��  "  v�@            ��    
@     �	      ��    J�@            ��    *�A     /       Æ  "  $/A     *       ��    ��@     ]       �    �A     �       !�    �=@     "       '�    ��A     3       /�  "  ��A            K�    Y�@     3       U�    @�B            b�    �@            l�  "  �M@     B       &r    ��@     �      ��    ��@            ��    L�@     U       ��  "  $"@            ��  "  �(@            ��  "  \�A            �    ��@     �       �  "  &�A            C�    ��@            K�  "  L�@     �       ƈ  "  �@     0       W�  "  ֲ@     4       ��  "  �o@            ��    �C            ��  "  &�A            ��    G�@     V       �    ~�A     3       
�  "  J�A     ,       :�  "  (p@     (       ��    m�@     /       ��    ��@     V       ��  "  �)@     #       ��  "  cj@            ��    v�@     +       L�    i�@     x       ��    I�@     V       ��  "  �@     -       ��  "  �@     -       ��    �@     "       Ռ    ?�A     g       �  "  "�A            �  "  �)@            5�  "  �o@     j       !�    QA     ;      0�  "  �,@     &       q�    ��A     r       x�  "  ��@     r       ��  "  ��A     P       ��  "  �aA     �       v�     �A     �       ��  "  �+@            ��  "  
�@            &�    �@     .       ;�  "  ��A     |       ��  "  �$A     Q       ��    �"@             ��  "  �A     U       �  "  \_@     #      )�    Q�A             /�  "  ��A     �      q�  "  4�A            ��  "  �V@     E       ܑ  "  �~A     �      D�  "  ��@     �       ��    k�@     D       ��  "  N|@     �      4�    ��@     �       3�    o�@     �       ��    ��A     ]       ��    V�@     �      Ó    9@     %       ʓ    �I@     3       ӓ  "  �j@            �x    �>@     )       ��   T�A     .       Ɣ    ��A     m       Δ  "  �@     R       �  "  C,@     C       F�  "  2�@     a       �  "  "&A     	      ��  "  �1@     U       c�    � A     [       m�  "  ��@            �    3�@     S       �  "  �@            �  "  bMA     )       7�  "  �@            H�    ��@     x       �    H C            �  "  D6A     �      l�  "  trA     �       �    �C            �    �=@     Z       
�  "  %-@     C       ]�  "  X�A     7       ��    ��A     R       ��  "  �,@     4       ��  "  DA            0�  "  e�A     �      r�  "  �%A     O       ��  "  F_A     �       �  "  �A            7�    5�@     $       �    ~B@     /       H�  "  c�A     d       �    5�@     +       ��  "  ܝA     �       /�  "  :M@     Q       R�  "  �g@     �       ��  "  �q@            ߝ  "  �%A     .       ��    ��@     "       ��  "  �$A     6       �  "  ��A     P       ��  "  �!@            ��    �A            ��  "  *�@     %       �    �@     >       �  "  |�A     �       ��  "  .�@     H       o�    ��@            ��  "  ��A     P       Ӡ  "  8IA     )       ��  "   m@     �      �    �@     .       �    �@     S       �    y&@           ��    d�@     h       �    �@     I       .�    @     (       Q�  "   )@     �       q�  "  �@     I       Ӣ  "  z�A     �      �    ��@     /       �  "  �(@     \       8�  "  �h@     L       e�  "  6�A     G      �    �A     ;      �    =�A     3       ��  "  HDA     )       !�  "  Ȗ@     �      �    �B@     /       �  "  �a@     2       @�  "  |@     1       �    ��A     3       $�  "  ��A            ��  "  ؉A     �       	�    �@     �       -�    �@     V       5�   M%@            R�    ;�@     2       Y�    ` C             `�  "  �0@     �       ۧ    r&@            ��    �C             ��  "  ��A     X      w�   �A     :       ��  "  �@     -       ��    (�B            ��  "  �@     <      �  "  ��A     �      F�    �@     `       N�  "  M@     6       ��    T�@     R       ��  "  0�@     P       �  "  �r@     a      ڪ  "  :M@     Q       ��    ��@     3       �  "  ��@     �      �  "  �A     W       -�    A     D       <�  "  ��@     (       ��  "  �)@            ��  "  F{@     K       �    ��@     .       ��  "  G/@     �       t�  "  ��@            �  "  �tA     �       zz    6?@            ��  "  �J@     �       ��    �@     �       �    �@     �       �    ��A            4�  "  ��A     �      w�  "  ǒA     �      ߯    R�@     *       �  "  �{@            ��    ��A     �       ܰ    -B@     +       �  "  ��@     1       ��  "  �,@     E       �   ��A     f       0�    ��@     2       7�  "  ��@           c�    ٝ@     S       R    7�@     x       l�    y�A     /       s�  "  ��@     G       ݲ  "  ��A     -       �    {8@     $       #�  "  �QA     )       I�    K�@     K       Q�    G@     �      j�  "  .b@     '       ��    �A            ��    ��@     +       ��  "  ��@     J       +�  "  N�A     �       ��    �@            ��    �A     2       ��  "  �*@     ,       �    ��@     �      �    F @     �       7�  "  @�A            g�  "  4+@     )       ��  "  �A            �    �A     /       �  "  n�A     %       �    (�A     m       �  "  ]u@            �  "  �1@     �      o�  "  �{@            N�  "  6@     �       ��    8@     <       ��  "  �,@     4       ۸  "  ^+@     (       "�  "   `A     �       ��    �C            ��  "  �@     *       ӹ    �@     Q       M�    �@     x       ۹  "  0�A            �    �8@     $       �    ��A           0�  "  �VA     ;       H�  "  !�A     W       ��  "  (+@            ĺ    
�A     3       ̺  "  *@     -      �    XB@     &       �  "  Vb@     �       ް    �A@     *       1�  "  ��A     �      ��    t�A     i       ��   �$@     6       ��  "  ��A     {       �    A�@     %       ��    g@     ,       �  "  s�@     O       �   �$@     �       >�  "  95@     (       X�    @�B            a�  "  a@     }       ͼ    �A     a       �  "  �+@            �    M�@     +       �    ��@     3       �  "  ˦A     J       2�    # A     �       <�    � C            C�    ��@     K       R�    ��A     \       \�  "  .b@     '       ��  "  ��@     �       ڽ  "  ´@     I       *�  "  �A     W       ��  "  .(A     *       ʾ  "  2"@            Ҿ    ��A     �       �    @"@             ��    ��A     �       �     >@     I       &�   
�A     J       :�    %I@     �       I�  "  4�@            n�  "  i@     �       ��  "  B�@     +       Ϳ    pC            տ  "  x"A     &       ��  !  �B             A�  "  z@     7      '�    ��@     E       U�    �C@     1      \�  "  ��@     6       ��  "  �A     �      ��    ��@     }       ��    J�A     n       �  "  ~�@            o�    � @     �       ��  "  DW@     h      ��  "  T�@     *        �    ��@     .       �  "  ~�A           ��    ��@     �      ��  "  �*@     (       ��    �F@     �       ��  "  ��@     0        crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.5415 dtor_idx.5417 frame_dummy object.5427 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/.local/share/lemon/sysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_keymap_us fb.cpp filesystem.cpp graphics.cpp ipc.cpp runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp syscall.c lemon.cpp _ZN3frgL8null_optE _ZN3frg15_to_string_implL12small_digitsE _ZN3frgL6endlogE _ZZN5mlibc17sys_anon_allocateEmPPvE8__func__ ensure.cpp essential.cpp stdlib-stubs.cpp _ZN3frgL9dont_lockE _ZN3frg9_redblack12_GLOBAL__N_1L15enable_checkingE _ZN3frg12_GLOBAL__N_1L15enable_checkingE _ZZN13AllocatorLock4lockEvE8__func__ _ZN12_GLOBAL__N_111mblen_stateE _ZZ6strtolE8__func__ _ZZ6rand_rE8__func__ _ZZ5abortE8__func__ _ZZ13at_quick_exitE8__func__ _ZZ10quick_exitE8__func__ _ZZ6systemE8__func__ _ZZ6mktempE8__func__ _ZZ7bsearchE8__func__ _ZZ3absE8__func__ _ZZ4labsE8__func__ _ZZ5llabsE8__func__ _ZZ4ldivE8__func__ _ZZ5lldivE8__func__ _ZZ5mblenE8__func__ _ZZ6mbtowcE8__func__ _ZZ6wctombE8__func__ _ZZ8mbstowcsE8__func__ _ZZ8wcstombsE8__func__ _ZZ14posix_memalignE8__func__ _ZZ8strtod_lE8__func__ _ZZN5mlibc7strtofpIdEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIfEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIeEET_PKcPPcE8__func__ _GLOBAL__sub_I_stdlib_stubs.cpp ctype-stubs.cpp _ZZN5mlibc20polymorphic_charcode7promoteEcRjE8__func__ _ZZ8iswctypeE8__func__ _ZZ8towlowerE8__func__ _ZZ8towupperE8__func__ environment.cpp _ZN12_GLOBAL__N_117empty_environmentE _ZN12_GLOBAL__N_118find_environ_indexEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_110get_vectorEvE6vector _ZGVZN12_GLOBAL__N_110get_vectorEvE6vector _ZN12_GLOBAL__N_110get_vectorEv _ZN12_GLOBAL__N_113update_vectorEv _ZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcb _ZZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcbE8__func__ _ZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEEE8__func__ _ZZ6getenvE8__func__ _ZZ6putenvE8__func__ _ZZ6setenvE8__func__ errno-stubs.cpp file-io.cpp _ZN5mlibc12_GLOBAL__N_1L24globallyDisableBufferingE _ZN5mlibc12_GLOBAL__N_116global_file_listE _ZZN5mlibc13abstract_file4readEPcmPmE8__func__ _ZZN5mlibc13abstract_file5writeEPKcmPmE8__func__ _ZZN5mlibc13abstract_file5ungetEcE8__func__ _ZZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeEE8__func__ _ZZN5mlibc13abstract_file4seekEliE8__func__ _ZZN5mlibc13abstract_file10_init_typeEvE8__func__ _ZZN5mlibc13abstract_file13_init_bufmodeEvE8__func__ _ZZN5mlibc13abstract_file11_write_backEvE8__func__ _ZZN5mlibc13abstract_file6_resetEvE8__func__ _ZZN5mlibc13abstract_file18_ensure_allocationEvE8__func__ _ZZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeEE8__func__ _ZN12_GLOBAL__N_110stdin_fileE _ZN12_GLOBAL__N_111stdout_fileE _ZN12_GLOBAL__N_111stderr_fileE _ZN12_GLOBAL__N_111stdio_guardC2Ev _ZN12_GLOBAL__N_111stdio_guardC1Ev _ZN12_GLOBAL__N_111stdio_guardD2Ev _ZN12_GLOBAL__N_111stdio_guardD1Ev _ZN12_GLOBAL__N_118global_stdio_guardE _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ5fopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ5fopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ6fdopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ6fdopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZSt7forwardIZ5fopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _ZSt7forwardIZ6fdopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _GLOBAL__sub_I_file_io.cpp stdio-stubs.cpp _ZZN13ResizePrinter6expandEvE8__func__ _ZZ6removeE8__func__ _ZZ6renameE8__func__ _ZZ8renameatE8__func__ _ZZ7tmpfileE8__func__ _ZZ6tmpnamE8__func__ _ZZ7freopenE8__func__ _ZZ6setbufE8__func__ _ZL9store_intPvjy _ZZ5scanfE8__func__ _ZZ6sscanfENUt_10look_aheadEv _ZZ6sscanfENUt_7consumeEv _Z8do_scanfIZ6sscanfEUt_EiRT_PKcP13__va_list_tag _ZZ7vfscanfENUt_10look_aheadEv _ZZ7vfscanfENUt_7consumeEv _Z8do_scanfIZ7vfscanfEUt_EiRT_PKcP13__va_list_tag _ZZ6vscanfE8__func__ _ZZ7vsscanfE8__func__ _ZZ8fwprintfE8__func__ _ZZ7fwscanfE8__func__ _ZZ9vfwprintfE8__func__ _ZZ8vfwscanfE8__func__ _ZZ8swprintfE8__func__ _ZZ7swscanfE8__func__ _ZZ9vswprintfE8__func__ _ZZ8vswscanfE8__func__ _ZZ7wprintfE8__func__ _ZZ6wscanfE8__func__ _ZZ8vwprintfE8__func__ _ZZ7vwscanfE8__func__ _ZZ5fgetsE8__func__ _ZZ6fgetwcE8__func__ _ZZ6fgetwsE8__func__ _ZZ6fputwcE8__func__ _ZZ6fputwsE8__func__ _ZZ5fwideE8__func__ _ZZ5getwcE8__func__ _ZZ8getwcharE8__func__ _ZZ5putwcE8__func__ _ZZ8putwcharE8__func__ _ZZ7ungetwcE8__func__ _ZZ7fgetposE8__func__ _ZZ7fsetposE8__func__ _ZZ8getdelimE8__func__ _ZZ14fgets_unlockedE8__func__ _ZZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ string-stubs.cpp _ZZ7strxfrmE8__func__ _ZZ8strtok_rE8__func__ _ZZ6strtokE5saved _ZZ6wcstodE8__func__ _ZZ6wcstofE8__func__ _ZZ7wcstoldE8__func__ _ZZ6wcstolE8__func__ _ZZ7wcstollE8__func__ _ZZ7wcstoulE8__func__ _ZZ8wcstoullE8__func__ _ZZ6wcscpyE8__func__ _ZZ7wcsncpyE8__func__ _ZZ7wmemcpyE8__func__ _ZZ8wmemmoveE8__func__ _ZZ6wcscatE8__func__ _ZZ7wcsncatE8__func__ _ZZ6wcscmpE8__func__ _ZZ7wcscollE8__func__ _ZZ7wcsncmpE8__func__ _ZZ7wcsxfrmE8__func__ _ZZ7wmemcmpE8__func__ _ZZ6wcschrE8__func__ _ZZ7wcscspnE8__func__ _ZZ7wcspbrkE8__func__ _ZZ7wcsrchrE8__func__ _ZZ6wcsspnE8__func__ _ZZ6wcsstrE8__func__ _ZZ6wcstokE8__func__ _ZZ6wcslenE8__func__ _ZZ7wmemsetE8__func__ allocator.cpp _ZZ12getAllocatorvE16virtualAllocator _ZGVZ12getAllocatorvE16virtualAllocator _ZZ12getAllocatorvE4heap _ZGVZ12getAllocatorvE4heap _ZZ12getAllocatorvE9singleton _ZGVZ12getAllocatorvE9singleton _ZZN16VirtualAllocator3mapEmE8__func__ _ZZN16VirtualAllocator5unmapEmmE8__func__ charcode.cpp _ZZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEEE8__func__ _ZZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEEE8__func__ _ZZN5mlibc16current_charcodeEvE15global_charcode _ZGVZN5mlibc16current_charcodeEvE15global_charcode _ZZN5mlibc22platform_wide_charcodeEvE20global_wide_charcode _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstateE8__func__ charset.cpp _ZZN5mlibc15current_charsetEvE14global_charset debug.cpp guard-abi.cpp _ZN12_GLOBAL__N_15Guard6lockedE _ZN12_GLOBAL__N_15Guard4lockEv _ZN12_GLOBAL__N_15Guard6unlockEv getwchar _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ stpcpy putchar _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13BufferPrinterEC1EPS0_PN3frg9va_structE _ZN5mlibc7charset8to_upperEj strcpy _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN3frg14format_optionsC2Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN5mlibc13abstract_file4tellEPl unsetenv _ZN3frg8optionalIiEC2ERKS1_ _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN5mlibc7charset8is_alnumEj _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ _ZN3frg8optionalIiEC2IRivEEOT_ _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev tmpfile mousePos _ZN5mlibc7charset8is_alphaEj _ZN3frg8optionalIiEaSES1_ vscanf _ZN13BufferPrinterC1EPc _ZTVN5mlibc20polymorphic_charcodeE strtok_r wcstok _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer stdout vsprintf _ZN3frg8optionalIiEC2Ev wcstof _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg17basic_string_viewIcEC2EPKc vswprintf _ZN5mlibc13abstract_file4readEPcmPm _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC1EPS3_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev _ZN11PrintfAgentI13BufferPrinterEclEPKcm _ZN5mlibc8code_seqIwEcvbEv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm ungetc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ _ZN3frg17basic_string_viewIcE10find_firstEcm strerror _ZN5mlibc10sys_accessEPKci _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _Z10lemon_readiPvm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN13StreamPrinterC1EP17__mlibc_file_base _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15_construct_slabEi _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi syscall _ZN5mlibc20polymorphic_charcodeC1Ebb _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN5mlibc8sys_openEPKciPi _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ fileno_unlocked _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg3maxImEERKT_S3_S3_ wcstoull _ZN5mlibc7fd_fileD1Ev atol _ZN5mlibc15current_charsetEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC1ENS3_10frame_typeEmm _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv _ZN5mlibc13wide_charcode7promoteEwRj _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg8optionalIiE13storage_unionC2Ev getenv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv wcslen iswcntrl _ZN13BufferPrinter6appendEc _Z12lemon_map_fbP6FBInfo iswpunct _Znwm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ strtold isblank wcstoll iswalpha iswblank bsearch _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ _ZN3frg14format_optionsC1ERKS0_ _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic vsscanf _ZN5mlibc13sys_clock_getEiPlS0_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZN5mlibc7strtofpIdEET_PKcPPc qsort _ZN5mlibc13utf8_charcode12decode_stateC2Ev wcsrchr _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10reallocateEPvm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ fgets _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ vwprintf _Z13AddNewWindowsv iswxdigit _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg8optionalIiEC1IRivEEOT_ _ZN5mlibc13abstract_file13_init_bufmodeEv _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC2Ev _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic _ZN5mlibc13abstract_fileD2Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic _ZN8ListNodeIP8Window_sEC2Ev _ZN5mlibc9PanicSinkclEPKc _ZplRK8Vector2iS1_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14size_to_bucketEm setvbuf __TMC_END__ _ZTVN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEE _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv renameat perror _ZN3frg10bitop_implImE3clzEm _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ __DTOR_END__ _ZN5mlibc7charset17is_ascii_supersetEv _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ _ZN3frg17basic_string_viewIwEC2EPKw _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC2Ev dragOffset _ZN5mlibc8sys_seekEiliPl islower _ZN5mlibc20polymorphic_charcodeD1Ev __fpurge tolower _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ _ZN5mlibc20polymorphic_charcodeD0Ev _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC2ERS1_ iswlower _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ system feof _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv fgetws wcspbrk _ZN5mlibc7strtofpIfEET_PKcPPc wcstol _ZN5mlibc13abstract_fileD1Ev _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE malloc remove iswspace _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE _ZN13AllocatorLockC2Ev mainFont _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic vsnprintf strtoll _ZN5mlibc13abstract_file18_ensure_allocationEv _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZN13ResizePrinter6appendEPKcm _ZN5mlibc7fd_file2fdEv wcsncmp _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ strtoul __dso_handle _ZN3frg8optionalIiEcvbEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED1Ev wcsstr _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _ZN5mlibc8code_seqIKwEcvbEv _ZN13BufferPrinterC2EPc _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE mktemp _ZN5mlibc13abstract_file5purgeEv ispunct _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC1Ev __mlibc_errno _ZN5mlibc20polymorphic_charcodeC2Ebb wctomb _ZN5mlibc12sys_libc_logEPKc _ZN13StreamPrinter6appendEc wcstombs _ZN8ListNodeIP8Window_sEC1Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ _ZN3frg8optionalIiEC1ERKS1_ _Z10lemon_openPKci _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD1Ev _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic _ZN4ListIP8Window_sE8add_backES1_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE _Z11SendMessagem13ipc_message_t clearerr_unlocked isspace vwscanf _ZN5mlibc13abstract_file7disposeEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic mempcpy fflush _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ _ZN13AllocatorLock6unlockEv _ZTVN5mlibc7fd_fileE _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ _ZN3frg6formatIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN14LimitedPrinter6appendEPKc _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE _ZN5mlibc7charset8is_digitEj _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ _ZN3frg11unique_lockI13AllocatorLockE6unlockEv _Z10lemon_seekili mbstowcs _ZN5mlibc22platform_wide_charcodeEv _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic putenv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED1Ev wmemcpy _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZdlPv _ZN13StreamPrinter6appendEPKcm _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ vswscanf _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ _Exit _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _ZN5mlibc13abstract_file5ungetEc _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8allocateEm drag _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv backgroundColor abort _ZN4ListIP8Window_sEixEj _ZN3frg8optionalIiEC2EOi fb _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ wcscoll _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frame8containsEPv _ZSt4moveIRN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ ftrylockfile isxdigit _init _ZN5mlibc10sys_getpidEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC1Ev _Z12getAllocatorv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ strtol _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC1Ev fsetpos __mlibc_rand_engine wcstod mblen iswprint _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZN5mlibc13abstract_file6_resetEv _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ lastKey active _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE rename _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm _ZNK3frg17basic_string_viewIcE4dataEv _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _Z22RemoveDestroyedWindowsv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1ES5_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic strrchr _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv _Z14ReceiveMessageP13ipc_message_t wcscpy calloc memcpy_sse2_unaligned _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv mouseData _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ strtod _ZN3frg15aligned_storageILm456ELm8EEC1Ev _ZN3frg7mt19937clEv _ZSt4swapIbEvRT_S1_ _ZN11PrintfAgentI13ResizePrinterEclEPKcm _ZN3frg7mt19937C2Ev wmemchr atof environ fputs_unlocked iswgraph _ZN13BufferPrinter6appendEPKcm _ZN3frg17basic_string_viewIcEC1EPKcm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ _ZN16VirtualAllocator3mapEm _Z16memcpy_optimizedPvS_m _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC1ES6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ strcat __ensure_warn _ZN13ResizePrinterC1Ev _ZN5mlibc7charset8is_printEj _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc rand_r _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv vprintf closeButtonSurface _ZN5mlibc8code_seqIcEcvbEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN5mlibc14sys_libc_panicEv _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE _ZN13ResizePrinter6appendEc _ZN5mlibc7fd_file5closeEv memset32_sse2 _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE fseek _ZN3frg8optionalIiEC1EOi _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev _ZN3frg7eternalI16VirtualAllocatorEC1IJEEEDpOT_ _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg8optionalIiE13storage_unionD2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev getdelim _ZN5mlibc7fd_file7io_readEPcmPm _ZN5mlibc13abstract_file4seekEli _ZTVN5mlibc13abstract_fileE wcstold _Z8DrawCharciihhhP7Surface _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev _ZN5mlibc14sys_futex_wakeEPi stdin _ZN13BufferPrinter6appendEPKc _ZN10win_info_tC1Ev _ZN5mlibc8InfoSinkclEPKc _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic _ZN5mlibc7charset8is_spaceEj _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC1Ev _ZN5mlibc8code_seqIjEcvbEv _ZN5mlibc13abstract_file10_init_typeEv _ZN3frg7eternalI16VirtualAllocatorE3getEv ferror strstr _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC1Emmi __cxa_pure_virtual _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZN11PrintfAgentI13StreamPrinterEC1EPS0_PN3frg9va_structE _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev iswctype _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic strcoll _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE isupper _ZN3frg15aligned_storageILm8ELm8EEC1Ev _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE strncmp _ZN4ListIP8Window_sE6get_atEj _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZN5mlibc7strtofpIeEET_PKcPPc library wmemset _ZdlPvm _Z18memset64_optimizedPvmm strncpy _ZN3frg15aligned_storageILm1ELm1EEC2Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ program_invocation_short_name _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic _ZN5mlibc7fd_file7io_seekEliPl _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic _ZN3frg17basic_string_viewIwEC1EPKw _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC1Ev funlockfile _ZN13ResizePrinter6appendEPKc _ZN5mlibc14sys_futex_waitEPii _ZN11PrintfAgentI13ResizePrinterEC1EPS0_PN3frg9va_structE isascii _ZN3frg4swapERNS_8optionalIiEES2_ realloc _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ windowCount towupper _ZN5mlibc7fd_fileD2Ev _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZN5mlibc7charset8is_graphEj __cxa_atexit _ZNK3frg17basic_string_viewIcE4sizeEv _Z8DrawRectiiii10RGBAColourP7Surface _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN13StreamPrinter6appendEPKc strtok _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC1Ev at_quick_exit _ZN3frg8optionalIiED2Ev mouseDown _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic fdopen _ZN3frg7mt19937C1Ev _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface isalpha _ZN5mlibc13utf8_charcode12decode_stateC1Ev wcscspn _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ wcstoul strncat _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEE3getEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ wcschr _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ _ZN3frg10escape_fmtC1EPKvm _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev _ZN3frg3minImEERKT_S3_S3_ _ZN3frg8optionalIiED1Ev fread _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ _ZN5mlibc7fd_fileC1EiPFvPNS_13abstract_fileEE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ strtoull _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN14LimitedPrinterC2EPcm fopen __bss_start wcsncat _Z8DrawRect4Rect10RGBAColourP7Surface _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm putwchar _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ main _ZN5mlibc13abstract_file9_save_posEv wcsspn _ZN11PrintfAgentI14LimitedPrinterEC1EPS0_PN3frg9va_structE ftell _ZN5mlibc7charset8is_lowerEj srand strxfrm _ZN5mlibc8code_seqIKcEcvbEv vfwprintf font_default _Z5floord _ZN13AllocatorLock4lockEv clearerr _ZN5mlibc7fd_file8io_writeEPKcmPm _ZdaPv _ZnwmPv _ZN3frg15aligned_storageILm1ELm1EEC1Ev fclose _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2EPNS_9slab_poolIS1_S2_EE getchar _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv _ZN5mlibc10infoLoggerE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC1EPNS_9slab_poolIS1_S2_EE isgraph wcsncpy _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ fgetpos isalnum _ZN3frg8optionalIiEC1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ tmpnam isprint _ZN4ListIP8Window_sED2Ev _ZN4ListIP8Window_sED1Ev _ZN5mlibc16current_charcodeEv _ZNK3frg17basic_string_viewIwE4sizeEv _ZN3frg14format_optionsD2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ fread_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc strcmp _ZN3frg17basic_string_viewIcE10sub_stringEmm _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC1IJRS2_EEEDpOT_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN5mlibc7charset9is_xdigitEj _ZN3frg8optionalIiE13storage_unionC1Ev _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ _Z11lemon_writeiPKvm _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE _ZN14LimitedPrinter6appendEc memset64_sse2 _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE7reallocEPvm _fini _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic _ZN13AllocatorLockC1Ev _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic fgetc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ strerror_r _ZN5mlibc13abstract_file11_write_backEv strtof strtod_l _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ __cxa_guard_release strcspn _ZN3frg17basic_string_viewIcEC1EPKc _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ _ZN13ResizePrinter6expandEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic flockfile _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ iswdigit _ZN4ListIP8Window_sE10get_lengthEv _ZN11PrintfAgentI13BufferPrinterEclEc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ stderr _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN5mlibc11panicLoggerE srandom _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC1Ev _ZN16VirtualAllocator5unmapEmm _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZN14LimitedPrinter6appendEPKcm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN3frg15aligned_storageILm8ELm8EEC2Ev putchar_unlocked _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg9_redblack11hook_structC2Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ _ZN13ResizePrinterC2Ev fputc _ZN14LimitedPrinterC1EPcm _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _Znam feof_unlocked _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _Z24CreateFramebufferSurface6FBInfoPv _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ getchar_unlocked _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ _ZN11PrintfAgentI14LimitedPrinterEclEc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ fwide iswupper __ensure_fail _ZN5mlibc13abstract_file5flushEv fflush_unlocked _Z13lemon_readdirimP12lemon_dirent _ZN3frg14format_optionsC2ERKS0_ _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic fputws _ZN3frg14format_optionsC1Ev _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate fwrite_unlocked wmemcmp _ZN11PrintfAgentI13StreamPrinterEclEc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ lldiv _ZN3frg11unique_lockI13AllocatorLockEC1ERS1_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ wmemmove _ZSt7forwardIPN3frg9slab_poolI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN5mlibc13abstract_fileC2EPFvPS0_E isdigit _ZN5mlibc13sys_anon_freeEPvm fwrite _edata _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _Z19__mlibc_do_finalizev _end _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _ZN5mlibc9sys_closeEi _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic vfscanf _ZN3frg14format_options15with_conversionENS_17format_conversionE rewind _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ES5_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ _ZN3frg9_redblack11hook_structC1Ev freopen _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic fgetc_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIiEERS4_T_ _ZN3frg14format_optionsD1Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm ungetwc _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg7mt199374seedEj _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc13abstract_fileC1EPFvPS0_E _ZN5mlibc20polymorphic_charcodeD2Ev _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE towlower _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ _ZN5mlibc7charset8is_upperEj llabs _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc9sys_writeEiPKvmPl setbuf _ZN5mlibc20polymorphic_charcode7promoteEcRj iswalnum wcscmp _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev atoi _ZN11PrintfAgentI13ResizePrinterEclEc iscntrl _Z10DrawWindowP8Window_s _ZN3frg11unique_lockI13AllocatorLockED2Ev ferror_unlocked _ZN5mlibc13abstract_fileD0Ev _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ fileno fgets_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE getline _Z10surfacecpyP7SurfaceS0_8Vector2i _ZN5mlibc13utf8_charcode12decode_state6cpointEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ wcscat _ZN3frg15aligned_storageILm456ELm8EEC2Ev strspn _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc strlen _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC1EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ program_invocation_name _ZN3frg10escape_fmtC2EPKvm toupper _ZN5mlibc13utf8_charcode12decode_state8progressEv atoll _ZN5mlibc7charset8is_punctEj _ZN3frg8optionalIiEdeEv _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD1Ev wcsxfrm _ZN4ListIP8Window_sE9remove_atEj _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11_find_frameEm _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE strchr _ZN5mlibc8sys_exitEi _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC1ERS1_ fputs _Z11lemon_closei _ZSt4swapIPcEvRT_S2_ _ZN5mlibc17sys_anon_allocateEmPPv _ZN3frg3maxIiEERKT_S3_S3_ font_old _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN5mlibc8sys_readEiPvmPl _ZN3frg8optionalIiE13storage_unionD1Ev fgetwc vfwscanf _ZSt4swapIiEvRT_S1_ vasprintf fbInfo fputc_unlocked strchrnul _ZN3frg11unique_lockI13AllocatorLockED1Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZdaPvm _ZN5mlibc7charset8is_blankEj memcpy_sse2 _ZN5mlibc7charset8to_lowerEj aligned_alloc __cxa_guard_acquire posix_memalign _ZNK3frg17basic_string_viewIcEeqES1_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE16_construct_largeEm _ZN5mlibc7fd_fileD0Ev windows _ZN13StreamPrinterC2EP17__mlibc_file_base _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10tiny_sizesE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE mbtowc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic vfprintf strpbrk _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEENSt16remove_referenceIT_E4typeEOS7_ _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE4freeEPv _ZN3frg17basic_string_viewIcEC2EPKcm fputwc _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13abstract_file5writeEPKcmPm _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ free _ZN5mlibc18generic_is_controlEj  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .tbss .init_array .ctors .dtors .data.rel.ro .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                � @     �                                     !              @            Q�                            '             Q�A     Q�                                   -             `�A     `�     ��                              5             `�B     `�     �[                             ?            8�B     8�                                   E             8�B     8�                                  Q             P�B     P�                                   X             `�B     `�                                   _             p�B     p�     x                             l              �B      �     `                              r             ` C     `�     `                              w      0               `�     +                             �                      ��     �1                             �                      ["                                   �                      m"     o�                            �                      �     �W                             �                      �Z     �\                            �                      �                                   �      0               �     7)                           �                      K�                                   �                      [�     p6                                                   �	     @h         0                	                      	     �                                                   (C
     �                              