ELF              ��4   `1      4    (  
         � ��%  �%           �%  ��   �                     �   ��U��S��D  ��������P�M  ��������f������fǅ����  fǅ����  �������� f������ǅ����   ��������P�  ���E�fǅd���� fǅf���,fǅ`���  ������f-Lf��b���ǅh���   �E� �E� ��hU�hW���  ���E܃�������P�  ����������   ��������u���   ��������u]�E� �}�~��}�~��}���}���u��}� t����`���P�R  ���E�눃}� t����u��'  ���E�    �h������������Y�����������f�Eڋ�����f�E��EډE��E؉E�}��*����}�� ����}������}������E������}� t���u���  ���E䍐�   ��Rh�   h�   h�   j Pj j �  �� �E䍐�   ��Rj j j jPj j �~  �� �E��   Pj j j j jj j �_  �� �E䍐�   ����Rj j j j jj P�8  �� �E䍐�   ��Rj j j jPjj �  �� �E��   Pj j j jjjj��  �� �E��   �}� t�@   ���   �}� t�@   ���   �}� t�@   ���   PSQRjjjj�  �� �E��   �E�@��j j j RPj�4  �� ����U��S���k  &2  ��h   ���.  ���E�}� u�    �%�E�U�P�E�   �E�P�E��@   �E�]���U��S���  ���1  ���u��u�N  ���E��}� y�    �$���u�u��b������E�}� t�E���    �]���U��S���   m1  �U�R�U���u���!  ����]���U��S���   =1  �U�R�U�U�U��R�u�u���  ����]���U��S���G   1  �} t&�U�R�U�U�U��R�u�u���  �����]���U���   �0  �]Ë$Ë$�U���������0  �E�    ��U�E�ЋU��E��E�;Er�E��U�������q0  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���E������/  �E���E�E���   �E�    ��Ѕ�u��   �E�    ���E����   �E�    �����E䋃   9E�s	��   �E���u��9  ���E��}� u%��h   ��l   ���� ��h   ��l   �    �l�E��     �E��@    �E��U�P��   �E�E��P�E��@   �E��@    �E��@�ƿ    ��(��P� ����(���Q�E��e�[^_]�U��WVS��L�������.  �E�    �E�    �E�    �E�    �E�E��E� �$  �}� u5��h   ��l   ���� ��h   ��l   �  ��j�������  ��`   ��u-���u��K�������`   ��`   ��u��
  �    �{  ��`   �E��E�    ��d   ���C  ��d   �P��d   �@)ЉE��E�    �E����    ;E؉�E��
  ��d   �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ�d   �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u��`   �E��E�    �|  ���u��9������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��0��P� ����0���Q��8��0�x��0��P� 9Ɖ��s�Ɖ���8��0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��0��P� ����0���Q��8��0�x��0��P� 9Ɖ��s�Ɖ���8��0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���O  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    ��0��P� ����0���Q��8��0�x��0��P� 9Ɖ��s�Ɖ���8��0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    ��0��P� ����0���Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u��`   �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������P  �    �e�[^_]�U��WVS��,������â'  �} u#��h   ��l   ���� ��h   ��l   �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx��p   ��t   ���� ��p   ��t   �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��x   ��|   ���� ��x   ��|   �Z  �  �E��@�E���0��P� �M��I�ο    )����0���Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ��`   9E�u�E܋@��`   ��d   9E�u
ǃd       �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋���(��P� �M܋I�ο    )����(���Q�E܋@��P�u��q  ���G��d   ��t=��d   �P��d   �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉�d   ��  �e�[^_]�U��S���k���&%  �U�U�U�U��R���%������E��E��Pj �u��?������E��]���U��S���$������$  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E���   �E���E�E�@=���tz��p   ��t   ���� ��p   ��t   �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��x   ��|   ���� ��x   ��|   �   �    �_�E�@�E�E�;Er�E�U�P�Y   �E�;�O   ���u��������E���u��u�u����������u��������E�]���U������y#  �    ]�U������e#  ��`��  �    ]�U��S������D#  �M�U��j j j QRj���   �� �E�]���U���W���#  �    ]�U��WVS�@����"  �E�]�M�U�u�}�i�[^_]�U��S�������"  �M�U��j j j QRj�������� �E�]���U��S��������"  �U�U�U�U���j j �u��u��uj���j����� ��]���U��S������["  �M�U��j j j QRj���6����� �E�]���U��S���j���%"  �U��j j j j Rj�������� ��]���U��S���8����!  �M�U��j j �uQRj��������� ��]���U��S�������!  �M�U��j j �uQRj�������� ��]���U���������!  �E�������E����	��E����	��E��	ЉE�E�@�E��E�    �E9E�}G�E�    �E9E�}2�U�E�E�@�M�U��Ѝ�    �E�E��E��ƃE�뱐��U��S���,����   �U��j j j j Rj ��������� ��E�]��� U���������   �M�U�E �M�U�E�} y�EE�E    �} y�EE�E    �E������E���	��E�	ЉE�E$�@�E��E�    �E�;E}k�U��EE$�@9�}Y�E�    �E�;E}D�U�E�E$�@9�}2�U��EE$�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��������  �} y�EE�E    �} y�EE�E    �E�������E����	��E��	ЉE�E�@�E��E�    �E�;E}k�U��EE�@9�}Y�E�    �E�;E}D�U�E�E�@9�}2�U��EE�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��� �-����  �E�E�E�E��E��}��E��f�E��m��]��m��E��E�������v�E�����E���U��S��4�7  ���  �U���������P��H����E��Eԃ��d$��$���l��������E��E�    �E�   �E�    �E�;E��   �E�    �E�;E��   �U�E�E�@�������U�E���E�ȉE��U���ЉE�E��E�P�E�����U���ЉE�ЍP�E��E�@�U�������U���ЉE�ЍP�E��E�@�U�������E��F����E�E�E��$�����]��Ë$�U��S������O  ���u���Y������]���U��S���n���)  ���u���3������]���U��S���H���  ���u���A�������]���U��S���!����  ���u����������]���U��S��������  ���u�����������]���U��S��������  ���u����������]���U��S������g  �M�U��j j j QRj���B����� �E�]���U��S���v���1  �U��j j j j Rj!�������� ��]���U��S���D����  �M�U��j j j QRj��������� ��]���U��WVS��,�������  ���u�E������E��h�   �J������Ɖ��    �*   ����V�  ���u��E��U�P�E��U���ֺ   �ǉ��E�@���EЋE�@���EԋUЋE�������P�O������E܋E��Uȉ��   �Ủ��   �UЉ��   �Uԉ��   �U؉��   �U܉��   �E��e�[^_]�U��VS�(������  �E�@��P�������u��t��V�?  ����h�   V��������e�[^]�U��S��������Ï  �E���   �E�@�ЋE�@����Q�M���   RPj j ������ �E�    �E��P�L  ��9E�����t0�U�E��RP�E  �����M���   ��QP�҃��E�뷋E���   �E�@��RP���������]���U��S��$�������  �E�    �E��P��  ��9E�������   �U�E��RP�  ���P�U�P�U�P�U�@�E��U�E9�}Y�U�E9�}O�U�E�E9�~@�U�E�E9�~1�U�E��RP�`  ��������P�҃��E�U􉐤   �	�E��L�����]���U��S���E���   �U���   �ыU��QR���  ��������P�҃���]���U��S�������  �U��R���Y   ���Eƀ�   ��Eƀ�   ��Eƀ�   ��Eƀ�   ���]���U��S������l  �U��R���-   ����]���U������H  �E�     �E�@    �]ÐU��S���i�����   �E� �E�E� ��t���u��N������琋]��ÐU���/����  �E�@]ÐU��������  �E�@9Er	�    � �+�E� �E��E�    �E�;Es�E�� �E��E���E��@��r /menu.txt           zR |�        ���'   A�BG�    8   ���]    A�BD�U��     \   G���\    A�BD�T��     �   ���0    A�BD�h��      �   ����;    A�BD�s��      �   ����C    A�BD�{��     �   ����    A�BL�       ����             ����          4  ����7    A�Bs�     T  ����r    A�Bn� ,   t  ����&   A�BF����A�A�A�   ,   �  ����4   A�BF���'�A�A�A�   ,   �  ����~   A�BF���q�A�A�A�         B���K    A�BD�C��     (  i���f   A�BD�^��   L  ����    A�BP�     l  ����    A�BY�      �  ����6    A�BD�n��     �  ����    A�BP�  (   �  ����*    A�BC���`�A�A�A�     �  ����6    A�BD�n��         ����?    A�BD�w��      D  ����6    A�BD�n��      h  ����2    A�BD�j��      �  ����5    A�BD�m��      �  ����5    A�BD�m��     �  ����    A�B��     �  ����7    A�BD�m��       �����    A�B��    8  m����    A�B��    X  -���Q    A�BM�     x  ^���C   A�BD�;��   �  }���           �  m���&    A�BD�^��      �  o���&    A�BD�^��      �  q���'    A�BD�_��        t���'    A�BD�_��      @  w���'    A�BD�_��      d  z���'    A�BD�_��      �  }���6    A�BD�n��      �  ����2    A�BD�j��      �  ����4    A�BD�l��      �  ����P    A�BD�H�� (     �����    A�BF�����A�A�A�    D  ����(    A�BD�`��  $   h  '���N    A�BB��F�A�A�    �  M����    A�BD����     �  �����    A�BD����     �  ����D    A�BD�|��     �  ,���#    A�B_�        0���9    A�BD�q��     @  F���    A�BQ�     `  <���Q    A�BM�                   GCC: (GNU) 8.2.0                        ��          U�          d�          �          �          ��                                ��~  ��                   ��            ���            ��   @�     '   D�     1   �     <   �     H   H�     W   P�     d   X�     w   -�7     �   d�r     �   օ&    �   ��4    �            ���            ���            ���            ���            ���            ��             ���   �        ��     *  (�     6  �7     H  m�6     g  8�     s  ��2     �  ڒ*     �  ��9   "  �  s�     �  �6     �  `�     �  ��&     �  �5     �  ��9   "  �  0�     �  :�?       y�6       E��     %  ��4    ,  %�     B  h�(   "  Q  ј'     X  ��     }  h�(   "  �  _�     �  ��#   "  �  ��K     �  �P   "  �  �P   "  �  �     �  �5     �  ��      �  ��6     �  ��       ��'       ��f      ��     8  )�     N  	��     l  ��]     s  >�C    �  $��     �  ��N     �  �Q   "  �  ��;     �  �\     �  ��      �  K��     !  �Q     +  �'     2  g�0     9  ՙ4     U  ƒ     c  ��'    i  ��&     o  ҄C     v  ��      }  d�      �  ԜD     �  �     �  ��#   "  �  ��2     �  F�'     �  �   "  ^  0�~     shell.asm main.cpp fileio.c l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 _liballoc.c syscall.c ipc.c filesystem.c graphics.cpp window.cpp _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx l_allocated _Z12GetVideoModev _Z13_CreateWindowP10win_info_t l_max_inuse _Z14_DestroyWindowPv syscall _ZN4ListIP6WidgetED2Ev liballoc_unlock ReceiveMessage _Znwm lemon_read _ZN4ListIP6WidgetED1Ev l_inuse SendMessage lemon_open _Z11PaintWindowP6Window malloc __x86.get_pc_thunk.ax _ZN6WindowD1Ev _ZdlPv _Z15HandleMouseDownP6Window8Vector2i _ZN6WindowD2Ev liballoc_lock _ZN4ListIP6WidgetEC1Ev calloc _ZN6WindowC1Ev _ZN6WindowC2Ev fseek lemon_write liballoc_alloc menuSurface _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx _Z12CreateWindowP10win_info_t fdopen _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window _ZN4ListIP6WidgetEixEj fread fopen __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface _Z5floord _ZdaPv fclose _Z12_PaintWindowPvP7Surface liballoc_free pmain _Znam fwrite _edata _end _Z13HandleMouseUpP6Window windowSurface _ZN4ListIP6WidgetEC2Ev lemon_close _ZdaPvm _ZN4ListIP6WidgetE10get_lengthEv  .symtab .strtab .shstrtab .text .rodata .eh_frame .got.plt .data .bss .comment                                                    ���   �                 !         U�U                    )         d�d  |                 3         ��%                   <         ��%                    B         ���%  l                  G      0       �%                                 &    	             	              ,  �                               1  P                  