ELF          >    � @     @       XC          @ 8  @                   @       @     �      �                              `       `     H
                    �+  �  �     H��    UUH��������7  ����    �H*` H=H*` t�    H��t	�H*` ��f��ff.�     @ �H*` H��H*` H��H��H��?H�H��t�    H��t�H*` ���ff.�     @ �=	)   uwUH�)  H��ATA� ` S� ` H�� ` H��H��H9�s%f.�     H��H��(  A��H��(  H9�r��0����    H��t
�(@ �<���[A\��(  ]��ff.�     @ �    H��tU��*` �(@ H������]����D  ����UH��H�� ��*` �Q  H��(  �(   �p  H�E�H�E��@    H�E��PH�E���f(  ��H�E��P�[(  ��H�E��P�R(  ��H�E��P�@(  ��H�E��P�E�    �&(  �&(  �ЋE�9�vH�(  �E�H�H��  �E����E�    H�E��PH�E��@��9E�}H��'  �E�H�H�� ��E���H�E�@ H�E�H���u�A�    A�    �    �(   �    H���g  H�����AW�B��A��AVAUE��ATU��SH��H��@$` �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�z  _AXA��@�w���A��AV�   ��RD�L$A��   D�D$�F  Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�  XZA���%���A��AVA��   RD�L$�   ��D�D$��  A[XA�������A��AVA��   RD�L$�   ��D�D$�  AYAZA�������A��AVA��   RD�L$�   ��D�D$�w  _AXA�������A��AV�   ��RD�L$A��   D�D$�C  A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃��	  XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_� L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A���$  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�SH���(   �R	  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     H��I��UD�>H�� I�� SE1҉�E����xA��A���yE� 1ۉ���L�A����   �	ǉЁ� �  ����	�	�E��~_;Y}Z��A�\�G�L�@ E��~9�iA9�}1D���fD  �i��9�~�A ��������H�A�<�D9�u�9�t��9q�[]� H���ff.�     �AWAVAUATUS��H���D$PL�l$X��y�1ۅ�y�1�E����E��M�eA��A��A	�E	�D�$��~dA;u}^�D�D�<Lc���D$Hc�H�D$�
���A9m~9A�E A�M�4$������)��Hc�D9�HOT$��L�I�<������;l$u�H��[]A\A]A^A_�ff.�     @ D��SE������AQ��A��P����XZ[�AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*�������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   D�CE9���   D��D��D�\$�UD  D�S L�[G��D��E��G�M��L�KD�A�HE�	D�A�HH�{D�D9�t?D�C����A9�~0���xD�L �HH�H�A��u��9u��?u�D9�u��    D�\$E)�9t$t��9s�>���H��[]A\A]A^A_�ff.�     @ AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�W���XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�����XZD9�u�H��8[]A\A]A^A_Ð�ff.�     @ �NA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      UH��H��H��L��fof H��H����H��]�UH��H��H��L���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo%`@ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo%`@ f��fs�f��f H����H��]Ð�����������                H��H��E1�E1�H�t$1ɿ   H�D$    �  H�D$H���f.�     D  �GP1�S�5�  �����9x  Cq  ��H���  f��H���*` @�X�R  H�     H�@    H�@     �X�@(   H[��     H���*` H��      H��      H�     H���*` ��     H�     H���*` ��      H�     H�y      H�f      H�S      �f.�     AWAVAUI��ATUSH���D  1�H�6  A�   �  M�e 1��  M��t�H�$  H����  H�  I�mHH����  �S�KA�   A��A)�I9���  ��)�L9�v
H��  I��H9�s$H�CH����   �P�HH�É�)�L9�w�H9�r�H�S H���@  H��H)�H��(H9���  H�J�rH��t%H��H)�H��(H)�H9���   H��H�J�rH��uۋCH�D�H)�H)�H9��8  H�CH���t���A��t#D�������H�CH����  H��Q���A��uH�  H����  E1��3���f�D������H�CH���r  H�H���(���H�T$�~D$H�H�L$H�F(H��`�F����D�f�D$D�n�F�H�JH�^�H�H�BA�D$(H��CH���*` L ��u<H���   �F�1���  H��H��[]A\A]A^A_ËP�HH��E1��[����    �   H)�Hƃ�H���D  �P�HH��E1�E1��(���@ H�2H�H(H�JH�P(A�T$(D�`DH�@0    �@@���H�X8D�hHSH���*` L"L�"H���*` L9"LC"H��`H��L�"��uH�ź   �P�1��  �2����   H)�HЃ�H����D���)���H�z  H���V���1�1���  �����H�C(�C@���f��H�C C(A�D$(CH���*` D�cDL D�kHH�[8L� H���*` L9 LC H��`H��L� ��u7H�ݸ   �C�1��t  ����H�C(H�H�S0H�C �C@���H�C(    닸   H)�HÃ�H���ff.�     �H����   SH�G�H��H)�H�� HC�1���  �C�H�s�=���u~�K�H�{�H���*` H��H)
�OH�S�)���H�K؃�(�G�C�ޭ�H��tH�
H�H����   H�QH�W H�+  H��tnH��t�w�Q+Q)�9�}H�=  1�[�   ��H��  ����� ���� t
f=��t<�u�H��  1�[�N  fD  H��  ��    H9=�  H�GtKH9�tVH�H��tH�BH�GH��tH�H���*` �W�wH)�9  1�[��  �H�W �5����    H�a  ��    H�E      � ��SHc�H�������H��t1�1��     � �QH��H9�w�[�ff.�     @ AUATUSH��H��H����  I��H����  H�G�H��H)�H�� HC�1��4  �E�H�U�=����2  D�e�M9��e  1��  L���6���H��I����  H�CI�L$�H9�H�E��H9������  H���v  H��1�H��H��H��H��H��fD  �oD H��H9�u�H��H���H��H��    H��L�H�I�<�H9�t'A��H�W�H��vA�PH���PH��vA�P�PH��H��H��   H��H�4L�$�H�M��t��I��t�V�PI��t�V�PH�������H��H��[]A\A]�f.�     ��H�f  ����� ���� tHf=��tB<�t>1�1���   H��H��[]A\A]��    D�j 1�H���   H��H��[]A\A]�@ H�   �fD  �[���1��l���@ H��H��[]A\A]����fD  H��H��H�4�   1��    ��T H��H9�u������ H�������I��SH��H��H��L��L��L���i[�fD  1��ff.�     f�H��+` �  1�� H��Hc�E1�E1�H�T$1ɿ   ����H�D$H����     1��f.�      H�)  H���t3UH��S�  ` H��D  ��H��H�H���u�H��[]�f.�     ��:����  trsteaf               zR x�        ����"   A�C       �   <   ����R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   �   ����m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        <  ����k       <   P  �����    B�A�D �G0U
 AABI[ AAB   �  ����3    A�q      �  ����           �  �����    G�M��A     �  P���       D   �  L����    B�B�B �B(�A0�A8�FP�8A0A(B BBB$   @  ����     D�LG FAA   H   h  ����Q   B�F�E �H(�G0�A8�GP"8A0A(B BBB   T   �  ����o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T     ����o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB     d  ���       0   x  ����    H�F�E �A(�� ABB     �  ����1    D l    �  ����h    F�a     �  ���v       H   �  �����   B�B�B �E(�A0�A8�DP�
8D0A(B BBBA,   @  ����m   J��
�Hm�[�B
�F    p  $���1    D�l   t   �  H���P   B�B�A �A(�G0_
(D ABBKo
(D ABBHR
(D ABBEd
(D ABBK            ���    D�U          $   ���          8  ���          L  ���(    D c    d  0���                                                                                                                                                                                                                                                                                                                                                                           ��������        ��������                                                                                                                                                                                                                                                                                                               <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o ,             @     "                      ,    �       �@     �                                       �       {         @     "          o   T  int 9  %  U   m   e  h   �   n  {   �   �   -  
�   N  o    �   o   bpp \   H  o   
 �   �   4  w  Q   e   (\  x ;    y 	;   N  ;   �   ;   H  ;   B  
I   ^  	\    

I     	I   G   �   3   �  x 	;    y ;    <   	n  v   
fb 
\  	�*`       �   	�*`     �   �  	�*`       ;   @     "      �~  c   ~  �`a #�  �Xbg (;   �  *;   �@     5       ^  i 
;   �l �@     5       i  
;   �h  	b  	�   N      �@     p@     �  src/gfx/sse2.asm NASM 2.14.02 ��@              %  $ >  $ >   :;9I  :;9   :;9I8   :;9I8  ;   	 I  
4 :;9I?  4 :;9I?  .?:;9I@�B  4 :;9I  4 :;9I  4 :;9I  4 :;9I       %  . @   �     �      /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/lemon /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx  main.cpp    stdint.h   fb.h   surface.h   graphics.h     	@     ��+v��tg�u�u�ut
� t* f" f < u	 � ;
j  t2 t& t < Y	 � ;i� 2 �    '   �       src/gfx/sse2.asm      	�@     !>==?LLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""��     /home/computerfido/Desktop/Lemon/Applications/Init Vector2i vector2i_t surface_t decltype(nullptr) fbSurface unsigned char GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions -fno-rtti fb_info_t long unsigned int short unsigned int mousePos height main.cpp main linePadding fbInfo uint8_t FBInfo long long int depth pitch width short int buffer uint16_t uint32_t long double size                                                   � @                   � @                   @                   @                   (@                     `                    `                     `                  	 `*`                  
                                                                                                                                                                                                     ��                       `                   `             (     (@             ;     � @             =     @             P     P@             f    	 `*`            u    	 h*`            �     �@             �    	 �*`     0           ��                �      `             �     �@             �     �@             �    ��                     � @                ��                   ��                   ��                (   ��                5   ��                F     �@             W     �@             r     @             �     @             �     E@             �     O@             �    `@            �   ��                @   ��                �    �@     h       �    D*`            �    @*`            �   	 +`            �   	  +`               	 �*`               	 �*`            "   	 �*`            5   ��                ?   ��                K   	 �*`            W    `@            i    0@     o      �   	 �*`            �   	 �*`            �    P@            �     @     v       �    �@            O   	 +`            �    �
@     o         	 �*`               H*`                 `             %    �@     �      ,     `             9    p@     1       C   	 �*`            �    � @             F    p@            T     @     k       o    �@     1       v    �@             �    �@             �    0@     R      o    � @            �    �@     (       �    p@     �       �     @     P      �    @	@                 `	@     Q      /    p@     �       K    �@     m       j   	 H*`             v    �@     �       �    @     "      �    @$`            �    �@            �    @             �    @             �    �@            �    @@     3            H*`                	 +`                 �@            0    @ `            9   	 �*`            @    �@             L    �@     �       �    P@     m       crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4699 dtor_idx.4701 frame_dummy object.4711 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp text.cpp font.cpp graphics.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero fb.c allocate_new_page l_pageSize l_pageCount l_memRoot l_bestBet l_warningCount l_errorCount l_possibleOverruns syscall.c _liballoc.c l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos l_max_inuse syscall liballoc_init liballoc_unlock _Z12DrawGradientiiii10RGBAColourS_P7Surface l_inuse __TMC_END__ __DTOR_END__ malloc __dso_handle lemon_map_fb liballoc_lock _Z18memset32_optimizedPvjm calloc memcpy_sse2_unaligned memset32_sse2 _Z8DrawCharciihhhP7Surface liballoc_alloc _Z18memset64_optimizedPvmm realloc _Z8DrawRectiiii10RGBAColourP7Surface _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface main font_default _Z5floord memset64_sse2 _fini liballoc_free _Z24CreateFramebufferSurface6FBInfoPv _edata _end _Z10surfacecpyP7SurfaceS0_8Vector2i font_old fbInfo memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc                                                                                  � @     �                                     !             � @     �       Q                             '             @                                         -             @                                         5             (@     (      x                             ?               `                                           F              `                                          M               `             (
                              S             `*`     H*      �                               X      0               H*      +                             a                      s*      `                              p                      �*                                    �                      �*      �                             �                      �-      -                             �                      �.      I                             �                      81                                    �      0               <1      �                            �                      �2                                                          �2      8
         <                 	                      =      {                                                   �B      �                              