ELF          >    � @     @       ��          @ 8  @                   @       @     A      A                   A      Q@     Q@     p                    �+  �v5  �     H��    UUH��������&
  ����    ��]@ H=�]@ t�    H��t	��]@ ��f��ff.�     @ ��]@ H��]@ H��H��H��?H�H��t�    H��t��]@ ���ff.�     @ �=I\   uwUH�G\  H��ATA�0Q@ S�8Q@ H��0Q@ H��H��H9�s%f.�     H��H�\  A��H�\  H9�r��0����    H��t
��6@ �<���[A\��[  ]��ff.�     @ �    H��tU��]@ ��6@ H������]����D  ����UH��H����^@ ��^@ A�    A�    �    H�ƿ   �s3  H�<\  H�\  H)�H��Hi��  H�\  H)�H�\  H�H�E�H�}��  v[H��[  H�E�H��H���S㥛� H��H��H��H�Ⱥ    H����[  H��[      H��[  H��[  H��[  H��[  ���UH��H��   H�E�A�    A�    �    �    H�ƿ   �2  �E��[  �E�    ��^@ ��  9E�������   �E� �E�    ��[  9E�}kH��`���H���S  �E�Hc�H��`���A�    A�    �    H�ƿ   �.2  H�E�H�E�E��ƿ�^@ �  H� H9E�����t�E���E���E�����t�E��ƿ�^@ �q  ��O  �E��=������UH��H��   H�E�A�    A�    �    �    H�ƿ   �1  �E܉�Z  �E�    ��Z  9E���  �E� H��`���H���f  �E�Hc�H��`���A�    A�    �    H�ƿ   �A1  H�E�H�E��E�    ��^@ �  9E�����t)�E�ƿ�^@ �{  H� H9E�����t�E���E����E�������   ��   �&  H�E�H�E�H��`���H��h���H�PH�HH��p���H��x���H�PH�H H�U�H�M�H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�U؉��   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�E�H�ƿ�^@ ��  ��M  �E��c������UH��AWAVAUATSH��   H�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸ ^@ A�    A�    H�ƿ   �/  ��  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H����  H��@���H�E��@����H��H���H�    ����H!�H	�H��H���H��H�����H�       H	�H��H���H��@���H��H���H��H��H�й ^@ ��H��H���  �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H���?  H��P���H��X���H�    ����H!�H��H��X���H�E��@������H�� H��X�����H	�H��X���H��P���H��X���H��H��H�й ^@ ��H��H���X  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H���{  H��`���H�E��@������H��h���H�    ����H!�H	�H��h���H��h�����H�       H	�H��h���H��`���H��h���H��H��H�й ^@ ��H��H���  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H���  H��p���H��x���H�    ����H!�H��H��x���H�E��@������H�� H��x�����H	�H��x���H��p���H��x���H��H��H�й ^@ ��H��H����  A�    A�*�2   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H����  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A� ^@ D���H��H���Q  H�E����   H�E��@��Ѓ���H�    ����L!�H	�I��H�E����   ����H�� D��H	�I��L����^@ � ^@ �$  H�E����   ����H�E����   ����H�E�H��H��h ^@ A��   A��   ��   H���  H���E�   �E�   H�E�H���   H�E�H��H���  H�E�H�E�H�U�H�� ^@ A�    A�    H���   ��*  H�e�[A\A]A^A_]�UH��H��@  �^@ ��  H��R  H��R  H��H��H��R  H���R  �H��R  f�HH���  H��H�E�H�E�H�H�HH��R  H��R  H�PH�HH��R  H��R  H�@ H��R  ��R  ��R  ��H�H���I  H��R  H�E��PH�E��@�u�h�   A�    A��   �щ¾    �    �M  H��A�    A�    �    �    �    �   �)  H��0���H���
  fǅ4���d fǅ6���d fǅ0���
 fǅ2���
 H��0���H��H�Test WinH�0�@dow ǅ8���    �    �y6@ ��  �E܋Eܺ   �    ���r  H��(����Eܺ    �    ���W  H��(���H�H���5  H�E�H��(���H�MЋE�H�Ή���  H�EЋ@��H��H��H�H��H��H�E�H�H�E���Q     ��Q     ��  ��  H��Q  ��Q  �{Q  H�M�A��^@ I�ȉщ¾    �    ��  H�Eȋ@H�H�U�H��A�    A�    �    H�¿    �5(  H��0���A�    A�    �    �    H�ƿ   �(  ��6@ A�    A�    �    �    H�ƿ   ��'  �    ��6@ �t  �EċEĺ   �H^@ ���  H�fP  H��H�[P  �����WE  ��t,�P  �P  A� ^@ D�;E  �щ¾    �    �  �E�    �zP  9E�}%�E��ƿ�^@ �  H�E�H�E�H���P����E�����D   �Eĺ   �H^@ ���  ��D  ��O  ��Љ�D  ��D  ��O  ��)Љ�D  ��O  ����   ��D  �D  �iO  H��O  )щʉ��   �fD  �PO  H��O  )щʉ��   H��O  ���   ��yH��O  ǀ�       H��O  ���   ��yH��O  ǀ�       ��N  �������5  ��N  �����#  ��N  ��^@ �y  ���E��}� �  �E��ƿ�^@ �l  H�E���C  H�E����   9���  ��C  H�E����   H�E��@���9���  �mC  H�E����   9���  �UC  H�E����   H�E��@���9��l  �E��ƿ�^@ �  H�ƿ�^@ �D  H�E�H��N  �C  H�E����   �P��B  9�|LH�E��@����u>��B  H�E����   )�B  H�E����   )��ȉ�M  ��M  ��M  ��   Hǅ ���   H�E��@����t0��B  H�E����   )ЉE�oB  H�E����   )ЉE��4�RB  H�E����   )Ѓ��E�<B  H�E����   )Ѓ��E��E�H�� H�E�H	�H�����H�E�H�@|H�����H�E�H�@tH�������������� ���������������H���|  H��0�	�m��������L  ����t��L  ��t��L   ��L  ����  �oL  ��������  �]L   �WL   H��L  H����  �UA  H��L  ���   9���  �:A  H��L  ���   H��L  �@���9��j  �A  H��L  ���   9��O  ��@  H�uL  ���   H�hL  �@���9��$  ��@  H�IL  ���   �P��@  9�|H�/L  �@������   Hǅ ���   H�L  �@����t6�w@  H��K  ���   )ЉE�a@  H��K  ���   )ЉE��:�A@  H��K  ���   )Ѓ��E�(@  H��K  ���   )Ѓ��E�E�H�� H�E�H	�H�����H�wK  H�@|H�����H�eK  H�@tH�������������� ���������������H���_  H��0H������H���  H�������%  H������H=�  ��   H=� u�H��J  H����   H������H����   H������H��H��t6H��������H��t'Hǅ ���   H����������`Q@ H�H������"Hǅ ���   H��������`Q@ H�H�����H�kJ  H�@|H�����H�YJ  H�@tH�������������� ���������������H���S  H��0�(H������H��u�����H������H��u�����������������h ^@ j A�    A�    �   �   �    �    �  H���KI  H�H��#����
   H��H���:  H��#���H��h ^@ A��   A��   ��   �    �    H���'  H���5�=  ��=  h ^@ j A�    A��   �   �   ���  H���QH  �OH  ������H�lH  H�E�H�@H��H���  �5=  �u=  A� ^@ D�q=  �   �   ����  �����UH��H���}��u��}�u'�}���  u��^@ �   �@Q@ ��^@ ��@ ��  ���UH����  �   ����]�UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]�UH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H��H�}��u�U�H�E���H���   ��UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H���;  H�E��ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �'
  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H�� H�}�H�E�H� H�E�H�E�@��tH�E�    H���'�������@ L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A����  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�AUI��H��ATA��H	�I��UH��SH��L)�H��H��H���t:��  M��uH��[]A\A]�D  H��I�4H�| L��[]A\A]��  D  �  �ĐSH���(   �  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     US�D$L�T$ ��y�1���y�1�E����E��M�ZA��A��A	�E	�A��   ���~OA;r}I��l��t�D  A�BA��D�ȅ�~9�~���
���A9B~A�E��9�u�9�t	��A9Z�[]�ff.�     D��SE������AQ��A��P�D���XZ[�H��I��H��A��H�� ��H�� ������� AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   �CA9���   D��D��D�\$�NfD  ��L�[�D��    G�L��L�KD��x��E�9E� H�{D�D9�t=�C����9�~0��D�BD�L= �zI�H�A��u��?u�A�8u�D9�u�D  D�\$E)�9t$t��9s�F���H��[]A\A]A^A_��    AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�w���XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_ÐH��H��A��H��APH�� A��H�� ����m���H����     �NH��H�� ��~zAVAUATUS�O��)���~^I��I����E1��f�A�F)�D9�~DA�EB�<#A�~��    A��Hc�A������4�    Hc�I~Hc�Iu�w���E9e�[]A\A]A^���    �NA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      H���   HD��  ff.�     @ ��  ff.�     �  ff.�     �����ff.�     �{  ff.�     �k  ff.�     1��f.�      UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo%0$@ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo%0$@ f��fs�f��f H����H��]Ð�����������                AW�B��A��AVAUE��ATU��SH��H�ÀW@ �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�*���_AXA��@�w���A��AV�   ��RD�L$A��   D�D$�����Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�����XZA���%���A��AVA��   RD�L$�   ��D�D$����A[XA�������A��AVA��   RD�L$�   ��D�D$�\���AYAZA�������A��AVA��   RD�L$�   ��D�D$�'���_AXA�������A��AV�   ��RD�L$A��   D�D$�����A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃�����XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_� H��H��E1�E1�H�t$1ɿ   H�D$    �y  H�D$H���f.�     D  H��H��E1�E1�H�T$1ɿ   �B  �D$H���f�     Hc�E1�E1�1�1ҿ   �  f�     H��H��H��Hc�L�D$H��E1ɿ   ��  �D$H���D  H��H��H��Hc�L�D$H��E1ɿ   �  �D$H���D  H��H��Hc�Hc�L�D$H��E1ɿ   �  H�D$H���@ H��H��E1�Hc�L�D$�!   �d  �D$H���ff.�     H���7���H��H��H���W���H��H���{���ff.�     ����ff.�     H�������1�H���H��1������   ��u��H���D  ������1�H�����H��H��E1�E1�H�T$1ɿ   �  H�D$H����     L�D$(H�L$ H��E1�H�T$�   �  ���~C�F�H�TA��A��A�A����~$1��    �
�4H��@�r�H��A9���@ H���� H��SHc�H��   H��tT@ H���H��H��	~+��W�T�H��H��u�Hc�H��� �l���H��[��    ��0�T�H��H��u���fD  �0   f�H��[�f.�     ��GP1�S�5x3  �����9h3  Ca3  ��H����  f��H�� _@ @�X�B3  H�     H�@    H�@     �X�@(   H[��     H�� _@ H��4      H��4      H�     H���^@ ��2     H�     H���^@ ��2      H�     H�I4      H�64      H�#4      �f.�     AWAVAUI��ATUSH���D  1�H�4  A�   ��
  M�e 1��
  M��t�H��3  H����  H��3  I�mHH����  �S�KA�   A��A)�I9���  ��)�L9�v
H��3  I��H9�s$H�CH����   �P�HH�É�)�L9�w�H9�r�H�S H���@  H��H)�H��(H9���  H�J�rH��t%H��H)�H��(H)�H9���   H��H�J�rH��uۋCH�D�H)�H)�H9��8  H�CH���t���A��t#D�������H�CH����  H��Q���A��uH��2  H����  E1��3���f�D������H�CH���r  H�H���(���H�T$�~D$H�H�L$H�F(H��`�F����D�f�D$D�n�F�H�JH�^�H�H�BA�D$(H��CH���^@ L ��u<H���   �F�1���  H��H��[]A\A]A^A_ËP�HH��E1��[����    �   H)�Hƃ�H���D  �P�HH��E1�E1��(���@ H�2H�H(H�JH�P(A�T$(D�`DH�@0    �@@���H�X8D�hHSH���^@ L"L�"H���^@ L9"LC"H��`H��L�"��uH�ź   �P�1��)  �2����   H)�HЃ�H����D���)���H�J1  H���V���1�1���  �����H�C(�C@���f��H�C C(A�D$(CH���^@ D�cDL D�kHH�[8L� H���^@ L9 LC H��`H��L� ��u7H�ݸ   �C�1��  ����H�C(H�H�S0H�C �C@���H�C(    닸   H)�HÃ�H���ff.�     �H����   SH�G�H��H)�H�� HC�1��  �C�H�s�=���u~�K�H�{�H���^@ H��H)
�OH�S�)���H�K؃�(�G�C�ޭ�H��tH�
H�H����   H�QH�W H��/  H��tnH��t�w�Q+Q)�9�}H�=�/  1�[�   ��H��/  ����� ���� t
f=��t<�u�H��/  1�[�^  fD  H��/  ��    H9=�/  H�GtKH9�tVH�H��tH�BH�GH��tH�H�� _@ �W�wH)�I  1�[�  �H�W �5����    H�1/  ��    H�/      � ��SHc�H�������H��t1�1��     � �QH��H9�w�[�ff.�     @ AUATUSH��H��H����  I��H����  H�G�H��H)�H�� HC�1��D  �E�H�U�=����2  D�e�M9��e  1��.  L���6���H��I����  H�CI�L$�H9�H�E��H9������  H���v  H��1�H��H��H��H��H��fD  �oD H��H9�u�H��H���H��H��    H��L�H�I�<�H9�t'A��H�W�H��vA�PH���PH��vA�P�PH��H��H��   H��H�4L�$�H�M��t��I��t�V�PI��t�V�PH�������H��H��[]A\A]�f.�     ��H�6-  ����� ���� tHf=��tB<�t>1�1���  H��H��[]A\A]��    D�j 1�H����  H��H��[]A\A]�@ H��,  �fD  �[���1��l���@ H��H��[]A\A]����fD  H��H��H�4�   1��    ��T H��H9�u������ H�������H��L�B�H����   I����   �t$�I��H��I���I�fnD$�f`�fa�fp� f�H��L9�u�H��H���H�8I)�H9���   @�1M����   @�qI��t|@�qI��tr@�qI��th@�qI��t^@�qI��tT@�qI��tJ@�qI��t@@�qI��t6@�q	I��	t,@�q
I��
t"@�qI��t@�qI��t@�qI��t@�q�H���e���ÐH��H���  H�NL�B�H9�H�H@��H9���@���   I����   M��1�I��I��L��H��H���oH��H9�u�M��I���J�<�    H�>H�M9�tH�	H�I����J��   H�H�H��v�>H��H��H���y�H��t)�<@�<H��H��tD�D�D�D�H��t�V�Q�f�L��H��L��   1��    H�<H�<H��L9�u��u���f�H���ff.�     H��t#�H�9�u��    �9�tH��H9�u���    H���ff.�     �H��t*D��A8�u'1�� D��A8�uH��H9�u�1��fD  1�A8�������)���    AU1�I��ATI��H��UH��SH������H��L��Hc�H���"���H��H��L������H��1��
���H��L��[]A\A]�f.�     f�I��SH��H��H��L��L��L���i[�fD  1��ff.�     f�H��0_@ �  1�� H��Hc�E1�E1�H�T$1ɿ   ����H�D$H����     1��f.�      H��  H���t3UH��S� Q@ H��D  ��H��H�H���u�H��[]�f.�     �������  /close.bmp /shell.lef /dev/mouse0             zR x�        ����I    A�CD     <   -����    A�C�     \   ����2    A�Cm      |   ����   A�C    �   �����   A�C� (   �   b���:   A�CP�����%     �   p���   A�C        4���-    A�Ch      $  B���    A�CL      D  4���"    A�C]      d  6���-   A�C(    �  D���"    A�C]       �  F����    A�CE��      �  �����    A�C�     �  ����>    A�Cy        8���8    A�Cs       (  ����    A�CP          L  0���k       <   `  �����    B�A�D �G0U
 AABI[ AABH   �  ���o    B�H�K �D(�M0V
(A ABBFD
(M ABBJ   �  @���3    A�q        d���             p����    A�A��A  $   @  ����     D�LG FAA      h  ����       H   |  ����I   B�F�E �H(�G0�A8�GP8A0A(B BBB   T   �  ����o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T      ���o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB     x  $���(    DK X  <   �  8����    P�B�B �A(�A0�j(A BBBA�����4   �  �����    H�F�E �A(�� ABB            ���             ,���          4  (���          H  $���          \   ���          p  ���          �  ���           �   �   ���R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   D  ����m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        �  ����1    D l    �  ����'    D b    �  ���          �  ���+    D f    �  4���+    D f      L���,    D g    (  d���%    D `    @  |���    DI    X  t���    DI    p  l���          �  h���          �  d���    DK     �  \���0    DV
FM          �  h���(    D c    �  ����                ����M             ����u    D�D
Hd       <   ���h    F�a     X  t���v       H   l  �����   B�B�B �E(�A0�A8�DP�
8D0A(B BBBA,   �  D���m   J��
�Hm�[�B
�F    �  ����1    D�l   t   	  ����P   B�B�A �A(�G0_
(D ABBKo
(D ABBHR
(D ABBEd
(D ABBK         |	  �����          �	  l���         �	  x���4          �	  ����I       4   �	  ����T    B�G�G �D(�D0r(D ABB    
  ���    D�U          $
  ���          8
  ���          L
   ���(    D c    d
  ���           L@     ��������        ��������                                               1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             @     T      a@     I       �@     2       �@     -       
@            @     "       >@     -      l@     "       �@     �       \@     �       �@     8                       ,    �       P#@     �                                       �       �  �  �                  b  
5   �  �    O   int O     a  n   �    �   �     �   T  G   �   O     �   ;  
�   �  �    �  �   bpp u   �  �   
 K  �      ��     v  	)  Y  (�  x O    y 	O   �  O   �  O   �  O   �  
b   m  	�  8  

b     
b   	  '  �  �  x 	O    y O    d  	�  �  D    r b    g b   b b   a b    �  �  "z  h  �  #h   �  $�   �  %�   �  &�   
 x  x  �    �  |  '&  ()�  (  �  *�    �  +
C   �  ,
C   �   -u   bpp .u   |  /�   �  0�   �  1
C   �  2
C   :  3�    o  4�   $ �  5�  �   	@  
�  |�  �  x u    y u   �  u   �  u   �  �   P   �  (  �   l  4  t�  D  �      x  �  �   _ �  H  �  
�  �  �  
  
�  "  
  �  
  (�   s  �  �      �   msg �   �  �   D  �     �   $  O   �  �    T    	`Q@     q  �<�    =4   ?  >�  pos ?�  ��  @�  �   fb C
�  	 ^@     o  D�   	^@     |  E�  	 ^@     )   ?  �      G/  	H^@     �  H�  	`S@         I�  	K^@     �  J�  	L^@     �   K�  	P^@     U  M�  	hS@     O  Ox  	X^@     1  T  	`^@     �  V
�   	h^@     �   W
�   	p^@     �  YO   	x^@     �  [
�   	�^@     �  \
�   	�^@     �  j  	iS@     8  k�  	�^@     p  mO   	�^@       b  �  V   �  �  b   �  �  �  �  b  O    �  !�  �    b   �  *%     "  b  m     ;J  7  B  b  m   M  L�  m  [  f  b  �    �  PQ  m    �  b  �    �  Zt  �  �  b  �   m   4  dm  O   �  �  b   �  h
  m  �  �  b  �    0  }�  m      b     ��  m  *  0  b     ��   �  ��  num ��   T m   
�  b  
�  �  �  �   	�   J  
�  obj m  �  �  �  �  �   T m   
s  �  t  n�  	�^@     �  om  	�^@       @  E  L@            ��  /	  P	   X  h   
   V   !"�  �    #!	  �  s	  �@     8       ��	  $/	  �X%A	  �	  &B	   'A	  �@     )       (B	  �h  )o   @     >       ��	  *�  vO   �l*�  vO   �h +f  
  \@     �       �N
  ,X  h  �X-pos P�   �T.   S�  �h/�@     8       0i U�   �d  1  m
  �@     �       ��
  ,X  h  �H-obj *m  �@.�  +�  �X 2�  �
  �
   X  �   3�
    �
  l@     "       ��
  $�
  �h 1�  �
  >@     -      �|  ,X  h  �H-pos h�   �D.   n�  �h0obj rm  �X4d@     	       \  .+  jm  �P /x@     8       0i p�   �d  1B  �  @     "       ��  ,X  h  �h-pos L�   �d +�  �  
@            ��  ,X  h  �h �  �  �   X  h   3�  �    �@     -       �'  $�  �h 5  �O   �
@           �$  .W  �B  �P.�   ��  ��~.9  �O   �L.  ��   ��~.]  ��  �@.(  �$  ��.�  �O   ��/�@           6msg Is  ��}7+  h*  ��~4A@     7       .  0i �O   �l/S@            0win �m  ��  4�@           �  6i O   �h/�@     �      6win m  ��/�@     �       7  s  ��}7  �   �d7-  �   �`   4�@     �       �  7  7s  ��}7  9�   �\7-  :�   �X /@     �       7>  Ns  ��}   
(  x  :  �    8i  �a  �@     :      �}  -win �m  ��~.$  ��  �� 8�  �%  �@     �      �R  .o  �O   �L/@     �      0j �
O   �l/1@     �      .X  ��  �k.�  ��  ��~.�  �4  �X4w@     D       .  0i �O   �d /�@     �       0win �m  �P    8�   q.  �@           �  .o  rO   �T/@     �       0i u
O   �l/2@     �       .X  v	�  �k/6@     }       0j wO   �d/H@     e       .�  x�  ��~.�  y4  �X     
�    2�  0  :   X     3  %  ]  �@     2       �f  $0  �h 8�  ^�  @     �       ��  .B  `�   �h 9G    �  a@     I       ��  -l 0�  �h-r E�  �` :�   N    t  P#@     @$@       src/gfx/sse2.asm NASM 2.14.02 �P#@              %U   :;9I  $ >  $ >  & I  :;9   :;9I8   :;9I8  	;   
 I  :;9n  I  ! I/     .?n4<d   I4   <  4 :;9I?<  4 :;9I?  4 :;9I?  :;9  .?:;9n2<d   I  .?:;9nI2<d   :;9I82   :;9I82  / I  .?n42<d  4 I?4<  . 4@�B  .Gd     I4  !  "4 :;9I  #.1nd@�B  $ 1  %1  &4 1  '1  (4 1  ).4@�B  * :;9I  +.Gd@�B  , I4  - :;9I  .4 :;9I  /  04 :;9I  1.Gd@�B  2.G:;9d   3.1nd@�B  4  5.?:;9I@�B  64 :;9I  74 :;9I  8.?:;9n@�B  9.?:;9nI@�B  : I   %  . @      �  �      /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx/window /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/lemon /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include  graphics.h   main.cpp    window.h   list.h   stdint.h   fb.h   stddef.h   surface.h   types.h   stdio.h   ipc.h    G 	a@     
�ff!.  tt!.�  	@     � 	�2(K�d�tu�'t��g���
<	�'
�' t �	�K t��+��<tKxfftK� ot�>	�'
� t�K
�+�( t ���<tKK +mt%����'��= jt�>vt<ZK
�H<
t&$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�XK�k�<B0B�4�B �<RJ�>�P.<_Ja�<8�:�<(.*�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9%������ �)!D<u/>Y�vT���.��u\,	tD.	J�*(!@![�, t � / �kv>f��f���u,fftJg,fftJg�& J( t��& J( t�tf � ��"u%�* f�/f�, �9 fG �; �  .Y �f fM �t �� f� �� �h .���u�<f5 J; t& <K+f �7.Df9�J�trX�t<K'f�J='f�JZ'f�)J<='f�)J<">4<;tf6u�u6 g.�� J	�w  �" t f�	u*ut �* f �8 �H fY �J �, .k �{ f_ �� �� f� �� �} .�!u�<f: J@ �( <���<K)f�J=)f�JZ)f�+J<=)f�+J<! >3 <: t f8 u � u9���t � t�tJ" X' t <Y$�)t/<��$�(t�.v�u90tg\+tgZy.mh X0�7C4RfIfY<<4.t��*[� f�}���<J  	�@     �*  	�@     ����  	
@     � 
�u  	@     � �  	>@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K  	l@     �  	�@     )�#���tY��Y����  	\@     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	�@     �	 � t J / �    '   �       src/gfx/sse2.asm      	P#@     !>==ALLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""��            mouseDown __in_chrg size_t uintptr_t _ZN4ListIP8Window_sE8add_backES1_ uint64_t title _ZN4ListIP8Window_sEC4Ev __static_initialization_and_destruction_0 dragOffset testWindow handle_t lastUptimeMilliseconds 13ipc_message_t colourPlanes next RemoveDestroyedWindows long long int mouseEventMessage closeInfoHeader closeButtonSurface fb_info_t redrawWindowDecorations _ZN4ListIP8Window_sE10get_lengthEv mouseDevice Vector2i lastUptimeSeconds active remove_at _ZN4ListIP8Window_sE9get_frontEv stdin _ZN8ListNodeIP8Window_sEC4Ev List<Window_s*> uint16_t _Z13AddNewWindowsv linePadding _ZN10win_info_tC4Ev this closeButtonBuffer _windowCount compression _Z15UpdateFrameRatev currentUptimeSeconds GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions reserved __initialize_p _ZN4ListIP8Window_sE9remove_atEj temp get_front colourNum RGBAColour long unsigned int _Z10DrawWindowP8Window_s 20bitmap_file_header_t width data size short unsigned int AddNewWindows UpdateFrameRate depth _ZN4ListIP8Window_sE8get_backEv _ZN4ListIP8Window_sEC2Ev recieverPID bool stdout decltype(nullptr) FBInfo difference operator[] windowFound vector2i_t fbInfo long double windowInfo 20bitmap_info_header_t pitch /home/computerfido/Desktop/Lemon/Applications/Init frameRate _ZN4ListIP8Window_sEixEj current _ZN8ListNodeIP8Window_sEC2Ev _ZN10win_info_tC2Ev closeButtonFd operator+ _ZN4ListIP8Window_sE6get_atEj importantColours unsigned char node _ZN4ListIP8Window_sED2Ev short int magic main.cpp 10win_info_t vres currentUptimeMilliseconds clear ListNode uint32_t surface_t mouseX _ZplRK8Vector2iS1_ mouseY get_length info data2 _ZN4ListIP8Window_sE9add_frontES1_ buffer _ZN4ListIP8Window_sE10replace_atEjS1_ _ZN4ListIP8Window_sE5clearEv hdrSize offset add_back drag IOFILE replace_at get_at stderr ListNode<Window_s*> closeButtonLength add_front renderPos _Z22RemoveDestroyedWindowsv prev lastKey fbSurface uint8_t DrawWindow windows renderBuffer flags windowHandle hres backgroundColor senderPID _ZN4ListIP8Window_sED4Ev mousePos ~List height rgba_colour_t __priority main mouseData __dso_handle get_back ownerPID frameCounter keyMsg _GLOBAL__sub_I_keymap_us                 @     a@     a@     �@     �@     �@     �@     	@     
@     @     @     >@     >@     k@     l@     �@     �@     \@     \@     �@     �@     @                                                         � @                   � @                   q6@                   y6@                   �6@                   Q@                    Q@                   0Q@                  	 @Q@                  
 �]@                                                                                                                                                                                                                                             ��                      Q@                  0Q@             (     �6@             ;     � @             =     @             P     P@             f    
 �]@            u    
 �]@            �     �@             �    
 �]@     0           ��                �     (Q@             �     A@             �     06@             �    ��                �    ��                     � @                ��                #    @     >       S    L@            l   ��                x   ��                �     ]#@             �     �#@             �     �#@             �     �#@             �     $@             �     $@             �    0$@               ��                   ��                   ��                   ��                +   ��                1   ��                �   ��                8     *@     h       J   	 �]@            U   	 �]@            a   
 (_@            k   
  _@            u   
 _@            �   
 _@            �   
 _@            �   ��                �   ��                �   ��                �   
  _@            �    � @             �    �@     o         	 `S@                @!@     (       T   
  ^@     (       a   
 �^@            m    P5@     T       u    �5@            }    0)@     M       �   
 `^@            �    p*@     v       �    �5@            �   
 p^@            �    �(@     (       c   
 0_@            �  "  �"@            �    �'@     +       �    `@     o          �@     �      &  "  l@     "       C    �3@           J  "  a@     I       ]   
 �^@            e  	 �]@             q    )@            }   8Q@             �   
 P^@            �    P'@     '       �    �*@     �      �  	 @Q@             �    �)@     u       �   
 �^@            �  "  l@     "       �  "  �@     �           '@     1           �(@            %  "   #@            ,   
 L^@            1   	 iS@            A  "  @     "          
  ^@            �    � @             Z    �5@            b   	 `Q@            h   
 X^@            p   
 �^@            w  "  �@     2       �     @     k       �    �@           �    0@     1       �    t#@             �   
 x^@            �   
 H^@            4    p(@            �    `@     o          
 �^@     (            �#@             .    �'@     +       :    �4@     4       A    @$@     R      \  "  �@     2       p   
 �^@            �    � @            �    `(@            �  "  \@     �       �    �5@     (       �  "  #@            �    �@     �       �    P0@     P      �   
 �^@            �    @#@            �    �@                  5@     I       "   
 K^@            ,    @     I      O    0@     �       k    �&@     m       �  "  �@     -       �   
 h^@            �   
 �]@             �    �@            �    �2@     �       �    �
@           �   	 �W@                 @            
  "   #@              "  �@     8       *  "  �@     8       C    �#@             Q    q6@             W  "  
@            z    @     �       �     6@            �  "  �"@            �    �@     3       �    �(@     0       �   	 �]@             �   
 8_@             �  "  �@     -       �   	 hS@            	     (@     ,       	    �@     :      1	    p!@     �       �    �(@            U	    �'@            a	  "  >@     -      �	   	 �S@            �	   
 ^@            �	  "  0#@            �	    0(@     %       �	    P#@             [	    �(@            �	   
 �^@            �	     "@     �       �    �.@     m       crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4699 dtor_idx.4701 frame_dummy object.4711 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux graphics.cpp /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_keymap_us runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp fb.c filesystem.c ipc.c itoa.c allocate_new_page l_pageSize l_pageCount l_memRoot l_bestBet l_warningCount l_errorCount l_possibleOverruns memory.c syscall.c _liballoc.c l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer l_max_inuse memmove syscall reverse frameCounter liballoc_init liballoc_unlock lastUptimeMilliseconds ReceiveMessage _Znwm lemon_read _Z12DrawGradientiiii10RGBAColourS_P7Surface _Z13AddNewWindowsv _ZN8ListNodeIP8Window_sEC2Ev memcpy _ZplRK8Vector2iS1_ l_inuse __TMC_END__ SendMessage __DTOR_END__ dragOffset lemon_open malloc __dso_handle itoa currentUptimeMilliseconds _ZN8ListNodeIP8Window_sEC1Ev _ZN4ListIP8Window_sE8add_backES1_ lemon_map_fb lseek _ZdlPv drag backgroundColor _ZN4ListIP8Window_sEixEj liballoc_lock lastKey active _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm _Z22RemoveDestroyedWindowsv calloc memcpy_sse2_unaligned frameRate mouseData _Z16memcpy_optimizedPvS_m closeButtonSurface memset32_sse2 lemon_write memchr _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev currentUptimeSeconds _ZN4ListIP8Window_sE6get_atEj liballoc_alloc _ZdlPvm _Z18memset64_optimizedPvmm realloc windowCount __cxa_atexit _Z8DrawRectiiii10RGBAColourP7Surface memcmp mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main font_default _Z5floord _ZdaPv _ZN4ListIP8Window_sED2Ev _ZN4ListIP8Window_sED1Ev memset64_sse2 _fini _ZN4ListIP8Window_sE10get_lengthEv _Z15UpdateFrameRatev liballoc_free _Znam _Z24CreateFramebufferSurface6FBInfoPv access _edata _end _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close _ZN4ListIP8Window_sE9remove_atEj font_old fbInfo _ZdaPvm lemon_readdir memcpy_sse2 windows _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                � @     �                                     !             � @     �       �5                             '             q6@     q6                                    -             y6@     y6      "                              5             �6@     �6      x
                             ?             Q@     A                                   K              Q@      A                                    R             0Q@     0A                                    Y             @Q@     @A      H                              _             �]@     �M      �                              d      0               �M      +                             m                      �M                                    |                      �N                                    �                      �N      2                             �                      �_      �                             �                      �c      �                             �                      0o                                    �      0               4o      ^                            �                      �w                                    �                      �w      �                                                    hx      X         E                 	                      ��      �	                                                   ��      �                              