ELF              ��4   �      4    (           � �x\  x\            `   � ��
  �        �W  ��?  �                 �    UU���*  VW�����_^�g  �    �i���f�f�f�f�f����=��t$�    ��tU���h���Ѓ��Í�&    f�Í�&    ��&    ����-�����������t(�    ��tU���Ph���҃��Í�&    �t& �Í�&    ��&    ��=�� ugU�����V��S���������9�s�v ����������9�r��'����    ��t��h���Q~��������e�[^]�Í�&    ��&    ��    ��t'U���h��h���~������	�����&    f������U��S��   ������L���Pj R��9  ���E��E�    �E�    �E�    �}� ��  �E����EԋE���E��E�`   �E�H   ��hp  �f  ���Ã��u��u��u��uԍ�L�����PS�\  �� �]�E�ƀ�   /�E�ƀ�    �E��   ����L�����RP�=4  ���E��   ��P��2  ���P��E����   <fuy�E��   ��P�2  ���P��E����   <euS�E��   ��P�2  ���P��E����   <lu-�E��   ��P�g2  ���P��E����   <.u�   ��    ��t�E��@a�E�ǀ�      �EЃ�u�E�ǀ�      ����P�u���"  ���E��E���у���L���RPQ�58  ���E�E�d�E��Pc�$���9��F����E�L�E�    �6�����]��ÍL$����q�U��VSQ��<�ȋ �E�f�$��f�&��f� �2 f�"�2 �(�    �,�File�0� Man�4�ager�8� ��h ��s  ������j h���L6  ������h��h���#  ���E���u��$  ���E����u���&  ��� �� ��u�j�u�P�5#  �����u���"  ����h��h���"  ���E���u��#  ���E����u��&  �������u�j�u�P��"  �����u��"  ����h��h���B"  ���E���u��A#  ���E����u��0&  �������u�j�u�P�u"  �����u��7"  ���4������E�P�7  ����������   �EЃ�u��y�EЃ�u����P��  ��뾋EЃ�u2�E���f�EދE�f�E��Eމ��E܉ơ���VSP�  ��넋EЃ��x�������P�  ���7  ���[�������P�  ����D���U����}u�}��  u��h ��!   �����U�����h��  j��������ÐU��Ef�   �Ef�@  �Ef�@  �Ef�@  �]ÐU����E���u�u�u�u�uP�%  �� ����E��Eǀ�       ���U����E�@ �E�@a��t�E�   ��j j j j Pj�u6  �� �E���   ��uP����P�3  ����    �E�   ��j P�F3  ��������t����P��  ����ÐU��VS�E�@���r  �E�@��������X��E�@�H��E�@�P�E�@���uh�   h�   h�   SQRP�D  �� �E�@��������X��E�@�H��E�P�E�@�������E�@���uh�   h�   h�   SQRP��  �� �E�@�H��E�@�U�R���uj`j`j`jQPR�  �� �E�@�H��E�P�E�@ЍP��E�@���uj`j`j`jQRP�  �� �E�@�H��E�@�P�E�@�uj`j`j`QjRP�V  �� �E�@�H��E�@�P�E�X�E�@؃��uj`j`j`QjRP�  �� �E���   ��u@� ��E�P�E�X�E�@�������؃����uQj0j0RP�  �� �   �E���   ��u=���E�P�E�X�E�@�������؃����uQj0j0RP�7  �� �I�E���   ��u;���E�P�E�X�E�@�������؃����uQj0j0RP��  �� �E�P�E�@Ѓ��ËE�P�E�@�������E�@X��)ЉE�����uj j j SRP�  �� ��e�[^]ÐU����E� �E�E� ��t�E� �E����u���$  ���E��E��ًE�     �E�@    �E�@    ���f�f��UWVS��
  �ÓU  ���D$(�|$$�ƃ�)����ŋD$ ��	��t>��QW�t$,��  ����u	��[^_]Ð���/VR�D$,�P�)  ����[^_]Ð��QW�t$,�r  ������&    ��    UWVS�P
  ��U  ���t$ �|$$�T$(��   t*�B���t�v ���>�����u��[^_]Í�&    �t& ������R��WV�=  ����tӉ>��t̉~��tĉ~��[^_]Í�&    �t& ���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���|$$�L$,�D$4�\$8�t$(�T$0�|$�L$��y��D$    �L$��y�1����ȁ�   ���	���% �  ���͉���	�k	ǅ�~u;s}p�D2��L$�D$�D$�D��$��&    �D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�  ��ES  ���t$j j j j Vj �|0  ��$��[^� f��`  S  UWVS��,�|$@�t$D�D$�L$L�D$P�\$T�T$X�l$\��y|$H1���y�1�����������	�	E�T$�D$��~\;u}W�D$H��D$�D��D$�
f���9u~9�]������)�;\$OT$H��R��t$�L$ ��P�\$�X�����;t$u���,[^_]Í�&    �  GR  UWVS��,�t$@�l$D�D$�L$L�D$P�|$T��yt$H1���y�1��؉������� �  ��	�	G�T$�D$��~i;o}d�D$H��D$�D��D$��t& ���9o~C�G�_������)����;\$OT$H��R�t$�L$ ���P�\$�~�����;l$u���,[^_]Í�&    ��    UWVS�  ��cQ  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$�������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�@  ���O  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�,����� 9t$h�_�����L[^_]Í�&    UWVS�p  ��#N  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�\����� 9t$l�_�����L[^_]Í�&    UWVS�  ��SL  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�)�����9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$Ë$�f��S�   ������áJ  ���D$��D�P��  ��[Í�&    �S�������vJ  ���t$�  ��[Ív S������VJ  ���t$�h  ��[Ív S������6J  ���t$�������[Ív S�c�����J  ���t$�(  ��[Ív S�C������I  ���t$�  ��[�f��UWVS� ������I  ���D$<�|$8�t$0�D$�G�D$�D$D�������D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�M����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�~����� 9|$�b�����[^_]Í�&    f�UWVS�������sG  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��Ð��&    ��&    Ð��&    ��&    �D$�@Ð��    �D$�@Ð��    �D$�@ Ð��    UW1�V1�S������ßF  ���l$0�t$4h�   h�   h�   �u�u�u�u�R����E�D$,�� �l$0���|$0�D$    ��t& �|7
t^�����t$�j  ��9�~S���t$8��  P��  P��  P�D$GP�G��P�D7P�����G�� ��9���D$1��f��|$0��l$0�O�t$4j j j jj�t$ Q������ �t$4h�   h�   h�   �ujj �E��P�r����� �t$4h�   h�   h�   jjj�E��P�J����� �t$4h�   h�   h�   jj�E��P�E��P������<[^_]Ð�t& U1�WV1�S�l�����E  ���|$0�D$    �G���&    f��<0
tN����P�  ��9�~G���t$8j j j �D$ GP�G��P�G�0P������G�� ��9�G��D$1�멍v ��[^_]Í�&    �UWVS������ÃD  ���t$ �l$$�F ��~J1���&    ��    �F����    ��R�V(��P�F�U��EF����P�  ��9~ Ń�[^_]Ð��&    �t& ���  ��D  �D$ǀ     ���(�����T$�P�T$�P�T$�P�T$�PÐ��&    ��&    WVS�|$������ðC  ��W��  �T$ ���r=   $��h   j V��  XZWV��  ��[^_Ít& ��W�  YZPV�  ���Ő��&    �WVS�t$������@C  �|$����<����W�V  �FXX�FZWP�w  �D$(�F�D$,�F�D$0�F�D$4���F[^_Ít& WVS�t$�-������B  �|$�F�N�P��F���|$ ��   Wh�   h�   h�   jRQP������ Wh�   h�   h�   j�F��P�FF��P�F��P�T����� Wh�   h�   h�   �F��Pj�F��P�v�)����� Wh�   h�   h�   �F��Pj�F��P�FF��P������� [^_�Wj`j`j`jRQP������� Wj`j`j`j�F��P�FF��P�F��P������ Wj`j`j`�F��Pj�F��P�v������ Wj`j`j`�o�����t& UWVS������ÓA  ���t$0�|$4�F�n�N�P��F���l$���~ ��   ���n\�L$�N�L$����  ����  ����  ��Wh����h�����t$RP�t$ �������j WV������Wj j j �V�������F��P�V����ЋVX��F��)�P�t$(�P����� ��[^_]Ít& ���W��h�   �h�   ��h�   ��QRP�t$ �x����V�� W��h�   ��h�   �h�   ���P�R�N�Q�RFP�F��P�>����� Wj`j`j`j�F��P�v�F��P������ Wj`j`j`j�F��P�FF��P�F��P������� Wj`j`j`�F��Pj�F��P�v������� Wj`j`j`�F��Pj�F��P�FF��P������ ��[^_]Í�&    ��    ��Wh--��h22���t$RP�t$ �c�����jWV������Wh�   h�   h�   �k�����&    ��&    ���Wh��-�hȠ2�뮃�Wh�77�h�<<��VS������5?  ���t$�T$,�V��P�����D$ �F�D$$�F�D$(�F����P�9
  �V�F(�F�V�F ��[^Ít& WVS�t$�������>  �|$����d����W��  �F�$��	  �FZYWP��  �D$(�F�D$,�F�D$0�F�D$4���F[^_Í�&    �t& ��G   ��g>  �D$�@    �@    �@    ��x�����T$�P�T$�P�T$�P�T$�PË$�S�c�����>  �� j j j �t$4�D$$Pj�K  �D$,��8[�f�S�3������=  ��j j j j �t$(j!�  ��([Í�&    f�S�����ö=  ��j j j �t$(�t$(j��  ��([Í�&    UWVS������Ã=  ��(�l$<U�T����$�   �D$�����+   �T$����1����FjtUPǆ�   ����ǆ�   �����V�  �}�m����    ���� ��f��� vf��� wd���   ������P�/  �����   ���   ���   ��ǆ�       ǆ�       Ɔ�    Ɔ�    ��[^_]Í�&    ��&    �ȃ���P��  ��롍�&    ��    S�������v<  ���D$�p�u�����[��7�����W<  UWVS���l$0�T$�Eu(�����   S�����   �EP�EPj j ������� �E���   ��~?1����   �v 9�v\�M ��t1��v ���	9�u��A�������WP��E��9�̋��   ��t	��S�Ѓ���S�u�\$�������,[^_]Ð�    ��&    f�UWVS���D$0�l$4�|$8�p��~G� 1ۉD$��&    ��&    9�t<�D$��t1�f���� 9�u��@�P�H9�~9�|&��9�uσ�[^_]Í�&    �    ��&    f�H9�~�P9�~̅�t�T$1���&    ����9�u��T$�D$���@�P�R�D$@�����   ��[^_]Í�&    ��&    S���\$���   ��xn;CsY���t1Ґ���	9�u��A���P�R���   ��;Ss-���t1��t& ����	9�u��A��[Í�&    ��&    ��    ��&    f�ǃ�   ������1�[Í�&    ��&    �VS�R�����:  ���t$ j�E����T$ ���     �P��@    ��t�V��P�F�F��[^Ív ��F�F��[^ÐU��E�]�Mfof ��������]�U��E�]�M�o� ��������]�U��E�]�M��~4fn�fop�f��fs�f��fs�f��fs�f��f ������]Ð������                S�S�����9  ��h   �7  ����t�T$�@   �P��   �P��[Ít& S�������8  ��j �t$�  ����1���x���t$R��������[Í�    S������Æ8  ���D$�p�  ��1�[Í�&    ��&    S������V8  ���D$�D$P�t$�D$(�p��  ��[�f�S�s�����&8  ���T$��t���D$�D$PR�D$(�p��  ����[Í�&    S�3������7  ���t$�t$�D$�p�  ��[Í�&    �S�����ö7  ��jj �D$�p��  ��[Í�&    �t& �1�Í�&    ��    1�Í�&    ��    S������f7  ���t$jj�D$P������[Í�&    �v WVS�|$�}�����07  ��W�U  �t$$j��PW������� 9�[^��_�����f�f��U��01�WVS�;������6  ��(��8
  �����9�4
  C�4
  P���8  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p�¨�1���8
  �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � �����4  ��8   �g�����&    �t& ����g5  ǀ@      �¨�ǀ<      �    �B    � �ǀ8
     �    �B    ��ǀ4
      �    �B    ǀ4      ǀ8      ǀ,      ǀ0      ǀ$      ǀ(      Í�&    �UWVS� ����ó4  ���|$0� ��&    ���4  �   ��8   ��  �w ��  ��t܋�@  �t$�|$0����  �|$0��<  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s��<  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ���@  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$���������B1ҋD$~Q��@�����   ��   �E���  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,�����E$���~�Ƙ�Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ�������������@  ���K�����  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~�ǘ��N,�����ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��t  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS� ������0  ���D$ ����   �P���)փ� C���  �N�A=����~   �y�Š�1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o��<  ����   ��t�J+J�ʋO)�9�|W�  ��[^_]Í�&    �v ��,  ��0   ����� ���� t
f=��t<�u���$  ��(   뱍�&    ���<  롍�&    ���4  ��8   ��[^_]Í�&    �v �G9�@  tU9�ta���t�B�G��t������G1�)Q���wW�  ���4�����&    �t& �o�������&    ���@  룍�&    �ǃ<      듍t& WVS�t$�m����� /  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS������3.  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��A  �G�P�������   �P9���   �T$�+  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ�,  ��0   %��� =�� tDf����t=���t8�s  1���[��^_]Í�&    �p���V  ����[^_]Í�&    �t& ���$  ��(   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ�����f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f��T$1��: t�t& ����< u�Í�    Í�&    ��&    �UWV1�S������Ñ*  ���|$ �l$$�f��D5 �7����U�����7��9��� ����[^_]Ít& �UWVS�t$�\$�L$��t}�A�S9���9���	ЍV�����tm��	Ȩue���ȉڃ��ύ�&    �v �(�����j�9�u����9�t'���B9�v�D�D�B9�v	�D�D�� [^_]Í�&    �ȉٍ<0��&    f�������Q�9�u��͍�&    ��&    VS�������u)  ���t$V����ZY�t$�P��������[^ËD$�L$��t& �����t	�8�u�Ð1�Í�&    ��    �D$�8 t��&    ���8 u�Í�&    U1�WVS�>������(  ���t$ �|$$���u�'��&    �t& ���.��t��PW�k�������u����[^_]Í�&    �v U1�WVS������Ñ(  ���t$ �|$$���u�'��&    �t& ���.��t��PW��������t����[^_]Í�&    �v WVS�t$�}�����0(  �|$��tV��D  ��WV�����XZWV�k��������D  9�t<1Ҁ8 u��D  ��[^_Í�&    f��  �P�㍴&    ���D  ��u�1���f�ǃD      1���f�VS�\$�t$��8�u"��t(�   ������t��8�t���)�[^Ít& �1�[^)�Í�&    f�UWVS�D$�\$�l$�0���8�u`��t@�<(��u�[��&    ��t,9�t8�����0���8�t�����[)�^_]Í�&    f�1�1�[)�^_]Ít& ���[��)�^_]�����������ōt& �UWVS�������&  ���t$ �|$$��t& ��t)�������P��  ����$�  ��9��t����[^)�_]Í�    UWVS������c&  ���l$0�D$8�t$4�D$���&    �v ��t1;l$t+�����E ��P�S  ����$�F  ��9��E t����[^)�_]Í�&    ��&    WVS�t$�-������%  ��V�������$�
����4$�����������Pj W�!���XZVW������[^_ÐS������Ö%  �� j j j �D$ P�t$8j��  �D$,��8[�f�S������f%  ��j j j j �t$(j�  ��([Í�&    f�S������6%  �� j �D$P�t$8�t$8�t$8j�g  �D$,��8[Í�&    ��&    S�C������$  �� j �D$P�t$8�t$8�t$8j�'  �D$,��8[Í�&    ��&    S�����ö$  �� j �D$P�t$8�t$8�t$8j��  �D$,��8[Í�&    ��&    S�������v$  �� j �D$P�t$4�t$<�t$8j�  �D$,��8[Í�&    ��&    S������6$  ���t$�t$�t$�������[Í�&    �t& S�S�����$  ���t$�t$�t$�������[Í�&    �t& S�#������#  ���t$�t$�t$� �����[Í�&    �t& S������æ#  ���t$�t$�������[Í�&    ��&    �S�������v#  ���t$�������1�[ÐS������V#  ��j �t$�������   ��u
����[Ív ��P������1҃���[�f�f�f�f�f��S�S�����#  �� j j j �D$ P�t$8j�;   �D$,��8[�f�S�#������"  ��j �t$0�t$0�t$0�t$(j�   ��([�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��S�������v"  ��j j j j j j������ ��&    ��    ���f�f�f�f�f�f���T$�   �JЃ�	v���1���A����ËD$��߃�A������Í�&    �t& �1��|$z��Ít& �1��|$@��Ít& ��D$��0��	����Í�&    ��&    ��T$�   �JЃ�	v���1���A�����Í�&    ��&    ��D$��!��]����Í�&    ��&    ��T$�� ����	��	���Í�&    �v Í�&    ��&    �1�Í�&    ��    VS�r�����%!  ���t$V��������u��[^Í�&    f���V��������������[^Í�    �D$��_Í�&    ��D$�� �f�f�f�f�1�Í�&    ��    ������   �����  1�Í�&    �v S������Æ   �� j j j �D$ P�t$8j�����D$,��8[�f�1��f�f�f�f�f�f�������t6U��S������&    �v �Ѓ�����u��[]Í�&    ��&    �������     / r /file.bmp /binfile.bmp /folder.bmp          Ї��8�       zR |�        ����)    A�Be�     <   ����>    A�Bz�     \   ����    A�B�� (   |   �����   A�BB����A�A�       �   ����   A�BG���(   �   {���z   D Gu Eutu|ux    �   ����U    A�BQ�      ����(    A�Bd�     8  ����    A�BV�  �   X  �����    A�A�A�A�N c$A(A,D0H G
A�A�A�A�BC$D(A,G0H C
A�A�A�A�BC$A(A,D0H    \   �  �����    A�A�A�A�N n
A�A�A�A�LC$F(D,A0H YA�A�A�A�   <  ���?    Cy 8   T  0����    A�A�A�A�C$�A�A�A�A�8   �  ����.    A�A�NFB B$B(A,B0HC�A� H   �  �����    K�A�A�A�C@�DAHFLHPL@IA�A�A�A� H     \����    K�A�A�A�C@�DAHDLJPL@IA�A�A�A� <   d  ����b   A�A�A�A�NPL@�A�A�A�A�X   �   ����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X      �����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   \  ����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   �  l����    A�A�A�A�C(�A�A�A�A�   �  %���          �  ���             ���(    A�SJ HA�     0  ���    A�ND HA�     T  ���    A�ND HA�     x  ���    A�ND HA�     �  ���    A�ND HA�     �  ���    A�ND HA�   �   ���W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   �  L���s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�     P  t���          d  p���          x  l���	          �  h���	          �  d���	       �   �  `���{   A�A�C�C�N0H4E8E<E@CDCHCLCPO0e<D@H0G4D8H<H@HDHHILFPK0c4B8B<B@BDBHDLAPH0D4E8E<E@CDBHBLGPH0D4E8E<E@BDBHBLGPH0D4E8E<E@BDBHGLGPHA�A�A�A� \   �  �����    A�C�A�C�N0f<A@H0G4D8B<B@BDHHILHPK0YA�A�A�A� H   �  <���s    A�A�A�A�N d$K(G,V0H HA�A�A�A�     D	  p���A       d   X	  ����g    A�A�A�RA LMEBA FAAA HA
�A�A�ECA FAAA H@   �	  ����\    A�A�A�VL IDAA aD�A�A�   �   
  ����K   A�A�A�nEEE B$A(A,A0HAEEE B$G(J,G0HAEEE G$B(G,C0HAEEE G$B(G,J0HA
�A�A�AABBB B$A(A,A0HABBB B$G(J,G0HABBB G$B(G,C0HABBB �  �
  (���`   A�A�A�A�N0Z4A8E<E@DDAHALDPH4B8A<A@H4A8B<B@BDSHXLDPH0C
A�A�A�A�FC4H8G<G@DDAHALDPK0A4G8H<G@FDGHDLGPH0A4B8B<B@BDGHCLGPH0A4B8B<B@BDGHJLGPH0A4B8B<B@GDBHGLCPH0A4B8B<B@GDBHGLJPH0C
A�A�A�A�NC4A8E<E@DDAHALDPH4B8A<A@H4A8E<E@EDT0C
4A8E<E@BC4A8E<E@ (   �   ���\    A�A�Nr WA�A�@   �  4���d    A�A�A�VL TAAA aD�A�A�      �  `���L            ����       0     ����.    A�N(B,B0B4D8E<B@LA�  0   P  ����'    A�NBB B$B(D,B0HA�  0   �  ����)    A�NBB B$D(D,B0HA�  `   �  |���   A�A�A�A�N<E@a4M8A<A@g0g<G@H0y
A�A�A�A�OE<D@H0        (���     A�NG HA� x   @  $����    L�A�A�A�C0Q8G<H@EDEHBLBPH0w8H<A@H0Q<A@E0C8A<C@LA�A�A�A�B0����X   �  x����    A�A�A�A�C0]
A�A�A�A�HD<F@J0IA�A�A�A�0     �����    A�CkC La
A�P]C� <   L  h���_    A�A�NF Lh
A�A�DLA�A�   $   �  (���<    A�NE H^A�  4   �  @���:    A�NBD HKDA HCA�       �  H���"    A�NG HC� (     T���.    A�NJDG HA�   ,   <  X���9    A�NKJAG HCA� (   l  h���(    A�NDDG HA�   (   �  l���$    A�NBBG HA�      �  p���          �  l���       (   �  h���&    A�NDBBE HA�@     l���;    A�A�A�RA I$B(C,A0HC�A�D�   D   \  h����   A�F�A�A�N<Z@J0�
A�A�A�A�M      �  �����       T   �  L����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `     �����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   t   ����    A�A�A�WA H��A�A�  �   �  �����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0<   <  ����   A�A�A�A�C �
C�A�A�A�A 8   |  �����    A�A�A�A��
�A�A�A�P      �  <���!       @   �  X���K    A�A�A�C�N Z,A0K JC�A�A�A�8     d����    A�A�A�A��
�A�A�A�H   4   L  ����0    A�A�NE FADC HC�A�   �  ����#          �  ���       D   �  ���V    A�C�A�A�N j(A,A0H GC�A�A�A� D   �  0���V    A�C�A�A�N j(A,A0H GC�A�A�A� D   <  H����    A�A�A�`AA HAAA H\
�A�A�J ,   �  ����G    A�A�w
�A�FC�A�  \   �  �����    A�A�A�A�M
�C�A�A�JE
�C�A�A�FD
�E�A�A�A @     ����Z    A�A�A�A�N ^,A0U MA�A�C�A�@   X  ����r    A�A�A�A�N0u<A@U0NA�A�C�A�L   �  8���O    A�A�A�RA ]DBA FAAA HA�A�A�   0   �  8���.    A�N(B,B0B4E8D<B@LA�  0      4���'    A�NBB B$B(D,B0HA�  0   T  0���2    A�N(B,E0D4D8D<B@LA�  0   �  <���2    A�N(B,E0D4D8D<B@LA�  0   �  H���2    A�N(B,E0D4D8D<B@LA�  0   �  T���2    A�N(B,E0D4D8D<B@LA�  (   $  `���%    A�NDDD HA�   (   P  d���%    A�NDDD HA�   (   |  h���%    A�NDDD HA�   $   �  l���!    A�NDD HA�      �  t���    A�ND HC� 8   �  p���E    A�NBD HL
C�DCA HEC�0   0  ����.    A�N(B,B0B4E8D<B@LA�  0   d  ����-    A�NBD D$D(D,B0HA�  (   �  |���!    A�A�A�[�A�A�,   �  ����3    A�NBB B$B(B,B0H     �  ����             ����            ����          0  ����          D  ����          X  ����           l  ����          �  ����          �  ����          �  ����          �  ����       D   �  ����J    A�A�NE HG
A�A�JCA HHD�A�       ����          ,  ����          @  ����          T  ����       0   h  ����.    A�N(B,B0B4E8D<B@LA�     �  ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ������    ����            ������        ������        ���Й         �����        `�����        ������                                                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              ��                           >        ���    src/gfx/sse2.asm NASM 2.14.02 ��     %  . @   l    '   �       src/gfx/sse2.asm      �!0==?LL==0/!$!0==?LL==0/!#!0==>=0K�KYKYKYMK>1/""u�                                               t�          ��          ��          ��          ��           �          �          �          �     	     ��     
     ��          ��                                                                                                                                  ��   �         �      (   ��      ;   ��      =    �      P   P�      f   ��     u   ��     �   Ё      �   ��                 ���   �      �   t�      �   @�      �            ��  ��                  ��  ��(     F  ��     d           ��q           ��}           ���           ���           ���           ���           ���  �       �  �       �  \�       �  e�         p�                ���           ��  ���    '  ��     2  ��     >  ��     M  ��     W  ��     a  ��     n  ��     �           ���           ���  ��     �           ���           ���           ���           ���           ���           ��             ���  ��     
 �  ��     �  �K     �  @�.       `��    A  ��     f  p�.     �  Ї�  "  �  �`    �  ��     �  ��'     �  �!     �   ��     �  �       ��.       ��       ��(   "    P�2     '  @�     /  ���    [  ��A     o  ��     v  @�\     �  ��     �  ��     �  ��-     �  �     �  �.     �  ��     �  ��     �  �     �  0��     �  Ы�    �   �t       Օ       ��     %  `�J     -  ��{    I   �     Q   �     X  ��K    �  <�   ! 	 �  ��%     �  �     �  0�   "  �  (�   ! 	 �   �r     �  l�     �   ��     �  ��U   "    о      �  t�        п     #  ��>   "  =  ��	     W  І)   "  k  ���     �  p�     �  @�\     �  `��     �   �      *  ��%     �  �     �  ���     �  `��       �0       �      ��(     $  ��2     0  ��W    K  І)   "  _  ��     y  �     9	  ��&     }  �     �  x�   ! 	 "  P�%     �  ��A     �  ��     �  0��     �  ��_     �   �.     �   �s       P�   "    @��       ��Z     &  P��    .  @��     S  P��     Z  ٕ     p   �    �  ��<     �   �b    �  p��     �  �      �  p�     �  �   ! 	 	  �s     !	  0�.     '	  ��O     .	  ��:     4	  ��      @	  P��     f	   �    m	  �z    r	  Ш$     x	  ��     �	  �?     �	  P�   ! 	 U   �     �	  p�   "  �	   �L     �	   �"     �	   �     �	  P�      �	  P�     �	  �G     �	  P�\     �	  ��   !  	
  ��      
  Мg     '
  �V     /
  Т)     K
  ��     f
  0�     t
  P�\     �
   �&     �
  �   "  �
  8��   "  �
  ��     �
  ��     �
  `�9     �
  0�E     �
  ��      �
  ��      �
  ��d     �
  ��       л2     !  �3     &  Й	     =  �     E  0��     i  ��V     p  ��!     �  �!     w  ��        �'     �  ��d     �  @�#     �  P�;     �  ��     �  d�   ! 	 �  ��	     �   �      �  ��   "  �  �2     �  �      �  �     	  ��>   "  #  ���     o
  ���    R   �L      crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_fileIconBuffer graphics.cpp runtime.cpp text.cpp widgets.cpp window.cpp font.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset_sse2.loop memset_sse2.ret bigzero fileio.c allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns memory.c string.c p.1056 filesystem.c ipc.c syscall.c exit.c ctype.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated strcpy _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN15ScrollContainer5PaintEP7Surface _Z13_CreateWindowP10win_info_t _ZN10FileButton5PaintEP7Surface _ZN6Button5PaintEP7Surface l_max_inuse _Z14_DestroyWindowPv syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm lemon_read isblank _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN7TextBoxC2E4Rect memcpy _ZN6ButtonC1EPc4Rect l_inuse __TMC_END__ SendMessage __DTOR_END__ lemon_open islower tolower feof _Z11PaintWindowP6Window malloc windowInfo __x86.get_pc_thunk.ax __dso_handle ispunct _ZN7TextBox5PaintEP7Surface isspace fflush _ZN6Button17DrawButtonBordersEP7Surfaceb _ZTV6Button lseek fd _ZdlPv _ZTV7TextBox strncasecmp __x86.get_pc_thunk.dx _Z15HandleMouseDownP6Window8Vector2i _ZN4ListIP6WidgetE5clearEv isxdigit liballoc_lock _ZN10FileButtonC2EPc4Rect _ZN6Button11OnMouseDownEv _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm strrchr _ZN6ButtonC2EPc4Rect calloc memcpy_sse2_unaligned folderIconBuffer _Z16memcpy_optimizedPvS_m _ZN5Label5PaintEP7Surface strcat _Z12RefreshFilesv fseek lemon_write _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev _ZN6Widget11OnMouseDownEv win exIconBuffer _ZTV15ScrollContainer _ZN7TextBoxC1E4Rect isupper strncmp _Z9AddWidgetP6WidgetP6Window liballoc_alloc _ZN6Bitmap5PaintEP7Surface _ZdlPvm strncpy strcasecmp realloc _Z8DrawRectiiii10RGBAColourP7Surface strtok __x86.get_pc_thunk.bx _Z12CreateWindowP10win_info_t fdopen _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window isalpha _ZTV6Widget _Z10DrawStringPcjjhhhP7Surface fread strdup fopen __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main ftell font_default _Z5floord _ZTV6Bitmap _ZdaPv _ZN15ScrollContainerC2E4Rect fclose isgraph isalnum isprint strcmp _ZN6BitmapC1E4Rect _ZTV10FileButton _fini _ZN7TextBox8LoadTextEPc strcspn _Z12_PaintWindowPvP7Surface _ZN6Widget5PaintEP7Surface liballoc_free _ZN6BitmapC2E4Rect fputc _Znam _ZN10FileButton9OnMouseUpEv _ZN6Widget9OnMouseUpEv isdigit fwrite access _edata _end _ZN5LabelC2EPc4Rect _Z13HandleMouseUpP6Window lemon_seek exit _ZN6Button9OnMouseUpEv iscntrl _Z10surfacecpyP7SurfaceS0_8Vector2i strspn strlen toupper lemon_close _ZN5LabelC1EPc4Rect strchr fputs font_old _ZTV5Label _ZN7TextBox11OnMouseDownEv memset_sse2 _ZdaPvm lemon_readdir memcpy_sse2 _ZN10FileButtonC1EPc4Rect _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN15ScrollContainerC1E4Rect  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .data.rel.ro .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                   t�t                     !         ���   �?                 '         ���@                    -         ���@  <                  5         ���@  �                 ?          � `                   K         �`                    R         �`                    Y         �`  x                  f         ���`                   o         ���`  (
                  u         ���j  �                   z      0       �j  +                 �              �j                     �              k                    �              %k  B                  �              gk                    �              �k  p                  �              �k                    �              �k                                  l  �     J         	              �z  o                               +�  �                  