ELF              ��4   d      4    (           � ��A  �A           �A  �����  �        �W  �24  �                 �    UU���s   VW�����_^�y  �    �i���f�f�f�f�f��(�=(�t$�    ��tU���h(��Ѓ��Í�&    f�Í�&    ��&    ��(�-(����������t(�    ��tU���Ph(��҃��Í�&    �t& �Í�&    ��&    ��=(� ugU�,���V���S����������9�s�v ���,����,�9�r��'����    ��t��h(��Q~�����(��e�[^]�Í�&    ��&    ��    ��t'U���h0�h(��~������	�����&    f���������t$�!  ��Ã��t$�~!  ��Ã��t$�(  ��Ã��t$�(  ��Ã��t$�(  ��Ã��t$�r(  ���UWVS���t$(�|$,�T$4�\$0�T$�F�D$�G�D$�~ ��   �G)Ѕ���   �T$�$    �[���F9�~4�O��)�9�~)�$Ћl$�l� ������v��L$���D$�,��$�$9F~*�D$�G+D$;$~�F��~܋O��)څ�~Ѻ    롃�[^_]�UWVS��8�l$L�|$P�D$T�D$�L$X�L$ �t$\�L$`�L$�\$d�\$$�T$h�T$(j�/   ���     �@    �@    ��9�
�D$�9�}R�L$9��D$�9���   t$9�|�D$�9���   �t$�T$�9�|�D$�9��  �؃�,[^_]Ã�j�  �     �@    �h�x��)���P�L$$�H��C�C   �����j�����j�h  �     �@    �h�x�L$ �H�T$)����P���; t�S��S�P�C�C�|$�-�������)�D$��j�	  �     �@    �p�x�T$ +T$(�P�L$$�H���; t�S��S�P�C�C�D$�D$���������j�  �     �@    �h�p�L$ �H)��T$$)�P���; t�S��S�P�C�C�������S��(�\$0�St�T$�Kx�L$�D$    �D$    �C|�D$���   �D$�Cu	�=�� u#��j �D$P�D$(P�sph��j�4-  ��H[�h��j j j ��PjQR�  �� h��j j j ���   ��Pj�sx�C|Ct��P��  �� h��j j j j�C|��P�sx�st��  �� h��j j j j�C|��P���   Cx��P�st�  �� 9���6  h��h�   h�   h�   j�s|�Cx��P�Ct��P�b  �� ��h��h�   h�   h�   �Cx��P�Ct��P�CP��  �Ct�Sx�H�L$8�J�L$<�� h��j2j2jdjj��RC|��P��  �� h��j2j2jdjj�Cx��P�C|Ct��P��  �� h��j2j2jdjj�Cx��P�C|Ct��P�  �� h��j2j2jdjj�Cx��P�C|Ct��P�  �K|Kt�A�Kx�Q�� RPh��h���  ��������h��h```�h   �j�s|�Cx��P�Ct��P�>  �� �����S��j j j hh�hl�j�+  �l��h���+x�i��  ��+t�Ѓ� =�  v,����̉��%|����p��|�    �x��t���[�ÍL$����q�U��WVSQ���   j j j h���E�Pj�~*  ����������P�5  ��������n  ���   ���   ��� ���j��  �     �@    �@    �H���j j j j h��j��)  ��j j j �E�Ph�j��)  ���   ���   ��j h��(  ���$   �  �����jj S�\(  �ǉ$�g  �ƃ�WPS��'  ��h��Vjjj j �  ��S�{(  ��j h��C(  �Ã�jj P�(  �ǉ$�  �ƃ�WPS�'  �T�   �X�   �$  0 ��  �`�����u%ǅ@���    ǅ8���    ǅD���    �  ����hL�Vh   h   j j �j  �� �ǅ<���    fǅl���  fǅn���  fǅp���  fǅr���  ��j j j ��l���P��<���j�z(  ��@����ǃ� ����   �uܻ    � �    �	��D����B;ppt/��9���   ��9�@���vօ�tً�D����    ���9�u���9�@���vQ���+	  ��D����    ���9�u��Bƀ�   ��D����    ���9�u��B��l����   ����   �    ƀ�   �    �ك�h�   �o  �Í�l����   �����l����Ct��n����Cx��p����C|��r������   ƃ�   ����$   �  �     �@    �X����D��� t=��8�����H��@��������8�����<�����<���9�T�����  �7�����D����������@���������  ��������<����  �5    �   ��D����  ��D����H��4������t�H��t�J�P��t���t�
��u���D�����@�����@���9�t��P�U  ����8�����H��8����ድ8�����j��  ��8����     �@    ��4����H����D��� ��   ��p��@�����@���9���   ����   ��D����    � ��9�u��@�������Wx����J9���   �G��  �5���Ot��<���O|�Y�9�}�Z9���9�|�J9�E+�<����5��)У�������  ��8�����D����E����    �o�����D����a���ǅt���   �Gp��|�����P��x���j��p�����l����wl�$  �� �m  ǅt���   �G�  ���+Ot����)��
  �������  ��9���������������D����    �6��9�u��v�Ft9�~�F|9�}��Fx9�<���~���   9�<���}�����@���������9��������������D���� ���(  �    ��9�@��������9��~�������  ���ۡ    ���    t���5    �\����    ���i  �    ;���_  ���    �    �K  ��D������t�Q��t�P�A��t���t���u���D�����9�t��Q�  ���    ��  �A��8����߉�@�����X�����S��"  ������   ��`���� uࡨ���t׋�d�������t �у�tǅt���   �� ���x����ǅt���   �� ���x����Pp��|�����R��x�����t�����p�����l����pl�}"  �� �^����5���5��h��h���5���h��j j j jjj j �  ��,j
��l���S�5p��#  ��h��h�   h�   h�   j j S�  ��j j j h���u�j�8"  �� �|�������j ��P���Pjh���u�j�"  �� ��P��� t>����Q����P���    H£���A�؋���B���    H£���=�� t3���������+���    HӉQt+���    HAx�����j j j j ��T���Pj�f!  �� ��T��� ������������t���S�������   �=�� t��� h��h�   h�   j@�����P�5��j j ��  �� �    ��@�����@��� �u  �y�����D����@���ǅt���   ���+Ot)�����ȉ�x����Wp��|�����RP��t�����p�����l����wl�@   �� �=�� �Q������� �C������ ��� ǅt���   �������������|�����x�����t�����p�����l����pl��  �� �������D����H��4����������    ��   ����D����s�F��������V��D����@��D������    ��   ��tȋ�D����    ���9�u����r� �������D����    ���9�u��Bƀ�    ��9�������9��R�����t���D����    ���9�u��B���    u���D����    ���9�u����9B�������R�����D�������(����    ��9��8���9��0�������Q������ߋ�D����Bƀ�   �����f�f�f�f��UWVS�
  �Ï=  ���|$$�D$ �l$(	��t��UW�t$,��  �������)�����RW�t$,�  ����u
��[^_]�f����VW�t$,�V�  ����[^_]�f���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���D$4�|$,�L$$�\$8�T$0�t$(�|$�ǉL$�ȁ�   ���	���% �  ���͉���	�k	ǅ�~o;s}j�L$�D$�T2��T$�D��$��D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�~  ��<  ���t$j j j j Vj �  ��$��[^� f�UWVS���|$�t$ �l$(�D$,�\$0�L$4�T$8��y|$$1���y�1�����������	�	��B�D$��~j;r}e�D.��$�D$$�\���&    f��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS���|$�t$ �\$(�D$,�T$0��y|$$1���y�1���������� �  ��	�	��B�D$��~m;r}h�D��$�D$$�\���&    �t& ��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS�  ��/:  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$��������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�<  �ÿ8  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�<����� 9t$h�_�����L[^_]Í�&    UWVS�l  ���6  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�l����� 9t$l�_�����L[^_]Í�&    UWVS�  ��5  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�������9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$�f�f�f��UWVS�������o3  ���D$<�|$8�t$0�D$�G�D$�D$D���� ��D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ�`����� ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�-����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�^����� 9|$�b�����[^_]Í�&    f�UWVS������1  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f���U����  �0  ǀX      ǀ\      ǀx     ǀ|      �����    �B    �����    �B    �����    �B    ǀ`      ǀd      ǀh      ǀl      ǀp      ǀt      �]�U����9  �/  �E�    ��U�E�ЋU��E��E�;Er�E��U����  �/  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS��������3/  �E���E�E���x  �E�    ��Ѕ�u��x  �E�    ���E����x  �E�    �����E䋃|  9E�s	��|  �E���u��q  ���E���jj �u���������}� u%��`  ��d  ���� ��`  ��d  �    �l�E��     �E��@    �E��U�P��x  �E�E��P�E��@   �E��@    �E��@�ƿ    �����P� ��������Q�E��e�[^_]�U��WVS��L�x������-  �E�    �E�    �E�    �E�    �E�E��E� �J  �}� u5��`  ��d  ���� ��`  ��d  �5  ��j�������  ��X  ��u-���u��9�������X  ��X  ��u��  �    �{  ��X  �E��E�    ��\  ���C  ��\  �P��\  �@)ЉE��E�    �E����    ;E؉�E��
  ��\  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ�\  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u��X  �E��E�    �|  ���u��'������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���u  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ���  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����	  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u��X  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������v	  �    �e�[^_]�U��WVS��,�D������&  �} u#��`  ��d  ���� ��`  ��d  �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx��h  ��l  ���� ��h  ��l  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��p  ��t  ���� ��p  ��t  �  �  �E��@�E������P� �M��I�ο    )��������Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ��X  9E�u�E܋@��X  ��\  9E�u
ǃ\      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋������P� �M܋I�ο    )��������Q�E܋@��P�u��  ���G��\  ��t=��\  �P��\  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉�\  ��  �e�[^_]�U��S���  K$  �U�U�U�U��R���%������E��E��Pj �u��-������E��]���U��S���}����� $  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E��  �E���E�E�@=���tz��h  ��l  ���� ��h  ��l  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��p  ��t  ���� ��p  ��t  �  �    �_�E�@�E�E�;Er�E�U�P�  �E�;�u  ���u��������E���u��u�u����������u��������E�]��Ë$�U���������"  �E�E���E��P�U��U��E�P��U��u�E��U��� ����_"  �E�E��E�E��E�E��"�E��P� �M���Q�E��E��m�E�E�}�w؋E�E���E���E���E��E��m�E�E��}�wދE�E���U��E�ЋM��U��� ��m�E�E�}� uۋE��U��S�������!  �M�U��j j j QRj���  �� �E�]���U��S��������!  �U��j j j j Rj���  �� ��]���U��S������N!  �]�M�U��j S�uQRj���T  �� �E�]���U��S���o���!  �]�M�U��j S�uQRj���  �� �E�]���U��S���6����   �]�M�U��j SQ�uRj����  �� �E�]���U��S��������   �]�M�U��j S�uQRj���  �� �E�]���U��S�������j   ���u�u�u����������]���U��S������>   ���u�u�u���������]���U��S���l���   ���u�u�u���������]���U��S���@����  ���u�u���������]���U��S�������  ���u���������    �]���U��S�������Ò  ��j �u�������E�}� t���u���������    ��   �]���U��S������H  �M�U��j j j QRj���Q   �� �E�]���U��S���l���  �U�U�U�U��U�U��j �u��u��u��uj���	   �� ��]���U��WVS�'����  �E�]�M�U�u�}�i�[^_]�U���������  �E�E��E�E��E�    ��E��E��E��9E�|��E�    �)�E�� �E�E���E��E��U��E��m��E��E�������9E�|Ɛ��U��S���   ��$  �E�    �} ua�E�P�U�E�� 0�U�E��  �E�e�E��}�U��}�	~
�E���W����E���0�ËE�P�U�EЈ�E��}�E�} u��U�E��  ���u��u����������E�]��Ë$�U�������x  �    ]�U������d  �� ��  �    ]�U��S������C  �M�U��j j j QRj���L����� �E�]���U���k���  �    ]�f�f�f�f�f�f��������t6U��S�������&    �v �Ѓ�����u��[]Í�&    ��&    ��Z����  /taskbar.lef /dev/mouse0 /close.bmp /bg1.bmp          zR |�        ����    CD H     8   ����    CD H     T   ����    CD H     p   ����    CD H     �   ����    CD H     �   ����    CD H  8   �   u����    A�A�A�A�C(�A�A�A�A�h      ���
   A�A�A�A�CLvP^@[
A�A�A�A�ACLBPx@JLBPn@oLBPm@kLBPm@   p  l  ����r   A�C0E8B<E@EDCHELBPHA�A0�E4B8B<B@DDBHALAPH0E4B8B<B@JDBHCLJPH0E4B8B<B@BDGHCLCPH0E4B8B<B@BDGHMLCPH0Q4E8E<E@BDCHGLGPH0C4E8E<E@EDGHGLDP\0E4B8B<B@BDBHDLGPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPW0A4A8E<E@H0H4E8E<E@BDCHGLGPH0 4   �  ����z    A�CBB B$E(E,B0lvA�        ����       ,   ,  �����   D Gu Fupu|uxut|   \  ����~    A�A�A�A�N U$A(A,D0H E$K(A,D0H G
A�A�A�A�CC$C(A,G0H CA�A�A�A�     �  ����?    Cy 8   �  �����    A�A�A�A�C$�A�A�A�A�8   0  D���.    A�A�NFB B$B(A,B0HC�A� 8   l  8����    A�A�A�A�C�A�A�A�A�8   �  �����    A�A�A�A�C�A�A�A�A�<   �  `���b   A�A�A�A�NPL@�A�A�A�A�X   $  �����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   �  ����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   �  x����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   (  �����    A�A�A�A�C(�A�A�A�A�   d  ����         x  ����W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   �  ����s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�     �  ����    A�B��      ����7    A�Bs�     $  ����r    A�Bn� ,   D  ����8   A�BF���+�A�A�A�   ,   t  ����4   A�BF���'�A�A�A�   ,   �  ���~   A�BF���q�A�A�A�       �  Q���K    A�BD�C��     �  x���f   A�BD�^��   	  ����          0	  ����8    A�Bt�     P	  �����    A�B��     p	  J���6    A�BD�n��      �	  \���2    A�BD�j��      �	  j���9    A�BD�q��      �	  ���9    A�BD�q��       
  ����9    A�BD�q��      $
  ����9    A�BD�q��      H
  ����,    A�BD�d��      l
  ����,    A�BD�d��      �
  ����,    A�BD�d��      �
  ����)    A�BD�a��      �
  ����+    A�BD�c��      �
  ����J    A�BD�B��        ���6    A�BD�n��      D  ���F    A�BD�~��  (   h  <���*    A�BC���`�A�A�A�    �  :���~    A�Bz�     �  �����    A�BD����    �   ���          �  ���    A�BP�       ���    A�BY�      ,  ���6    A�BD�n��     P  ���    A�BP�      ����    ����                                                              @  �                          �             �   �            �����   �           ���������   �          �������������   �         �����������������   �        ���������������������   �       �������������������������   �      �����������������������������   �     ���������������������������������   �    �������������������������������������   �   ���������������������   �   �   �   �   �   ���������   ���������   �����      �����   �    ���������   �      �   �     ���������   �����      ����   ���������   �          ���������   �       ����   �   �����                 1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                                                                                                                                                                                                                                                                                            <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              �                           >        ��    src/gfx/sse2.asm NASM 2.14.02 ��     %  . @   :    '   �       src/gfx/sse2.asm      �                                         t�          ��          �          ��          (�          ��          ��          ��          ��     	     (�     
                                                                                                                             ��   ��         ��      (   (�      ;   ��      =    �      P   P�      f   (�    
 u   ,�    
 �   Ё      �   0�    
             ���   ��      �   ��      �   ��      �            ��  ��                  ��           ��#           ��,           ��5           ��           ��F   �    
 P  �    
 Z   �    	 e  $�    	 q  �    
 �  �    
 �  �    
 �  ��7     �  ��r     �  g�8    �  ��4    �           ���           ���           ��           ��           ��           ��             ��  ��      5  $�     K  ��    
 W  ��.     i  ���    �  ��    	 �  ��    
 �  в*     �  ��~     �  |�    
 �  ��     �  <�     �  t�    
   T�6     >   �    
   �       N�9     $  H�    
 0  ���    �  >��     \  ��    
 d  (�    	 p  ��F     |  ��     �  ��    
 �  �6     �  e��     �  ��4    �  �     �  ��    
 �  ��    	 �  x��       h�    
   ��,     !  ��    
 )  %�     0  ��    
 �  t�      5  (�     C   �    	 M  ��    
 T  Q�K     [  p�    
 e  ��    
 �  ^�,     o  �~     �  ��    
 �  ��9     �  0�W    �  $�     �  l�    
 �  ��&       2�,        �   	    Y�6     /  5�     7  ��f    ?  ���     d  %�     z  ��    
 �  p�b    �  Е�     �  ��s     �  x�    
 �  (�     
    Д�     �  �8     &  %��    +  ��    	 3   �    	 @  ��?     J  L�    
 T  E�     [  �      a  ��z     v  ��     �  �     �  
�J     �  (�     	 �  $�     
 �  ��    	 �  .�
    �  ��9     �  8�r    �  ���     �  ��)       �2     #   �    	 ,  U�     4  ��9     B  �        ߱+     N  0��       Ӫ~     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp graphics.cpp text.cpp font.cpp src/gfx/sse2.asm l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 memory.c filesystem.c ipc.c syscall.c itoa.c _liballoc.c _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos l_max_inuse syscall reverse frameCounter liballoc_init liballoc_unlock lastUptimeMilliseconds ReceiveMessage _Znwm lemon_read bgClipRects _Z12DrawGradientiiii10RGBAColourS_P7Surface l_inuse __TMC_END__ SendMessage __DTOR_END__ dragOffset lemon_open _Z12surfacecpy_tP7SurfaceS0_8Vector2i malloc __x86.get_pc_thunk.ax mouseSurface __dso_handle itoa currentUptimeMilliseconds lseek surface _ZdlPv drag liballoc_lock keymap_us active calloc frameRate mouseData _Z16memcpy_optimizedPvS_m closeButtonSurface lemon_write _Z8DrawCharciihhhP7Surface _Z30RecalculateBackgroundClipRectsP4ListIP8Window_sE currentUptimeSeconds mouseSurfaceBuffer liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface main testKey font_default _Z5floord bgSurface _ZdaPv _fini _Z15UpdateFrameRatev liballoc_free _Znam access _edata _end redrawWindowDecorations _Z14SplitRectangle4RectS_ lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close font_old _ZdaPvm lemon_readdir memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                  t�t                     !         ���   a4                 '         ��4                    -      2   ���4  -                 5         (�(5  p                 ?         ���A                    F         ���A                    M         ���A                   V         ���A  h                  \         (�(Q  �                  a      0       (Q  +                 j              SQ                     y              sQ                    �              �Q  B                  �              �Q                    �              �Q  >                  �               R                    �              $R                                  4R  �	     =         	              �[  }                               Qc  �                  