ELF              ��4   HC      4    (           � ��,  �,            0   � ��  �                    �   ��U��WVS��L  fǅL����fǅN���,fǅH���2 fǅJ���2 ǅP���    ����H���P��  ���E؍�D����أ��j j j PRj�  �� ��������������D�����j Qj RPj�  �� �E�
   �E�
   �E�    ����������  �E�E��E��E��E�x   �E�   ��hd  ��  ���ǃ��u��u��u��u���������PW��  �� �}ԋE�ƀ�   /�E�ƀ�    �E��   ����������RP��!  ���E��   ��P�H!  ���P��E����   <fuy�E��   ��P�"!  ���P��E����   <euS�E��   ��P��   ���P��E����   <lu-�E��   ��P��   ���P��E����   <.u�   ��    ��t�E��@]���u��u���   ���������E��M܍�������D�����j WQRPj��  �� �m䀁}�  �r����E� �E�
   �b�����������P�.  ��������tl��������u��Y��������u���u��w  ��뼋�������u���������f�Eҋ�����f�E��E҉��EЉƃ�VS�u��d  ���y������u��  ���f����U����E���uP�   ����ÐU����E���u�u�u�u�uP�Q  �� ���E���ÐU����E�@ �E�@]��t�E�   ��j j j j Pj�   �� ��ÐU��E�     �E�@    �]ÐU�����j�  ���E��E�    �E�    �E�    ���E�P�������E�U��U�P�U��P�E�U�P�E� ��u
�E�U���E�@�U��E�P�E�P�E�U�P�E�@�P�E�P���U��WVS�   �+  �E�]�M�U�u�}�i�[^_]Ë$�U��������[+  �E�    ��U�E�ЋU��E��E�;Er�E��U�������$+  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���{  �ï*  �E���E�E���$   �E�    ��Ѕ�u��$   �E�    ���E����$   �E�    �����E䋃(   9E�s	��(   �E���u��8  ���E��}� u%��d  ��h  ���� ��d  ��h  �    �l�E��     �E��@    �E��U�P��$   �E�E��P�E��@   �E��@    �E��@�ƿ    �����P� ��������Q�E��e�[^_]�U��WVS��L�U  �É)  �E�    �E�    �E�    �E�    �E�E��E� �#  �}� u5��d  ��h  ���� ��d  ��h  �  ��j�������  ��\  ��u-���u��K�������\  ��\  ��u��  �    �{  ��\  �E��E�    ��`  ���C  ��`  �P��`  �@)ЉE��E�    �E����    ;E؉�E��
  ��`  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ�`  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u��\  �E��E�    �|  ���u��9������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���N  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u��\  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������O  �    �e�[^_]�U��WVS��,�!  ��U"  �} u#��d  ��h  ���� ��d  ��h  �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx��l  ��p  ���� ��l  ��p  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��t  ��x  ���� ��t  ��x  �Y  �  �E��@�E������P� �M��I�ο    )��������Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ��\  9E�u�E܋@��\  ��`  9E�u
ǃ`      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋������P� �M܋I�ο    )��������Q�E܋@��P�u��p  ���G��`  ��t=��`  �P��`  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉�`  ��  �e�[^_]�U��S���o����  �U�U�U�U��R���%������E��E��Pj �u��?������E��]���U��S���Z  �Î  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E���  �E���E�E�@=���tz��l  ��p  ���� ��l  ��p  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��t  ��x  ���� ��t  ��x  �~  �    �_�E�@�E�E�;Er�E�U�P�X  �E�;�N  ���u��������E���u��u�u����������u��������E�]��Ë$�U��S������$  �M�U��j j j QRj���q����� �E�]���U��S�������  �U�U�U�U���j j �u��u��uj���0����� ��]��ÐU���H����  �]�U���8����  �]�U���(����  �]�U��S���J�����~  �E��P�H  ������P�E���]��ÐU�������L  �]�U��S��������8  �E��P�  ���� ��P�E����u��  ���E�PX�E�����uP��  ���E�U�P�U�P�U�P�U�P��]��ÐU��WVS�������ú  �E�@���w  �E�@��������p��E�@�H��E�@�P�E�@���uh�   h�   h�   VQRP�|
  �� �E�@��������p��E�@�H��E�P�E�@�������E�@���uh�   h�   h�   VQRP�#
  �� �E�@�H��E�@�U�R���uj`j`j`jQPR��	  �� �E�@�H��E�P�E�@ЍP��E�@���uj`j`j`jQRP�	  �� �E�@�H��E�@�P�E�@�uj`j`j`QjRP�	  �� �E�@�H��E�@�P�E�p�E�@����uj`j`j`QjRP�U	  �� �r  �E�@��������p��E�@�H��E�@�P�E�@���uh�   h�   h�   VQRP�	  �� �E�@��������p��E�@�H��E�P�E�@�������E�@���uh�   h�   h�   VQRP�  �� �E�@�H��E�@�U�R���uj`j`j`jQPR�~  �� �E�@�H��E�P�E�@ЍP��E�@���uj`j`j`jQRP�E  �� �E�@�H��E�@�P�E�@�uj`j`j`QjRP�  �� �E�@�H��E�@�P�E�p�E�@����uj`j`j`QjRP��  �� �E�P�E�@�������Ѓ��ƋE�P�E�@�������E�@X��)ЉE�����uj j j VRP�  �� ��e�[^_]�U�������L  �E�@�]ÐU�������4  �E�@ �]ÐU������  ��(��P�E��]�U��S�������  ���u���Q������]���U��S���j����  ���u���+������]���U��S���D����  ���u���9�������]���U��S�������  ���u����������]���U��S�������`  ���u�����������]���U��S�������9  ���u����������]���U��S������  �M�U��j j j QRj���_����� �E�]���U��S���r����  �U��j j j j Rj!���+����� ��]���U��S���@����  �M�U��j j j QRj��������� ��]���U��WVS��,�@�����t  ���u�E������E��h�   �J������Ɖ��    �*   ����V��  ���u��E��U�P�E��U���ֺ   �ǉ��E�@���EЋE�@���EԋUЋE�������P�G������E܋E��Uȉ��   �Ủ��   �UЉ��   �Uԉ��   �U؉��   �U܉��   �E��e�[^_]�U��VS�V����Ê  �E�@��P�������u��t��V�@  ����h�   V��������e�[^]�U��S��������:  �E���   �E�@�ЋE�@����Q�M���   RPj j �  �� �E�    �E��P�M  ��9E�����t0�U�E��RP�F  �����M���   ��QP�҃��E�뷋E���   �E�@��RP���������]���U��S��$�J�����~  �E�    �E��P��  ��9E�������   �U�E��RP�  ���P�U�P�U�P�U�@�E��U�E9�}Y�U�E9�}O�U�E�E9�~@�U�E�E9�~1�U�E��RP�a  ��������P�҃��E�U􉐤   �	�E��L�����]���U��S���A����  �U���   �ыU��QR���  ��������P�҃���]��ÐU��S�������f  �U��R���Y   ���Eƀ�   ��Eƀ�   ��Eƀ�   ��Eƀ�   ���]���U��S������  �U��R���-   ����]���U�������  �E�     �E�@    �]ÐU��S���������  �E� �E�E� ��t���u��E������琋]��ÐU���*����  �E�@]ÐU�������{  �E�@9Er	�    � �+�E� �E��E�    �E�;Es�E�� �E��E���E��@��U�������-  �    ]�U������  �����  �    ]�U��S�������  �M�U��j j j QRj���E����� �E�]���U���\����  �    ]�U����E����  �E�������E����	��E����	��E��	ЉE�E�@�E��E�    �E9E�}G�E�    �E9E�}2�U�E�E�@�M�U��Ѝ�    �E�E��E��ƃE�뱐��U��S������  �U��j j j j Rj ���[����� ��E�]��� U����l����  �M�U�E �M�U�E�} y�EE�E    �} y�EE�E    �E������E���	��E�	ЉE�E$�@�E��E�    �E�;E}k�U��EE$�@9�}Y�E�    �E�;E}D�U�E�E$�@9�}2�U��EE$�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��������  �} y�EE�E    �} y�EE�E    �E�������E����	��E��	ЉE�E�@�E��E�    �E�;E}k�U��EE�@9�}Y�E�    �E�;E}D�U�E�E�@9�}2�U��EE�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��� ����  �E�E�E�E��E��}��E��f�E��m��]��m��E��E�������v�E�����E���U��S��4�7  ���  �U���������P��H����E��Eԃ��d$��$���l��������E��E�    �E�   �E�    �E�;E��   �E�    �E�;E��   �U�E�E�@�������U�E���E�ȉE��U���ЉE�E��E�P�E�����U���ЉE�ЍP�E��E�@�U�������U���ЉE�ЍP�E��E�@�U�������E��F����E�E�E��$�����]��Ë$�U��WVS��<�>�����r  �u�M�U�}���EԈMЈỦ��E��E�    �}���   �U�������E��� ���E��E�    �}�]�E�   �����#E܉E������Ѕ�t7�}��u��MЋE� �EE�EċE�E��u WVQjjRP������� �E�띃E��f�����e�[^_]�U��WVS��,�.����  �EȋM�U�E�MԈUЈE��E�    �E� ��tC�}��u��]ԋM�U�EЉE� �����u WVSQRP�]������� �E��E볐�e�[^_]�U�������  �E�    ��E��U��E�� ��u�E���U��S���������  �E�    ��U�EЋM�U�� ��E����u������9E�|Ԑ�]���U��S���c����×  ���u�e������EЃ��uP�������E�]��� /           t����       zR |�        Z���    A�BW�     <   V���1    A�Bm�     \   h���9    A�Bu�     |   ����   A�BI���   �   b���    A�BU�     �   \����    A�B�� (   �   ����*    A�BC���`�A�A�A�      ����            ����7    A�Bs�     <  ����r    A�Bn� ,   \  /���&   A�BF����A�A�A�   ,   �  %���4   A�BF���'�A�A�A�   ,   �  )���~   A�BF���q�A�A�A�       �  w���K    A�BD�C��       ����f   A�BD�^��   4  ����           H  ����6    A�BD�n��      l  ����?    A�BD�w��     �  ����    A�BL�     �  ����    A�BL�     �  ����    A�BL�     �  4���    A�BZ�        ����5    A�BD�m��     4  ����    A�BL�      T  ����{    A�BD�s�� ,   x  ���t   A�BF���g�A�A�A�      �  L���    A�BS�     �  D���    A�BS�      �  Z���&    A�BD�^��        \���&    A�BD�^��      0  ^���'    A�BD�_��      T  a���'    A�BD�_��      x  d���'    A�BD�_��      �  g���'    A�BD�_��      �  j���6    A�BD�n��      �  |���2    A�BD�j��        ����4    A�BD�l��      ,  ����P    A�BD�H�� (   P  v����    A�BF�����A�A�A�    |  ����(    A�BD�`��  $   �  ���N    A�BB��F�A�A�    �  :����    A�BD����     �  �����    A�BD����       ����D    A�BD�|��     4  ���#    A�B_�      T  ���9    A�BD�q��     x  4���    A�BQ�     �  *���Q    A�BM�    �  [���    A�BP�     �  O���    A�BY�      �  L���6    A�BD�n��       ^���    A�BP�     <  R����    A�B��     \  ����7    A�BD�m��     �  �����    A�B��    �  �����    A�B��    �  p���Q    A�BM�     �  ����C   A�BD�;��     ����       (     �����    A�BF�����A�A�A�(   D  ^����    A�BF���x�A�A�A�   p  ����1    A�Bm�      �  ����M    A�BD�E��     �  ����>    A�BD�v��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      t�� �        �����        ������                                                                                                                                                                                                                                                                                                                                         <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;              GCC: (GNU) 8.2.0                        ��          أ          �           �          <�          `�          ��                                ��p  ��                   ��            ���            ��   ��     %   ��     /   `�     :   d�     F   ��     U   ��     b   ��     u   ք7     �   �r     �   �&    �   ��4    �            ���            ���            ���            ���            ���            ���            ��             ��  <�        ��     /  ��     ;  $�7     M  L�M     T  �6     s  t�t    �  ��     �  �   "  �  T�2     �  ��   "  �  ��*     �  f�9   "  �  �       �6     �  ��       6�&     "  f�9   "  9  ��5     M  �   "  h  ��{     }  ��     �  B�?     �  ���     �  ��4    �  j�   "  �  ҄     �  �        �   "    �(   "  *   �   !  6  ��'     =  �   !  J  ���     o  �(   "  ~  �     �  ��1   "  �  �     �  B�#   "  �  ��{     �  W�K     �  ʛP   "    ��>     	  ʛP   "    �   "  '  ���     B  ��     �  ��      \  ��5     p  8�6       ��'     �  ��f    �  D��     �  �     �  ���     �  u�C      [��     '  ��N     A  ��Q   "  X  (�   !  d  ���     �  ��      �  ���     �  ��     �  $�Q     �  З'     �  ܣ   !  �  ��4        ��       n�     )  ���    /  \�&     5  ��9   "  Q  ��     h  ��      o  ��      t  ��D     �   �     �  �1     �  B�#   "  �  ��'     �  ��   "  �  ��1   "  $  ٍ~     fm.asm main.cpp syscall.c l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 ipc.c widgets.cpp window.cpp _liballoc.c graphics.cpp text.cpp string.c _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx l_allocated _Z12GetVideoModev strcpy _Z13_CreateWindowP10win_info_t _ZN6Button5PaintEP7Surface l_max_inuse _ZN6WidgetC1Ev _Z14_DestroyWindowPv _ZN4ListIP6WidgetE8add_backES1_ syscall _ZN4ListIP6WidgetED2Ev liballoc_unlock ReceiveMessage _Znwm _ZN4ListIP6WidgetED1Ev _ZN7TextBoxC2E4Rect _ZN8ListNodeIP6WidgetEC2Ev _ZN6ButtonC1EPc4Rect l_inuse SendMessage _Z11PaintWindowP6Window malloc _ZN6Window9AddWidgetEP6Widget __x86.get_pc_thunk.ax _ZN7TextBox5PaintEP7Surface _ZN8ListNodeIP6WidgetEC1Ev _ZN6WindowD1Ev _ZTV6Button _ZdlPv _ZTV7TextBox _Z15HandleMouseDownP6Window8Vector2i _ZN6WindowD2Ev liballoc_lock _ZN10FileButtonC2EPc4Rect _ZN6Button11OnMouseDownEv _ZN4ListIP6WidgetEC1Ev _ZN6ButtonC2EPc4Rect calloc _ZN6WindowC1Ev strcat _ZN6WindowC2Ev _ZN6WidgetC2Ev _Z8DrawCharciihhhP7Surface _ZN6Widget11OnMouseDownEv _ZN7TextBoxC1E4Rect liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx _Z12CreateWindowP10win_info_t _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window _ZN4ListIP6WidgetEixEj _ZTV6Widget _Z10DrawStringPcjjhhhP7Surface __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface font_default _Z5floord _ZdaPv _ZTV10FileButton _Z12_PaintWindowPvP7Surface _ZN6Widget5PaintEP7Surface liballoc_free pmain _Znam _ZN10FileButton9OnMouseUpEv _ZN6Widget9OnMouseUpEv _edata _end _Z13HandleMouseUpP6Window _ZN6Button9OnMouseUpEv strlen _ZN4ListIP6WidgetEC2Ev _ZdaPvm _ZN4ListIP6WidgetE10get_lengthEv _ZN10FileButtonC1EPc4Rect  .symtab .strtab .shstrtab .text .rodata .eh_frame .data.rel.ro .got.plt .data .bss .comment                                                   ���   W#                 !         أ�#                    )         ��#  �                 3          � 0  <                  @         <�<0                   I         `�`0                     O         ���4  <                  T      0       �4                                 �4  P  
   "         	              �;                                 �B  ]                  