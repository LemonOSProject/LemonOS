ELF              ��4   _      4    (           � ��@  �@           �@  �����
          �W  �R3  �                 �    UU���#  VW�����_^�  �    �i���f�f�f�f�f���=�t$�    ��tU���h��Ѓ��Í�&    f�Í�&    ��&    ���-����������t(�    ��tU���Ph��҃��Í�&    �t& �Í�&    ��&    ��= � ugU�$���V���S����������9�s�v ���$����$�9�r��'����    ��t��h@��Q~����� ��e�[^]�Í�&    ��&    ��    ��t'U���h(�h@��~������	�����&    f������U����i�mN�A90  ��������%�  ]�U��S���T����9�sz�U��E��j j j RPj�0  �� �E���    �H��L�)�Ӊȉ�i��  �M��P�)щ�¡T�УT��E��    �H��L��E�P��w����T�    ��]���U��WVS����j�  ���ǃ�W�/  ���=\��\��E�   �E�   ���u��u�P�B  ���\��	   �   ��VSP�%  ���@�    ��������������e�[^_]ÍL$����q�U��WVSQ���  �ȋ ��T�������p���P�c
  ��fǅt��� fǅv��� fǅp���@ fǅr���  ǅx���    ��j�  ���Ã�S�D
  ���\��\��   �   ��WVP�_
  ���\�ǅ���	   ǅ���   ������������P�.
  ���E�    �}�.�E�    �}��E����E��`��  �E��߃E��̃���p���P�7  ���E������@���tR�`���t+�`����`�������� ��� ������@�    ����������������\���P�-  ����������   ��d�����ui�X���t�X� ������h���=  t)=  w	=
  t�=  t=  t��E�    �>�E�   �5�E�   �,�E�   ��"��d������^������u��4  ���-  �F����X����C  �E�    �}�.�E�    �}��E����E��`��  �E��߃E��̡d���t�   ��   ���������`���E�    �\���P��  ��9E�����t[�\��EЍ�������PQR�  ���������\��EЍ�������PQR�  �������������`�� �E���E�    �}���   �E�    �}���   �Eč��   �E����E��`�� ���������E����E��`�� �������؋E����E��`�� �������ЋE������E���WVSRjjQP��  �� �E��[����E��A����}���   �}��}� t�  �}��W  �}���  �  �\��\���P�`  ������������RSP��  ���\��\���������j RP�2  ���������� ����\��������j RP�  �����������$�������$����� ���S�  ����  �\��\���P�  �����������RSP�9  ���\��\��������j RP�  �����������(����\��������j RP�d  ���� �����,�������,�����(���S��  ���D  �\��\���P�  ������$�����RSP�  ���\��\���,�����j RP��  ����,�������0����\���4�����j RP��  ����8�����4�������4�����0���S�<  ���   �\��\���P�t  ������<�����RSP��  ���\��\���D�����j RP�F  ����D�����8����\���L�����j RP�  ����P�������<�������<�����8���S�  ����\���T�����j RP��  ����T����\���\�����j RP�  ����`��������`�� <��   �\���d�����j RP�  ����h�����xq�\���l�����j RP�^  ����l�����xL�\���t�����j RP�9  ����x�����&�\���|�����j RP�  ����|�����~�   ��    ��t]�X��E��   ��Ph�   h�   h�   j j h��_  �� �E��   �Eċ@��j j j RPj�'  �� �~  �\��E���j RP�  ���]��\��E���j RP�h  ���U������`�� <������   �\��E���j RP�1  ���]��\��E���j RP�  ���U������`��  �����������������������������������t�d�   �
�d�    �\�ǅ@���    ǅD���    ����D�����@���P��  ���B  �\��E���j RP�r  ���]��\��E���j RP�W  ���U������`�� <������   �\��E���j RP�   ���]��\��E���j RP�  ���U������`��  �@�   ����`���������������������������������������������������)Ѕ�����t�d�   �
�d�    �\�ǅH���    ǅL���    ����L�����H���P�   ���E��   �Eċ@��j j j RPj�%  �� ����������U��Ef�   �Ef�@  �Ef�@  �Ef�@  �]ÐU��E�     �E�@    �E�@    �]ÐU��E�     �E�@    �]ÐU��S����j�  �����    �C    �C    �C    ��S�������]�E��     �M�E�U�A�Q�E� ��u
�E�U���E�@�U��E�P�E�P�E�U�P�E�@�P�E�P��]���U��E�@]ÐU����E�@��t�E�@9Es	�E� ��u�E� �M�P�@��Q�J�E� �E��E�    �E�;Es"�E�@9E�s�E�� ��t�E�� �E��E��֋M�E��P�@��Q�E�� U���(�E�@��t�E�@9Er�M�E��U��Q��   �E� �E��E�    �E�;Es"�E�@9E�s�E� ��t�E� �E�E��֋E�P�@�E�U�E� ��t�E�@��t�E� �U�R�P�E�@��t�E� ��t�E�@�U���} u
�E��E��E�@�P��E�P�E�@9E����t�E�P�E�P���u���  ���M�E�U��Q�E�� �U��S����j�
  �����    �C    �C    �C    ��S�`������]�E��     �M�E�U�A�Q�E�@��u�E�U�P��E� �U�P�E��E��E�U��E�@�P�E�P��]���f�f�f�f�f��UWVS�
  ��??  ���|$$�D$ �l$(	��t��UW�t$,�L   �������)�����RW�t$,�  ����u
��[^_]�f����VW�t$,�V�   ����[^_]�f���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���D$4�|$,�L$$�\$8�T$0�t$(�|$�ǉL$�ȁ�   ���	���% �  ���͉���	�k	ǅ�~o;s}j�L$�D$�T2��T$�D��$��D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�~  �ñ=  ���t$j j j j Vj ��  ��$��[^� f�UWVS���|$�t$ �l$(�D$,�\$0�L$4�T$8��y|$$1���y�1�����������	�	��B�D$��~j;r}e�D.��$�D$$�\���&    f��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS���|$�t$ �\$(�D$,�T$0��y|$$1���y�1���������� �  ��	�	��B�D$��~m;r}h�D��$�D$$�\���&    �t& ��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS�  ���;  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$��������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�<  ��o:  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�<����� 9t$h�_�����L[^_]Í�&    UWVS�l  �ß8  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�l����� 9t$l�_�����L[^_]Í�&    UWVS�  ���6  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�������9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$�f�f�f��S�   �������5  ���D$��D�P�
  ��[Í�&    �S�������4  ���t$�w
  ��[Ív S�������4  ���t$�  ��[Ív S�����ò4  ���t$�������[Ív S�_����Ò4  ���t$�K  ��[Ív S�?�����r4  ���t$�+  ��[�f��UWVS������O4  ���D$<�|$8�t$0�D$�G�D$�D$D���� ��D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������� ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�]����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ�*����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��������t$H���t$�t$�D$PjjW�D$P����P������ 9|$�b�����[^_]Í�&    f�UWVS�������1  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��S�?�����r1  �� j j j �t$4�D$$Pj�  �D$,��8[�f�S������B1  ��j j j j �t$(j!�  ��([Í�&    f�S�������1  ��j j j �t$(�t$(j�N  ��([Í�&    UWVS�������0  ��(�l$<U�T����$�   �D$�����+   �T$����1����FjtUPǆ�   ����ǆ�   �����V�  �}�m����    ���� ��f��� vf��� wd���   ������P��  �����   ���   ���   ��ǆ�       ǆ�       Ɔ�    Ɔ�    ��[^_]Í�&    ��&    �ȃ���P�  ��롍�&    ��    S�������/  ���D$�p�u�����[��  �³/  UWVS���l$0�T$�Eu(�����   S�����   �EP�EPj j ������ �E���   ��~?1����   �v 9�v\�M ��t1��v ���	9�u��A�������WP��E��9�̋��   ��t	��S�Ѓ���S�u�\$�������,[^_]Ð�    ��&    f�UWVS���D$0�l$4�|$8�p��~G� 1ۉD$��&    ��&    9�t<�D$��t1�f���� 9�u��@�P�H9�~9�|&��9�uσ�[^_]Í�&    �    ��&    f�H9�~�P9�~̅�t�T$1���&    ����9�u��T$�D$���@�P�R�D$@�����   ��[^_]Í�&    ��&    S���\$���   ��xn;CsY���t1Ґ���	9�u��A���P�R���   ��;Ss-���t1��t& ����	9�u��A��[Í�&    ��&    ��    ��&    f�ǃ�   ������1�[Í�&    ��&    �VS�.�����a-  ���t$ j�%����T$ ���     �P��@    ��t�V��P�F�F��[^Ív ��F�F��[^Ë$�f�f�f�f�f�f���U����  �,  ǀ�      ǀ�      ǀh
     ǀl
      ��h��    �B    ��p��    �B    ��x��    �B    ǀ�      ǀ�      ǀ�      ǀ�      ǀ       ǀ      �]�U����9  ?,  �E�    ��U�E�ЋU��E��E�;Er�E��U����  ,  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���`����Ó+  �E���E�E���h
  �E�    ��Ѕ�u��h
  �E�    ���E����h
  �E�    �����E䋃l
  9E�s	��l
  �E���u��  ���E���jj �u���������}� u%���  ���  ���� ���  ���  �    �l�E��     �E��@    �E��U�P��h
  �E�E��P�E��@   �E��@    �E��@�ƿ    ��h��P� ����h���Q�E��e�[^_]�U��WVS��L�(�����[*  �E�    �E�    �E�    �E�    �E�E��E� ��  �}� u5���  ���  ���� ���  ���  ��  ��j�������  ���  ��u-���u��9��������  ���  ��u�  �    �{  ���  �E��E�    ���  ���C  ���  �P���  �@)ЉE��E�    �E����    ;E؉�E��
  ���  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ��  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u���  �E��E�    �|  ���u��'������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��p��P� ����p���Q��x��0�x��p��P� 9Ɖ��s�Ɖ���x��0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���J
  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��p��P� ����p���Q��x��0�x��p��P� 9Ɖ��s�Ɖ���x��0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���	  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    ��p��P� ����p���Q��x��0�x��p��P� 9Ɖ��s�Ɖ���x��0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ���  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    ��p��P� ����p���Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ���  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u���  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������  �    �e�[^_]�U��WVS��,�������'#  �} u#���  ���  ���� ���  ���  �9  �E��� ���E�}�w	�E+E�E�  �E���E��E��@=���tx���  ���  ���� ���  ���  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��   ��  ���� ��   ��  �  �  �E��@�E���p��P� �M��I�ο    )����p���Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ���  9E�u�E܋@���  ���  9E�u
ǃ�      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋���h��P� �M܋I�ο    )����h���Q�E܋@��P�u��(  ���G���  ��t=���  �P���  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉��  �  �e�[^_]�U��S���  �   �U�U�U�U��R���%������E��E��Pj �u��-������E��]���U��S���-�����`   �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E��  �E���E�E�@=���tz���  ���  ���� ���  ���  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��   ��  ���� ��   ��  �6  �    �_�E�@�E�E�;Er�E�U�P�  �E�;�  ���u��������E���u��u�u����������u��������E�]��Ë$�U���������  �E�E���E��P�U��U��E�P��U��u�E��U��� �����  �E�E��E�E��E�E��"�E��P� �M���Q�E��E��m�E�E�}�w؋E�E���E���E���E��E��m�E�E��}�wދE�E���U��E�ЋM��U��� ��m�E�E�}� uۋE��U��S������  �M�U��j j j QRj���Q   �� �E�]���U��S��������  �U�U�U�U��U�U��j �u��u��u��uj���	   �� ��]���U��WVS�����  �E�]�M�U�u�}�i�[^_]�U��S���j���p  ��j j j j j j�������� ���U���A���G  �    ]�U���-���3  �����  �    ]�U��S������  �M�U��j j j QRj���M����� �E�]���U��������  �    ]�f�f�f�f�f�f�������t6U��S�������&    �v �Ѓ�����u��[]Í�&    ��&    ��:����     Game Over, Press any key to Reset          zR |�        ����'    A�Bc�      <   �����    A�BD���� (   `   (����    A�BF�����A�A�A�   �   "���)    A�Be�  ,   �   o����
   D Gu Fupu|uxut   �   ����#    A�B_�     �    ���    A�BU�        �����    A�BD����    @  v���    A�BG�     `  b����    A�B��    �  ����   A�B�    �  �����    A�BD���� |   �  H���~    A�A�A�A�N U$A(A,D0H E$K(A,D0H G
A�A�A�A�CC$C(A,G0H CA�A�A�A�     D  H���?    Cy 8   \  p����    A�A�A�A�C$�A�A�A�A�8   �  ���.    A�A�NFB B$B(A,B0HC�A� 8   �  �����    A�A�A�A�C�A�A�A�A�8     �����    A�A�A�A�C�A�A�A�A�<   L   ���b   A�A�A�A�NPL@�A�A�A�A�X   �  P����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   �  �����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   D  8����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   �  �����    A�A�A�A�C(�A�A�A�A�   �  U���           �  L���(    A�SJ HA�       X���    A�ND HA�     (  T���    A�ND HA�     L  P���    A�ND HA�     p  L���    A�ND HA�     �  H���    A�ND HA�   �  D���W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   �  ����s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�  0   $  ����.    A�N(B,B0B4D8E<B@LA�  0   X  ����'    A�NBB B$B(D,B0HA�  0   �  ����)    A�NBB B$D(D,B0HA�  `   �  ����   A�A�A�A�N<E@a4M8A<A@g0g<G@H0y
A�A�A�A�OE<D@H0      $  X���     A�NG HA� x   H  T����    L�A�A�A�C0Q8G<H@EDEHBLBPH0w8H<A@H0Q<A@E0C8A<C@LA�A�A�A�B0����X   �  �����    A�A�A�A�C0]
A�A�A�A�HD<F@J0IA�A�A�A�0    	  ,����    A�CkC La
A�P]C� <   T	  ����_    A�A�NF Lh
A�A�DLA�A�      �	  ����          �	  �����    A�B��    �	  B���7    A�Bs�     �	  Y���r    A�Bn� ,   
  ����8   A�BF���+�A�A�A�   ,   8
  ����4   A�BF���'�A�A�A�   ,   h
  ����~   A�BF���q�A�A�A�       �
  ���K    A�BD�C��     �
  ,���f   A�BD�^��   �
  n���          �
  ^���8    A�Bt�       v����    A�B��     4  ����6    A�BD�n��      X  ���F    A�BD�~��  (   |  2���*    A�BC���`�A�A�A�    �  0���-    A�BD�   �  A���    A�BP�     �  5���    A�BY�        2���6    A�BD�n��     (  D���    A�BP�      ����    ����                                                `�`�@@@�@@@�@@ �`�`�S   S      d                                                                                                                                                                                                                                                                                                <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              ��                           >        ����    src/gfx/sse2.asm NASM 2.14.02 ���     %  . @   :    '   �       src/gfx/sse2.asm      ��                                         t�          ��          �          �          @�          ��          ��          ��          ��     	      �     
                                                                                                                             ��   ��         ��      (   @�      ;   ��      =    �      P   P�      f    �    
 u   $�    
 �   Ё      �   (�    
             ���   ��      �   ��      �   г      �            ��  ��                  ��           ��#           ��/           ��8           ��C           ��L           ��           ��]  ��    
 g  ��    
 q   �    	 |  �    	 �  ��    
 �  ��    
 �  ��    
 �  N�7     �  ��r     �  ��8    �  /�4    �           ��           ��           ��           ��           ��             ��)  ��      ?  h�    
 K  ��.     ]  ��    �  \�    
 �   �.     �  ���   "  �  @�   "  �  x�    
    P�'       `�    
 "  �*     *  ���     8  ]�     H  v�6     �  ��    
 W  p�(   "  ]  ��    	 m   ��    �  α�     �  p�    
 �  �    	 �  ��F     �  ��     �  ��     �  /�4    �  ��    	 �  Z��   "    ��     1  ��    	 >  P�    
 K  ��   "  R  ,��     [  ��     q  ���     2  t�      �  I�     �  ��    	 �  @�   "  �  @�    
 �  �)   "  �  �K     �  P�~       X�    
   �#   "  ,  @�W    G  �)   "  �  ��&     [  0�_     x  ��    	 �  z�6     �  ��   "  �  ,�f    �  ���     �  e�     �  `�    
 �  ��      ��    	   ��b    >  ��     Z  ��      t  ��    	 ~  ��s     �  ��  "  �  ̂�     �  H�    
 �  �     
 �  ��     �  ��8       _��
       �    	   Б?     '   �   "  .  T�    
 8  �      >  �#   "  V  ��)     r  �'     {  ��     �  d�    
 �  ��   "  �  ��    	 �  ��   "  �  �     	 �  ��     
 �  ���     �  �-     �  ��   "    ���     8   �    	 A   �   "  I  ��      U  p��     �  c�~     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp graphics.cpp runtime.cpp text.cpp window.cpp font.cpp src/gfx/sse2.asm l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 memory.c ipc.c syscall.c exit.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface snake _Z13_CreateWindowP10win_info_t _ZN4ListI8Vector2iE9add_frontES0_ _ZN8ListNodeI8Vector2iEC1Ev l_max_inuse _Z14_DestroyWindowPv powerUpTimer syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm bgColourDefault _Z12DrawGradientiiii10RGBAColourS_P7Surface l_inuse __TMC_END__ SendMessage __DTOR_END__ _Z11PaintWindowP6Window malloc frameWaitTimeDefault _ZN4ListI8Vector2iE8add_backES0_ __x86.get_pc_thunk.ax __dso_handle lastUptimeMs _ZdlPv _Z4Waitv __x86.get_pc_thunk.dx _Z15HandleMouseDownP6Window8Vector2i liballoc_lock frameWaitTime _ZN8ListNodeI8Vector2iEC2Ev powerUp _ZN10win_info_tC2Ev calloc _Z16memcpy_optimizedPvS_m gameOver _ZN4ListI8Vector2iEC2Ev _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev _Z9AddWidgetP6WidgetP6Window applePos liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx snakeMapCells _Z12CreateWindowP10win_info_t powerUpTimerDefault _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window rand_next _Z10DrawStringPcjjhhhP7Surface _ZN4ListI8Vector2iE9remove_atEj _Z5Resetv lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface main font_default _Z5floord _ZdaPv msCounter _fini _ZN4ListI8Vector2iEC1Ev _Z12_PaintWindowPvP7Surface _Z4randv liballoc_free fruitType _Znam snakeCellColours _ZN4ListI8Vector2iE6get_atEj _edata _end _Z13HandleMouseUpP6Window exit _ZN4ListI8Vector2iE10get_lengthEv _Z10surfacecpyP7SurfaceS0_8Vector2i font_old _ZdaPvm memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                   t�t                     !         ���   �3                 '         �4                    -         �4  "                  5         @�@4  H                 ?         ���@                    F         ���@                    M         ���@                   V         ���@  H
                  \          �K  �                  a      0       K  +                 j              3K                     y              SK                    �              eK  B                  �              �K                    �              �K  >                  �               L                    �              L                                  L  �	     >         	              �U  �                               H^  �                  