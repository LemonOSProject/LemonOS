ELF          >    � @     @       Ȇ          @ 8  @                   @       @     �:      �:                    @       @@      @@     h      �             �+  �v0  �     H��    UUH��������
  ����    �hL@ H=hL@ t�    H��t	�hL@ ��f��ff.�     @ �hL@ H��hL@ H��H��H��?H�H��t�    H��t�hL@ ���ff.�     @ �=)K   uwUH�'K  H��ATA�@@ S�@@ H��@@ H��H��H9�s%f.�     H��H��J  A��H��J  H9�r��0����    H��t
��1@ �<���[A\��J  ]��ff.�     @ �    H��tU��L@ ��1@ H������]����D  ����UH��AVAUATSH��   H�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸ M@ A�    A�    H�ƿ   �J.  �h  ��?  ���  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H���,  H��P���H�E��@����H��X���H�    ����H!�H	�H��X���H��X�����H�       H	�H��X���H��P���H��X���H��H��H�й M@ ��H��H���  �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H���p  H��`���H��h���H�    ����H!�H��H��h���H�E��@������H�� H��h�����H	�H��h���H��`���H��h���H��H��H�й M@ ��H��H����  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H���  H��p���H�E��@������H��x���H�    ����H!�H	�H��x���H��x�����H�       H	�H��x���H��p���H��x���H��H��H�й M@ ��H��H���  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H����  H�E�H�U�H�    ����H!�H��H�E�H�E��@������H�� H�U���H	�H�E�H�E�H�U�H��H��H�й M@ ��H��H���h  A�    A�@�@   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H���  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A� M@ D���H��H����  H�E����   ����H�E����   ����H�E�H��H��h M@ A��   A��   ��   H����  H���E�   �E�   H�E�H���   H�E�H��H���D  H�E�H�E�H�U�H�� M@ A�    A�    H���   ��)  H�e�[A\A]A^]�UH��SH���  ��L@ ��  H��E  H��E  H��H��H��E  H���E  �H��E  f�HH���  H��H�E�H�E�H�H�HH��E  H��E  H�PH�HH��E  H��E  H�@ H��E  ��E  ��E  ��H�H���d  H��E  H�E��PH�E��@�u�h�   A�    A��   �щ¾    �    �X  H��A�    A�    �    �    �    �   �(  H��`���H���f  H������H���%  fǅ����d fǅ����d fǅ����
 fǅ����
 H������H��H�Test WinH�0�@dow ǅ����    H������A�    A�    �    �    H�ƿ   �*(  �y1@ A�    A�    �    �    H�ƿ   �(  �    ��1@ �c  �E��E��   �(M@ ���  H������A�    A�    �    �    H�ƿ   �'  ������9E���  �������E��E�    �E�;E���  �E� H��`���H����	  �E�Hc�H��`���A�    A�    �    H�ƿ   �I'  H������H�E��E�    H��`���H���
  9E�����t.�U�H��`�����H��� 
  H� H9E�����t�E���E���Eۃ����  ��   �  H�E�H�E�H��`���H��h���H�PH�HH��p���H��x���H�PH�H H������H������H�P(H�H0H������H������H�P8H�H@H������H������H�PHH�HPH������H������H�PXH�H`H������H������H�PhH�HpH������H�Px���������   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�U�H��`���H��H���A	  �d7  �E��0����T7  ��t,�B  �B  A� M@ D�87  �щ¾    �    �  �E�    �E�;E�}*�U�H��`�����H���_  H�E�H�E�H�������E�����6   �E��   �(M@ ����  ��6  ��A  ��Љ�6  ��6  ��A  ��)Љ�6  �xA  ��u�nA  ��t��6  �^A  ��to�o6  �a6  �KA  )�H�E����   �M6  �7A  )�H�E����   H�E����   ��yH�E�ǀ�       H�E����   ��yH�E�ǀ�       ��@  �������J  ��@  �����8  ��@  H��`���H���  ���Ẽ}� �  �U�H��`�����H���  H�E���5  H�E����   9���  �|5  H�E����   H�E��@���9���  �[5  H�E����   9���  �C5  H�E����   H�E��@���9��w  �U�H��`�����H���  H��H��`���H��H����  H�E�H�E���4  H�E����   �P��4  9�|LH�E��@����u>��4  H�E����   )�4  H�E����   )��ȉ�?  ��?  �v?  ��   Hǅp���   H�E��@����t0�f4  H�E����   )ЉEȋS4  H�E����   )ЉE��4�64  H�E����   )Ѓ��Eȋ 4  H�E����   )Ѓ��Eĺ    �Eȉ���Eĉ�H��x���H�E�H�@|H������H�E�H�@tH����������x�����p�����h�����`���H���O  H��0�	�m��������>  ����t�w>  ��t�l>   �d>  ����  �R>  ��������  �@>   �:>   H�}� ��  �=3  H�E����   9��l  �%3  H�E����   H�E��@���9��G  �3  H�E����   9��/  ��2  H�E����   H�E��@���9��
  ��2  H�E����   �P��2  9�|H�E��@������   Hǅp���   H�E��@����t0�z2  H�E����   )ЉE��g2  H�E����   )ЉE��4�J2  H�E����   )Ѓ��E��42  H�E����   )Ѓ��E��    �E�����E���H��x���H�E�H�@|H������H�E�H�@tH����������x�����p�����h�����`���H���c  H��0�E�    H��`���H����  9E�������   �E� �E�    �E�;E�}|H��`���H���m  �E�Hc�H��`���A�    A�    �    H�ƿ   �  H������H��x����U�H��`�����H���  H� H9�x�������t�E��	�E��|����E�����t�U�H��`�����H���  ��0  �E��%���H��0���H���>  H��������   H��@���H=� u�H�}� ��   H��H���H����   H��H���H��H��t6H��H�����H��t'Hǅp���   H��H�������@@@ H�H��x����"Hǅp���   H��H�����@@@ H�H��x���H�E�H�@|H������H�E�H�@tH����������x�����p�����h�����`���H���  H��0������5�/  ��/  h M@ j A�    A��   �   �   ���  H��H�    ����H!�H�É�H��H�E�H�ھ M@ H���
  �5�/  �y/  A� M@ D�u/  �   �   ����  �����UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]ÐUH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H�}�u�H�E�@9E�r
�    H� �3H�E�H� H�E��E�    �E�;E�sH�E�H� H�E��E���H�E�H�@]�UH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �w
  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��H�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]ÐUH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H���  H�E��� L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A���  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�AUI��H��ATA��H	�I��UH��SH��L)�H��H��H���t:��  M��uH��[]A\A]�D  H��I�4H�| L��[]A\A]��  D  �c  �ĐSH���(   �"  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     SD�\$L�T$��y�1���y�1�A��E��E��M�J��A��D	�A	���~LA;r}F�\�D�\�D  ��~'A�B9�}���A�B��9�~���H�E��D9�u�9�t	��A9r�[�fD  D��SE������AQ��A��P�T���XZ[�H��I��H��A��H�� ��H�� ������� AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*�������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   �CA9���   D��D��D�\$�NfD  ��L�[�D��    G�L��L�KD��x��E�9E� H�{D�D9�t=�C����9�~0��D�BD�L= �zI�H�A��u��?u�A�8u�D9�u�D  D�\$E)�9t$t��9s�F���H��[]A\A]A^A_��    AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_ÐH��H��A��H��APH�� A��H�� ����m���H����     �NH��H�� ��~zAVAUATUS�O��)���~^I��I����E1��f�A�F)�D9�~DA�EB�<#A�~��    A��Hc�A������4�    Hc�I~Hc�Iu����E9e�[]A\A]A^���    �NA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      H���   HD��/  ff.�     @ �  ff.�     �
  ff.�     �����ff.�     �
  ff.�     �
  f.�     �UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo%  @ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo%  @ f��fs�f��f H����H��]Ð�����������                AW�B��A��AVAUE��ATU��SH��H��`F@ �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�J���_AXA��@�w���A��AV�   ��RD�L$A��   D�D$����Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�����XZA���%���A��AVA��   RD�L$�   ��D�D$����A[XA�������A��AVA��   RD�L$�   ��D�D$�|���AYAZA�������A��AVA��   RD�L$�   ��D�D$�G���_AXA�������A��AV�   ��RD�L$A��   D�D$����A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃������XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_� H��H��E1�E1�H�t$1ɿ   H�D$    �  H�D$H���f.�     D  H��H��E1�E1�H�T$1ɿ   �r  �D$H���f�     Hc�E1�E1�1�1ҿ   �I  f�     H��H��H��Hc�L�D$H��E1ɿ   �  �D$H���D  H��H��H��Hc�L�D$H��E1ɿ   ��  �D$H���D  H��H��Hc�Hc�L�D$H��E1ɿ   �  H�D$H���@ H����E1�Hc�L�D$1��  �D$H���ff.�     @ H���7���H��H��H���W���H��H���{���ff.�     ����ff.�     H�������1�H���H��1������   ��u��H���D  ������1�H�����H��H��E1�E1�H�T$1ɿ   ��  H�D$H����     L�D$(H�L$ H��E1�H�T$�   �  ��GP1�S�5X'  �����9H'  CA'  ��H����  f��H��PM@ @�X�"'  H�     H�@    H�@     �X�@(   H[��     H��PM@ H��'      H��'      H�     H��HM@ ��&     H�     H��@M@ ��&      H�     H��'      H��'      H�s'      �f.�     AWAVAUI��ATUSH���D  1�H�V'  A�   ��
  M�e 1��
  M��t�H�D'  H����  H�,'  I�mHH����  �S�KA�   A��A)�I9���  ��)�L9�v
H��&  I��H9�s$H�CH����   �P�HH�É�)�L9�w�H9�r�H�S H���@  H��H)�H��(H9���  H�J�rH��t%H��H)�H��(H)�H9���   H��H�J�rH��uۋCH�D�H)�H)�H9��8  H�CH���t���A��t#D�������H�CH����  H��Q���A��uH�+&  H����  E1��3���f�D������H�CH���r  H�H���(���H�T$�~D$H�H�L$H�F(H��`�F����D�f�D$D�n�F�H�JH�^�H�H�BA�D$(H��CH��HM@ L ��u<H���   �F�1���  H��H��[]A\A]A^A_ËP�HH��E1��[����    �   H)�Hƃ�H���D  �P�HH��E1�E1��(���@ H�2H�H(H�JH�P(A�T$(D�`DH�@0    �@@���H�X8D�hHSH��HM@ L"L�"H��@M@ L9"LC"H��`H��L�"��uH�ź   �P�1��)  �2����   H)�HЃ�H����D���)���H��$  H���V���1�1���  �����H�C(�C@���f��H�C C(A�D$(CH��HM@ D�cDL D�kHH�[8L� H��@M@ L9 LC H��`H��L� ��u7H�ݸ   �C�1��  ����H�C(H�H�S0H�C �C@���H�C(    닸   H)�HÃ�H���ff.�     �H����   SH�G�H��H)�H�� HC�1��  �C�H�s�=���u~�K�H�{�H��HM@ H��H)
�OH�S�)���H�K؃�(�G�C�ޭ�H��tH�
H�H����   H�QH�W H�K#  H��tnH��t�w�Q+Q)�9�}H�=+#  1�[�   ��H�#  ����� ���� t
f=��t<�u�H��"  1�[�^  fD  H��"  ��    H9=�"  H�GtKH9�tVH�H��tH�BH�GH��tH�H��PM@ �W�wH)�I  1�[�  �H�W �5����    H��"  ��    H�e"      � ��SHc�H�������H��t1�1��     � �QH��H9�w�[�ff.�     @ AUATUSH��H��H����  I��H����  H�G�H��H)�H�� HC�1��D  �E�H�U�=����2  D�e�M9��e  1��.  L���6���H��I����  H�CI�L$�H9�H�E��H9������  H���v  H��1�H��H��H��H��H��fD  �oD H��H9�u�H��H���H��H��    H��L�H�I�<�H9�t'A��H�W�H��vA�PH���PH��vA�P�PH��H��H��   H��H�4L�$�H�M��t��I��t�V�PI��t�V�PH�������H��H��[]A\A]�f.�     ��H��   ����� ���� tHf=��tB<�t>1�1���  H��H��[]A\A]��    D�j 1�H����  H��H��[]A\A]�@ H�    �fD  �[���1��l���@ H��H��[]A\A]����fD  H��H��H�4�   1��    ��T H��H9�u������ H�������H��L�B�H����   I����   �t$�I��H��I���I�fnD$�f`�fa�fp� f�H��L9�u�H��H���H�8I)�H9���   @�1M����   @�qI��t|@�qI��tr@�qI��th@�qI��t^@�qI��tT@�qI��tJ@�qI��t@@�qI��t6@�q	I��	t,@�q
I��
t"@�qI��t@�qI��t@�qI��t@�q�H���e���ÐH��H���  H�NL�B�H9�H�H@��H9���@���   I����   M��1�I��I��L��H��H���oH��H9�u�M��I���J�<�    H�>H�M9�tH�	H�I����J��   H�H�H��v�>H��H��H���y�H��t)�<@�<H��H��tD�D�D�D�H��t�V�Q�f�L��H��L��   1��    H�<H�<H��L9�u��u���f�H���ff.�     H��t#�H�9�u��    �9�tH��H9�u���    H���ff.�     �H��t*D��A8�u'1�� D��A8�uH��H9�u�1��fD  1�A8�������)���    AU1�I��ATI��H��UH��SH������H��L��Hc�H���"���H��H��L������H��1��
���H��L��[]A\A]�f.�     f�I��SH��H��H��L��L��L���i[�fD  1��ff.�     f�H���M@ �  1�� H��Hc�E1�E1�H�T$1ɿ   ����H�D$H����     1��f.�      H��  H���t3UH��S� @@ H��D  ��H��H�H���u�H��[]�f.�     �������  /shell.lef /dev/mouse0        zR x�        :���I    A�CD  $   <   =����   A�CN�����   d   <���2    A�Cm      �   ����
   A�CH�   �   2���-    A�Ch      �   @���    A�CL      �   2���V    A�CQ        h���"    A�C]          j����    A�CE��      D  ���-   A�C(    d  ���k       <   x  t����    B�A�D �G0U
 AABI[ AABH   �  ���o    B�H�K �D(�M0V
(A ABBFD
(M ABBJ     (���3    A�q         L���          4  X����    A��  $   P  ����     D�LG FAA      x  ����       H   �  ����I   B�F�E �H(�G0�A8�GP8A0A(B BBB   T   �  ����o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T   0  ����o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB     �  ���(    DK X  <   �  ����    P�B�B �A(�A0�j(A BBBA�����4   �  h����    H�F�E �A(�� ABB            ���          0  ���          D  ���          X  ���          l   ���          �  ����       �   �  ����R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   <  ����m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        �  ����1    D l    �  ����'    D b    �  ����          �  ���+    D f    �  ���+    D f      4���,    D g       L���!    D \    8  d���    DI    P  \���    DI    h  T���          |  P���          �  L���    DK     �  D���0    DV
FM          �  P���(    D c    �  h���              �  p���h    F�a       ����v       H   ,  0����   B�B�B �E(�A0�A8�DP�
8D0A(B BBBA,   x  ����m   J��
�Hm�[�B
�F    �  ����1    D�l   t   �  ����P   B�B�A �A(�G0_
(D ABBKo
(D ABBHR
(D ABBEd
(D ABBK         <  �����          P  ����         d  ����4          x  ����I       4   �  0���T    B�G�G �D(�D0r(D ABB    �  X���    D�U          �  X���          �  T���          	  P���(    D c    $	  h���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��������        ��������                                               1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             @     �      �@     I       4@     2       f@     -       �@            �@     V       �@     "       @     �       �@     -                      ,            @     �                                              �    #                  Q  
5   �  �  int �   P  ]   �  i  p   _  6  �   .  6   �   )  
   �   �  
�   T  w    �  w   bpp d     w   
 �   �   �     �  H  (|  x C    y 	C   T  C   �  C     C   r  
Q   �  	|  r  

Q     	Q   �  
  �   �  x 	C    y C    �  	�  
�    �  r Q    g Q   b Q   a Q    �  �  �  n     	�  |#  �  x d    y d   T  d   �  d   x  w     �  �  �   l�    t%  ~  �  ;    	  �  �   _ %  $  �  	�  �  
  	�  	�  �  	�  6  	�  (
w   O  �  
�    �  
�   msg 
�   Z  
�   p  
�     y   
   C   k  �    �  [  	@@@     K  �<�  �  =   k  >�  pos ?�  �  @�  � �  fb C
|  	�L@       D�   	�L@     k  E�  	 M@     )     �    �  G  	(M@     �  H�  	@B@         I�  	+M@     �  J�  	,M@     X   K�  	0M@     �   M�  	HB@     >  O	  	8M@     ~  j�  	IB@     Y  �  �  ?   �  �  �   �  �      �  C    0  !�  (  .  �   �  *   C  N  �  �   %  ;v  c  n  �  �   �  LV  �  �  �  �  �      V�  �  �  �  �  �    �  `�  �  �  �  �   �   `  j�  C   �  �  �     n�  �      �  �      �  �  7  =  �   �  �x  �  V  \  �   )  ��   �  ��  num ��   T �   	�  
�  	�    �  �   	�   9  
�  obj �  �   <  �  �  �   T �   	�  
�  �     �@     -      ��  �  �  �Hpos n�   �D o  t�  �h!obj x�  �X"@     	       ~     p�  �P #@     8       !i v�   �d  .  �  @     �       ��  �  �  �Hobj *�  �@ �  +�  �X $�  �    %�  �   &�  w  &  �@     "       �/  '�  �h (n  N  �@     V       ��  �  �  �Xpos L�   �T o  O�  �h#�@             !i Q�   �d  (�  �  �@            ��  �  �  �h )�  �  �  %�  �   &�  �  �  f@     -       �	  '�  �h *�  �C   �@     
      �;   F  �  �� �  �C   �\ c  ��  ��~   ��  �P c   ��  ��} �   �C   ��#�@     
       �  �C   ��}+msg 2O  ��|"	@     �      c
  !j �C   �L#)	@     �       �  �
�  �K �   ��  ��| �   �  ��"r	@     N       ?
  !i �C   �D #�	@           !win ��  ��   "$@     9       �
  !i �C   �@#3@     $       !win ��  ��~  "o@     1      0  !i �C   ��#�@     	      !win ��  ��~#�@     �        �   �O  ��| ?  �w   �� Y  �w   ��   "�@     �       y  ,�   O  ��|,?  w   ��,Y  w   �� "�@     �         +i C   ��#�@     �       ,�  	�  ��#�@     �       +j C   ��#�@     s       ,�    �  ��|,�   !  ��~    #�@     �       ,�  7O  ��|   	�  
;  $�  W  a  %�  A   &F  �  �  4@     2       ��  'W  �h -X  l;  @     �      ��  win l�  �� /  ~�  �� .�  F  �  �@     I       �  l 0  �hr E  �` /�   N    �   @      @     7	  src/gfx/sse2.asm NASM 2.14.02 � @              %U   :;9I  $ >  $ >  :;9   :;9I8   :;9I8  ;   	 I  
& I     :;9n  .?n4<d   I4  I  ! I/   <  4 :;9I?<  4 :;9I?  4 :;9I?  :;9  .?:;9n2<d   I  .?:;9nI2<d   :;9I82   :;9I82  / I  .?n42<d  .Gd@�B   I4   :;9I   4 :;9I  !4 :;9I  "  #  $.G:;9d   % I4  &.1nd@�B  ' 1  (.Gd@�B  ).Gd   *.?:;9I@�B  +4 :;9I  ,4 :;9I  -.?:;9n@�B  ..?:;9nI@�B  / I   %  . @   3	   |  �      /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx/window /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/lemon  graphics.h   main.cpp    window.h   list.h   stdint.h   fb.h   surface.h   types.h   stdio.h   ipc.h    G 	�@     
�ff!.  tt!.�  	@     � Zt<ZK
�H<
t&�$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�.K�k�<60B�4�B �8R:�<(.*�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9%�������	�*(!
	<*f�� t
�K�+�* t ��<<tKK +mt'����)��=Z jt��, t � u �kv>f��f��t! J t< Jv�u,ff.�,ff.��( J��( J�tf � ��"u%�* f�uf�, �9 fG �; �  .Y �f fM �t �� f� �� �h .�)�u�<f5 J; t& <K+f �7.Df9�J�trX�t<K'f�J='f�JZ'f�)J<='f�)J<(>/�X6u�u6 g.�� J	�w  �" t f�	uu �* f �8 �H fY �J �, .k �{ f_ �� �� f� �� �} .�!u�<f: J@ t( <��t<K)f�J=)f�JZ)f�+J<=)f�+J<' >. � X8 u � u6( t �	�K t��+�<<�Kxf�tK= ot���t� � t�tJ" X' t <Y$�)t/<��$�(t�.v�u6o X4)*  	4@     �*  	f@     ����  	�@     � 
�u  	�@     � �t* X�� t* � �h�  	�@     �  	@     )�#���tY�����  	�@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K �    '   �       src/gfx/sse2.asm      	 @     !>==?LLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""��      mouseDown uintptr_t _ZN4ListIP8Window_sE8add_backES1_ uint64_t _ZN4ListIP8Window_sEC4Ev dragOffset testWindow handle_t 13ipc_message_t next long long int mouseEventMessage windowHandle windowInfo fb_info_t redrawWindowDecorations ListNode mouseDevice Vector2i active remove_at _ZN4ListIP8Window_sE9get_frontEv stdin _ZN8ListNodeIP8Window_sEC4Ev List<Window_s*> uint16_t linePadding _ZN10win_info_tC4Ev this _windowCount keymap_us GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions _ZN4ListIP8Window_sE9remove_atEj temp get_front RGBAColour long unsigned int _Z10DrawWindowP8Window_s width data short unsigned int depth _ZN4ListIP8Window_sE8get_backEv _ZN4ListIP8Window_sEC2Ev recieverPID bool stdout decltype(nullptr) FBInfo operator[] windowFound vector2i_t fbInfo long double title pitch /home/computerfido/Desktop/Lemon/Applications/Init _ZN4ListIP8Window_sEixEj current _ZN8ListNodeIP8Window_sEC2Ev _ZN10win_info_tC2Ev operator+ _ZN4ListIP8Window_sE6get_atEj surface_t unsigned char node short int _ZN4ListIP8Window_sE10get_lengthEv main.cpp 10win_info_t clear uint32_t mouseX _ZplRK8Vector2iS1_ mouseY get_length info data2 _ZN4ListIP8Window_sE9add_frontES1_ buffer _ZN4ListIP8Window_sE10replace_atEjS1_ _ZN4ListIP8Window_sE5clearEv add_back drag IOFILE replace_at get_at stderr ListNode<Window_s*> add_front renderPos prev lastKey fbSurface uint8_t DrawWindow windows renderBuffer flags backgroundColor handle senderPID _ZN4ListIP8Window_sED4Ev mousePos ~List height rgba_colour_t main mouseData get_back ownerPID keyMsg                 @     �@     �@     3@     4@     f@     f@     �@     �@     �@     �@     �@     �@     @     @     �@     �@     @                                                   � @                   � @                   q1@                   y1@                   �1@                    @@                   @@                    @@                  	 �L@                  
                                                                                                                                                                                                                           ��                      @@                  @@             (     �1@             ;     � @             =     @             P     P@             f    	 �L@            u    	 �L@            �     �@             �    	 �L@     0           ��                �     @@             �     �:@             �     01@             �    ��                �    ��                     � @                ��                #   ��                /   ��                @     -@             Q     Q@             l     �@                  �@             �     �@             �     �@             �      @            �   ��                �   ��                �   ��                �   ��                �   ��                h   ��                �     %@     h       �    dL@                `L@               	 xM@               	 pM@            %   	 hM@            4   	 `M@            A   	 XM@            T   ��                ]   ��                g   ��                s   	 PM@                � @             �    �@     o      �    @B@            �     @     (          	  M@     (          	 @M@                P0@     T       %    �0@            -    p%@     v       ;    �0@            K    �$@     (       �   	 �M@            Z  "  �@            `    p#@     +       k    @@     o      �  "  �@     "       �    �.@           �  "  �@     I       �   	 HM@            �   hL@             �    �$@            �   @@             �   	 0M@                 #@     '           �%@     �          @@             %  "  �@     "       B  "  @     �       d    �"@     1       q    P$@            w  "  �@            ~   	 ,M@            �    IB@            �  "  �@     V       n   	 �L@            5    � @             �    �0@            �    @@@            �   	 8M@            �  "  4@     2       �    @     k       �    +@     1           D@                	 (M@            P    @$@            "    P@     o       <    h@             J    �#@     +       V    �/@     4       ]     @     R      x  "  4@     2       x    � @            f    0$@            �    �0@     (       �  "  �@            �    �@     �       �    P+@     P      �    �@             �     0@     I       �   	 +M@            �    �@     I           @     �       ;    p"@     m       Z  "  f@     -       s   	 hL@                 �@            �    �-@     �       �    �@     
      �    `F@            �     @            �  "   @            �    �@             �    q1@             �  "  �@                 1@              "  �@                �@     3       @    �$@     0       G    hL@             N   	 �M@             S  "  f@     -       l    HB@            �    �#@     ,       �    @     �      �    P@     �           `$@            �    P#@            �  "  �@     -      �    `B@               	 �L@            	  "  @                 $@     !            @             �    p$@            +    �@     �           �)@     m       crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4699 dtor_idx.4701 frame_dummy object.4711 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux graphics.cpp /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp fb.c filesystem.c ipc.c allocate_new_page l_pageSize l_pageCount l_memRoot l_bestBet l_warningCount l_errorCount l_possibleOverruns memory.c syscall.c _liballoc.c l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer l_max_inuse memmove syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm lemon_read _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN8ListNodeIP8Window_sEC2Ev memcpy _ZplRK8Vector2iS1_ l_inuse __TMC_END__ SendMessage __DTOR_END__ dragOffset lemon_open malloc __dso_handle _ZN8ListNodeIP8Window_sEC1Ev _ZN4ListIP8Window_sE8add_backES1_ lemon_map_fb lseek _ZdlPv drag backgroundColor _ZN4ListIP8Window_sEixEj liballoc_lock keymap_us lastKey _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm calloc memcpy_sse2_unaligned mouseData _Z16memcpy_optimizedPvS_m memset32_sse2 lemon_write memchr _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev liballoc_alloc _ZdlPvm _Z18memset64_optimizedPvmm realloc _Z8DrawRectiiii10RGBAColourP7Surface memcmp mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main font_default _Z5floord _ZdaPv memset64_sse2 _fini _ZN4ListIP8Window_sE10get_lengthEv liballoc_free _Znam _Z24CreateFramebufferSurface6FBInfoPv access _edata _end _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close _ZN4ListIP8Window_sE9remove_atEj font_old fbInfo _ZdaPvm lemon_readdir memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                     � @     �                                     !             � @     �       �0                             '             q1@     q1                                    -             y1@     y1                                    5             �1@     �1      8	                             ?              @@      @                                    F             @@     @                                    M              @@      @      H                              S             �L@     hL                                    X      0               hL      +                             a                      �L      �                              p                      sM                                    �                      �M      j                             �                      �Z      �                             �                      �]      �	                             �                      �g                                    �      0               �g                                  �                      �m                                    �                      �m      �                                                    `n      0         A                 	                      �}      Z                                                   �      �                              