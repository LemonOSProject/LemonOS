ELF              ��4   ,g      4    (           � ��C  �C           �C  �����  �        �W  �R3  �                 �    UU���B$  VW�����_^�y  �    �i���f�f�f�f�f��(�=(�t$�    ��tU���h(��Ѓ��Í�&    f�Í�&    ��&    ��(�-(����������t(�    ��tU���Ph(��҃��Í�&    �t& �Í�&    ��&    ��=(� ugU�,���V���S����������9�s�v ���,����,�9�r��'����    ��t��hH��Q~�����(��e�[^]�Í�&    ��&    ��    ��t'U���h0�hH��~������	�����&    f���������t$�#  ��Ã��t$�o#  ��Ã��t$�?'  ��Ã��t$�/'  ��Ã��t$�'  ��Ã��t$�'  ���UWVS���t$(�|$,�T$4�\$0�T$�F�D$�G�D$�~ ��   �G)Ѕ���   �T$�$    �[���F9�~4�O��)�9�~)�$Ћl$�l� ������v��L$���D$�,��$�$9F~*�D$�G+D$;$~�F��~܋O��)څ�~Ѻ    롃�[^_]�UWVS��8�l$L�|$P�D$T�D$�L$X�L$ �t$\�L$`�L$�\$d�\$$�T$h�T$(j� "  ���     �@    �@    ��9�
�D$�9�}R�L$9��D$�9���   t$9�|�D$�9���   �t$�T$�9�|�D$�9��  �؃�,[^_]Ã�j�!  �     �@    �h�x��)���P�L$$�H��C�C   �����j�����j�Y!  �     �@    �h�x�L$ �H�T$)����P���; t�S��S�P�C�C�|$�-�������)�D$��j��   �     �@    �p�x�T$ +T$(�P�L$$�H���; t�S��S�P�C�C�D$�D$���������j�   �     �@    �h�p�L$ �H)��T$$)�P���; t�S��S�P�C�C�������S��(�\$0�St�T$�Kx�L$�D$    �D$    �C|�D$���   �D$�Cu	�=�� u#��j �D$P�D$(P�sph��j��,  ��H[�h��j j j ��PjQR��  �� h��j j j ���   ��Pj�sx�C|Ct��P�  �� h��j j j j�C|��P�sx�st�y  �� h��j j j j�C|��P���   Cx��P�st�M  �� 9���6  h��h�   h�   h�   j�s|�Cx��P�Ct��P�  �� ��h��h�   h�   h�   �Cx��P�Ct��P�CP�  �Ct�Sx�H�L$8�J�L$<�� h��j2j2jdjj��RC|��P�  �� h��j2j2jdjj�Cx��P�C|Ct��P�  �� h��j2j2jdjj�Cx��P�C|Ct��P�[  �� h��j2j2jdjj�Cx��P�C|Ct��P�3  �K|Kt�A�Kx�Q�� RPh��h����  ��������h��h```�h   �j�s|�Cx��P�Ct��P��  �� �����S��j j j hh�hl�j�*  �l��h���+x�i��  ��+t�Ѓ� =�  v,����̉��%|����p��|�    �x��t���[�ÍL$����q�U��WVSQ���   j j j h���E�Pj�*  ����������P�&  ��������n  ���   ���   ��� ���j��  �     �@    �@    �H���j j j j h�j�)  ��j j j �E�Ph&�j�)  ���   ���   ��j h2��b(  ���$   �t  �����jj S�(  �ǉ$�X  �ƃ�WPS�'  ��h��Vjjj j ��  ��S�<(  ��j h=���'  �Ã�jj P�'  �ǉ$�  �ƃ�WPS�G'  �T�   �X�   �$  0 ��  �`�����u%ǅ@���    ǅ8���    ǅD���    �  ����hL�Vh   h   j j �*  �� �ǅ<���    fǅl���  fǅn���  fǅp���  fǅr���  ��j j j ��l���P��<���j�(  ��@����ǃ� ����   �uܻ    � �    �	��D����B;ppt/��9���   ��9�@���vօ�tً�D����    ���9�u���9�@���vQ���+	  ��D����    ���9�u��Bƀ�   ��D����    ���9�u��B��l����   ����   �    ƀ�   �    �ك�h�   �`  �Í�l����   �����l����Ct��n����Cx��p����C|��r������   ƃ�   ����$   �  �     �@    �X����D��� t=��8�����H��@��������8�����<�����<���9�T�����  �7�����D����������@���������  ��������<����  �5    �   ��D����  ��D����H��4������t�H��t�J�P��t���t�
��u���D�����@�����@���9�t��P��  ����8�����H��8����ድ8�����j��  ��8����     �@    ��4����H����D��� ��   ��p��@�����@���9���   ����   ��D����    � ��9�u��@�������Wx����J9���   �G��  �5���Ot��<���O|�Y�9�}�Z9���9�|�J9�E+�<����5��)У�������  ��8�����D����E����    �o�����D����a���ǅt���   �Gp��|�����P��x���j��p�����l����wl�h$  �� �m  ǅt���   �G�  ���+Ot����)��
  �������  ��9���������������D����    �6��9�u��v�Ft9�~�F|9�}��Fx9�<���~���   9�<���}�����@���������9��������������D���� ���(  �    ��9�@��������9��~�������  ���ۡ    ���    t���5    �\����    ���i  �    ;���_  ���    �    �K  ��D������t�Q��t�P�A��t���t���u���D�����9�t��Q�!  ���    ��  �A��8����߉�@�����X�����S�"  ������   ��`���� uࡨ���t׋�d�������t �у�tǅt���   �� ���x����ǅt���   �� ���x����Pp��|�����R��x�����t�����p�����l����pl�3"  �� �^����5���5��h��h���5���h��j j j jjj j �8  ��,j
��l���S�5p��"  ��h��h�   h�   h�   j j S��  ��j j j h���u�j��!  �� �|�������j ��P���Pjh���u�j�!  �� ��P��� t>����Q����P���    H£���A�؋���B���    H£���=�� t3���������+���    HӉQt+���    HAx�����j j j j ��T���Pj�!  �� ��T��� ������������t���S�������   �=�� t��� h��h�   h�   j@�����P�5��j j �  �� �    ��@�����@��� �u  �y�����D����@���ǅt���   ���+Ot)�����ȉ�x����Wp��|�����RP��t�����p�����l����wl��  �� �=�� �Q������� �C������ ��� ǅt���   �������������|�����x�����t�����p�����l����pl�  �� �������D����H��4����������    ��   ����D����s�F��������V��D����@��D������    ��   ��tȋ�D����    ���9�u����r� �������D����    ���9�u��Bƀ�    ��9�������9��R�����t���D����    ���9�u��B���    u���D����    ���9�u����9B�������R�����D�������(����    ��9��8���9��0�������Q������ߋ�D����Bƀ�   �����f�f�f�f��UWVS��  �Û?  ���|$$�D$ �l$(	��t��UW�t$,�  �������)�����RW�t$,�q  ����u
��[^_]�f����VW�t$,�V�M  ����[^_]�f��T$�D$�Í�    �T$�Í�&    �v S�3  ���>  ��h�  ��������� [��Í�&    �t& �VS�  ���>  ���t$��&    �t& �������t�������Vh�  �t�����[^Í�&    ��&    VS�
  ��}>  ���t$�> t-��&    �[�����t����F���Ph�  �"������> uڃ�[^Ít& UWVS�`
  ��+>  ���t$ �|$$�T$(��   t*�B���t�v ���>�����u��[^_]Í�&    �t& ������R��WV�  ����tӉ>��t̉~��tĉ~��[^_]Í�&    �t& ���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�Ð�	  _=  UWVS��,�T$H�|$@�D$�t$T�D$P�l$D�L$L�T$��y�1��T$��y�1���Ё�   ���	ډ�% �  ����	�	ËF�\$�D$��~v;n}q�D$�t$T����D$�D)��l$T�D$���&    ���9u~C�]��)�;\$OD$��P�t$�E�L$ ����������P�\$�N�����;t$u���,[^_]Í�&    ��    VS�  ��]<  ���t$j j j j Vj ��  ��$��[^� f��`  /<  UWVS��,�|$@�t$D�D$�L$L�D$P�\$T�T$X�l$\��y|$H1���y�1�����������	�	E�T$�D$��~\;u}W�D$H��D$�D��D$�
f���9u~9�]������)�;\$OT$H��R��t$�L$ ��P�\$�H�����;t$u���,[^_]Í�&    �  _;  UWVS��,�t$@�l$D�D$�L$L�D$P�|$T��yt$H1���y�1��؉������� �  ��	�	G�T$�D$��~i;o}d�D$H��D$�D��D$��t& ���9o~C�G�_������)����;\$OT$H��R�t$�L$ ���P�\$�n�����;l$u���,[^_]Í�&    ��    UWVS�  ��{:  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$�������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�@  ��9  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�,����� 9t$h�_�����L[^_]Í�&    UWVS�p  ��;7  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�\����� 9t$l�_�����L[^_]Í�&    UWVS�  ��k5  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�9�����9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$Ë$�f��UWVS������û3  ���D$<�|$8�t$0�D$�G�D$�D$D���� ��D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������ ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ�P����� ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�N����� 9|$�b�����[^_]Í�&    f�UWVS������[1  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��U��E�]�Mfof ��������]�U��E�]�M��~4fn�fo@�f��fs�f��fs�f��fs�f��f ������]Ð������                U��01�WVS������V0  ��(��p  �����9�l  C�l  P���  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p����1���p  �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � �����\  ��`   �g�����&    �t& � ����.  ǀh      ����ǀd      �    �B    ����ǀp     �    �B    ����ǀl      �    �B    ǀ\      ǀ`      ǀT      ǀX      ǀL      ǀP      Í�&    �UWVS�P�����.  ���|$0� ��&    ���\  �   ��`   �  �w �  ��t܋�h  �t$�|$0����  �|$0��d  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s��d  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ���h  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$���������B1ҋD$~Q��@�����   ��   �E��  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,�����E$���~����Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ�������������h  ���K�����
  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~�����N,�����ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��D
  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS�p�����;*  ���D$ ����   �P���)փ� C��	  �N�A=����~   �y����1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o��d  ����   ��t�J+J�ʋO)�9�|W�R	  ��[^_]Í�&    �v ��T  ��X   ����� ���� t
f=��t<�u���L  ��P   뱍�&    ���d  롍�&    ���\  ��`   ��[^_]Í�&    �v �G9�h  tU9�ta���t�B�G��t������G1�)Q���wW��  ���4�����&    �t& �o�������&    ���h  룍�&    �ǃd      듍t& WVS�t$�����È(  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS������Û'  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��  �G�P�������   �P9���   �T$��  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ�T  ��X   %��� =�� tDf����t=���t8�C  1���[��^_]Í�&    �p���&  ����[^_]Í�&    �t& ���L  ��P   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ�����f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f�S�c�����.$  �� j j j �D$ P�t$8j��  �D$,��8[�f�S�3������#  ��j j j j �t$(j�  ��([Í�&    f�S�������#  �� j �D$P�t$8�t$8�t$8j�g  �D$,��8[Í�&    ��&    S������Î#  �� j �D$P�t$8�t$8�t$8j�'  �D$,��8[Í�&    ��&    S������N#  �� j �D$P�t$8�t$8�t$8j��  �D$,��8[Í�&    ��&    S�C�����#  �� j �D$P�t$4�t$<�t$8j�  �D$,��8[Í�&    ��&    S�������"  ���t$�t$�t$�������[Í�&    �t& S������Þ"  ���t$�t$�t$�������[Í�&    �t& S������n"  ���t$�t$�t$� �����[Í�&    �t& S�s�����>"  ���t$�t$�������[Í�&    ��&    �S�C�����"  ���t$�������1�[ÐS�#������!  ��j �t$�������   ��u
����[Ív ��P������1҃���[�f�f�f�f�f��S������Þ!  �� j j j �D$ P�t$8j�;   �D$,��8[�f�S������n!  ��j �t$0�t$0�t$0�t$(j�   ��([�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��WVS�D$�L$���ƍT�N��������~&1���&    �t& �:����Z�����9�|�[^_Ív W1�VS�D$������ö   �|$�t$��t@�������	~%��W�T���u��� QW�l�������[^_Ív ��0�T���u��ٍv �0   f���[^_�f�1�Í�&    ��    �p���?   �� ��  1�Í�&    �v S�S�����   �� j j j �D$ P�t$8j�����D$,��8[�f�1��f�f�f�f�f�f��������t6U��S�������&    �v �Ѓ�����u��[]Í�&    ��&    ��:����  /taskbar.lef /dev/mouse0 /close.bmp /bg1.bmp          zR |�        ����    CD H     8   ����    CD H     T   ����    CD H     p   y���    CD H     �   m���    CD H     �   a���    CD H  8   �   U����    A�A�A�A�C(�A�A�A�A�h      ����
   A�A�A�A�CLvP^@[
A�A�A�A�ACLBPx@JLBPn@oLBPm@kLBPm@   p  l  ����r   A�C0E8B<E@EDCHELBPHA�A0�E4B8B<B@DDBHALAPH0E4B8B<B@JDBHCLJPH0E4B8B<B@BDGHCLCPH0E4B8B<B@BDGHMLCPH0Q4E8E<E@BDCHGLGPH0C4E8E<E@EDGHGLDP\0E4B8B<B@BDBHDLGPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPH0E4B8B<B@BDBHGLJPW0A4A8E<E@H0H4E8E<E@BDCHGLGPH0 4   �  ~���z    A�CBB B$E(E,B0lvA�        ����       ,   ,  �����   D Gu Fupu|uxut|   \  h���~    A�A�A�A�N U$A(A,D0H E$K(A,D0H G
A�A�A�A�CC$C(A,G0H CA�A�A�A�     �  h���
          �  d���             `���$    A�NE HD� 0   (  l���B    A�A�N^DE HA�A�  4   \  ����L    A�A�NcAE HHA�A�   \   �  �����    A�A�A�A�N n
A�A�A�A�LC$F(D,A0H YA�A�A�A�   �  ����?    Cy H     �����    K�A�A�A�C@�DAHDLYPL@IA�A�A�A� 8   X  ����.    A�A�NFB B$B(A,B0HC�A� H   �  �����    K�A�A�A�C@�DAHFLHPL@IA�A�A�A� H   �  $����    K�A�A�A�C@�DAHDLJPL@IA�A�A�A� <   ,  ����b   A�A�A�A�NPL@�A�A�A�A�X   l  �����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   �  \����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   $  �����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   p  4����    A�A�A�A�C(�A�A�A�A�   �  ����          �  ����         �  ����W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   �  ���s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�  D   @	  �����   A�F�A�A�N<Z@J0�
A�A�A�A�M      �	  ����       T   �	  �����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `   �	  0����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   X
  |����    A�A�A�WA H��A�A�  �   �
  4����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0<      T���   A�A�A�A�C �
C�A�A�A�A 8   `  $����    A�A�A�A��
�A�A�A�P   0   �  ����.    A�N(B,B0B4E8D<B@LA�  0   �  ����'    A�NBB B$B(D,B0HA�  0     ����2    A�N(B,E0D4D8D<B@LA�  0   8  ����2    A�N(B,E0D4D8D<B@LA�  0   l  ����2    A�N(B,E0D4D8D<B@LA�  0   �  ����2    A�N(B,E0D4D8D<B@LA�  (   �  ����%    A�NDDD HA�   (      ����%    A�NDDD HA�   (   ,  ����%    A�NDDD HA�   $   X  ����!    A�NDD HA�      �  ����    A�ND HC� 8   �  ����E    A�NBD HL
C�DCA HEC�0   �  ����.    A�N(B,B0B4E8D<B@LA�  0     ����-    A�NBD D$D(D,B0HA�  (   H  ����!    A�A�A�[�A�A�,   t  ����M    A�A�A�G�A�A�   D   �   ���n    A�C�A�tEA HC
�A�A�D[�A�A�    �  (���             $���       0     0���.    A�N(B,B0B4E8D<B@LA�     H  ,���           ����    ����                                                  @  �                          �             �   �            �����   �           ���������   �          �������������   �         �����������������   �        ���������������������   �       �������������������������   �      �����������������������������   �     ���������������������������������   �    �������������������������������������   �   ���������������������   �   �   �   �   �   ���������   ���������   �����      �����   �    ���������   �      �   �     ���������   �����      ����   ���������   �          ���������   �       ����   �   �����                 1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                                                                                                                                                                                                                                                                                            <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              Т�                           >        ТP�    src/gfx/sse2.asm NASM 2.14.02 �Т     %  . @   _    '   �       src/gfx/sse2.asm      Т!0==?LL==0/!#!0==>=0K�KYKYKYMK>1/""u�                                            t�          ��          �          �          H�          ��          ��          ��          ��     	     (�     
                                                                                                                             ��   ��         ��      (   H�      ;   ��      =    �      P   P�      f   (�    
 u   ,�    
 �   Ё      �   0�    
             ���   ��      �   ��      �   г      �            ��  ��                  ��           ��#           ��,           ��5           ��F  ܢ       W  ,�       h  5�       x  @�                ���  P��    �  $�    	 �   �    	 �  �    
 �  �    
 �  �    
 �  �    
 �   �    
 �           ���           ��           ��           ��           ��           ��             ��%  ��      ;  ��    
 G  P�.     Y  p��    �  ��     �  ��    	 �  ��    
 �  p�!     �  ��M     �  |�    
 �  ��     �  p�     �  t�    
    �.     S   �    
   �       �2        H�    
 ,  ���    X  ��B     j  Ю�     q  ��    
 y  (�    	 �  @�-     �  ��     �  ��    
 �  ��.     �  e��     �  ���    �  �     �  ��    
   ��    	   �n       h�    
 0  @�%     6  ��    
 >  %�     E  ��    
 �  t�      J  `�     X   �    	 b  ��    
 i  ���     �   ��     �  p�    
 �  ��    
 �  �%     �  �~     �  ��    
 �   �2     �  �W    �  $�     (  l�    
 7  ��&       �%     =   �   	 P  ��.     _  5�     g  ��    o  ��
     }  P��     �  �     �  ��    
 �  0�b    �  ���       P�s        x�    
 2  (�     
 >  P��     d  ��    k  %��    p  ��    	 x   �    	 �  �?     �  L�    
 �  E�     �  ��$     �  �      �  ��z     �  ��     �  �     �  0�L     �  ��E        (�     	   $�     
   ��    	 $  .�
    >  `�2     I  8�r    b  @��     �  p�!     �  ��'     �   �    	 �  �      �  U�     �  ��2     �  Т      �  ��     �  ��     �  p��     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp graphics.cpp text.cpp font.cpp src/gfx/sse2.asm memcpy_sse2.loop memset_sse2.loop memset_sse2.ret bigzero allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns memory.c filesystem.c ipc.c syscall.c itoa.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _Z7inportbt mousePos l_max_inuse syscall reverse frameCounter liballoc_init liballoc_unlock lastUptimeMilliseconds ReceiveMessage _Znwm lemon_read bgClipRects _Z12DrawGradientiiii10RGBAColourS_P7Surface _Z12write_serialc memcpy l_inuse __TMC_END__ SendMessage __DTOR_END__ dragOffset lemon_open _Z12surfacecpy_tP7SurfaceS0_8Vector2i malloc __x86.get_pc_thunk.ax mouseSurface __dso_handle itoa currentUptimeMilliseconds lseek surface _ZdlPv drag liballoc_lock keymap_us active _Z18memset32_optimizedPvjm calloc frameRate mouseData _Z16memcpy_optimizedPvS_m closeButtonSurface lemon_write _Z8DrawCharciihhhP7Surface _Z30RecalculateBackgroundClipRectsP4ListIP8Window_sE currentUptimeSeconds mouseSurfaceBuffer liballoc_alloc _ZdlPvm realloc _Z8outportbth _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main testKey font_default _Z5floord bgSurface _ZdaPv _Z17is_transmit_emptyv _fini _Z15UpdateFrameRatev liballoc_free _Znam _Z12write_serialPc access _edata _end redrawWindowDecorations _Z14SplitRectangle4RectS_ lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close font_old memset_sse2 _ZdaPvm lemon_readdir memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                   t�t                     !         ���   �3                 '         �4                    -      2   �4  -                 5         H�H4  \                 ?         ���C                    F         ���C                    M         ���C                   V         ���C  h                  \         (�(S  �                  a      0       (S  +                 j              SS                     y              sS                    �              �S  B                  �              �S                    �              �S  c                  �              HT                    �              LT                                  \T  
     >         	              l^  �                               df  �                  