ELF          >     @     @       ؘ
         @ 8  @                   @       @     ��     ��                           C       C     �      `                            C       C                           �3  �>� �             H��    UUH��������	  ����    ��C H=�C t�    H��t	��C ��f��ff.�     @ ��C H���C H��H��H��?H�H��t�    H��t��C ���ff.�     @ �=)  uwUH�' H��ATA�( C S�0 C H��( C H��H��H9�s%f.�     H��H�� A��H�� H9�r��0����    H��t
�șB �����[A\�� ]��ff.�     @ �    H��tU��C �șB H�������]����D  ����UH��H����C ��C A�    A�    �    H�ƿ   �t%  H� H�� H)�H��Hi��  H�� H)�H�� H�H�E�H�}��  v[H�� H�E�H��H���S㥛� H��H��H��H�Ⱥ    H���� H��     H�� H�� H�� H�{ ���UH��H��   H�E�A�    A�    �    �    H�ƿ   �$  �E�� �E�    ��C �  9E�������   �E� �E�    �e 9E�}kH��`���H���  �E�Hc�H��`���A�    A�    �    H�ƿ   �/$  H�E�H�E�E��ƿ�C �=  H� H9E�����t�E���E���E�����t�E��ƿ�C �+  �t� �E��=������UH��H��   H�E�A�    A�    �    �    H�ƿ   �#  �E܉�
 �E�    ��
 9E���  �E� H��`���H���   �E�Hc�H��`���A�    A�    �    H�ƿ   �B#  H�E�H�E��E�    ��C �<  9E�����t)�E�ƿ�C �5  H� H9E�����t�E���E����E�������   ��   �5  H�E�H�E�H��`���H��h���H�PH�HH��p���H��x���H�PH�H H�U�H�M�H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�U؉��   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�E�H�ƿ�C �  ��� �E��c������UH��AVAUATSH��   H�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸@C A�    A�    H�ƿ   �!  �Y  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H���  H��P���H�E��@����H��X���H�    ����H!�H	�H��X���H��X�����H�       H	�H��X���H��P���H��X���H��H��H�й@C ��H��H����  �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H����  H��`���H��h���H�    ����H!�H��H��h���H�E��@������H�� H��h�����H	�H��h���H��`���H��h���H��H��H�й@C ��H��H���  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H���6  H��p���H�E��@������H��x���H�    ����H!�H	�H��x���H��x�����H�       H	�H��x���H��p���H��x���H��H��H�й@C ��H��H���Q  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H���m  H�E�H�U�H�    ����H!�H��H�E�H�E��@������H�� H�U���H	�H�E�H�E�H�U�H��H��H�й@C ��H��H���  A�    A�*�2   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H���  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A�@C D���H��H���(  H�E����   ����H�E����   ����H�E�H��H��h@C A��   A��   ��   H���0  H���E�   �E�   H�E�H���   H�E�H��H����
  H�E�H�E�H�U�H��@C A�    A�    H���   �8  H�e�[A\A]A^]�UH��H���   �(C �T  H�> H�7 H��H��H�1 H��0 �H�* f�HH���  H��H�E�H�E�H�H�HH� H� H�PH�HH�
 H� H�@ H� �� �� ��H�H���G/  H�� H�E��PH�E��@�u�h�   A�    A��   �щ¾    �    �  H��A�    A�    �    �    �    �   �  �    ���A �  �E܋Eܺ   �    ����  H�E��Eܺ   �    ����  H�E�H�H���.  H�E�H�U�H�MЋE�H�Ή��1  H�EЋ@��H��H��H�H��H��H�E�H�H�E��]    �W    ��  �9.  H�R �@ �6 H�M�A��C I�ȉщ¾    �    �^  H�Eȋ@H�H�U�H��A�    A�    �    H�¿    �  ���A A�    A�    �    �    H�ƿ   ��  �    ���A ��  �EċEĺ   �hC ���?  H�K H��H�@ �����<� ��t,��  ��  A�@C D� � �щ¾    �    �T  �E�    �_ 9E�}%�E��ƿ�C �y  H�E�H�E�H���U����E������  �Eĺ   �hC ���  ��� ��  ��Љ�� ��� �w  ��)Љ�� �e  ����   �r� �d� �N  H��  )щʉ��   �K� �5  H��  )щʉ��   H��  ���   ��yH��  ǀ�       H��  ���   ��yH�~  ǀ�       ��� �������#  ��� �����  ��� ��C �8  ���E��}� ��  �E��ƿ�C �+  H�E���� H�E����   9���  �s� H�E����   H�E��@���9���  �R� H�E����   9��  �:� H�E����   H�E��@���9��Z  �E��ƿ�C ��  H�ƿ�C �  H�E�H�x� ��� H�E����   �P��� 9�|LH�E��@����u>��� H�E����   )�� H�E����   )��ȉ�� ��� �w� ��   H�E�   H�E��@����t0�j� H�E����   )ЉE�W� H�E����   )ЉE��4�:� H�E����   )Ѓ��E�$� H�E����   )Ѓ��E��E�H�� H�E�H	�H�E�H�E�H�@|H�E�H�E�H�@tH���u��u��u���x�����p���H����  H��0�	�m�������� ����t��� ��t���  �x� ����  �f� ��������  �T�  �N�  H��� H����  �L� H��� ���   9���  �1� H��� ���   H��� �@���9��X  �
� H��� ���   9��=  ��� H�l� ���   H�_� �@���9��  ��� H�@� ���   �P��� 9�|H�&� �@������   H�E�   H�	� �@����t6�q� H��� ���   )ЉE�[� H��� ���   )ЉE��:�;� H��� ���   )Ѓ��E�"� H��� ���   )Ѓ��E�E�H�� H�E�H	�H�E�H�t� H�@|H�E�H�e� H�@tH���u��u��u���x�����p���H����  H��0H��@���H���  H�������  H��P���H=�  ��   H=� u�H��� H����   H��X���H����   H��X���H��H��t0H��X�����H��t!H�E�   H��X��������C H�H�E��H�E�   H��X������C H�H�E�H��� H�@|H�E�H�q� H�@tH���u��u��u���x�����p���H����  H��0�(H��X���H��u�D����H��X���H��u�8����������������h@C j A�    A�    �   �   �    �    �  H���l� H�H�M��
   H��H���  H�E�H��h@C A��   A��   ��   �    �    H���  H���5� ��� h@C j A�    A��   �   �   ���  H���x� �v� ������H��� H�E�H�@H��H���  �5�� ��� A�@C D��� �   �   ����  �'���UH��H���}��u��}�u'�}���  u��C �   �`C ��C ��@ 襐 ���UH����  �   ����]�UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]ÐUH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H��H�}��u�U�H�E���H���   ��UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H���]"  H�E��ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �-
  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H�� H�}�H�E�H� H�E�H�E�@��tH�E�    H���'�������f.�     L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A����  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�H��H	�t�  �AUI��ATA��I��UH��SH��L)�H��H��H���  M��uH��[]A\A]��    H��I�4H�| L��[]A\A]�E  D  SH���(   ��  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     US�D$L�T$ ��y�1���y�1�E����E��M�ZA��A��A	�E	�A��   ���~OA;r}I��l��t�D  A�BA��D�ȅ�~9�~���
���A9B~A�E��9�u�9�t	��A9Z�[]�ff.�     D��SE������AQ��A��P�D���XZ[�H��I��H��A��H�� ��H�� ������� AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   �CA9���   D��D��D�\$�NfD  ��L�[�D��    G�L��L�KD��x��E�9E� H�{D�D9�t=�C����9�~0��D�BD�L= �zI�H�A��u��?u�A�8u�D9�u�D  D�\$E)�9t$t��9s�F���H��[]A\A]A^A_��    AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�w���XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_ÐH��H��A��H��APH�� A��H�� ����m���H����     �NH��H�� ��~zAVAUATUS�O��)���~^I��I����E1��f�A�F)�D9�~DA�EB�<#A�~��    A��Hc�A������4�    Hc�I~Hc�Iu�w���E9e�[]A\A]A^���    �NA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      H���   HD���  ff.�     @ ��  ff.�     �  ff.�     �����ff.�     �  ff.�     �  f.�     �UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo% #@ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo% #@ f��fs�f��f H����H��]Ð�����������                AW�B��A��AVAUE��ATU��SH��H�àC �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�:���_AXA��@�w���A��AV�   ��RD�L$A��   D�D$����Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�����XZA���%���A��AVA��   RD�L$�   ��D�D$����A[XA�������A��AVA��   RD�L$�   ��D�D$�l���AYAZA�������A��AVA��   RD�L$�   ��D�D$�7���_AXA�������A��AV�   ��RD�L$A��   D�D$����A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃������XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_�UH��H�� H�}�u�H�U�H�E�A�    A�    �    H�ƿ   �  �E���UH��H���}��E�H�A�    A�    �    �    H�ƿ   �  ���UH��H��0�}�H�u�H�U�H�u�H�U��E�H�H�M�A�    I��H�ƿ   �J  �E���UH��H��0�}�H�u�H�U�H�u�H�U��E�H�H�M�A�    I��H�ƿ   �  �E���UH��H�� �}�H�u��U�H�u��E�Hc�H�U��E�H�A�    I��H�ƿ   ��   H�E���UH��H��0�}�H�u�H�U�H�u�H�U؋E�H�H�M�A�    I��H�ƿ!   �   H�E���UH��H�� H�}�H�U�H�E�A�    A�    �    H�ƿ   �S   H�E���UH��H��0H�}�H�E H�E�H�E(H�E�H�E0H�E�H�u�H�M�H�U�H�E�A�    I��H�ƿ   �   ���UH��SH�}�H�u�H�U�H�M�L�E�L�M�H�E�L�E�H�M�H�U�H�u�H�}�L���i�[]�UH��H�� H�}�H�E�    H�U�H�E�A�    A�    �    H�ƿ   ����H�E���UH��H�}؉u�H�E�H�E�H�E�H�E��E�    �	H�E��E��Eԃ�9E�|��E�    �/H�E�� �E�H�E��H�E�H�E��U�H�E�H�m��E��Eԉ������9E�|��]�UH��H��0H�}�H�u��U��E�    H�}� ��   �E��P�U�Hc�H�E�H�� 0�E�Hc�H�E�H��  H�E��   �E�Hc�H�E�H�H��H�ЉE��}�	~
�E���W����E���0���E��P�U�Hc�H�E�HЈ�E�Hc�H�E�H�H��H�E�H�}� u��E�Hc�H�E�H��  �U�H�E���H������H�E���UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�sH�U�H�E�HЋU�H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�H;E�s"H�U�H�E�H�H�M�H�U�H�� �H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H;E�s4H�E�    H�E�H;E�sgH�U�H�E�H�H�M�H�U�H�� �H�E���H�E�    H�E�H;E�s3H�E�H+E�H�P�H�E�H�H�E�H+E�H�P�H�E�H���H�E���H�E�]�UH��H�}�H�E�    H�E�    H�U�H�E�H�� ��tH�E�H�E���H�E�]�UH��H��H�}�H�E��    H���|   fH~�H�E��E���UH��H��H�}�H�E��
   �    H����   ��UH��H��H�}�H�E��
   �    H���   ��UH��H��H�}�H�E��
   �    H����  ��UH��H�� H�}�H�u�H�U�H�E�H��H���+  fH~�H�E��E���UH��H��H�}�H�u�H�U�H�E�H��H���E  ��UH��H�� H�}�H�u�H�U�H�E�H��H���l  �}�H�E��U�H�E��U��m���UH��H��0H�}�H�u��U�H�E�� ��t"H�E�� �����e  ������uH�E��ԐH�E�� <+uH�=� �:   H�59� H�=[� 蒖 �E� H�E�� <-u	�E�H�E��}�
t@�}� tH��� �B   H�5�� H�='� �O� �U�H�M�H�E�H��H���   �   H�E�    H�E�� ��tGH�E�� </~<H�E�� <91H�U�H��H��H�H�H��H�E�� ����0H�H�H�E�H�E��H�}� tH�E�H�U�H��}� t	H�E�H���H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H��`H�}�H�u��U�H�E�����H�E�H�E��E�    H�E�H�PH�U�� ���E�E���d  ������t�փ}�-u�E�   H�E�H�PH�U�� ���E���}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��E�Hc�H�������    H��H�E؋E�Hc�H�������    H��H�ЉE�H�E�    �E�    �E���a  ������t�m�0�4�E���`  ��������   �E����c  ��t�7   ��W   )E�E�;E�}r�}� xH�E�H9E�rH�E�H9E�u�E�;E�~	�E������*�E�   �E�Hc�H�E�H��H�EȋE�Hc�H�E�H�H�E�H�E�H�PH�U�� ���E��<�������}� y
H�E�������}� tH�E�H��H�E�H�}� t�}� t
H�E�H���H�E�H�U�H�H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H�� C H����  %���]�UH��H��H�}�H��� ��   H�5w� H�=�� �В UH��H���}��E���H�� C H����  ���UH��H��   ��\���H��`���H�ªC H��H����  H��`���H�5f� H���  H���=  H��`���H����  ���UH��H�� H�}�H�u�H�U�H�M�H�E�H��H����
  �E��}� tdH�%    H������H�E���    �H�E���UH��H�� H�}�H�u�H�E�H�E�H���!	  H�E�H�}� u�    �!H�E�H�E�H��H�E��    H������H�E���UH��H�?� ��   H�5-� H�=h� 膑 UH��H��H�}�H�E��    �    H����s �    ��UH��H��H�}�H��� ��   H�5�� H�=� �2� UH��H���}���s �E����w UH��H���}��E����w UH��H���}�H��� ��   H�5�� H�=�� �ِ UH��H��H�}�H��� ��   H�5U� H�=�� 讐 UH��H��H�}�H�h� ��   H�5*� H�=e� 胐 UH��H��`H�}�H�u�H�U�H�M�L�E�H�E�    H�E�H�E�H�E�H;E�s|H�E�H+E�H��H�E�H�U�H�E�H�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���ЉE܃}� yH�U�H�E�H�H�E�뛃}� ~H�U�H�E�H�H��H�E��H�E��.H�E�H;E�tH��� ��   H�5O� H�=�� 訏 �    ��UH��H��`H�}�H�u�H�U�H�M�H�E�    H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�E�H��H�E�H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���Ѕ�����ufH�E�H�E�H�E�H�E�H�E�    H�E�H;E�sEH�U�H�E�H�� �E�H�U�H�E�H�H�M�H�U�H�� �H�U�H�E�H��EǈH�E�벐H�E��M���H�E��������UH��H���}�H�a� �  H�5� H�=H� �f� UH��H��H�}�H�:� �  H�5�� H�=� �;� UH��H��H�}�H�� �  H�5�� H�=�� �� UH��}�u�E��}�E��E��}�ЉE�H�E�]�UH��H��H�}�H�u�H��� �'  H�5b� H�=�� 軍 UH��H��H�}�H�u�H��� �+  H�53� H�=n� 茍 UH��SH��HH�}�H�u��
x H�E�H�E�H�E�H�U�H�E�H�H�E�H�E�H�E�H�E�H��H�E�H�}� uOdH�%    H������f�   dH�%    H������f�@  dH�%    H�������@    H�E��@	���bH�E�H� H��H�dH�%    H������H��H�U�H�u�H�E�H���ӉE�}� tH��� �;  H�5>� H�=�� 藌 H�E�H+E�H��H[]�UH��H���   H��X���H��P���H��H���H��`���H�ªC H��H����  H��`���H�5�� H����  H���  H��`���H����  H��X���H��uH�� �@  H�5�� H�=[� ��� H��P���H��uH��� �A  H�5s� H�=3� �̋ H��H���H��uH��� �B  H�5H� H�=� 衋 H��P���� ��uH��� �C  H�5� H�=�� �t� H��P����H��X����҉�   ��UH��H��H�}��u�H�K� �H  H�5�� H�=� �)� UH��H��pH�}�H�u�H�U��u H�E�f�E�  f�E�  �E�    H�E�    H�E�    H�E�H�E�H�E�H�E�H�E�H��    H�E�H�H�E�H�}� uNH�E�H� H�� H� H�M�H�U�H�u�H�}��ЉE�}� tH��� �U  H�5� H�=�� �s� H�E��H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� tH�P� �Z  H�5�� H�==� �%� H�E�H+E�H��H�E�H�E�H;E�sH�E�H��    H�E�H��     H�E���UH��H�� H�}�H�u�H�U�H��� �e  H�5`� H�=�� 蹉 UH��H��P  H������H�=� ��j  H��������   H������H�ªC H��H����  H������H�5�� H���  H��H������H��H���L  H���  H������H����  H��������H��tIH��`���H�ªC H��H���  H�EH��H��`���H��H����  H����  H��`���H���{  �o H��H������H��H����  ���UH��H��   H��X����o H��H��X���H��H���&  H�E�H�=�� �i  H������tXH��`���H�ªC H��H����  H��`���H�5�� H����  H��H�E�H��H���9  H���  H��`���H����  H�E���UH��H��   H��X���H��P�����n H��H��P���H��X���H��H���$  H�E�H�=H� ��h  H������t|H��`���H�ªC H��H���#  H��`���H�5b� H���C  H��H��X���H��H���  H�5[� H���  H��H�E�H��H���c  H���/  H��`���H����  H�E���UH��SH��8H�}�H�u�H�U�H�E�H��w
�  �   H�E�H�P�H�E�H!�H��t�  �~��m H��H�U�H�E�H��H���L  H� H��H���k  H�E�H�}� u�  �CH�E�H�P�H�E�H!�H��tH��� ��  H�58� H�=�� 葆 H�E�H�U�H��    H��8[]�UH��H�� H�}�H�u�H�U�H��� ��  H�5� H�=)� �G� UH��H���}��u��}�u�}���  uH�� C H���   ���UH����  �   ����]�UH��H��H�}�H�E��q  H���   ���UH��H�}��u�H�E��U�H�E�ǀ�	     H�E����	  =o  wH�E����	  �P�H�E�Hcҋ�H�E����	  �P�H�E�Hcҋ���1�i�e�lH�E����	  ��H�E����	  �H�E�Hc҉�H�E����	  �PH�E����	  �x����]ÐUH��H�}��E�    �E�߰�H�E؋��	  =o  �N  �E�    �}��   kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE�E����  H�E�Hcҋ��U���1E�����D����1�H�E؋U�Hc҉��E���E��   �}�n  kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE��E������H�E�Hcҋ��U���1E������D����1�H�E؋U�Hc҉��E��H�E؋��	  %   ���H�E؋ %���	ЉE�H�E؋�0  �U���1E�����D��1�H�E؉��	  H�E�ǀ�	      H�E؋��	  �HH�U؉��	  H�U�H����E�E���1E�E���%�V,�1E�E���%  ��1E�E���1E�E�]�UH��H�}�H�u�H�E�]ÐUH��H��H�}�H�E��     H�E��@    H�E�H��H���M  H�E��@ H�E��@ H�E��@ H�E��@ H�E��@ ���UH��H��H�}�H�u�H�E��H�E��H�E��PH�E��PH�E�H��H�U�H��H��H���  H�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��P��ÐUH��H��H�}�H�E�H��H���  ��ÐUH��H�� H�}�H�u��U�H�U�H�E�H��H���&���H�E��U��H�E���UH��H�}�H�E�H�     H�E�H�@    H�E�H�@    H�E�H�@    H�E�H�@     H�E��@(    �]�UH��H�}�H�E�H��?]�UH��H��H�}�H�U��   �������tH��� �   H�5�� H�=� �j� ���UH��H�}�H�E��    ��]�UH��}�H�E�   �E�H9E�vH�� B �U�H���U�E�   �E�H+E�H��H�E�E�H+E�H�P�E��H�H!�H�E�H�E�H��H�E؋E�Hc�H�E�H�H�E؉�H��H��]�UH��H��@H�}�H�E�   H�E������_���H9E�����tG�E�    �E�H�U�H��H9�s#�E����3���H9E�����t�E��   �E���H�E�H���   H�E�H������H��?   H)�H��H�E�H�E�H�E�H�E�H��H�E�H�E�   ��H��H�E�H)�H��H�E�   ��H��H��H�H�P�H�E���H��H��H�E�H�U�H�E�H�H�E�H�H����UH��H��H�}�H�E�H���P  H�E��@ ��ÐUH��H��H�}�H�E�H���8  ��ÐUH��H��H�}�H�u�H�E�H���  H�E��PH�E��PH�E��@��tH�E�H�ƿ   �����H��H�E�� ����UH��H��PH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH�P� �   H�5� H�=� �~ f���E�H�E��.   H���U H�E�H�E�H���1���H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� ����� K  �������  �M���� �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   �?� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH�&� �&   H�5�� H�=� �} H�E�H;E�sbH�E�H�E�� �����KJ  ������uBH�E�� ����0�*��^E��M��X��E��M���� �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E��~]� fW��E��E���UH��H��@H�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH�� �   H�5�� H�=�� �p| f���E�H�EȾ.   H���rS H�E�H�E�H�������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� ������H  �������  �M��L� �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   �
� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�5m� H�=�� �F{ H�E�H;E�sbH�E�H�E�� ������G  ������uBH�E�� ����0�*��^E��M��X��E��M��W� �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E��0� W��E��E���UH��H��pH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH��� �   H�5K� H�=t� �$z ���}�H�E��.   H���*Q H�E�H�E�H������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sNH�E�� �����F  ��������   �m��-(� ���}�H�E�� ����0�E��E��m����}�H�E��H�}� ��   �-�� �}�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�55� H�=^� �y H�E�H;E�sVH�E�H�E�� ������E  ������u6H�E�� ����0�E��E��m����m����}��m��-G� ���}�말����H�}� tH�E�H�U�H��}� t�m����}��m���UH��H��H�}�H�u�H�U�H�E�H��H���  H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���  H�E��ÐUH��H��H�}�H�E�H� H�U�H��H��H���(  H�E���UH��H��H�}�H�u�H�U�H�E�H��H���%  H�E��ÐUH��SH��xH�}�H�u�H�}� �D  H�E�H�E�H�E�H�PH�E�H��H���)  H�U�H�E�H��H���p  H�E�H�}� uH��    H��uH�=� �볿�H�E�� ����   H�E�H�@H9E�tH��    H��uH�=� 贳��H�E�H�PH�E�H��H����  H�E�H�P H�E�H�@H   H��H)�H�E�H�P H�E�H���P  H�E�H� H�U�H�RH��   H�U�H�RH�� ���H��H��H���^ �    �   H�E�� ��tH��    H��uH�=ϱ �
���H�E�H����  H�E�H�E�H�E�H%  ��H��H�E�H9�tH��    H��uH�=� �Ʋ��H�E؋@HH�H��H��H��H�E�H�H��H�E�H�E؋@H������H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=	� �T���H�U�H�E�H��H���G	  H�E�H�@PH�����E�H�E؋@L��uH��    H��uH�=0� ����H�E�H�ƿ   �	���H��H���#  H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H���  ����t�   ��    ��tH��    H��uH�=� 薱��H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H����
  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���
  H�E�H���L  �   H�E�H���;  ����H��x[]�UH��SH��   H��x���H��p���H��p��� uHǅp���   H��p��� �  ��  H��p���H���J����E�}�~H��    H��uH�=y� 脰���E�H�H��H��H��H��x���H�H��H�E�H�U�H�E�H��H���U  H�E�H�@H���*  H�E�H�@H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=P� ����H�E�H�U�H��H���:	  ����tH��    H��uH�=l� �ϯ��H�E�H� H��t$H�E�H�U�H�H��H����  ����t�   ��    ��tH��    H��uH�=y� �|���H�E�H�H�E�H�PPH�E؋@L�PH�E؉PLH�E�H�@PH���$  H�E�H�PH�E�H��H���	  H�E�H��H���h
  H��H�E�H�P��  H�E�H����  �U�H��x�����H���
  H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=F� �����H�E�H�U�H��H����  ����tH��    H��uH�=b� 荮��H�E�H� H��t$H�E�H�U�H�H��H���  ����t�   ��    ��tH��    H��uH�=o� �:���H�E�H�H�E�H�PPH�EЋ@L�PH�EЉPLH��x���H�PH�E�H��H���  H��x���H�PH�E�H��H����
  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H���  H�E�H���w  H�E�H�@PH��uH��    H��uH�=9� �|���H�E�H�PH�E�H��H����  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���_  H�E�H����  H�]�H�E�H���C  �   H��p���H�  H% ���H�E�H�U�H��x���H��H����
  H�E�H��x���H�PH�E�H��H����  H��x���H�PH�E�H��H���	  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H���N  H�E�H�@H��H�E�H���  H��H�Ĉ   []�UH��SH��hH�}�H�u�H�U�H�}� uH�U�H�E�H��H���!���H����  H�}� uH�U�H�E�H��H�������    �  H�E�H�E�H�E�H�PH�E�H��H����  H�U�H�E�H��H���  H�E�H�E�H���  H�}� uH��    H��uH�=�� 舫��H�E�� ����   H�E�H�E�H�E؋@H������H�E�H�E�H;E�w	H�]��  H�U�H�E�H��H���C���H�E�H�}� u
�    ��   H�U�H�M�H�E�H��H������H�U�H�E�H��H������H�]��   H�E�� ��tH��    H��uH�=Q� �̪��H�E�H�@H9E�tH��    H��uH�=�� 褪��H�E�H�@H9E�sH�]��WH�U�H�E�H��H������H�E�H�}� u�    �2H�E�H�PH�M�H�E�H��H���`���H�U�H�E�H��H�������H�]�H�E�H���e  H��H��h[]�UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]�UH��H�}��]ÐUH��H�}��]ÐUH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H������H�E�H� H�U�H�M�H��H���2  H�E�H���|�����ÐUH��H��H�}�H�u�H�E�H�U�H��H���wl ���UH��H��0H�}�H�u�H�E�H���F���H�E�H� H�U�H�M�H��H����  H�E�H��������ÐUH��H��H�}�H�u�H�E�H�U�H�H�E��@ H�E�H���  ���UH��H��H�}�H�E��@��tH�E�H���  ��ÐUH��H�� H�}�H�u�H�E�H��H����  H�E�H�}� ��   H�E�H�@H9E�sH�E�H����  H�E���H�E�H�PH�E�H�@H�H9E�rH�E�H���  H�E��H�E�H�@H9E�rH�E�H�PH�E�H�@H�H9E�rH��    H��uH�=2� �姿�H�E���    ��UH��H��0H�}�H�u�H�E�H���1  H�E�H�E�H���?  H�E�H�}� uH�U�H�M�H�E�H��H���<  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���o	  H�E�H�E�H����  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���Q	  ���UH��H��H�}�H�E��@����tH��    H��uH�=Ĭ �禿�H�E�H� H�������H�E��@ ��ÐUH��H�}�H�E�H�     �]�UH��H�}�H�u�H�E�H�E�H�E�H�@H9E�r H�E�H�PH�E�H�@H�H9E�s�   ��    ]ÐUH��H�� H�}�H�u�H�E�H���  H������tH�E�H�U�H��H���  �   H�E�H����
  H�E�H�E�H�HH�U�H�E�H��H���=  ��tAH�E�H���U  H������tH�E�H�U�H�M�H��H���R  �VH�E�H���&  H�E��H�E�H���i  H������tH�E�H�U�H�M�H��H���g  �H�E�H���:  H�E��\�����UH��H��0H�}�H�u�H�E�H���
  H�E�H�E�H���  H�E�H�}� uH�U�H�M�H�E�H��H���8  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���k  H�E�H�E�H���N
  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���M  ���UH��H�� H�}�H�E�H���b	  H�E�H�}� u�    �,H�E�H����	  H������tH�E�H����	  H�E���H�E���UH��SH��XH�}��u�H�E�H� �   H���6O H�E�H�E�H�� H%  ��H�EЋE����B���H�E�H�E�    H�}�   w
H�E�HE���H�}��� vH��    H��uH�=� �ڣ��H�E�H�ƿ�   �����H�ø   H+E�H�M�H�U�H�4�U���H��H���  H�]�H�E�    H�E�    H�E�H�@H9E�sHH�E�H�PH�E�H�H�ƿ   �r���H��H������H�]�H�E�H�U�H�H�E�H�E�H�E�HE��H�E�H�U�H�PPH�E�H��X[]�UH��H�� H�}�H�u�H�E�H���h  H������tH�E�H�U�H��H���e  �   H�E�H���:  H�E�H�E�H�HH�U�H�E�H��H����  ��tAH�E�H���  H������tH�E�H�U�H�M�H��H���n  �VH�E�H����  H�E��H�E�H����  H������tH�E�H�U�H�M�H��H���e  �H�E�H����  H�E��\�����UH��H��H�}�H�E��@��tH��    H��uH�=� �����H�E�H� H������H�E��@���UH��SH��(H�}�H�u�H�E�%�  H��tH��    H��uH�=|� 觡��H�E�H� H�U�H��   H��H���L H�E�H�E�H�ƿH   ����H��H�E�H��   H�E�H���   H���  H�]�H�E�H��([]�UH��H�� H�}�H�u�H�U�H�U�H�E�H��H����  ���UH��H��`H�}�H�u�H�U�H�E�H�5-� H���  H�E�H���	���H�E�H�M�   H��H������H�E�H�U�H�M�H��H���-  H�E�H������H�E�H��������ÐUH��H�}�H�E�H� ]�UH��H��H�}�H�E�H���  H�@��UH��H��H�}�H�E�H���i  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���G  H�E�H�}� tH�]�H�E�H���  H�X H�}� tH�]�H�E�H����  H�XH�E�H����  �@(������t8H�E�H���  ��tH�E�H����  �@(   �H�U�H�E�H��H���  H�E�H�������H��uH�E�H������H9E�t*H�E�H�������H9E�uH�E�H�������H��t�   ��    ��tH��    H��uH�=_� �"���H�E�H���S  H�E�H�}� uH�E�H�U�H��rH�E�H���g���H9E�����tH�]�H�E�H����  H�X�EH�E�H���X���H9E�����tH��    H��uH�=�� 蠞��H�]�H�E�H���  H�XH�}� tH�]�H�E�H���  H�H�E�H���z  H�@    H�E�H���f  H�@    H�E�H���R  H�     H�E�H���?  H�@    H�E�H���+  H�@     H�}� tH�U�H�E�H��H���O  �H��H[]�UH��H��H�}�H�E�H����  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H��� ���H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���b  H�X�EH�E�H�������H9E�����tH��    H��uH�=\� ����H�]�H�E�H���  H�XH�]�H�E�H���  H�H�E�H����  �X(H�E�H����  �X(H�]�H�E�H����  H�XH�}� tH�]�H�E�H���  H�H�]�H�E�H���  H�XH�}� tH�]�H�E�H���  H�H�E�H���}���H������tH�]�H�E�H���c���H���\  H�X H�E�H���K���H��H�E�H���=  H�XH�E�H���C  H��H�E�H���  H�X H�E�H���$  H������tH�]�H�E�H���
  H����  H�XH�E�H����  H�@    H�E�H����  H�@    H�E�H���  H�     H�E�H���  H�@    H�E�H���  H�@     H�U�H�E�H��H���   H�U�H�E�H��H���  �H��H[]ÐUH��H�}�H�E�H� ]ÐUH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=�� �����H�E�H�U�H�H�U�H�E�H��H���  H�U�H�E�H��H���  ���UH��H�}�H�u�H�U�H�E�H�PH�E�H�@H9���]�UH��H��H�}�H�E�H���  H�@��UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�==� �H���H�E�H������H������tH��    H��uH�=]� ����H�]�H�E�H���@  H�XH�]�H�E�H���,  H�H�E�H���T  H�E�H�}� tH�]�H�E�H���  H�X H�]�H�E�H����  H�XH�]�H�E�H����  H�X H�]�H�E�H����  H�XH�U�H�E�H��H���9  H�U�H�E�H��H���  H�U�H�E�H��H���3  �H��8[]�UH��H��H�}�H�E�H���i  H�@�ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=�� ���H�E�H������H������tH��    H��uH�=�� ���H�]�H�E�H����  H�XH�]�H�E�H����  H�H�E�H���%  H�E�H�]�H�E�H���  H�X H�]�H�E�H���  H�XH�]�H�E�H���  H�X H�}� tH�]�H�E�H���p  H�XH�U�H�E�H��H����  H�U�H�E�H��H���\  H�U�H�E�H��H����  �H��8[]ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���W  H�E�H�}� tH�]�H�E�H����  H�X H�}� tH�]�H�E�H����  H�XH�E�H���  �@(������t8H�E�H���  ��tH�E�H���  �@(   �H�U�H�E�H��H���  H�E�H������H��uH�E�H�������H9E�t*H�E�H���i���H9E�uH�E�H������H��t�   ��    ��tH��    H��uH�=� �Ɩ��H�E�H���c  H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���  H�X�EH�E�H��� ���H9E�����tH��    H��uH�=)� �D���H�]�H�E�H���l  H�XH�}� tH�]�H�E�H���Q  H�H�E�H���B  H�@    H�E�H���.  H�@    H�E�H���  H�     H�E�H���  H�@    H�E�H����  H�@     H�}� tH�U�H�E�H��H����  �H��H[]�UH��H��H�}�H�E�H���  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H�������H�E�H�}� uH�E�H�U�H��rH�E�H���o���H9E�����tH�]�H�E�H���*  H�X�EH�E�H������H9E�����tH��    H��uH�= � 軔��H�]�H�E�H����  H�XH�]�H�E�H����  H�H�E�H����  �X(H�E�H���  �X(H�]�H�E�H���  H�XH�}� tH�]�H�E�H���  H�H�]�H�E�H���p  H�XH�}� tH�]�H�E�H���U  H�H�E�H���}���H������tH�]�H�E�H���c���H���$  H�X H�E�H���K���H��H�E�H���  H�XH�E�H���S  H��H�E�H����  H�X H�E�H���4  H������tH�]�H�E�H���  H���  H�XH�E�H���  H�@    H�E�H���  H�@    H�E�H���|  H�     H�E�H���i  H�@    H�E�H���U  H�@     H�U�H�E�H��H����  H�U�H�E�H��H���=  �H��H[]ÐUH��H�� H�}�H�u�H�U�M�H�E�H�M�H�U�   H���  H�E��U�PHH�E��@L    H�E�H�@P    H�E�H��XH����������UH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=� �L���H�E�H�U�H�H�U�H�E�H��H����
  H�U�H�E�H��H����  ���UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=՚ �����H�E�H���I���H������tH��    H��uH�=�� 谑��H�]�H�E�H���  H�XH�]�H�E�H���  H�H�E�H������H�E�H�}� tH�]�H�E�H���v  H�X H�]�H�E�H���b  H�XH�]�H�E�H���N  H�X H�]�H�E�H���:  H�XH�U�H�E�H��H���	  H�U�H�E�H��H���V	  H�U�H�E�H��H���  �H��8[]ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=E� 訐��H�E�H���/���H������tH��    H��uH�=e� �x���H�]�H�E�H���|  H�XH�]�H�E�H���h  H�H�E�H���o  H�E�H�]�H�E�H���E  H�X H�]�H�E�H���1  H�XH�]�H�E�H���  H�X H�}� tH�]�H�E�H���  H�XH�U�H�E�H��H���y  H�U�H�E�H��H���  H�U�H�E�H��H���w  �H��8[]ÐUH��H�� H�}��u�H�U�H�M�H�E��U�H�E�H�U�H�PH�E�H�U�H�PH�E�H��H���������ÐUH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=W� ����H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���b  �UH�E�� ��t%H�E�� ��tH��    H��uH�=�� ����H�u�H�E�A�    A�   �    �
   H���  ���UH��H�}��   H�E�H�]�UH��H��H�}�H�E�H�������H�@ ��UH��H��H�}�H�}� u�    �H�E�H�������@(�����ÐUH��SH��XH�}�H�u�H�E�H���}����@(������tH��    H��uH�=�� �B���H�E�H���s  H�E�H�}� �\  H�E�H������H9E�������   H�E�H������H������tH��    H��uH�=�� �܌��H�E�H���c���H��������@(��������   H�E�H���>���H�E�H�E�H���.���H��H�E�H��H���-  H�E�H�������H9E�����tH��    H��uH�=]� �X���H�E�H���`����@(   H�E�H���M����@(   H�E�H������H�E��  H�E�H������H9E�����tH��    H��uH�=Q� �싿�H�E�H���U���H������tH��    H��uH�=�� 輋��H�E�H���%���H�������@(������tzH�E�H������H�E�H�U�H�E�H��H���  H�E�H�������H9E�����tH��    H��uH�=d� �G���H�E�H���O����@(   H�E�H���<����@(   H�E�H������H�E�H�E�H���z���H���p  ��tH�E�H������H���X  ��t�   ��    ��toH�E�H��������@(������t+H�E�H��������@(   H�U�H�E�H��H��������  H�E�H�������@(   H�E�H�������@(   �  H�E�H���j����@(�E�H�E�H������H9E������  H�E�H������H���i�����tH�E�H������H���|  ��t�   ��    ��tQH�E�H���^���H�E�H�U�H�E�H��H���  H�E�H��������@(   H�E�H��������@(   H�E�H�E�H�E�H���+���H�����������tH��    H��uH�=� �o���H�U�H�E�H��H���   H�E�H���d����@(   �]�H�E�H���N����X(H�E�H������H���7����@(   �M  H�E�H������H9E�����tH��    H��uH�=Ö �房�H�E�H���m���H��������tH�E�H���7���H���-  ��t�   ��    ��tQH�E�H���-���H�E�H�U�H�E�H��H���'  H�E�H�������@(   H�E�H���x����@(   H�E�H�E�H�E�H������H����������tH��    H��uH�=]� � ���H�U�H�E�H��H���Q  H�E�H�������@(   �]�H�E�H��������X(H�E�H���Q���H��������@(   ��H��X[]�UH��H��H�}�H�E�H������H� ��UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H���_  ����uH�E�H������H�E��Ԑ���UH��H��H�}�H�u�H�E�H���&  ��ÐUH��H��H�}�H�u�H�E�H���  ��ÐUH��H�� H�}�H�u�H�E�H���	  H�E�H�}� uH�E�H���#  �@(   �  H�E�H���  �@(   H�E�H����  �@(��������  H�E�H���L	  H�E�H�}� tH�E�H����  �@(��t�   ��    ��tH��    H��uH�=� �Z���H�E�H������H9E�uH�E�H�������H����  ��t�   ��    ��tYH�E�H���L  �@(   H�E�H���9  �@(   H�E�H������H���  �@(   H�U�H�E�H��H��������  H�E�H���r���H9E�uH�E�H������H���U  ��t�   ��    ��tYH�E�H���  �@(   H�E�H���  �@(   H�E�H������H���  �@(   H�U�H�E�H��H�������j  H�E�H������H9E�������   H�E�H�������H9E�����t;H�U�H�E�H��H����  H�U�H�E�H��H���~  H�E�H���  �@(   �&H�U�H�E�H��H���V  H�E�H����   �@(   H�E�H����   �@(   �   H�E�H���4���H9E�����tH��    H��uH�=e� �X���H�E�H������H9E�����t;H�U�H�E�H��H����  H�U�H�E�H��H���  H�E�H���G   �@(   �&H�U�H�E�H��H����  H�E�H���   �@(   H�E�H���   �@(   ����UH��H�}��X   H�E�H�]�UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H���z  ����uH�E�H���  H�E��Ԑ���UH��H��H�}�H�E�H������H�@ ��UH��H��H�}�H�}� u�    �H�E�H���^����@(�����ÐUH��SH��XH�}�H�u�H�E�H���5����@(������tH��    H��uH�=� �ւ��H�E�H���s  H�E�H�}� �\  H�E�H������H9E�������   H�E�H���K���H������tH��    H��uH�=� �p���H�E�H������H�������@(��������   H�E�H�������H�E�H�E�H�������H��H�E�H��H���  H�E�H���s���H9E�����tH��    H��uH�=� �쁿�H�E�H�������@(   H�E�H�������@(   H�E�H���q���H�E��  H�E�H���\���H9E�����tH��    H��uH�=� 老��H�E�H�������H������tH��    H��uH�=� �P���H�E�H������H���t����@(������tzH�E�H������H�E�H�U�H�E�H��H���  H�E�H������H9E�����tH��    H��uH�=�� �ۀ��H�E�H�������@(   H�E�H��������@(   H�E�H������H�E�H�E�H�������H����  ��tH�E�H���8���H���  ��t�   ��    ��toH�E�H�������@(������t+H�E�H���x����@(   H�U�H�E�H��H��������  H�E�H���M����@(   H�E�H���:����@(   �  H�E�H���"����@(�E�H�E�H���:���H9E������  H�E�H������H���i�����tH�E�H���\���H����  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���  H�E�H�������@(   H�E�H�������@(   H�E�H�E�H�E�H�������H�����������tH��    H��uH�=�� ���H�U�H�E�H��H����  H�E�H�������@(   �]�H�E�H�������X(H�E�H���v���H��������@(   �M  H�E�H���V���H9E�����tH��    H��uH�=W� �z~��H�E�H���%���H��������tH�E�H������H���  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���  H�E�H���C����@(   H�E�H���0����@(   H�E�H�E�H�E�H���?���H����������tH��    H��uH�=� �}��H�U�H�E�H��H���C	  H�E�H��������@(   �]�H�E�H�������X(H�E�H�������H�������@(   ��H��X[]�UH��H��H�}�H�E�H���w���H� ��UH��H�� H�}�H�u�H�E�H���[���H�E�H�}� uH�E�H�������@(   �  H�E�H�������@(   H�E�H��������@(��������  H�E�H�������H�E�H�}� tH�E�H�������@(��t�   ��    ��tH��    H��uH�=� �v|��H�E�H�������H9E�uH�E�H�������H��������t�   ��    ��tYH�E�H���D����@(   H�E�H���1����@(   H�E�H������H�������@(   H�U�H�E�H��H��������  H�E�H���j���H9E�uH�E�H���:���H��������t�   ��    ��tYH�E�H�������@(   H�E�H�������@(   H�E�H�������H�������@(   H�U�H�E�H��H�������j  H�E�H������H9E�������   H�E�H������H9E�����t;H�U�H�E�H��H���  H�U�H�E�H��H���<  H�E�H��� ����@(   �&H�U�H�E�H��H���  H�E�H��������@(   H�E�H��������@(   �   H�E�H���,���H9E�����tH��    H��uH�=�� �tz��H�E�H�������H9E�����t;H�U�H�E�H��H���  H�U�H�E�H��H����   H�E�H���?����@(   �&H�U�H�E�H��H���   H�E�H�������@(   H�E�H�������@(   ����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H��H�}�H�}� u�   �H�E�H���{����@(������UH��SH��8H�}�H�u�H�E�H���|���H�E�H�}� tH�E�H������H9E�t�   ��    ��tH��    H��uH�=e� ��x��H�E�H���a���H�E�H�E�H������H�E�H�}� tH�]�H�E�H�������H�H�]�H�E�H�������H�XH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H������H�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���I���H�X�EH�E�H������H9E�����tH��    H��uH�=Ӈ ��w��H�]�H�E�H������H�XH�U�H�E�H��H���y���H�U�H�E�H��H���f����H��8[]�UH��SH��8H�}�H�u�H�E�H�������H�E�H�}� tH�E�H�������H9E�t�   ��    ��tH��    H��uH�=�� �Xw��H�E�H�������H�E�H�E�H���y���H�E�H�}� tH�]�H�E�H���5���H�H�]�H�E�H���"���H�XH�]�H�E�H������H�H�]�H�E�H�������H�XH�]�H�E�H�������H�H�}� uH�E�H�U�H��rH�E�H���%���H9E�����tH�]�H�E�H������H�X�EH�E�H������H9E�����tH��    H��uH�=� �^v��H�]�H�E�H���b���H�XH�U�H�E�H��H�������H�U�H�E�H��H��������H��8[]�UH��H�}��    ]�UH��H�}��    ]�UH��SH��8H�}�H�u�H�E�H������H�E�H�}� tH�E�H������H9E�t�   ��    ��tH��    H��uH�=� �u��H�E�H�������H�E�H�E�H���'���H�E�H�}� tH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H���t���H�H�]�H�E�H���a���H�XH�]�H�E�H���M���H�H�}� uH�E�H�U�H��rH�E�H���T���H9E�����tH�]�H�E�H������H�X�EH�E�H���|���H9E�����tH��    H��uH�=u� �t��H�]�H�E�H�������H�XH�U�H�E�H��H���;���H�U�H�E�H��H���(����H��8[]�UH��SH��8H�}�H�u�H�E�H�������H�E�H�}� tH�E�H������H9E�t�   ��    ��tH��    H��uH�='� ��s��H�E�H������H�E�H�E�H������H�E�H�}� tH�]�H�E�H�������H�H�]�H�E�H�������H�XH�]�H�E�H�������H�H�]�H�E�H�������H�XH�]�H�E�H������H�H�}� uH�E�H�U�H��rH�E�H������H9E�����tH�]�H�E�H���o���H�X�EH�E�H�������H9E�����tH��    H��uH�=�� � s��H�]�H�E�H���(���H�XH�U�H�E�H��H������H�U�H�E�H��H�������H��8[]�UH��H��H�}�H�}� u�   �H�E�H��������@(������UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�I� H�E��E�    �E���~H��    H��uH�=2� �5r���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=� ��q���E��P�U�H��D�-H�U�H�E�H��H���   � 9E�����tE�E�    H�U�H�E�H��H���   � �U�)�9E�����t�U�H�E���H���   �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���b   �E��ڋE����E�}� x!�E�H��D���H�E���H���2   �m��ِ��UH��H�}�H�u�H�E��H�E�� 9�}H�E��H�E�]ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=� �p��H�E�H���   H��u)H�E�H� H�U�H��H��H�������H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ���UH��H�� �}�� H�E��E���H�U�H�E���H����  �E�}� t�    ��2 H�E���H���' ����UH��H�� �}�� H�E��E���H�U�H�E���H���  �E�}� t�    ��,2 H�E���H���' ����UH��H�� �}��V H�E��E���H�U�H�E���H���5  �E�}� t�    ���1 H�E���H����' ����UH��H�� �}��  H�E��E���H�U�H�E���H����  �E�}� t�    ��1 H�E���H���~( ����UH��H�� �}�� H�E��E���H�U�H�E���H���  �E�}� t�    ��*1 H�E���H���) ����UH��H�� �}��T H�E��E���H�U�H�E���H���3  �E�}� t�    ���0 H�E���H����* ����UH��H�� �}��� H�E��E���H�U�H�E���H����
  �E�}� t�    ��~0 H�E���H���$+ ����UH��H�� �}�� H�E��E���H�U�H�E���H���
  �E�}� t�    ��(0 H�E���H���+ ����UH��H�� �}��R H�E��E���H�U�H�E���H���1
  �E�}� t�    ���/ H�E���H���$, ����UH��H�� �}��� H�E��E���H�U�H�E���H����	  �E�}� t�    ��|/ H�E���H���, ����UH��H�� �}�� H�E��E���H�U�H�E���H���	  �E�}� t�    ��&/ H�E���H����, ����UH��H�� �}��P H�E��E���H�U�H�E���H���/	  �E�}� t�    ��E����!
  ����UH��H�� �}�� H�E��E���H�U�H�E���H����  �E�}� t�    ��E���������UH��H�� �}��A H�E��M�H�U�H�E���H���	 �E�}� t�    ��>. H�E���H����" ����UH��H�� �}��� H�E��M�H�U�H�E���H��� �E�}� t�    ���- H�E���H���Q# ����UH��H�� �}�� H�E��M�H�U�H�E���H���c �E�}� t�    ��- H�E���H���# ����UH��H�� �}��H H�E��M�H�U�H�E���H��� �E�}� t�    ��E- H�E���H���C$ ����UH��H�� �}��� H�E��M�H�U�H�E���H��� �E�}� t�    ���, H�E���H����$ ����UH��H�� �}�� H�E��M�H�U�H�E���H���j �E�}� t�    ��, H�E���H���& ����UH��H�� �}��O H�E��M�H�U�H�E���H��� �E�}� t�    ��L, H�E���H����& ����UH��H�� �}��� H�E��M�H�U�H�E���H���� �E�}� t�    ���+ H�E���H���m' ����UH��H�� �}�� H�E��M�H�U�H�E���H���q �E�}� t�    ��+ H�E���H����' ����UH��H�� �}��V H�E��M�H�U�H�E���H��� �E�}� t�    ��S+ H�E���H���_( ����UH��H�� �}�� H�E��M�H�U�H�E���H���� �E�}� t�    �� + H�E���H����( ����UH��H�� �}�� H�E��M�H�U�H�E���H���x �E�}� t�    ��E�����  ����UH��H��  H������H������H������H��H����  H������H�5O{ H����  H������H������H������H��H���  ��t
�   �X  H������H�5{ H���  H������H������H������H��H����  ��t
�   �  H������H�5�z H���`  H������H������H������H��H���  ��t
�   ��  H������H�5�z H���  H������H������H������H��H���N  ��t
�   �  H������H�5Wz H����  H������H������H������H��H���
  ��t
�   �H  H������H�5z H���  H������H������H������H��H����  ��t
�   �  H�� ���H�5�y H���P  H�� ���H�����H������H��H���  ��t
�   ��  H�����H�5�y H���  H�����H�����H������H��H���>  ��t
�   �|  H�� ���H�5_y H����  H�� ���H��(���H������H��H����  ��t
�	   �8  H��0���H�5!y H���  H��0���H��8���H������H��H���  ��t
�
   ��   H��@���H�5�x H���@  H��@���H��H���H������H��H���r  ��t
�   �   H��P���H�5�x H����  H��P���H��X���H������H��H���.  ��t�   �oH��`���H�ªC H��H���d���H��`���H�5Rx H��脯��H��H������H��H���o���H�5>x H���`���H��肯��H��`���H���=����    ��UH��H���}�H�u�H��x �  H�5x H�=/x �g' UH��H�� �}��� H�E��E���H�U�H�E���H����   �E�}� t�E���m& H�E���H����$ ��UH��H�� �}�� H�E��E���H�U�H�E���H���y   �E�}� t�E���& H�E���H���T% ��UH��H���}�H��w �  H�5Bw H�=cw �& UH��H���}�H��w �$  H�5w H�=9w �q& UH��H��`H�}���H�U��E��E��E��E���x H�E��@��t�U�H�E���    ��   H�E�H�E�H�E�H��H�E�H�E�H�E�H�E�H��H�E�f�E�  f�E�  �E�    H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� t�E��]H�U�H�E�H9�tH��v �>   H�5wu H�=�u �% H�U�H�E�H9�tH��v �?   H�5Ku H�=�u �l% �    ��UH��}��}�v�}�t�}�v�}��   w�   ��    ]�UH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�PH�E�H�� ��tH�E�H�@H�PH�E�H�P�Ԑ]�UH��H�}�H��H��H��H�E�H�U�H�E�H�PH�E�H9�t�    �LH�E�    H�E�H�@H9E�s1H�E�H�H�E�H��H�M�H�E�H�� 8�t�    �H�E����   ]�UH��ATSH���   H��H��H��H�� ���H�����H�E�    H���C H� H�U�H��H�H� H���F  H���C H� H�U�H��H�H�H�����H��H������H������    �=   H����  H�E�H�}����   H�� ���H�ªC H��H���"���H�� ���H�5gu H���B���H��H�����H����  I��H�����H����  H��H�E�L��H���8  H�U�H�E�H��H��H����  H�5-u H������H���	���H�� ���H���Ī���GH�U�H������    H���  H�E�H�U�H�� ���H�����H�E�H��H��������tH�E��H�E�����H������H���   [A\]�UH���}x ������tRH�=mx �+ ������t=�t	 H��H�=0x �  H�=Dx ��+ H�X` H�5x H��֩@ H���� H��w ]�UH��H�� ����H�E�H�E�H����  H��H���C H� H9�������   H�E�H����  H�E�    H���C H� H�U�H��H�H� H��t+H���C H� H�U�H��H�H�E�H��H���  H�E��H�E�    H�U�H�E�H��H���	  H�E�H���:  H��H���C H�����UH��SH��HH��H��H��H��H��H�u�H�}�H�U��ȈE�����H�E�H�E�H����  H��H���C H� H9�����tH� � �>   H�5,s H�=Ms �! H�U�H�E�H��H������H�E�H�}��t&�}� ��   H�]�H�U�H�E�H��H���  H��fH�E�H����  H� H������tH��� �F   H�5�r H�=�r �  H�]�H�E�H���  H�H�E�    H�U�H�E�H��H����  H�E�H����  H��H���C H��H��H[]�UH��SH��(H��H��H��H�E�H�U��f���H�E�H�E�H���  H��H���C H� H9�����tH� � �Q   H�5�q H�=r �� H�U�H�E�H��H���f���H�E�H�}��uH��    H��uH�=r �0\��H�E�H����  H��vH�E�H���  H� H��t�   ��    ��tH�s� �W   H�5oq H�=r �P H�E�H���w  H�P�H�E�H��H���  H��H�U�H�E�H��H���  H��H���f  H�E�H���  H�E�H���  H�     H�E�H���  H��H���C H��H��([]�UH��H��@H�}�H�U�H�E�H��H���|���H�U�H�E�H��H���:���H�E�H�}��u
�    �   H���C H� H�U�H��H�H�H�E�H��H���-���H�Eк    �=   H���O  H�E�H�}��uH�W� �i   H�5Ap H�=�p �" H�E�H���m  H��H�E�H��H���UH��SH��8H�}�H�U�H�E�H��H������H�Eк    �=   H����  H�E�H�}��uH�� �q   H�5�o H�=�p � �S���H�U�H�Eо    H���=  H�u�H��H��H��H�й   H��H��������    H��8[]�UH��ATSH��  H������H������������H������H�����H��H�������H������    �=   H���  H�E�H�}����   H�� ���H�ªC H��H���[���H�� ���H�5�o H���{���H��H�����H���  I��H�����H���  H��H�E�L��H���q  H�U�H�E�H��H��H����  H�5�o H��� ���H���B���H�� ���H�������dH�%    H�������   �������   H������H������H�����H�5yo H�Ǹ    ��#  ������tH�.� ��   H�5
n H�=So �� H�����H��uH�� ��   H�5�m H�=To �� �m��������� ��D��H�����H������H�E�H��H���[���H�u�H�E�D��H��H��H��������    H��  [A\]�UH��H�� H�}�����H�U�H�E�H��H������H�U�H�E�H��H��������    �ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H�}��H�U؈E�H�E�H�E�H�E�H�@H9E�s#H�E�H�H�E�H�� 8E�uH�E��H�E���H������]ÐUH��H�}�H�E�H� ]ÐUH��H�}�H�E�H�@]�UH��H�� H�}�H��H��H��H�E�H�U�H�U�H�E�H��H���C  H�E���UH��H��0H�}�H�u�H�U�H�U�H�E�H�H�E�H�@H9�vH��    H��uH�=�m �V��H�E�H�H�E�H�H�U�H�E�H��H���  H�E�H�U���UH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�@    H�E�H�@    �]�UH��H�� H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H� H�U�H�RH��H��艡�����UH��H�}�H�E�H�@]�UH��H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H�@    �]�UH��H�� H�}�H�u�H�E�H�@H�PH�E�H��H���I  H�E�H�PH�E�H�@H��H�H�ƿ   �^���H�U�H�H�H�E�H�E�H�@H�PH�E�H�PH�E��ÐUH��SH��(H�}�H�u�H�E�H�@H�PH�E�H��H����  H�E�H���   H��H�E�H�PH�E�H�@H��H�H�ƿ   �֔��H�H�E�H�E�H�@H�PH�E�H�PH�E�H��([]ÐUH��H�}�H�u�H�E�H�@H�U�H��H�]ÐUH��H�}�H�E�H�PH�E�H�@H��H��H�]ÐUH��H�}�H�E�H�@]�UH��H�}�H�E�H� ]�UH��H�� H�}�H�u�H�E�H�������H�E�H�E�H�������H��H�E�H�H�E�H������H��H�E�H����UH��H�� H�}�H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��H�H���a���H�E�H�E���UH��H��0H�}�H�u�H�E�H��裓��H�M�H�U�H�E�H�0H�@H��H���<  H�E�H���i������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��SH��8H�}�H�u�H�E�H�@H9E���   H�E�H�H�E�H�E�H� H�U�H��H��H������H�E�H�E�    H�E�H�@H9E�sHH�E�H�@H�U�H��H�H���g���H��H�E�H��    H�E�H�H�ƿ   虒��H�H�E��H�E�    H�E�H�@H9E�sH�E���H�E�H� H�U�H�RH��H������H�E�H�U�H�PH�E�H�U�H�P��H��8[]�UH��H��PI��H��L��L��H��H�u�H�}�H�U�H�M�H�E�H�E�H�E�    H�E�H9E���  H�U�H�E�H�� �E�}�`v�}�zv�}�@v �}�Zw�E���H�E���H��������q  �}�/v �}�9w�E���H�E���H��������K  �}� uH�E��    H�������/  �E��H�=�k ���  H������t�E���H�E���H���p�����   �}�\uH�E�H�5�k H��������   �}�"uH�E�H�5�k H�������   �}�'uH�E�H�5jk H���v����   �}�
uH�E�H�5Ok H���X����   �}�	uH�E�H�54k H���:����fH�E�H�5"k H���%���H�E�H�M��   H��H��蛑���E�E�H�U�H�M�H�E�H��H���*   H�E�H���Q���H�E��}   H���r���H�E��4������UH��H��@H�}�H�u�H�U�H�U�H�E�H��H���x���H�E؋ H�U�H�M�H�Ή��   H�E�H���������UH��H��@�}�H�u�H�U�H�U�H�E�H��H���+���H�U�H�M��E�H�Ή��   H�E�H��螐�����UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=�v �O���u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�%x H�E��E�    �E���~H��    H��uH�=x �AN���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�w ��M���E��P�U�H��D�-H�U�H�E�H��H�������� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H�������E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���v����E��ڋE����E�}� x!�E�H��D���H�E���H���F����m��ِ�ÐUH��H��H�}�H�~� ��   H�5�w H�=x �B UH��H�� H�}�H�u�H��    H��u<H�J� ��   H�5�w H�=�w � dH�%    H�������   ������@H�U�H�E�H��H���bL���E��}� tdH�%    H������H�E���������    ��UH��H�� �}�H�u��U�H�M�H��� ��   H�5w H�=Lw �s UH��H��� ��   H�5�v H�=)w �P UH��H��H�}�H��� ��   H�5�v H�=�v �% UH��H�� H�}�H�u�H�U�H�]� ��   H�5�v H�=�v �� UH��H��H�}�H�u�H�6� ��   H�5bv H�=�v �� ���UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���#  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L�����UH��H���   H��(���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H���C H� H��0���H��(���H��H���  ��L�����L�����UH��H�}��u�H�U�}���   �E�H��    H��t �H�H��t H���H�E��H�E���]H�E��H�E�f��NH�U�H�E�H��AH�U�H�E�H��4H�U�H�E�H��'H�U�H�E�H��H�E�H�U�H��H�E��H�E����]�UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��� �p  H�5s H�=Xs � UH��H���   H��(���H�� ���H�����H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�����H�� ���H��(���H����  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L�����UH��H�}�H�E�H� � ]�UH��H�}�H�E��@�PH�E��PH�E�H� H�HH�U�H�
� ]�UH��H��   H�����H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�Hǅ0���    Hǅ8���    H�����H��0���ǅ���   ǅ���0   H�EH�� ���H��P���H��(���H�����H�� ���H��0���H��H���I  ��L�����L�����UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���u3  H�U�H�M�H�E�H��H���9  H�M�H�U�H�u�H�E�H��H���#9  H�E��ÐUH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H���o H�E�H��tH�E�H� �U��҉�H��� H�E�H��t�E���    ��UH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H��� H�E�H��tH�E�@�PH�E�PH�E�H��t�E���    ��UH��H��@H�}�H�u�H�U�H�}� t
H�E�H����    H�E�H�E�    H�E�    H�E�H�E�H�U�H�M�H�E�H��H���b$  ���UH��H��H�}�H�u�H���C H� H�U�H�M�H��H���8�����UH��H��H�}�H�u�H��� ��  H�5�n H�=�n �� UH��SH��   H�}�H�u�H��x���H��p���H�}� u
�    �   H�M�H��p���H�H�VH�H�QH�FH�AH�E�H�P�H�M�H�E�H��H���3  H�U�H�M�H�E�H��H����=  H�M�H��x���H�u�H�E�H��H����=  H�]�H�E�H��H�E�H�E�H�PH�E�H��H���D  H� H��  H�E�H�Ĉ   []�UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���1  H�U�H�M�H�E�H��H���QD  H�M�H�U�H�u�H�E�H��H���`D  H�U�H�E�H��  H�E���UH��H�� H�}�H�u�H�U�H�� ��  H�5�l H�=7m �^ UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��� ��  H�5�l H�=&m �� UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�A� ��  H�5l H�=�l �n UH��H�� H�}�H�u�H�U�H�� ��  H�5�k H�={l �; UH��H�� H�}�H�u�H�U�H�� ��  H�5�k H�=Hl � UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��� ��  H�5/k H�=�k � UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�#� ��  H�5�j H�=Xk � UH��H�� H�}�H�u�H�U�H�M�H��� ��  H�5�j H�=!k �� UH��H�� H�}�H�u�H�U�H�M�H�͒ ��  H�5Ij H�=�j � UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�e� ��  H�5�i H�=rj �2 UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��� ��  H�5Yi H�=�i � UH��H��H�}�H�u�H�Α ��  H�5*i H�=�i � UH��H��H�}�H�u�H��� ��  H�5�h H�=�i �\ UH��H�� H�}�H�U�H�E�H�Ѻ   �   H���u  H�E�H�}�t�������E�����UH��H��0H�}�H�u�H�U�H�}� uH�9� ��  H�5}h H�=?i ��  H�E�    H�E�H��H9E�uH�U�H�E�H��  H�E��oH�E�H���L����E�}��u"H�}� tH�U�H�E�H��  H�E��?�    �8H�U�H�E�HЋU��}�
uH�E�H�PH�E�H��  H�E��
H�E��o�����UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���  H������t�������   ��UH��H���}�H�u�H�U��E�H�։�������UH��H��H�}�H�u�H�E�H���Xg��H��H�U�H�E�H�Ѻ   H���  H������t�������   ��UH��H��H�}�H�u�H�U�H�E�H��H��������UH��H��H�}�H�E�H���	  ��UH��H��H�}�H�E�H���������UH��H���C H� H���o	  ]�UH��H���C H� H������]�UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���?  H������t�������E���UH��H���}�H�u�H�U��E�H�։�������UH��H���}�H���C H��E�H�։��s�����UH��H���}��E����������UH��H��@H�}�H���C H� H��tH���C H� H����    H�E�H�E�    H�E�H���e��H�E�H�E�H;E�sQH�E�H+E�H��H�M�H�E�H�4H�M�H�E�H��� ������t������NH�E�H��u������>H�E�HE��H�U�H�E�H�Ѻ   H�5f H���N ������t�������   ��UH��H��H�}�H��� �f  H�5�d H�=�e �O�  UH��H�� H�}��u�H�U�H��� �g  H�5�d H�=]e ��  UH��H���}�H�u�H�^� �h  H�5�d H�=/e ���  UH��H��H�}�H�u�H�6� �i  H�5_d H�= e ���  UH��H��H�}��u�H�� �j  H�51d H�=�d ��  UH��H��H�}�H�� �k  H�5d H�=�d �g�  UH��H�ό �l  H�5�c H�=�d �D�  UH��H���}�H�u�H��� �m  H�5�c H�=Vd ��  UH��H���}�H��� �n  H�5�c H�=,d ���  UH��H���}�H�u�H�i� �o  H�5]c H�=�c ��  UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���*  ��UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���3  ��UH��H��H�}�H�u�H�ދ �z  H�5�b H�=c �+�  UH��H��H�}�H�u�H��� �  H�5�b H�=�b ���  UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�dH�%    H������� �E�H�}� t-H�E�� ��t"H���C H� H�U�H�5�b H�Ǹ    �����E����^�  H��H���C H� H�5�b H�Ǹ    �~������UH��SH���   H�����H�����H�����H����� t
H����� u"dH�%    H�������   H�������^  H�E�    H�E�    H�����H� H��tH�����H� H�E�H�����H� H�E�H�}� u��  �   H���%���H�E�H�E�   H�����H�M�H�E�H��H���R���H������tH��������   H�E�H����`��H�E�H�U�H�E�H�� 
H�E�H�PH�E�H��  H�� ���H�ªC H��H��肀��H�� ���H�5qa H��袀��H��H�E�H�PH�M�H�E�H��H������H�U�H�E�H��H��H���<���H��萀��H�� ���H���K���H�����H�U�H�H�����H�U�H�H�E�H��H���   []�UH��H�� H�}�H�u��U�H�M�H�� ��  H�5�_ H�=` �F�  UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���   ��L�����L�����UH��H��pH�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�E�H���%  H�U�H�M�H�E�H��H����<  H�M�H�U�H�u�H�E�H��H����<  H�E�H���%  H�U�H�E�H��  H�U�H�E�H�H�E���UH��H��   H��X���H��`���H�ªC H��H���C~��H��`���H�5A_ H���c~��H���~��H��`���H���@~�����UH��H��   H��X���H��`���H�ªC H��H����}��H��`���H�5_ H���~��H���*~��H��`���H����}�����UH��H��   H��X���H��`���H�ªC H��H���}��H��`���H�5�^ H���}��H����}��H��`���H���}�����UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�H�U�H�E�H�Ѻ   �   H�������H������t�������E�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H���� ������tHH������H�ªC H��H����{��H������H�5�] H���|��H���?|��H������H����{���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H���� ������tHH��@���H�ªC H��H���{��H��@���H�5�\ H���2{��H���T{��H��@���H���{���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H���* ������tHH������H�ªC H��H����y��H������H�5�[ H����y��H���z��H������H���y���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H���? ������tHH��@���H�ªC H��H����x��H��@���H�5�Z H����x��H���y��H��@���H����x���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H�� H�}��u�H�U�H��� �b  H�5[X H�=�X ��  UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� �����K���������tbH�� ���H��� �����*���������t
H�� �����H�����H�����������������������  H�����H��������H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� �����U�����tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H�ªC H��H���v��H�� ���H�5�W H���4v��H���Vv��H�� ���H���v��H�� ����T  H�� ���� <muSH������H�ªC H��H���u��H������H�5�W H����u��H����u��H������H���u��H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H�W �H�H��V H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H��V �H�H��V H����E�
   H�E�    H�����H��������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���[����E�륀}�0uHH�����H���U���H�����H���2����E׀}�xu!H�����H���.���H�����H�������E׀}�/~2�}�9,H�����H������H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H�������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H������H�E�H��H���E׃�AH�H�H�E�H�����H���K����E��;����}�/~S�}�7MH�����H���<���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H��������E�뭐����H�}� ��  H�U؋M�H�E���H���;����  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���\����E��H�}� �/  H�UȋM�H�E���H�������  H�E�    H�����H�������E��}�0uHH�����H������H�����H��������E��}�xu!H�����H�������H�����H��������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H���S���H�E�H��H���E���AH�H�H�E�H�����H�������E��C���H�}� ��  H�U��M�H�E���H���_�����  H�E�H�E�H�����H��������E��E�    �}� t�E���襶����u�   ��    ��tPH�����H������H�}� t�E�Hc�H�E�H��E��H�����H���j����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H�������E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H�������H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H����L��ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H�������E��}� te�E�;E�}]H�����H�������E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H�������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H���s����E��}�0uHH�����H���o���H�����H���L����E��}�xu!H�����H���H���H�����H���%����E��}�/~2�}�9,H�����H������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H�������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H������H�E�H��H���E���AH�H�H�E�H�����H���m����E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E���UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� ����茱��������tbH�� ���H��� �����k���������t
H�� �����H�����H������������?�����������  H�����H���0�����H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� ����薮����tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H�ªC H��H���Uh��H�� ���H�5>J H���uh��H���h��H�� ���H���Rh��H�� ����T  H�� ���� <muSH������H�ªC H��H����g��H������H�5�I H���h��H���6h��H������H����g��H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H�}P �H�H�qP H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H�]P �H�H�QP H����E�
   H�E�    H�����H�������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H�������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���6����E�륀}�0uHH�����H���~���H�����H�������E׀}�xu!H�����H���W���H�����H��������E׀}�/~2�}�9,H�����H���*���H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H�������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H������H�E�H��H���E׃�AH�H�H�E�H�����H���&����E��;����}�/~S�}�7MH�����H���e���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H��������E�뭐����H�}� ��  H�U؋M�H�E���H���|����  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H�������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���7����E��H�}� �/  H�UȋM�H�E���H��������  H�E�    H�����H��������E��}�0uHH�����H���@���H�����H��������E��}�xu!H�����H������H�����H�������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H���|���H�E�H��H���E���AH�H�H�E�H�����H��������E��C���H�}� ��  H�U��M�H�E���H��������  H�E�H�E�H�����H�������E��E�    �}� t�E���������u�   ��    ��tPH�����H�������H�}� t�E�Hc�H�E�H��E��H�����H���E����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H��������E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H������H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H���?��ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H��������E��}� te�E�;E�}]H�����H���;����E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H�������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H���N����E��}�0uHH�����H������H�����H���'����E��}�xu!H�����H���q���H�����H��� ����E��}�/~2�}�9,H�����H���D���H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H�������H�E�H��H���E���AH�H�H�E�H�����H���H����E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H��H�}����E�H�E�H�H�E�H�Ѻ   �   H���Z���H�E�H�@H�PH�E�H�P���UH��SH��H�}�H�u�H�E�H�H�E�H���I<��H��H�E�H�ٺ   H������H�E�H���&<��H��H�E�H�@H�H�E�H�P�H��[]ÐUH��H�� H�}�H�u�H�U�H�E�H�H�u�H�E�H�Ѻ   H������H�E�H�PH�E�H�H�E�H�P��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H�}����E�H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]�UH��H�}�H�u�H�E�    H�U�H�E�H�� ��t>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�밐]ÐUH��H�}�H�u�H�U�H�E�    H�E�H;E�s>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�븐]ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�PH�E�H�@    �]�UH��H�}����E�H�E�H�PH�E�H�@H9�sH�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]ÐUH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���e���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E�H�     H�E�H�@    H�E�H�@    �]�UH��H��0H�}�H�E�H�PH�E�H�@H9���   H�E�   H�E�H�@H�H�E�H�U�H�E�H��H���c��H� H�E�H�E�H���tH��H�E�H�E�H��uH��a ��   H�5�8 H�=�8 ��  H�E�H�PH�E�H�H�E�H��H���7��H�E�H� H���G��H�U�H�E�H�H�E�H�U�H�PH�E�H�PH�E�H�@H9�rH�sa ��   H�5,8 H�=X8 ��  ��ÐUH��H��H�}����E�H�E�H�������H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P���UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���k���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E��@]�UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���G  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=�9 ���H��x���� <%uH�E��%   H���  H��x����  H�E�H����J��H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�9 �
���H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�9 �G
���u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�9 ��	���*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�9 �	�������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�9 �f	��������E���tH��    H��uH�=�9 �>	���E���tH��    H��uH�=1: �	��H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=[: ����H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�= : �3��돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=: ����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=: ���H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H���K����   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�9 ����H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�9 ����H�U�H�E�H��H���N  H�E�H�U�H��H��H���  H�E�H���J���E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=y9 ���H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�9 �����N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�9 �w��H�U�H�E�H��H����E��H��x���� ���M�H�U�H�E�H���h  H�E�H���JF��H��x���H�E�H���6F���g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���K  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=�2 ���H��x���� <%uH�E��%   H���  H��x����  H�E�H����C��H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�2 ����H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�2 �Q���u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�2 ����*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�2 ��������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�2 �p��������E���tH��    H��uH�=�2 �H���E���tH��    H��uH�=;3 �&��H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=e3 ����H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=
3 �=��돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=3 �� ��H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=3 � ��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H����  H�E�H�U�H��H��H���   H�E�H���D����   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�2 � ��H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�2 �����H�U�H�E�H��H���X  H�E�H�U�H��H��H���  H�E�H���#C���E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=�2 ����H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�2 ������N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�2 ����H�U�H�E�H��H����>��H��x���� ���M�H�U�H�E�H���  H�E�H���T?��H��x���H�E�H���@?���g������UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���]  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=�+ �����H��x���� <%uH�E��%   H���0  H��x����  H�E�H����<��H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�+ �s����H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�+ �/����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�+ ������*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�+ ���������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�+ �N���������E���tH��    H��uH�=�+ �&����E���tH��    H��uH�=, ����H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=C, �����H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�+ ����돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=�+ �����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=�+ ����H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���	  H�E�H�U�H��H��H����	  H�E�H����<����   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�+ �����H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�+ �u����H�U�H�E�H��H���6	  H�E�H�U�H��H��H����  H�E�H���<���E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=a+ �����H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=l+ �����N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=l+ �_���H�U�H�E�H��H����7��H��x���� ���M�H�U�H�E�H���  H�E�H���28��H��x���H�E�H���8���g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=�$ �����H��x���� <%uH�E��%   H���n  H��x����  H�E�H����5��H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�$ �}����H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�$ �9����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�$ ������*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�$ ���������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�$ �X���������E���tH��    H��uH�=�$ �0����E���tH��    H��uH�=#% ����H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=M% ����H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�$ �%��돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=�$ ����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=% ���H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H����5����   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�$ ����H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�$ ����H�U�H�E�H��H���@  H�E�H�U�H��H��H����  H�E�H���5���E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=k$ ����H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=v$ ����N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=v$ �i��H�U�H�E�H��H����0��H��x���� ���M�H�U�H�E�H����  H�E�H���<1��H��x���H�E�H���(1���g������UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���������ÐUH��H��H�}����E�H�E�H� �U��H��������ÐUH��SH��H�}�H�u�H�E�H���E��H�E��@H�E�H���c�����H�E�H�ƿ   �m/����H��[]�UH��H��H�}�H�u�H�U�H�E�H��H����  H�E��ÐUH��SH��H�}�H�u�H�E�H���E��H�E��@H�E�H���  �H�E�H�ƿ   ��.����H��[]�UH��SH��(  H��������H��������������������������E��3�	  ��H��    H��B �H�H��B H���H������H�XH������H������H��H����.��������H������H� ������H������I��H���  H������H���5/���  H������H�XH������H�����H��H���x.��������H������H� ������H�����I��H���7  H�����H����.���  H������H�XH������H��0���H��H���.��������H������H� ������H��0���I��H���#  H��0���H���s.���L  H�������@��tH�&@ �*   H�5B H�=U& 裰  H�������@��tH��? �+   H�5 H�=8& �u�  H�������@��tH��? �,   H�5� H�=& �G�  H�������@��tH��? �-   H�5� H�=& ��  ������ tH�u? �.   H�5� H�=�% ��  H������H��H���F�����tH�?? �/   H�5[ H�=�% 輯  H������H�dH�%    H������� ��蘏  H��H�������  ������ tH��> �3   H�5  H�=i% �a�  H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ªC H��H���k6��H��P���H�5)% H���6��H����������H����!  H�5.% H���h6��H���6��H��P���H���E6��H�> �;   H�5$ H�=�$ 腮  �H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���:�����ÐUH��H��H�}����E�H�E�H� �U��H���j�����ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H��? �H�H��? H���H������H�XH������H������H��H���*��������H������H� ������H������I��H���   H������H���+���  H������H�XH������H�����H��H���D*��������H������H� ������H�����I��H����+  H�����H���*���  H������H�XH������H��0���H��H����)��������H������H� ������H��0���I��H���#3  H��0���H���?*���L  H�������@��tH�
< �*   H�5 H�=!" �o�  H�������@��tH��; �+   H�5� H�=" �A�  H�������@��tH��; �,   H�5� H�=�! ��  H�������@��tH��; �-   H�5� H�=�! ��  ������ tH�Y; �.   H�5] H�=�! 辫  H������H��H��������tH�#; �/   H�5' H�=�! 舫  H������H�dH�%    H������� ���d�  H��H��������  ������ tH��: �3   H�5� H�=5! �-�  H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ªC H��H���72��H��P���H�5�  H���W2��H����������H���  H�5�  H���42��H���V2��H��P���H���2��H��9 �;   H�5� H�=�  �Q�  �H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���������ÐUH��H��H�}����E�H�E�H� �U��H���������ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H�(< �H�H�< H���H������H�XH������H������H��H���q&��������H������H� ������H������I��H���0  H������H����&���  H������H�XH������H�����H��H���&��������H������H� ������H�����I��H���=;  H�����H���l&���  H������H�XH������H��0���H��H���%��������H������H� ������H��0���I��H���B  H��0���H���&���L  H�������@��tH��7 �*   H�5� H�=� �;�  H�������@��tH��7 �+   H�5� H�=� ��  H�������@��tH��7 �,   H�5~ H�=� �ߧ  H�������@��tH�]7 �-   H�5Q H�=� 貧  ������ tH�57 �.   H�5) H�=� 芧  H������H��H���������tH��6 �/   H�5� H�=� �T�  H������H�dH�%    H������� ���0�  H��H���m����  ������ tH��6 �3   H�5� H�= ���  H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ªC H��H���.��H��P���H�5� H���#.��H����������H���m  H�5� H��� .��H���".��H��P���H����-��H��5 �;   H�5� H�=� ��  �H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���������ÐUH��H��H�}����E�H�E�H� �U��H���0�����ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H��8 �H�H��8 H���H������H�XH������H������H��H���="��������H������H� ������H������I��H���?  H������H���"���  H������H�XH������H�����H��H����!��������H������H� ������H�����I��H���J  H�����H���8"���  H������H�XH������H��0���H��H���{!��������H������H� ������H��0���I��H����Q  H��0���H����!���L  H�������@��tH��4 �*   H�5� H�=� ��  H�������@��tH��4 �+   H�5x H�=� �٣  H�������@��tH��4 �,   H�5J H�=� 諣  H�������@��tH�Y4 �-   H�5 H�=i �~�  ������ tH�14 �.   H�5�
 H�=^ �V�  H������H��H��������tH��3 �/   H�5�
 H�=T � �  H������H�dH�%    H������� �����  H��H�������  ������ tH��3 �3   H�5d
 H�=� �Ţ  H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H�ªC H��H����)��H��P���H�5� H����)��H����������H���9  H�5� H����)��H����)��H��P���H���)��H��2 �;   H�5�	 H�=` ��  �H��(  []�UH��SH��(H�}�H�u�H�E��@��t$H�E��@��tH�U�H�E�H��H���O  �   H�E��@��tAH�E��@����t2H�E�H��������E�H�E�H���������H�E�H�ƿ   ������KH�E��@����t<H�E��@��t0H�E�H�������E�H�E�H��������H�E�H�ƿ   ����H�E�H�PH�E�H��H��H���_O  �H��([]�UH��H�}�H�E�]ÐUH��H��H�}�H�E��@����tH��    H��uH�=� �)ݾ�H�E���UH��H�ĀH�}���H�U��M�L�E��E��E���pt��s�8  ��c�  �  H�E��@��tH��    H��uH�=~ ��ܾ�H�E��@��tH��    H��uH�=� �ܾ�H�E��@��tH��    H��uH�=� �uܾ�H�E��@��tH��    H��uH�=- �Pܾ�H�E�H�5~ H�������H�E����/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���N  �7  H�E��@��tH��    H��uH�= �۾�H�E��@��tH��    H��uH�=> �۾�H�E��@��tH��    H��uH�=x �s۾�H�E��@��tH��    H��uH�=� �N۾��}� tH��    H��uH�=� �.۾�H�E�H��H���������tH��    H��uH�== � ۾�H�E����/wH�P���Hʋ����H�PH�JH�H���H�E���H��� ����  H�E��@��tH��    H��uH�=4 �ھ�H�E��@��tH��    H��uH�=n �qھ��}� ��  H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�} H�E�H�U�H�E�H��H���Px��H�E�H�������E�H�E�H��H���������tH�E�H��H������� 9E�~�   ��    ��tH�E�H��H���X���� �E�H�E��@��tw�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H�������E�뽋E�E�H�E��@9E���  H�E��    H�������E��ًE�E�H�E��@9E�}H�E��    H���i����E����E�    �E�;E��C  �E�Hc�H�E�H�� ���+  �E�Hc�H�E�H�� ��H�E���H�������E�뵃}�tH��    H��uH�=� �ؾ�H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�# H�E�H�U�H�E�H��H����J  H�E�H���K  �E�H�E�H��H���������tH�E�H��H������� 9E�~�   ��    ��tH�E�H��H������� �E�H�E��@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H��������E�뱋EԉE�H�E��@9E���   H�E��    H�������E��ًEԉE�H�E��@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���/����E��H��    H��uH�=� �־�����ÐUH��SH��H�}�H�u�H�E�H� H��H���b�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��� �����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���H  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H���8���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���(�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���H  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H���a���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���P�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���]F  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���������t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���x�����tH�E�H� H��H���'������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����F  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���O������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���D  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���)�����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���w������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���9E  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H��( �H�H��( H���H�E��@��tH��    H��uH�=� �%Ѿ�H�E��@��tH��    H��uH�=� ��о��}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=H �+о�H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H���������t$H�E�H��H���v���� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���g�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���BB  �W  H�E��@��tH��    H��uH�=� �Ͼ�H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���P����}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=w �ξ�H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=� �$ξ�H�E��@��tH��    H��uH�=� ��;�H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=� �;�H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=� � ;�H�E��@��tH��    H��uH�=� ��̾�H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=� �<̾�H�E��@��tH��    H��uH�=� �̾�H�E�H��H��������tH��    H��uH�=� ��˾��}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���g?  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���==  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����<  �   �}� tH��    H��uH�=� �rʾ�H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���=  �H��    H��uH�=� ��ɾ����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5� H���F����H��    H��uH�=� �ɾ���ÐUH��H��H�}����E�H�U�H�E�H��H���=  H�E���UH��H�ĀH�}���H�U��M�L�E��E��E���pt��s�8  ��c�  �  H�E��@��tH��    H��uH�=� ��Ⱦ�H�E��@��tH��    H��uH�=� ��Ⱦ�H�E��@��tH��    H��uH�=% �Ⱦ�H�E��@��tH��    H��uH�=` �Ⱦ�H�E�H�5� H��耹��H�E����/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���<  �7  H�E��@��tH��    H��uH�=7 ��Ǿ�H�E��@��tH��    H��uH�=q ��Ǿ�H�E��@��tH��    H��uH�=� �Ǿ�H�E��@��tH��    H��uH�=� �Ǿ��}� tH��    H��uH�=. �aǾ�H�E�H��H���-�����tH��    H��uH�=p �3Ǿ�H�E����/wH�P���Hʋ����H�PH�JH�H���H�E���H��賷���  H�E��@��tH��    H��uH�=g ��ƾ�H�E��@��tH��    H��uH�=� �ƾ��}� ��  H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�� H�E�H�U�H�E�H��H���d��H�E�H���o���E�H�E�H��H��� �����tH�E�H��H������� 9E�~�   ��    ��tH�E�H��H������� �E�H�E��@��tw�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���R����E�뽋E�E�H�E��@9E���  H�E��    H���%����E��ًE�E�H�E��@9E�}H�E��    H��������E����E�    �E�;E��C  �E�Hc�H�E�H�� ���+  �E�Hc�H�E�H�� ��H�E���H��誵���E�뵃}�tH��    H��uH�=+ ��ľ�H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�V H�E�H�U�H�E�H��H����6  H�E�H���I7  �E�H�E�H��H���,�����tH�E�H��H�������� 9E�~�   ��    ��tH�E�H��H������� �E�H�E��@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���n����E�뱋EԉE�H�E��@9E���   H�E��    H���A����E��ًEԉE�H�E��@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���³���E��H��    H��uH�=� ��¾������UH��SH��H�}�H�u�H�E�H� H��H��薶����t'H�E�H� H��H���E���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���4�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���6  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��轵����t&H�E�H� H��H���l���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���\�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���6  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��脴����tH�E�H� H��H���3������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H����4  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��謳����tH�E�H� H��H���[������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���5  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���6�����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���Բ����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���73  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���]�����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���V3  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�� �H�H�� H���H�E��@��tH��    H��uH�=��  �Y���H�E��@��tH��    H��uH�=��  �3����}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=|�  �_���H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H���������t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H��蛯����tH�E�H��H���M������   H�E��PH�u�H�E�A��A�ȉѺ
   H���_0  �W  H�E��@��tH��    H��uH�=��  �S���H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H�������}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  辺��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=��  �X���H�E��@��tH��    H��uH�=��  �2���H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  躹��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=��  �T���H�E��@��tH��    H��uH�=�  �.���H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=��  �p���H�E��@��tH��    H��uH�=��  �J���H�E�H��H��������tH��    H��uH�=)�  �����}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���-  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����+  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���U+  �   �}� tH��    H��uH�=�  覶��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H����+  �H��    H��uH�=�  �$������H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5�  H�������H��    H��uH�=�  踵�����UH��H�ĀH�}���H�U��M�L�E��E��E���pt��s�8  ��c�  �  H�E��@��tH��    H��uH�=�  �S���H�E��@��tH��    H��uH�=J�  �-���H�E��@��tH��    H��uH�=��  ����H�E��@��tH��    H��uH�=��  �ⴾ�H�E�H�5�  H��苤��H�E����/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���*  �7  H�E��@��tH��    H��uH�=��  �Q���H�E��@��tH��    H��uH�=��  �+���H�E��@��tH��    H��uH�=
�  ����H�E��@��tH��    H��uH�=E�  �೾��}� tH��    H��uH�=��  �����H�E�H��H��茧����tH��    H��uH�=��  蒳��H�E����/wH�P���Hʋ����H�PH�JH�H���H�E���H���Ԣ���  H�E��@��tH��    H��uH�=��  �)���H�E��@��tH��    H��uH�= �  �����}� ��  H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��  H�E�H�U�H�E�H��H����P��H�E�H���t[���E�H�E�H��H���_�����tH�E�H��H������� 9E�~�   ��    ��tH�E�H��H�������� �E�H�E��@��tw�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���s����E�뽋E�E�H�E��@9E���  H�E��    H���F����E��ًE�E�H�E��@9E�}H�E��    H�������E����E�    �E�;E��C  �E�Hc�H�E�H�� ���+  �E�Hc�H�E�H�� ��H�E���H���ˠ���E�뵃}�tH��    H��uH�=��  �%���H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH���  H�E�H�U�H�E�H��H���Z#  H�E�H���#  �E�H�E�H��H��苤����tH�E�H��H���=���� 9E�~�   ��    ��tH�E�H��H������� �E�H�E��@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H��菟���E�뱋EԉE�H�E��@9E���   H�E��    H���b����E��ًEԉE�H�E��@9E�}H�E��    H���9����E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H�������E��H��    H��uH�=8�  �C�������ÐUH��SH��H�}�H�u�H�E�H� H��H���������t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��蒢����tH�E�H� H��H���A������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���$  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��躡����tH�E�H� H��H���i������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���$  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���D�����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H����"  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���k�����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���
�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���#  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��蔟����t'H�E�H� H��H���C���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���2�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���7!  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��軞����t&H�E�H� H��H���j���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���Z�����tH�E�H� H��H���	������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���V!  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�� �H�H�� H���H�E��@��tH��    H��uH�=�  跩��H�E��@��tH��    H��uH�=N�  葩���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=��  轨��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H���V�����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���������tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���_  �W  H�E��@��tH��    H��uH�=>�  豧��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H�������}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=	�  ����H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=�  趦��H�E��@��tH��    H��uH�=M�  萦��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=5�  ����H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=?�  貥��H�E��@��tH��    H��uH�=y�  茥��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=�  �Τ��H�E��@��tH��    H��uH�=U�  訤��H�E�H��H���t�����tH��    H��uH�=��  �z����}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���U  �   �}� tH��    H��uH�=q�  ����H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H����  �H��    H��uH�=_�  肢�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5y�  H�������H��    H��uH�=c�  �������UH��H�ĀH�}���H�U��M�L�E��E��E���pt��s�8  ��c�  �  H�E��@��tH��    H��uH�=n�  象��H�E��@��tH��    H��uH�=��  苡��H�E��@��tH��    H��uH�=��  �e���H�E��@��tH��    H��uH�=�  �@���H�E�H�5n�  H���e���H�E����/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���  �7  H�E��@��tH��    H��uH�=��  诠��H�E��@��tH��    H��uH�=.�  艠��H�E��@��tH��    H��uH�=h�  �c���H�E��@��tH��    H��uH�=��  �>����}� tH��    H��uH�=��  ����H�E�H��H��������tH��    H��uH�=-�  ���H�E����/wH�P���Hʋ����H�PH�JH�H���H�E���H��螒���  H�E��@��tH��    H��uH�=$�  臟��H�E��@��tH��    H��uH�=^�  �a����}� ��  H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�m�  H�E�H�U�H�E�H��H���@=��H�E�H����G���E�H�E�H��H��轒����tH�E�H��H���o���� 9E�~�   ��    ��tH�E�H��H���H���� �E�H�E��@��tw�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���=����E�뽋E�E�H�E��@9E���  H�E��    H�������E��ًE�E�H�E��@9E�}H�E��    H�������E����E�    �E�;E��C  �E�Hc�H�E�H�� ���+  �E�Hc�H�E�H�� ��H�E���H��蕐���E�뵃}�tH��    H��uH�=��  胝��H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��  H�E�H�U�H�E�H��H���  H�E�H���  �E�H�E�H��H��������tH�E�H��H��蛿��� 9E�~�   ��    ��tH�E�H��H���t���� �E�H�E��@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���Y����E�뱋EԉE�H�E��@9E���   H�E��    H���,����E��ًEԉE�H�E��@9E�}H�E��    H�������E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H��譎���E��H��    H��uH�=��  衛������ÐUH��SH��H�}�H�u�H�E�H� H��H���R�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H��蟽�����   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���y�����t&H�E�H� H��H���(���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���Ǽ�����   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��袍����t'H�E�H� H��H���Q���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���@�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H����  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���Ɍ����t&H�E�H� H��H���x���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���h�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H��衺��� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��萋����tH�E�H� H��H���?������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���7  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H���ȹ��� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��踊����tH�E�H� H��H���g������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���V  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�x�  �H�H�l�  H���H�E��@��tH��    H��uH�=r�  ����H�E��@��tH��    H��uH�=��  ���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=8�  ����H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��贈����t$H�E�H��H���f���� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���W�����tH�E�H��H���	������   H�E��PH�u�H�E�A��A�ȉѺ
   H���_  �W  H�E��@��tH��    H��uH�=��  ����H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���Ά���}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=g�  �z���H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=q�  ����H�E��@��tH��    H��uH�=��  ��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=��  �v���H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=��  ����H�E��@��tH��    H��uH�=��  �ꑾ�H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=y�  �,���H�E��@��tH��    H��uH�=��  ����H�E�H��H���҄����tH��    H��uH�=��  �ؐ���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���	  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���U  �   �}� tH��    H��uH�=��  �b���H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H����  �H��    H��uH�=��  ��������H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5��  H���ȁ���H��    H��uH�=��  �t������UH��H�� H�}�H�u�H�E�H���G����E�H�E�H���8�����H�E�H�E�H���$�����H�E�����UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�E�H��������E�H�E�H���������H�E�H�E�H��������H�E�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����  H����ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�@H��    H�E�HЋ ��tH�E�H�@H�PH�E�H�P�͐]ÐUH��H�}�H�E�H�@]�UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���#
  H�����UH��H��0H�}�H�u�H�E�H�������H�E�� ��H�U�H�M�H�Ή��  H�E�H���������UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���w  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���l  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���u  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���a  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H����  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���j  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�'�  H�E��E�    �E���~H��    H��uH�=�  �8����E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �ƅ���E��P�U�H��D�-H�U�H�E�H��H������ 9E�����tE�E�    H�U�H�E�H��H������ �U�)�9E�����t�U�H�E���H���s���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���s���E��ڋE����E�}� x!�E�H��D���H�E���H���Os���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=m�  萄���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=K�  �����E��P�U�H��D�-H�U�H�E�H��H������ 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���r���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����q���E��ڋE����E�}� x!�E�H��D���H�E���H���q���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  �邾��M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=��  �����E��P�U�H��D�-H�U�H�E�H��H���w��� 9E�����tE�E�    H�U�H�E�H��H���Q��� �U�)�9E�����t�U�H�E���H���op���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���8p���E��ڋE����E�}� x!�E�H��D���H�E���H���p���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�8�  H�E��E�    �E���~H��    H��uH�=&�  �I����E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  �׀���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H������ �U�)�9E�����t�U�H�E���H����n���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���n���E��ڋE����E�}� x!�E�H��D���H�E���H���`n���m��ِ��UH��H��@�}�H�u�H�U�H�U�H�E�H��H���Q���H�U�H�M��E�H�Ή���  H�E�H����������UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�F�  H�E��E�    �E���~H��    H��uH�=4�  �W���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�  ��~���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H������ �U�)�9E�����t�U�H�E���H���5o���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����n���E��ڋE����E�}� x!�E�H��D���H�E���H����n���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  �}���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=j�  �=}���E��P�U�H��D�-H�U�H�E�H��H���5��� 9E�����tE�E�    H�U�H�E�H��H������ �U�)�9E�����t�U�H�E���H���m���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���Vm���E��ڋE����E�}� x!�E�H��D���H�E���H���&m���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  �|���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=��  �{���E��P�U�H��D�-H�U�H�E�H��H���
��� 9E�����tE�E�    H�U�H�E�H��H���p
��� �U�)�9E�����t�U�H�E���H����k���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���k���E��ڋE����E�}� x!�E�H��D���H�E���H���k���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�W�  H�E��E�    �E���~H��    H��uH�=E�  �hz���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=#�  ��y���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���Fj���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���j���E��ڋE����E�}� x!�E�H��D���H�E���H����i���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  ��x���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�={�  �Nx���E��P�U�H��D�-H�U�H�E�H��H���F��� 9E�����tE�E�    H�U�H�E�H��H��� ��� �U�)�9E�����t�U�H�E���H���`g���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���)g���E��ڋE����E�}� x!�E�H��D���H�E���H����f���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=��  �w���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �v���E��P�U�H��D�-H�U�H�E�H��H������ 9E�����tE�E�    H�U�H�E�H��H���x��� �U�)�9E�����t�U�H�E���H���e���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���e���E��ڋE����E�}� x!�E�H��D���H�E���H���Qe���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�`�  H�E��E�    �E���~H��    H��uH�=N�  �qu���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=4�  �u���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���d���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����c���E��ڋE����E�}� x!�E�H��D���H�E���H���c���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=��  ��s���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �_s���E��P�U�H��D�-H�U�H�E�H��H���W��� 9E�����tE�E�    H�U�H�E�H��H���1��� �U�)�9E�����t�U�H�E���H���qb���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���:b���E��ڋE����E�}� x!�E�H��D���H�E���H���
b���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=�  �)r���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  �q���E��P�U�H��D�-H�U�H�E�H��H��� ��� 9E�����tE�E�    H�U�H�E�H��H��� ��� �U�)�9E�����t�U�H�E���H���5d���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����c���E��ڋE����E�}� x!�E�H��D���H�E���H����c���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�p�  H�E��E�    �E���~H��    H��uH�=^�  �p���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=<�  �p���E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H�������� �U�)�9E�����t�U�H�E���H���b���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���Vb���E��ڋE����E�}� x!�E�H��D���H�E���H���&b���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�ɾ  H�E��E�    �E���~H��    H��uH�=��  ��n���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=��  �pn���E��P�U�H��D�-H�U�H�E�H��H���h���� 9E�����tE�E�    H�U�H�E�H��H���B���� �U�)�9E�����t�U�H�E���H����`���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���`���E��ڋE����E�}� x!�E�H��D���H�E���H���`���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�)�  H�E��E�    �E���~H��    H��uH�=�  �:m���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=��  ��l���E��P�U�H��D�-H�U�H�E�H��H�������� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���F_���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���_���E��ڋE����E�}� x!�E�H��D���H�E���H����^���m��ِ��UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=s�  �vk���u�H�E�A�    A�   �    �
   H���   ���UH��H��0H�}�u�U��M�D�E�D�ȈEԃ}� y=�E��؉E��M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ   H���Z��H���3�M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�N�  H�E��E�    �E���~H��    H��uH�=<�  �_j���E���}���Hc�H�E�H���E��H�M�H��T��E���}��E��}� t맀}� t2�E���~H��    H��uH�=-�  � j���E��P�U�H��D�-H�U�H�E�H��H�������� 9E�����tE�E�    H�U�H�E�H��H�������� �U�)�9E�����t�U�H�E���H��������E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H�������E��ڋE����E�}� x!�E�H��D���H�E���H���o����m��ِ��UH��H�}�H�u�H�E�H�E�H�E�H�E�H�E�� ��tH�E�H�PH�U��H�E�H�HH�M����H�E��  H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E�H;E�sH�E�H�PH�U��  H�E���H�E�]�UH��H��H�}�H�u�H�E�H���?���H��H�E�H�H�E�H��H�������H�E���UH��H��@H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H������HE�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E��  H�E���UH��H�}�H�u�H�U�H�E�    H�E�H;E�sIH�U�H�E�H�� �E�H�U�H�E�H�� �E��E�:E�s�������E�:E�v�   �H�E�뭸    ]�UH��H�}�H�u�H�E�    H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H��H�}�H�u�H�U�H�E�H��H���k�����UH��H�}�H�u�H�U�H�E�    H�E�H;E�r�    �\H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H�� H�}�H�u�H�U�H�(�  �g   H�5��  H�=��  �=)  UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s)H�U�H�E�H�� �U�8�uH�U�H�E�H��H�E��͸    ]�UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E��ă}� uH�U�H�E�H���    ]�UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H���N���H��t�   ��    ��tH�E��H�E����UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t=H�U�H�E�H�� ��H�E���H�������H������tH�U�H�E�H��H�E�뱸    ��UH��H�� H�}�u�H�E�H���#���H�E�H�E�    H�E�H;E�w8H�E�H+E�H��H�E�H�� ��9E�uH�E�H+E�H��H�E�H��H�E�뾸    ��UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H������H��u�   ��    ��tH�E��H�E����UH��H�}�H�u�H�E�    H�U�H�E�H�� ����   �E�H�E�    H�U�H�E�H�� ��tGH�U�H�E�H�� ��t-H�U�H�E�H�H�E�H��H�M�H�E�H�� 8�t�E� ��H�E�맀}� tH�U�H�E�H��H�E��h����    ]�UH��H��H�}�H�u�H�Կ  ��   H�5(�  H�=J�  ��%  UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E���H�U�H�E�H�]�UH��H��H�}�H�u�H�P�  ��   H�5��  H�=ֻ  �V%  UH��H��H�}�H�u�H�(�  ��   H�5n�  H�=��  �'%  UH��H��H�}�H�u�H��  ��   H�5?�  H�=x�  ��$  UH��H�� H�}�H�u��U�H�پ  ��   H�5�  H�=F�  ��$  UH��H�� H�}�H�u��U�H���  ��   H�5ۺ  H�=�  �$  UH��H�� H�}�H�u��U�H���  ��   H�5��  H�=�  �b$  UH��H�� H�}�H�u��U�H�[�  ��   H�5w�  H�=��  �0$  UH��H��H�}�H�u�H�5�  ��   H�5H�  H�=��  �$  UH��H�� H�}�H�u�H�U�H�	�  ��   H�5�  H�=N�  ��#  UH��H�� H�}�H�u�H�U�H�޽  ��   H�5�  H�=�  �#  UH��H�� H�}�H�u�H�U�H���  ��   H�5��  H�=�  �h#  UH��H��H�}�H�u�H���  ��   H�5��  H�=��  �9#  UH��H�� H�}�H�u�H�U�H�a�  ��   H�5M�  H�=��  �#  UH��H��H�}�H�u�H�:�  ��   H�5�  H�=W�  ��"  UH��H��H�}�H�u�H��  ��   H�5�  H�=(�  �"  UH��H�� H�}�H�u�H�U�H��  ��   H�5��  H�=��  �u"  UH��H�� H�}�H�u�H�U�H���  ��   H�5��  H�=¸  �B"  UH��H�� H�}�H�u�H�U�H���  ��   H�5V�  H�=��  �"  UH��H��H�}��u�H�l�  ��   H�5(�  H�=a�  ��!  UH��H��H�}�H�u�H�E�  ��   H�5��  H�=2�  �!  UH��H��H�}�H�u�H��  ��   H�5ʷ  H�=�  �!  UH��H��H�}��u�H���  ��   H�5��  H�=շ  �U!  UH��H��H�}�H�u�H�ѻ  ��   H�5m�  H�=��  �&!  UH��H��H�}�H�u�H���  ��   H�5>�  H�=w�  ��   UH��H�� H�}�H�u�H�U�H�}�  ��   H�5�  H�=D�  ��   UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s6H�E�H��    H�E�HЋ 9E�uH�E�H��    H�E�H��H�E����    ]�UH��H��H�}�H��  ��   H�5z�  H�=��  �3   UH��H�� H�}��u�H�U�H�̺  ��   H�5H�  H�=��  �   UH��}�E�-�  ��C�  ��H��    H���  �H�H���  H���H�c�  H�E���   H�r�  H�E���   H�z�  H�E���   H���  H�E���   H���  H�E��   H���  H�E��   H���  H�E��   H���  H�E��   H���  H�E��sH�ζ  H�E��fH��  H�E��YH���  H�E��LH��  H�E��?H�2�  H�E��2H�F�  H�E��%H�M�  H�E��H�[�  H�E��H�p�  H�E�H�E�]�UH��H��0�}�H�u�H�U؋E������H�E�H�U�H�M�H�E�H��H���E���H�E�H������H9E�����t�   ��    ��UH��H�� H�}�H�u�H�U�H�U�H�M�H�E�H��H���Ԅ��H��H�E�H���UH��H�� H�}�H�u�H�E�H��诅��H�E�H�E�H�PH�M�H�E�H��H��荄��H�U�H�E�H���UH����s ������t5H�=�s ��&  ������t �  H��H�=�s ��   H�=�s ��&  H�=�s �  ]�UH��H��@H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H�E��x���H��H�E�H��H����   �    ��UH��H�� �R���H�E�H�E�H���@  H�E�H�}� t6H�E�H�P�H�E�H��H���0  H�E�H�E�H� H�U�H�RH����H�m��Ð��UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H���  H�E�H�������H��H�E�H�ƿ    �2���H��H���  �H��[]�UH��H�}�H�E�]�UH��H�� H�}�H�u�H�E�H�@H�PH�E�H��H���  H�E�H�HH�E�H�PH��H�H�H��H�H�ƿ   蹘��H�u�H�H�NH�H�HH�VH�PH�E�H�E�H�@H�PH�E�H�PH�E���UH��H�}�H�E�H�@]�UH��H�}�H�u�H�E�H�HH�U�H��H�H�H��H�]�UH��H�}�H�E�H�     H�@    H�@    H�@    �]�UH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�@    H�E�H�@    �]�UH��H��0H�}�H�u�H�E�H�@H9E���   H�E�H�H�E�H�E�H�H�U�H��H�H�H��H��H��脦��H�E�H�E�    H�E�H�@H9E�sVH�U�H��H�H�H��H��H�E�H�H�ƿ   �G���H��H�E�H�HH�U�H��H�H�H��H�H���[   H�E��H�E�    H�E�H�@H9E�sH�E���H�E�H� H�U�H�RH��H���u���H�E�H�U�H�PH�E�H�U�H�P����UH��H�}�H�u�H�M�H�u�H�H�VH�H�QH�FH�AH�E�]�UH��H���}�A�    A�    �    �    �    �   �G~�����UH��H��H�}�H�u�H�E�%�  H��tH���  �   H�5��  H�=��  �  H�E�H�U�H��H��A�    A�    �    H�¿   ��}��H�E�H� H��u�������    ��UH��H�}�H�u�    ]�UH��H��ޭޭ����    ��UH���Co ������t-H�=3o ��!  ������tH�=o �!  H�=o �'"  ��p ������t<H�=�p ��!  ������t'H�=�n �  H��H�=�n �  H�=�p ��!  H�=�n �U  ]ÐUH��H�� H�}�H�u�H�U�H�E�H��H������������tH��  �   H�5��  H�=��  �4  H�E��ÐUH��H�� H�}�H�u�H�U�H�E�H�U�H��H�������������tH���  �    H�55�  H�=��  ��  ���UH��H�}�H�E��     �]ÐUH��H��H�}�H�E�H���   H�E�H�ƿ   �6������UH��H�}�H�E�]�UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H���S   H�E�H�������H��H�E�H�ƿ�  �ړ��H��H���N   �H��[]�UH��H�}�H�E�]�UH��H�}�H�E��  �]�UH��H�}�H�E�H�Ƹ    �9   H��H���H��]ÐUH��ATSH��H�}�H�u�H�E�H�U�H�H�E�H��H�������H�E�H��H���>   H�E�H�@     H�E�H��(�   I��H��xL���9   I�� H����H��[A\]ÐUH��H��H�}�H�E�H���N   H�}�:   ���UH��H��H�}�H�E�H���T���H�E�H�@    H�E�H��H���$   ���UH��H�}�]ÐUH��H�}�H�E�H�     �]�UH��H��H�}�H�E�H���   H�}�������UH��H�}�H�E�H�     �]�UH��H�}�H��x C H�PH�E�H��]ÐUH��H��H�}�H�E�H�������H�E��   H���	t����UH����m ������tJH�=|m �O  ������t5H�=Wm ��  H�=[m �x  H�S H�58m H��Z�A H������H�"m ]�UH��H�}��u�H�U�U�H�E��    ]�UH��H�m ]�UH��H�}����E�ЈE�H��x C H�PH�E�H�H�E��U�PH�E��U��P	�]ÐUH��H�}�H�E��     H�E��@    �]�UH��H�}�H�E�� ]�UH��H�}�H�E��@]ÐUH��H�� H�}�H�u�H�E�H� � �E�H�E� ����   �E���x�U�H�E�P�-  �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    �   �E�%�   =�   t/�E�%�   =�   tH���  �'   H�5I�  H�=r�  �J  �   �q�E�%�   =�   tH�w�  �,   H�5�  H�=��  �  H�E�@�����E���?	�H�E�PH�E� �P�H�E�H�E�H� H�PH�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�E�H� � �E��}�vH���  �>   H�5��  H�="�  �  H�E�H� �U��H�E�H� H�PH�E�H�H�E�H� H�PH�E�H��    ��UH��H��H�}�H�E��    �   H���X���H��8 C H�PH�E�H���ÐUH��H��H�}�H��8 C H�PH�E�H�H�E�H���<�����ÐUH��H��H�}�H�E�H������H�E��   H���_p���ÐUH��SH��XH�}�H�u�H�U�H�M�H�E�� f��tH��  �W   H�5|�  H�=U�  �}  H�E�H�PH� H�E�H�U�H�E�H�������H�E�H���  ��tH�E�H���  ��t�   ��    ����   H�U�H�E�H��H�������E�}� t�E��   H�E�H������������t�H�U�H�E�H�H�E�H���o���������t�    �MH�E�H�H�E�H���L����H�E�H� H�PH�E�H��@���H�E�H������������t�   ��    H��X[]ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH���  �s   H�51�  H�=
�  �2  H�E�H�PH� H�E�H�U�H�E�H���x���H�E�H���F  ��tH�E�H���v  ��t�   ��    ����   H�U�H�E�H��H���s����E��}� t�E��   H�E�H���4���������t�H�U�H�E�H�H�E�H���$���������t�    �OH�E�H��������H�E�H� �H�E�H� H�PH�E�H��>���H�E�H�������������t�   ��    �ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH�-�  ��   H�5�  H�=¼  ��  H�E�H�PH� H�E�H�U�H�E�H���0���H�E�H�     H�E�H����  ��ttH�U�H�E�H��H���D����E��}� t�E��tH�E�H������������t�H�U�H�E�H�H�E�H�������������t�    �8H�E�H� H�PH�E�H��|���H�E�H������������t�   ��    ��UH��H��`H�}�H�u�H�U�H�M�H�E�� f��tH��  ��   H�5պ  H�=��  ��  H�E�H�PH� H�E�H�U�H�E�H���V  ��tH�E�H���f  ��t�   ��    ����   H�E�H� � �E؋E؅�u
�    �   H�E�H�E�H�E�H��H�E�H�U�H�M�H�E�H��H���x����E��}�tY�}� t�E��pH�U�H�E�H9�tH��  ��   H�5�  H�=�  �  H�E�H� H�PH�E�H�H�U�H�E�H��"��������H�U�H�E�H� H9�t�   ��    ��UH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}��   ]ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t2��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ªC H��H������H��`���H�5�  H������H���2���H��`���H�������    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t ��T���/v��T���9w�   �[�    �T��T���vFH��`���H�ªC H��H���6���H��`���H�5��  H���V���H���x���H��`���H���3����    ��UH��H��   H��X�����T�����T���wH��X���H���:�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���fv��T���@v��T���Fw�   �[�    �T��T���vFH��`���H�ªC H��H���X���H��`���H�5��  H���x���H��蚑��H��`���H���U����    ��UH��H��   H��X�����T�����T���wH��X���H���\�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ªC H��H���z���H��`���H�5h�  H��蚐��H��輐��H��`���H���w����    ��UH��H��   H��X�����T�����T���wH��X���H���~�����t�   ��    ���r  ��T���!�W  ��T���"�J  ��T���#�=  ��T���$�0  ��T���%�#  ��T���&�  ��T���'�	  ��T���(��   ��T���)��   ��T���*��   ��T���+��   ��T���,��   ��T���-��   ��T���.��   ��T���/��   ��T���:��   ��T���;��   ��T���<t~��T���=tu��T���>tl��T���?tc��T���@tZ��T���[tQ��T���\tH��T���]t?��T���^t6��T���_t-��T���`t$��T���{t��T���|t��T���}t	��T���~u�   �[�    �T��T���vFH��`���H�ªC H��H���j���H��`���H�5��  H��芎��H��謎��H��`���H���g����    ��UH��H��   H��X�����T�����T���wH��X���H���n�����t�   ��    ��t ��T��� v��T���~w�   �[�    �T��T���vFH��`���H�ªC H��H��谍��H��`���H�5>�  H���Ѝ��H������H��`���H��譍���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T��� t	��T���	u�   �n�    �g��T���vYH��`���H�ªC H��H�������H��`���H�5Ե  H������H��T�����H���  H���%���H��`���H��������    �ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��tD��T��� t-��T���	t$��T���
t��T���t��T���t	��T���u�   �[�    �T��T���vFH��`���H�ªC H��H������H��`���H�52�  H���$���H���F���H��`���H�������    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���v��T���~w�   �[�    �T��T���vFH��`���H�ªC H��H���J���H��`���H�5ȴ  H���j���H��茋��H��`���H���G����    ��UH��H��   H��X�����T�����T���wH��X���H���N�����t�   ��    ��t ��T���`v��T���zw�   �[�    �T��T���vFH��`���H�ªC H��H��萊��H��`���H�5�  H��谊��H���Ҋ��H��`���H��荊���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���@v��T���Zw�   �[�    �T��T���vFH��`���H�ªC H��H���։��H��`���H�5T�  H�������H������H��`���H���Ӊ���    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t��T���@v��T���Zw��T����� �U��T���vFH��`���H�ªC H��H������H��`���H�5�  H���?���H���a���H��`���H��������T�����UH��H��   H��X�����T�����T���wH��X���H���"�����t�   ��    ��t��T���`v��T���zw��T����� �U��T���vFH��`���H�ªC H��H���g���H��`���H�5��  H��臈��H��詈��H��`���H���d�����T�����UH��H��X ]ÐUH��H��H�}��u�H�U�H�E�H��H���   H�E���UH��H��0H�}�H�u�H�E�H���}��H�E؋ H�U�H�M�H�Ή��	���H�E�H����}����ÐUH��H��H�}�H�u�H�E�H����7  ��ÐUH��H��H�}�H�u�H�E�H���7  �����UH��H���   H��X���H��P�����L���H��@���H��`���H�«C H��H����  H��`���H�5��  H����  H��H��@���H��H����  H�5��  H����  H��H��P���H��H����  H�5}�  H���  H��L�����H����  H�5]�  H���  H�5P�  H���  H��H��X���H��H���l  H�56�  H���]  H���  H��`���H���:  ���UH��H���   H��X���H��P�����L���H��@���H��`���H�ªC H��H���,���H��`���H�5��  H���L���H��H��@���H��H���7���H�5��  H���(���H��H��P���H��H������H�5q�  H������H��L�����H������H�5Q�  H������H�5D�  H���Ӆ��H��H��X���H��H��辅��H�5*�  H��诅��H���х��H��`���H��茅����ÐUH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H��H�}��u�H�U�H�E�H��H���   H�E���UH��H��H�}�H�E�H� H�U�H��H��H����   H�E���UH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H���y��H�E�H� H�U�H�M�H��H���x   H�E�H���Zz�����UH��H��0H�}�H�u�H�E�H���Ky��H�E؋ H�U�H�M�H�Ή��_   H�E�H���z�����UH��H��H�}�H�u�H�E�H�U�H��H���3������UH��H�� H�}�H�u�H�U�H�U�H�E�H��H���M   ���UH��H��@�}�H�u�H�U�H�U�H�E�H��H���
y��H�U�H�M��E�H�Ή���   H�E�H���}y�����UH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=ï  �8��H�E�H���   H��u)H�E�H� H�U�H��H��H�������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�= �  �#7���u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��  H�E��E�    �E���~H��    H��uH�=�  �O6���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�  ��5���E��P�U�H��D�-H�U�H�E�H��H�������� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H���q   �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���:   �E��ڋE����E�}� x!�E�H��D���H�E���H���
   �m��ِ�ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=�  ��4��H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ��ÐUH��H�� H�}��E�    H�E�H�pH�U���   ��������u�
��uH�=­  �0/  ���UH��H�}�H�E�H���    ��]�UH��H��   H��`���H�«C H��H���X���H��`���H�5��  H���x���H��H�EH��H���   H������H��`���H���C������UH��H�� H�}�H�E�H�E�H�E�H������H�E�� ������tH�E�H���D����    ��   ��UH��H��H�}�H�E�H�E�H�E��   �H�E�H���������UH��H��H�}�H�u�H�U�H�E�H��H���   H�E���UH��H��0H�}�H�u�H�E�H����r��H�E�H� H�U�H�M�H��H���   H�E�H���s�����UH��H��`H�}�H�u�H�U�H�E�H�5��  H������H�E�H���r��H�E�H�M�   H��H���s��H�E�H�U�H�M�H��H���   H�E�H���Fs��H�E�H���:s�����UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���Z   �UH�E�� ��t%H�E�� ��tH��    H��uH�=�  �1��H�u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���   H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H���  H�E��E�    �E���~H��    H��uH�=�  ��0���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=ʫ  �e0���E��P�U�H��D�-H�U�H�E�H��H���]���� 9E�����tE�E�    H�U�H�E�H��H���7���� �U�)�9E�����t�U�H�E���H��������E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H�������E��ڋE����E�}� x!�E�H��D���H�E���H�������m��ِ�ÐUH��H��H�}�H�u�H��C H�PH�E�H�H�E��@H    H�E��@L    H�E�H�U�H�PPH�E�H��XH���  H�E�H�@    H�E�H�@�   H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�@0    H�E�H�@8    H�E��@@    H�E��@D    H�E�H��H�=zJ ��  ���UH��H���   H��H���H��C H�PH��H���H�H��H���H�P0H��H���H�@8H9�tFH��`���H�ªC H��H���Cy��H��`���H�5��  H���cy��H���y��H��`���H���@y��H��H���H�@H��t�o���H��H��H���H�@H��H���y��H��H���H��H�=�I �  H��X���H��X���H��H�=�I ��  ���UH��H��H�}�H�E�H�������H�E��p   H���O���ÐUH��H��H�}�H�E�H�@PH��tH�E�H�@PH�U�H�������ÐUH��H���   H��(���H�� ���H�����H�����H�����H��uH�W�  �W   H�5̩  H�=�  ����H��(���H���'  ������t
������%  H��(����@L����   H��(���H� H��(H� H�����H��8���H�� ���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��  H��8���H��uH��(����@D����H��(����PDH��8���H�����H��    �y  H��(����@@��tVH��(���H�@(H��tFH��@���H�«C H��H������H��@���H�5ݨ  H�������H������H��@���H������H��(����@@    H��(���H�PH��(���H�@(H9��  H��(���H���J
  �E��}� t�E���  H��(���H���  �E�}� t�E��  H��(���H����  H��(���H� H��(H� H��(���H�RH��(���H�qH��0���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��8  H��0���H��u1H��(����@D����H��(����PDH�����H�     �    ��   H��0���H��(���H�P H��0���H��(���H�P(H��(���H�PH��(���H�@(H9�rH���  ��   H�5"�  H�=}�  �����H��(���H�P(H��(���H�@H)�H��H�E�H�����H�E�H��H���,��H� H�E�H��(���H�PH��(���H�@H�H�U�H�� ���H��H���T��H��(���H�PH�E�H�H��(���H�PH�����H�U�H��    �ÐUH��H��   H�����H�����H�����H�� ���H�����H��uH���  ��   H�50�  H�=M�  �����H�����H���  ������t
������Q  H������@L����   H�����H�P0H�����H�@8H9�tH�Q�  ��   H�5��  H�=5�  ����H�����H� H��0H� H�����H�� ���H�����H������ЉE��}� t!H������@D����H������PD�E��  H�� ���H��uH���  ��   H�5=�  H�=Υ  �����H�� ���H�� ���H��    �e  H�����H�PH�����H�@H9�u@H�����H����  �E�}� t�E��*  H�����H���  �E��}� t�E��
  H������@@��uVH�����H�@(H��tFH��0���H�«C H��H���j���H��0���H�5��  H������H�������H��0���H���g���H������@@   H�����H�PH�����H�@H9�rH���  ��   H�5�  H�=��  �����H�����H�PH�����H�@H)�H��H�E�H�����H�E�H��H���)��H� H��(����E� H������@L��u@H��(���H������
   H���1���H�E�H�}� tH�E�H��H+����H��(����E�H��(���H��uH��  ��   H�5]�  H�=Q�  ����H�����H����  H��(���H�����H�HH�����H�@H�H�����H��H���xP��H�����H�P0H�����H�@8H9�trH�����H�PH�����H��0H��H���(��H�H�����H�P0H�����H�PH��(���H�H�E�H�����H�P8H�E�H��H����{��H�H�����H�P8�6H�����H�PH�����H�P0H�����H�PH��(���H�H�����H�P8H�����H�P(H�����H�HH��(���H�H�E�H�E�H��H���O{��H�H�����H�P(H�����H�PH��(���H�H�����H�P�}� tH�����H����  ������t������H��(���H�� ���H��    �ÐUH��H��H�}����E�H�E�H�@H��uH��  ��   H�5}�  H�=w�  �>���H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��E���ÐUH��H��H�}��u�H�E�H�P0H�E�H�@8H9�tH���  ��   H�5	�  H�=�  �����H�E��U�PL�    ��UH��H�}�H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�P0H�E�H�P8�]ÐUH��H��H�}�H�E�H���  ��UH��H�� H�}�H�u�H�E�H� H��8H� H�U�H�}�H�Ѻ   �    �ЉE��}� t�E��)H�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H��    ��UH��H��@H�}�H�uЉU�H�E�H����  �E��}� t�E���   �}�ueH�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� ��   H�E؋@D����H�E؉PD�E��|�}�t%�}�tH��  �
  H�5j�  H�=Ӡ  �+���H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� tH�E؋@D����H�E؉PD�E��H�E�H���&����    �ÐUH��H�� H�}�H�E�@H��t�    �_H�E�H� H��H� H�U�H�JHH�U�H��H���ЉE��}� t�E��/H�E�@H��uH�R�  �  H�5��  H�=0�  �_����    �ÐUH��H��H�}�H�E��@L��t�    �aH�E�H� H�� H� H�U�H�JLH�U�H��H���Ѕ�����t������/H�E��@L��uH��  �(  H�5�  H�=͟  ������    �ÐUH��H��0H�}�H�E�H��������E��}� t�E���  H�E�H�P0H�E�H�@8H9�u
�    �  H�E؋@H��u\H�E�H� H��8H� H�U�H�R0H��H�U�H�R H��H)�H�U�H�}�H�Ѻ   �ЉE��}� t�E��S  H�E�H�P0H�E�H�P �_H�E؋@H��tH��  �;  H�59�  H�=�  �����H�E�H�P H�E�H�@0H9�tH�ٹ  �<  H�5�  H�=��  �����H�E�H�P H�E�H�@8H9���   H�E�H� H��0H� H�U�H�J8H�U�H�R H)�I��H�U�H�JH�U�H�R H�4H�U�H�}�H��L���ЉE�}� tH�E؋@D����H�E؉PD�E��`H�E�H��uH�/�  �F  H�5[�  H�=�  ����H�E�H�P H�E�H�H�E�H�P H�E�H�P0H�E�H�H�E�H�P0�#����    �ÐUH��H�� H�}�H�E�H��������E��}� t�E��   H�E�@H��u4H�E�H�PH�E�H�@(H9�tH���  �U  H�5��  H�=͝  �x���H�E�H�P0H�E�H�@8H9�tH�c�  �W  H�5��  H�=��  �D���H�E�H�@    H�E�H�@     H�E�H�@(    �    ��UH��H�� H�}�H�E�H�@H��uH��  �`  H�5 �  H�=P�  �����H�E�H�@H��u-����H��H�E�H�@H��H���Nm��H�E�H�E�H�U�H�P���ÐUH��H�� H�}��u�H�U�H�E�H�U�H��H������H��� C H�PH�E�H�H�E��U�Pp��ÐUH��H�}�H�E��@p]ÐUH��H��   H��X���H��X���H�P0H��X���H�@8H9�tFH��`���H�ªC H��H���|h��H��`���H�5r�  H���h��H���h��H��`���H���yh��H��X����@p���  �E��}� t�E���    �ÐUH��H�� H�}�H�u�H�E�@pH�U�H�Ѻ   �    ���@  �E��}� uH�E��    �    ��}�-  uH�E��    �    ��E���UH��H��   H��X���H��P���H��    H��u6H�X�  ��  H�5D�  H�=��  ����H��P����    �    �   H��X����@p���h���E��}� uH��P����    �    �h�}�"  uH��P����    �    �KH��`���H�ªC H��H���g��H��`���H�5_�  H���!g��H���Cg��H��`���H����f��������ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u����  �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u�����  �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u��U�H�M�H�E�@pH�MЋU�H�u����7  �E��}� t�E���    �ÐUH��H�}��]ÐUH��H���   H��8���H��6 H�E�H�E�H���  H��H���H�E�H����  H��@���H��@���H��H���H��H����  ����   H��H���H���  H�E�H�E�H���[����E�}� tFH��P���H�ªC H��H���)e��H��P���H�5י  H���Ie��H���ke��H��P���H���&e��H��H���H���s  �]������UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���������UH��H��H�}�H�E�H�������ÐUH��H��H�}�H�u������H��H�E�H��H���8  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��p  H������H������H�������+   H��賳��H�����E�H������� <ru�}� t�E�   �   �E�   �   H������� <wu�}� t	�E�   ��E�   �M�  �oH������H�ªC H��H���c��H������H�5s�  H���c��H��H������� ����H����N��H�5a�  H���c��H���c��H������H���gc��H������H������� ����   H������� <+u
H��������H������� <bu
H�������H������� <eu�M� @  H�������H��P���H�ªC H��H���b��H��P���H�5��  H����b��H��H������H��H����b��H�5��  H���b��H����b��H��P���H���b��H�������(���H�������M�H��������H����  �E�}� tdH�%    H������H�E��    �.����H��H�U�H������H��H���  H��tH����    ��UH��H��H�}�H�u��C���H��H�E�H��H���  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��   ��\���H��P���H��`���H�ªC H��H���^a��H��`���H�5t�  H���~a��H�5��  H���oa��H���a��H��`���H���La������H��H�U�H��\���H��H���S  H��tH����    ��UH��H�� H�}�H�}� t
H�E�H����    H�E��E�    H�E�H�������������t�E�����H�E�H� H��H� H�U�H���Ѕ�����t�E�����H�E�H��������E���UH��H��0H�}�H�u��U�H�}� t
H�E�H����    H�E��U�H�M�H�E�H��H��������E�}� tdH�%    H������H�E��������    ��UH��H��0H�}�H�}� t
H�E�H����    H�E�H�U�H�E�H��H��������E�}� t!dH�%    H������H�E�H�������H�E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���t���������t�������    ��UH��H��H�}�H�E�H��������UH��H��@H�}�H�uЉU�H�M�H�}� t
H�E�H����    H�E��}�u@H�E��   H���g����E�}� ��   dH�%    H������H�E�������   �}�u9H�E��   H���!����E��}� t{dH�%    H������H�E��������a�}�u9H�E��   H��������E�}� t<dH�%    H������H�E�������"dH�%    H�������   �������    ��UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E��   �    H���v���H�E�@<�����H�E�P<���UH��H�� �}�H�u�H�}� t
H�E�H����    H�E��E���H�E���H�������E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���$������UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H���7a��H�E�H�E�H���4��D� H�E�H������H������I��H�E�H�ƿx   �R��H��L��D��H������H��H��8[A\A]]�UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H���`��H�E�H�E�H���4��D� H�E�H������H�������I��H�E�H�ƿx   �oQ��H��L��D��H���!���H��H��8[A\A]]�UH��H���}��u��}���   �}���  ��   H�=�, ��   �    �    H�=�, �����H�S H�5�, H��6�A H���Ķ���    �   H�=,- ����H�  H�5- H��6�A H��葶���    �   H�=y- �f���H�� H�5f- H��6�A H���^���H�=�- �}���H�� H�5�- H�=t����8������UH����  �   �����]ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@ �]�UH��SH��(H�}�H�u�H�E�H��uH��    H��uH�=�  ���H�E�H���  H�E�H�U�H�E�H��H���  �@��tH��    H��uH�=�  �s��H�U�H�E�H��H���j  H� H������tH��    H��uH�=.�  �9��H�U�H�E�H��H���0  H�@H������tH��    H��uH�=K�  ����H�E�H�@H��uH�E�H���  H��H�E�H��HH�E�H�XH�U�H�E�H��H����  H�XH�E�H����  H��H�E�H�PH�E�H��H���  H�H�E�H�U�H�PH�U�H�E�H��H���|  �@H�U�H�E�H��H���  H�E�H��([]�UH��H�� H�}�H�u�H�U�H�E�H��H���7  �@����tH��    H��uH�=��  ���H�U�H�E�H��H���A  H�E��ÐUH��SH��8H�}�H�u�H�E�H��uH��    H��uH�=��  ���H�U�H�E�H��H���  �@����tH��    H��uH�=ϒ  ���H�U�H�E�H��H���y  H���  H�E�H�U�H�E�H��H���Z  H�@H�E�H�E�H��u9H�E�H�PH�E�H9�tH��    H��uH�=��  ���H�E�H�U�H�P�pH�E�H����  H��H�E�H��H����  H�PH�E�H9�����tH��    H��uH�=��  ���H�]�H�E�H���  H��H�E�H��H���  H�XH�}� ueH�E�H� H���|  H��H�E�H9�����tH��    H��uH�=Ғ  �U��H�E�H���  H�E�H�E�H���s  H��H�E�H��   H�U�H�E�H��H���!  H� H���  H��H�E�H9�����tH��    H��uH�=ƒ  ����H�U�H�E�H��H����  H���   H�E�H�E�H����  H��H�U�H�E�H��H���  H�H�E�H���  H��H�E�H9�����tH��    H��uH�=Ò  �f��H�U�H�E�H��H���]  H�     H�U�H�E�H��H���C  H�@    H�U�H�E�H��H���(  �@ H�E�H��8[]ÐUH��H�� H�}�H�E�H� H����   H��H�E�H��H���-  H�E��ÐUH��H�� H�}�H�E��    H���	  H�E��ÐUH��H��H�}�H�u�H�U�H�E�H��H����   ����UH��H��H�}�H�E�H�H�E�H��H����   H�H�E�H�H�E���UH��H�}�H�E�H� ]�UH��H��H�}�H�u�H�}� t-H�E�H� H� H�U�H����H�M�H�E��p   H��H����   ����UH��H�}�H�E�]�UH��H��H�}�H�u�H�E�H����  H��H�E�H��H����  ��UH��H�}�H�E�H� ]ÐUH��H�}�H�u�H�E�H�U�H��]�UH��H�}�H�u�H�E�H�H�E�H� H9���]�UH��H��H�}�H�u�H�E�H���P  H��H�E�H��H���X  ��UH��SH��hH�}�H�u�H�U�H�}� �  H�}� �  vH�U�H�E�H��H���T����  H�E�H�E�H�E�H%  ��H�E�H�E�H�U�H��H���'b������tH��    H��uH�=��  ���H�E��@HH�H��H��H��H�E�H�H��H�E�H�E��@H���J��H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=�  �J��H�U�H�E�H��H���=_��H�E�H�@PH�����E�H�E��@L��uH��    H��uH�=��  ���H�E�H�ƿ   ��G��H��H���a��H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H���a������t�   ��    ��tH��    H��uH�=��  ���H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H����`��H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���N^����H��h[]�UH��H��H�}�H�E�H���   ��UH��H�}�H�u�X   H�E�H�]�UH��H�}�H�E�]�UH��H��H�}�H��� C H�PH�E�H�H�E�H���������ÐUH��H��H�}�H�E�H������H�E��x   H���(����UH��H��0�}�H�u�H�U�H�M�H�U�H�M��E�H�Ή���,��H�H�E�H�}��u������H�E�H�U�H��    ��UH��H��0�}�H�u�H�U�H�M�H�U�H�M��E�H�Ή��`,��H�H�E�H�}��u������H�E�H�U�H��    ��UH��H��0�}�H�u��U�H�M؋U�H�M��E�H�Ή��,��H�E�H�}��u������H�E�H�U�H��    ��UH��H��0H�}�u�H�U؋U�H�E��H���X+���E�H�}� u������H�E؋U���    ��UH��H���}��E����\+���    ��UH��H�� H�}�u�H�E�    H����*���E��}� t�E����"+���    ��   ��UH��H�}��]�f�H�� H���t3UH��S� C H��D  ��H��H�H���u�H��[]�f.�     �����         /close.bmp /shell.lef /dev/mouse0                       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    ../options/ansi/generic/stdlib-stubs.cpp *string != '+' !negative !"Not implemented" mlibc: srandom() is a no-op i == j !"decode_wtranscode() errors are not handled" mlibc: Broken mbtowc() called wc mbs max_size *mbs MLIBC_DEBUG_MALLOC mlibc (PID ?): free() on    mlibc (PID ?): malloc() returns  mlibc (PID ?): realloc() on   returns  !(reinterpret_cast<uintptr_t>(p) & (align - 1)) ../options/internal/include/mlibc/strtofp.hpp   !"hex numbers in strtofp are unsupported"       ../subprojects/frigg/include/frg/slab.hpp:393: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:399: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:417: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:425: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:432: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:435: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/slab.hpp:252: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:262: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:263: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:265: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:280: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:281: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:283: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:295: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:344: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:361: Assertion 'fra->type == frame_type::large' failed!       ../subprojects/frigg/include/frg/slab.hpp:362: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:504: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:525: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:550: Assertion '!(area_size & (page_size - 1))' failed! 0x    ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! 0123456789abcdef ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       strtofp strtofp strtofp strtol rand_r abort     at_quick_exit   quick_exit system mktemp        bsearch abs labs llabs ldiv lldiv mblen mbtowc wctomb   mbstowcs        wcstombs lock   posix_memalign  strtod_l              $@       �           A               �                   �@                                            @               ../options/internal/include/mlibc/charcode.hpp nseq.it == nseq.end wseq.it == wseq.end alnum alpha blank cntrl digit graph lower print punct space upper xdigit mlibc: wctype(" ") is not supported     ../options/ansi/generic/ctype-stubs.cpp !"Not implemented"      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       promote iswctype        towlower        towupper                ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"   mlibc: environment string "      " does not contain an equals sign (=)   ../options/ansi/generic/environment.cpp environ == vector.data() !vector.back() ../options/ansi/generic/environment.cpp:84: Assertion 'k != size_t(-1)' failed! vector.size() >= 2 && !vector.back() s != size_t(-1)    !"Environment strings need to contain an equals sign" mlibc: environment variable " " contains an equals sign %s=%s     asprintf(&string, "%s=%s", name, value) > 0 string      ../subprojects/frigg/include/frg/string.hpp:71: Assertion 'from + size <= _length' failed!      ../subprojects/frigg/include/frg/slab.hpp:393: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:399: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:417: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:425: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:432: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:435: Assertion '!slb->available || slb->contains(slb->available)' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{    ../subprojects/frigg/include/frg/slab.hpp:504: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:252: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:262: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:263: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:265: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:280: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:281: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:283: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:295: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/slab.hpp:525: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/slab.hpp:550: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! 0123456789abcdef ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed! lock     assign_variable unassign_variable getenv putenv setenv          ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    ../options/ansi/generic/stdio-stubs.cpp new_buffer count < limit !"Not implemented"     Library function fails due to missing sysdep    ��������������������ċ��ы��    Functionality is not implemented max_size > 0 
 %s:  %s
 returns:       mlibc: File locking (flockfile) is a no-op      mlibc: File locking (funlockfile) is a no-op    mlibc: File locking (ftrylockfile) is a no-op   mlibc: fread() I/O errors are not handled       mlibc: fwrite() I/O errors are not handled do_scanf: ' not implemented! do_scanf: m not implemented!    թ������������������������������������������������������������������������������������������������������������������������������������������������������������������������	������C������W��������������������������������������������ĩ�����������u���������������������������)���������������0���������������̱��R�������������.������)������������../subprojects/frigg/include/frg/formatting.hpp:200: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:213: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:217: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:221: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:225: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:229: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:235: Assertion '!opts.always_sign' failed!      ../subprojects/frigg/include/frg/formatting.hpp:236: Assertion '!opts.plus_becomes_space' failed!       ../subprojects/frigg/include/frg/formatting.hpp:240: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:247: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:254: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:258: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:262: Assertion '*s >= '0' && *s <= '9'' failed! ../subprojects/frigg/include/frg/formatting.hpp:266: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:275: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:279: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:286: Assertion '*s' failed! `��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������ί�������������������������-�����������>�����������������������O���o����������� �������������������������������r�������������������������������������������W���ݱ���������������������������������o���    ../subprojects/frigg/include/frg/slab.hpp:252: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:262: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:263: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:265: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:280: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:281: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:283: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:295: Assertion 'slb->available' failed! !opts.fill_zeros !opts.left_justify !opts.alt_conversion opts.minimum_width == 0      szmod == frg::printf_size_mod::default_size !opts.precision     [31mmlibc: Unknown printf terminator ' '[39m !"Illegal printf terminator"     ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:525: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:550: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/optional.hpp:97: Assertion '_non_null' failed! ../subprojects/frigg/include/frg/formatting.hpp:299: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:300: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:301: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:302: Assertion 'opts.minimum_width == 0' failed! 0x     ../subprojects/frigg/include/frg/formatting.hpp:307: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:308: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:309: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:310: Assertion 'opts.minimum_width == 0' failed!        ../subprojects/frigg/include/frg/formatting.hpp:311: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:312: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:316: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:317: Assertion '!opts.alt_conversion' failed! (null)    ../subprojects/frigg/include/frg/formatting.hpp:340: Assertion 'szmod == printf_size_mod::long_size' failed!    (   n   u   l   l   )           ../subprojects/frigg/include/frg/formatting.hpp:363: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/formatting.hpp:373: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:374: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:383: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:395: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:412: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:418: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:419: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:431: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:436: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:437: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:453: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:454: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:455: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:469: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:476: Assertion '!"Unexpected printf terminal"' failed! %f       ../subprojects/frigg/include/frg/formatting.hpp:493: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed! 0123456789abcdef      ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed! remove rename  renameat        tmpfile tmpnam  freopen setbuf scanf    operator() vscanf       operator()      operator()      vsscanf fwprintf        fwscanf vfwprintf       vfwscanf        swprintf        swscanf vswprintf       vswscanf        wprintf wscanf  vwprintf        vwscanf fgets fgetwc fgetws fputwc fputws fwide getwc   getwchar putwc  putwchar        ungetwc fgetpos fsetpos lock    getdelim        operator() expand       fgets_unlocked  �������������������������������������������������������������������������������������������!��������������������������������D�����������!���������!��������������������G���G���G���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l���l�������l���l���l���l���l���l���l���l���l���l�����������G���G���G���l�������l���l���l�������������������l���l�������l�������l���l�����������������������������������������������������������������������������������J�����������������������������������������������J�������������������J������������������T���J�����������������������J�����������J������������4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4�������4���4���4���4���4���4���4���4���4���4���M����������������4�������4���4���4���p�����������M���4���4���M���4�������4���4����������V���V���V���V���V���V���V���V���V���V���V������V���V���V���V������V���V���V���V���V������V���V���V���V���V�������V���V������b�����������������������������������������������]�������������������]�����������������������c�����������������������F�����������^���������������������������������������{���������������{�������������������������������������d��������| �����������������������������������������������������������������������������������������������������../options/ansi/generic/string-stubs.cpp !"Not implemented"     Functionality is not implemented        Operation would block (EAGAIN) Access denied (EACCESS) Bad file descriptor (EBADF) File exists already (EEXIST) Access violation (EFAULT) Operation interrupted (EINTR) Invalid argument (EINVAL) I/O error (EIO)       Resource is directory (EISDIR)  No such file or directory (ENOENT) Out of memory (ENOMEM)       Expected directory instead of file (ENOTDIR)    Operation not implemented (ENOSYS)      Operation not permitted (EFAULT) Broken pipe (EPIPE) Seek not possible (ESPIPE) No such device or address (ENXIO) Unknown error code (?)    �G��oH��oH��oH��zG��oH���G��oH��oH��oH��oH��oH��oH��oH��oH��oH��oH���G���G��oH��oH��oH��oH���G���G���G��oH���G��oH��oH��oH��oH��oH��oH��oH��oH��oH��oH��oH��oH��oH��H��oH��oH��oH��H��oH��oH��oH��.H��oH��!H��oH��oH��oH��oH��oH��bH��oH��oH��oH��;H��HH��oH��oH��oH��oH��UH��    strxfrm strtok wcstod wcstof    wcstold wcstol  wcstoll wcstoul wcstoull wcscpy wcsncpy wmemcpy wmemmove wcscat wcsncat wcscmp  wcscoll wcsncmp wcsxfrm wmemcmp wcschr  wcscspn wcspbrk wcsrchr wcsspn wcsstr wcstok wcslen     wmemset         ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    ../subprojects/frigg/include/frg/slab.hpp:252: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:262: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:263: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:265: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:280: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:281: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:283: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:295: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:393: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:399: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:417: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:425: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:432: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:435: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:525: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:550: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/slab.hpp:504: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! lock             ../sysdeps/lemon/generic/lemon.cpp !(size & 0xFFF)              sys_anon_allocate               ../options/internal/generic/allocator.cpp       !mlibc::sys_anon_allocate(length, &ptr) !mlibc::sys_anon_free((void *)address, length) map unmap                        ../options/internal/generic/charcode.cpp        (uc & 0b1100'0000) == 0b1000'0000 || (uc & 0b1111'1000) == 0b1111'1000  (uc & 0b1100'0000) == 0b1000'0000       wc <= 0x7F && "utf8_charcode cannot encode multibyte chars yet" !st.__progress cps.it == cps.end        encode_wtranscode       operator()              decode_wtranscode_length        operator()      decode_wtranscode decode                mlibc: charset::is_alpha() is not implemented for the full Unicode charset      mlibc: charset::is_digit() is not implemented for the full Unicode charset      mlibc: charset::is_xdigit() is not implemented for the full Unicode charset     mlibc: charset::is_alnum() is not implemented for the full Unicode charset      mlibc: charset::is_punct() is not implemented for the full Unicode charset      mlibc: charset::is_graph() is not implemented for the full Unicode charset      mlibc: charset::is_blank() is not implemented for the full Unicode charset      mlibc: charset::is_space() is not implemented for the full Unicode charset      mlibc: charset::is_print() is not implemented for the full Unicode charset      mlibc: charset::to_lower() is not implemented for the full Unicode charset      mlibc: charset::to_upper() is not implemented for the full Unicode charset      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed! 0123456789abcdef       ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!         In function  , file  : 
 __ensure( ) failed   ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed! 0123456789abcdef       ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!              __cxa_guard_acquire contention  mlibc: Pure virtual function called from IP  0x ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed! 0123456789abcdef       ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!                       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    mlibc warning: File is not flushed before destruction   ../options/ansi/generic/file-io.cpp max_size    mlibc: Cannot read-write to same pipe-like stream __offset < __valid_limit __dirty_begin == __dirty_end io_size > 0 && "io_write() is expected to always write at least one byte" __offset < __buffer_size chunk __offset       __dirty_begin == __dirty_end && "update_bufmode() must only be called before performing I/O"    whence == SEEK_SET || whence == SEEK_END _type != stream_type::unknown  _bufmode != buffer_mode::unknown        _type == stream_type::pipe_like __io_offset == __dirty_begin __offset == __valid_limit __buffer_size    mlibc warning: File is not flushed before closing       Library function fails due to missing sysdep    mlibc: sys_isatty() failed while determining whether stream is interactive      mlibc warning: Failed to flush file before exit() Illegal fopen() mode ' ' Illegal fopen() flag '       [31mmlibc: fdopen() ignores the file mode [39m        ../subprojects/frigg/include/frg/list.hpp:104: Assertion 'element' failed!      ../subprojects/frigg/include/frg/list.hpp:106: Assertion '!h(borrow).in_list' failed!   ../subprojects/frigg/include/frg/list.hpp:107: Assertion '!h(borrow).next' failed!      ../subprojects/frigg/include/frg/list.hpp:108: Assertion '!h(borrow).previous' failed!  ../subprojects/frigg/include/frg/slab.hpp:393: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:399: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:417: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:425: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:432: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:435: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/list.hpp:79: Assertion 'h(ptr).in_list' failed!        ../subprojects/frigg/include/frg/list.hpp:164: Assertion 'it._current' failed!  ../subprojects/frigg/include/frg/list.hpp:165: Assertion 'h(it._current).in_list' failed!       ../subprojects/frigg/include/frg/list.hpp:170: Assertion '_back == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:173: Assertion 'h(traits::decay(next)).previous == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:179: Assertion 'traits::decay(_front) == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:183: Assertion 'traits::decay(h(previous).next) == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:188: Assertion 'traits::decay(erased) == it._current' failed! ../subprojects/frigg/include/frg/slab.hpp:252: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:262: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:263: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:265: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:280: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:281: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:283: Assertion '!"slab_allocator corruption. Possible write to unallocated object"' failed!   ../subprojects/frigg/include/frg/slab.hpp:295: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:504: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:525: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:550: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/slab.hpp:467: Assertion 'slb->contains(pointer)' failed!       ../subprojects/frigg/include/frg/slab.hpp:471: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:478: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:481: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! 0123456789abcdef ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed! lock read write unget update_bufmode seek     _init_type      _init_bufmode   _write_back _reset              _ensure_allocation              determine_bufmode              zR x�        r{��I    A�CD     <   Eh���    A�C�     \   |{��2    A�Cm      |   �h��   A�C    �   �i���   A�C� $   �   zk���   A�CN�����   �   p��A
   A�C         
{��-    A�Ch         {��    A�CL      @  
{��"    A�C]      `  {��-   A�C(    �  |��"    A�C]       �  |���    A�CE��      �  �|���    A�C�     �  Wy��>    A�Cy        }��8    A�Cs      $  Uy��    A�CP      D  }��k       <   X  l}���    B�A�D �G0U
 AABI[ AABL   �  �}��k    R�E�H �D(�M0R
(A ABBHD(M� A�B�B�      �  ~��3    A�q        @~��             L~���    A�A��A  $   <  �~��     D�LG FAA      d  �~��       H   x  �~��I   B�F�E �H(�G0�A8�GP8A0A(B BBB   T   �  ���o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T     ���o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB     t   ���(    DK X  <   �  ����    P�B�B �A(�A0�j(A BBBA�����0   �  d����    H�F�E �A(�� ABB        ���            ���          ,  ���          @  ���          T   ���          h  ����       �   |  ���R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   $  ����m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        |  ����:    A�Cu      �  υ��6    A�Cq      �  ���?    A�Cz      �  ���?    A�Cz      �  #���A    A�C|        D���@    A�C{      <  d���8    A�Cs      \  |���M    A�CH     |  ����>    A�CA�x   �  ǆ��@    A�C{      �  ����    A�C     �  K����    A�C�     �  ���F    A�CA       (���Z    A�CU     <  b����    A�C�     \  ���<    A�Cw      |  *���     A�C[      �  *����    A�C�     �  �����   A�C�    �  g���    A�CM      �  Z���\    A�CW     	  �����    A�C�     <	  
���    A�CZ      \	  
���6    A�Cq      |	   ���Q    A�CL     �	  Q���    A�CN      �	  D���B    A�C}      �	  f���    A�CQ      �	  ����-    A�Ch      
  ����$    A�C_      <
  ����$    A�C_      \
  ����$    A�C_      |
  ����3    A�Cn      �
  ����%    A�C`      �
  ����9    A�Ct      �
  ч��J   A�CE    �
  ����+    A�Cf        ���G   A�CB    <  -���+    A�Cf      \  8���    A�CU      |  2���+    A�C      �  A���"    A�C]      �  C���Z    A�CU     �  }���U    A�CP     �  ����V    A�CQ       ���#    A�C      4  ���)    A�Cd      T  ����+    A�C      p  ���    A�C      �  ���    A�C      �  ����*    A�C      �  ���+    A�C      �  ���+    A�C      �  *����    A�C�       ���   A�C    <  ݍ��*    A�C      X  ���+    A�C      t  ����+    A�C      �  	���&    A�Ca      �  ���/    A�C      �  "���/    A�C       �  5���   A�CE��        ���1   A�C,    ,  &���.    A�C      H  8���=   A�C8    h  U���3    A�C      �  ԙ��    A�Cz     �  3����    A�C�     �  ,����    A�C�     �  ����    A�C�       �����    A�C�      $  B����    A�CE��      H  ���3    A�C      d  p���#    A�C^      �  t���    A�CV      �  p���V    A�CQ     �  ����M   A�CH    �  Ӝ��L   A�CG      ����   A�C    $  ����)    A�Cd      D  ���    A�CF      d  ���)    A�Cd      �  ����,    A�Cg      �  ���)    A�Cd       �  ���h   A�CE�^      �  V����   A�CH��        ���#   A�CE�     0  ���+    A�Cf      P  ���    A�CF      p  ت��    A�CF      �  Ī��4    A�Co      �  ت��E    A�C@     �  ����&    A�Ca      �  ���E    A�C@       *���2    A�Cm      0  <���'    A�Cb      P  D����    A�C�     p  ����    A�C�     �  ����O    A�CJ     �  ����    A�CQ      �  ����I    A�CD     �  ج���    A�C�       �����    A�C�     0  H���X    A�CS      P  ����D   A�CE�:     t  �����    A�C�     �  t���L    A�CG      �  �����    A�CE��      �  ���*    A�Ce      �  "���}    A�Cx       ����    A�CL      8  q���    A�CY      X  o���    A�CY       x  n���a   A�CE�W     �  ����    A�CY       �  �����   A�CE��     �  ���    A�CL         ���j    A�Ce        N���(    A�Cc      @  V���    A�CY       `  T���7   A�CE�-     �  g���    A�CY       �  f���7   A�CE�-      �  z���a   A�CE�W     �  ����    A�CY         �����   A�CE��     0  ���d    A�C_     P  b���j    A�Ce      p  ����7   A�CE�-      �  ����7   A�CE�-     �  Կ��K    A�CF     �   ����    A�C�     �  �����    A�C�       0���    A�CQ      8  &���    A�CY      X  $���1    A�Cl       x  6����   A�CE��     �  ����    A�CX      �  ����H    A�CC     �  ����    A�CZ      �  ����    A�CZ        ����V   A�CQ    <  0���    A�CQ      \  &���H    A�CC     |  N���    A�CY      �  L���1    A�Cl       �  ^����   A�CE��     �  ����    A�CX         ����V   A�CQ       0���W    A�CR     @  g���1    A�Cl       `  x����   A�CE��      �  �����   A�CE��     �  p���    A�CJ      �  _���    A�CJ       �  N����   A�CE��        �����   A�CE��     0  F���1    A�Cl      P  W����   A�C�    p  ����(    A�Cc      �  �����    A�C�     �  ����/    A�Cj       �  ����    A�CP          �  D���   A�C      0���0    A�Ck      4  ����V    A�CQ     T  -���V    A�CQ     t  c���V    A�CQ     �  ����V    A�CQ     �  ����V    A�CQ     �  ���V    A�CQ     �  ;���V    A�CQ       q���V    A�CQ     4  ����V    A�CQ     T  ����V    A�CQ     t  ���V    A�CQ     �  I���K    A�CF     �  t���J    A�CE     �  ����S    A�CN     �  ����S    A�CN       ���S    A�CN     4  7���S    A�CN     T  j���S    A�CN     t  ����S    A�CN     �  ����S    A�CN     �  ���S    A�CN     �  6���S    A�CN     �  i���S    A�CN       ����S    A�CN     4  ����H    A�CC     T  �����   A�C�    t  ����.    A�C      �  ����Q    A�CL     �  ����Q    A�CL     �  ���*    A�C      �  "���*    A�C        l���R    A�CM      (  ����    A�Cz         L  6���*    A�Ce       l  �����   A�CJ���   �  \���o    A�Cj     �  �����    A�C�      �  X���?   A�CE�5      �  s���r   A�CE�h        �����    A�C�      8   k����    A�CE��       \   �����   A�CJ���   �   ����>    A�Cy      �   ���S    A�CN     �   @���    A�CL      �   2���    A�CM       !  $���6    A�Cq       !  :���r    A�Cm     @!  ����>    A�Cy      `!  ����F    A�CA     �!  ����    A�CM      �!  ����4    A�Co      �!  ����w    A�Cr      �!  .����    A�CE�{      "  ����!    A�C\      $"  ����%    A�C`      D"  ����    A�CM      d"  ����    A�CL      �"  {���O    A�CJ     �"  ����I    A�CD     �"  ����I    A�CD     �"  ����*    A�Ce       #  ���   A�CE��      (#  ����   A�C    H#  ����N    A�CI     h#  ����J    A�CE     �#  #����    A�C�     �#  ����U    A�CP      �#  �����   A�C�        �#  �0��&    A�Ca      $  �0��H    A�CC      ,$  �0��e    A�CE�[      P$  �0��M    A�CH     p$  1��&    A�Ca      �$  $1��<    A�Cw      �$  @1��g    A�Cb     �$  �1��c    A�C^     �$  �1��6    A�Cq      %  �1��Q    A�CL     0%  2��S    A�CN     P%  H2��O    A�CJ     p%  x2��.    A�Ci      �%  �2��	   A�C    �%  p3��L    A�CG     �%  �3��S    A�CN     �%  �3��O    A�CJ     &  ,���+    A�C      ,&  ;����    A�C�     L&  ����5    A�C      h&  ����#    A�C      �&  ����+    A�C      �&  ����3    A�C      �&  ����2    A�Cm      �&  ����    A�C�     �&  �����    A�C�     '  5����    A�C�     <'  �����    A�C�     \'  V���x    A�C      x'  �����    A�C�     �'  J����    A�C�     �'  ����    A�CO      �'  ����0    A�Ck      �'  �����    A�C�     (  ����}    A�Cx     8(  ����b    A�C]     X(  :���[    A�CV     x(  u���`    A�C[     �(  ����/    A�Cj      �(  ����/    A�C       �(  �����    A�CH��      �(  �����    A�C�     )   ���3    A�C      4)  ���x    A�C      P)  s���x    A�C      l)  ����3    A�C      �)  ����3    A�C      �)  ����x    A�C      �)  Y���x    A�C      �)  ����7    A�C      �)  ����7    A�C      *  ����x    A�C      0*  G���x    A�C      L*  ����/    A�C      h*  ����/    A�C      �*  ����D    A�C      �*  �����    A�C�     �*  ����K    A�CF     �*  ����"    A�C]      +  ����P    A�CK     $+  ����%    A�C`      D+  ���    A�CU      d+  ����    A�CU      �+  ����    A�CS      �+  ����    A�CS      �+  ����I    A�CD     �+  ���"    A�C]      ,  ���$    A�C_      $,  ���    A�CR      D,  ����    A�C�     d,  ����+    A�C      �,  ����2    A�C      �,  ����.    A�C      �,   ��/    A�C      �,   ��.    A�C      �,  ' ��+    A�C      -  6 ��#    A�C      (-  = ��.    A�C      D-  O ��*    A�C      `-  ] ��.    A�C      |-  o ��2    A�Cm      �-  � ��2    A�Cm      �-  � ��/    A�C      �-  � ��/    A�C      �-  � ��    A�CQ      .  � ��    A�CO      4.  � ��    A�CO      T.  � ���    A�C~      t.  � ���   A�CH��     �.  ���6    A�C      �.  ����    A�C�     �.  C���    A�C�     �.  ���[    A�CV     /  ���[    A�CV     4/  4��[    A�CV     T/  o��    A�CQ      t/  e��    A�CO      �/  Y��    A�CO      �/  M��D    A�C      �/  q��;   A�C6    �/  ���;   A�C6    0  ���2    A�C      00  �)��    A�CM      P0  ����   A�C�    p0  �)��*    A�Ce      �0  �)���   A�C�    �0  ����   A�C�    �0  H0��*    A�Ce      �0  R0���   A�C�    1  �6��+    A�Cf      01  
7��*    A�Ce      P1  7���   A�C�    p1  �=��*    A�Ce      �1  �=���   A�C�    �1  vD��    A�CK      �1  fD��1    A�Cl      �1  xD��)    A�Cd       2  �D��N    A�CE�D      42  �D��)    A�Cd       T2  �D��N    A�CE�D       x2  �D���   A�CH��     �2  �H��1    A�Cl      �2  �H��)    A�Cd       �2  �H���   A�CH��      3  dL��1    A�Cl       3  vL��)    A�Cd       @3  �L���   A�CH��     d3  4P��1    A�Cl      �3  FP��)    A�Cd       �3  PP���   A�CH��      �3  T���    A�CE��      �3  �T��    A�CI      4  �T��;    A�Cv      ,4  �T��x   A�Cs     L4  >[���    A�CE��       p4  �[���    A�CE��       �4  �\���    A�CE��       �4  \]���    A�CE��       �4  ^���    A�CE��        5  �^���    A�CE��       $5  v_���   A�CE��     H5  g��d    A�C_     h5  Lg��*    A�Ce      �5  Vg��x   A�Cs     �5  �m���    A�CE��       �5  dn���    A�CE��       �5  o���    A�CE��       6  �o���    A�CE��       86  ~p���    A�CE��       \6  4q���    A�CE��       �6  �q���   A�CE��     �6  wy��d    A�C_     �6  �y��x   A�Cs     �6  ����    A�CE��       7  ʀ���    A�CE��       ,7  |����    A�CE��       P7  2����    A�CE��       t7  ����    A�CE��       �7  �����    A�CE��       �7  L����   A�CE��     �7  ݋��d    A�C_      8  !���x   A�Cs      8  z����    A�CE��       D8  0����    A�CE��       h8  ����    A�CE��       �8  �����    A�CE��       �8  J����    A�CE��       �8   ����    A�CE��       �8  �����   A�CE��     9  C���d    A�C_     <9  ����J    A�CE     \9  ����    A�CL      |9  ����J    A�CE     �9  ̞��W    A�CR     �9  ���Y    A�CT     �9  >���    A�CM      �9  0����    A�C�     :  ����U    A�CP     <:  ���W    A�CR     \:  ���G    A�CB     |:  B���W    A�CR     �:  y����    A�C�     �:  ����U    A�CP     �:  -���W    A�CR     �:  d���W    A�CR     ;  �����    A�C�     <;  ���U    A�CP     \;  O���W    A�CR     |;  ����W    A�CR     �;  �����    A�C�     �;  <���U    A�CP     �;  q���W    A�CR     �;  �����   A�C�    <  0����   A�C�    <<  �����   A�C�    \<  7����   A�C�    |<  ����J    A�CE     �<  ����   A�C�    �<  q����   A�C�    �<  �����   A�C�    �<  x����   A�C�    =   ����   A�C�    <=  �����   A�C�    \=  ����   A�C�    |=  �����   A�C�    �=  ����   A�C�    �=  �����   A�C�    �=  '����   A�C�    �=  �����   A�C�    >  .����    A�C�     <>  �����    A�C�     \>  "����   A�C�    |>  ����S    A�CN     �>  ɾ���    A�C�     �>  0���;    A�Cv      �>  K����    A�C}     �>  ����r    A�Cm     ?  ����r    A�Cm     <?  Q���%    A�C`      \?  V����    A�C�     |?  ����3    A�C      �?  ����Y    A�CT     �?  ���i    A�Cd     �?  V���m    A�Ch     �?  ����n    A�Ci     @  ����p    A�Ck     8@  A���m    A�Ch     X@  �����    A�C�     x@  !���/    A�C      �@  4���\    A�CW     �@  p���/    A�C      �@  ����/    A�C      �@  ����/    A�C      A  ����2    A�C      $A  ����2    A�C      @A  ����2    A�C      \A  ����2    A�C      xA  ���/    A�C      �A  ���3    A�C      �A  +���3    A�C      �A  B���3    A�C      �A  Y���/    A�C      B  l���3    A�C       B  ����/    A�C      <B  ����/    A�C      XB  ����3    A�C      tB  ����3    A�C      �B  ����3    A�C      �B  ����.    A�C      �B   ���/    A�C      �B  ���/    A�C       C  &���.    A�C      C  8���/    A�C      8C  K���/    A�C      TC  ^���3    A�C      pC  u���f    A�Ca     �C  ����+    A�C      �C  ����2    A�C      �C  ����@   A�C;    �C   ���]    A�CX     D  =���7    A�Cr       (D  T���H    A�CC         LD  x���W    A�CR     lD  ����J    A�CE     �D  ����a    A�C\     �D  ���    A�CI       �D  ���P    A�CE�F      �D  4���    A�CI      E  "����    A�C�     0E  ����    A�CM      PE  ����*    A�Ce      pE  ����.    A�Ci      �E  ����>    A�Cy      �E  ����   A�C     �E  ����0    A�Ck          �E  ����3    A�Cn      F  �����    A�C     4F  1���    A�CN      TF  $���    A�C          tF  Z���    A�CP      �F  �����    A�C�     �F  v���Q    A�CL     �F  ����R    A�CM     �F  ����,    A�Cg      G  ����    A�CI      4G  ����    A�CI       TG  ����P    A�CE�F      xG  ���    A�CI      �G  ����    A�CM      �G  ����%    A�C`       �G  ����{    A�CG��o    �G  B���$    A�C_      H  F���7    A�Cr      <H  ]���
    A�CE      \H  H���    A�CQ      |H  >���$    A�C_      �H  B���    A�CQ      �H  ���=    A�Cx      �H  2���     A�C[      �H  2���    A�CK      I  "���    A�CL      <I  ����   A�C�    \I  ~���|    A�Cw     |I  x���    A�CX      �I  v���+    A�Cf      �I  ����g    A�Cb     �I  ����    A�CZ      �I  ����    A�CH      J  :���7    A�Cr      <J  R���-    A�Ch      \J  `���+    A�Cf       |J  l���K   A�CE�A     �J  ����G   A�CB    �J  ����   A�C    �J  ����X   A�CS     K  ����    A�CZ       K  ����    A�CZ      @K  ����    A�CZ      `K  ����    A�CZ       �K  ����    A�CZ          �K  ����    A�CJ      �K  �����    A�C�     �K  �����    A�C�     L  ����    A�C�     $L  �����    A�C�     DL  ����   A�C    dL  �����    A�C�     �L   ����    A�C�     �L  �����    A�C�     �L  �����    A�C�     �L  &����    A�C�     M  �����    A�C�     $M  Z����    A�C�     DM  �����    A�C�     dM  ����    A�CH      �M  x���(    A�Cc      �M  ����C    A�C~      �M  ����    A�CZ      �M  ����!    A�C          N  ����   A�C    $N  ����   A�C    DN  ~���)    A�Cd      dN  ����    A�CF      �N  t���)    A�Cd      �N  ~���(    A�Cc      �N  ����,    A�Cg      �N  ����4    A�Co      O  ����E    A�C@     $O  ����C    A�C~      DO  ����&    A�Ca      dO  ����*    A�Ce      �O  ����J    A�CE     �O  (����    A�C�     �O  �����    A�C�     �O  U���U    A�CP     P  �����   A�C�    $P  
����    A�C�     DP  ����J    A�CE     dP  ����    A�CU      �P  ����f    A�Ca     �P  ���J    A�CE     �P  2���.    A�Ci      �P  @���)    A�Cd      Q  I���E    A�C@     $Q  n���}    A�Cx     DQ  �����    A�C�     dQ  J���W    A�CR     �Q  �����   A�C�    �Q  
����    A�C�     �Q  �����    A�C�     �Q  ����+    A�Cf      R  ����/    A�Cj      $R  �����   A�C�    DR  "����   A�C�    dR  ����m    A�Ch     �R  ���T    A�CO     �R  L���?    A�Cz      �R  l���    A�CU      �R  f���n    A�Ci     S  ����   A�C    $S  ����    A�Cz     DS  ����    A�C|     dS  p����   A�C�    �S  D����    A�C�     �S  ����u    A�Cp     �S  B���E    A�C@     �S  h���    A�CL      T  Z����    A�C�     $T  ����h    A�Cc     DT  ����    A�C�     dT  ����U    A�CP     �T  &���U    A�CP     �T  \���E    A�C@     �T  ����    A�CF      �T  n����    A�C�     U  7���4    A�Co      $U  K���    A�CU      DU  F���*    A�Ce      dU  P���    A�CZ      �U  P���    A�CL      �U  A���Q   A�CL    �U  r���*    A�Ce      �U  |���    A�CZ      V  |���    A�CL      $V  m����    A�C�     DV  �����    A�C|     dV  K���r    A�Cm     �V  ����i    A�Cd     �V  ����I    A�CD     �V  ���    A�CU      �V  	���   A�C    W  ���R    A�CM     $W  4���B    A�C}      DW  V���5    A�Cp      dW  ����"    A�C]      �W  ����*    A�Ce       �W  �����   A�CE��     �W   ��a    A�C\      �W  ^ ���   A�CE��     X  ��3    A�Cn      ,X  .��#    A�C^      LX  2��(    A�Cc      lX  :��2    A�Cm      �X  L��    A�CL      �X  =��G    A�CB     �X  ���    A�CI   $   �X  �����    A�CI���v      Y  M���    A�CI   $   4Y  ;����    A�CI���v      \Y  ���    A�CI      |Y  ���0    A�Ck      �Y  ���    A�CL      �Y  ���    A�CU      �Y  ���"    A�C]      �Y  ���0    A�Ck       Z  ���<   A�CE�2     @Z  ���    A�CU      `Z  ���    A�CU      �Z  ���    A�CI      �Z  ���-    A�Ch      �Z  ���+    A�Cf      �Z  ����    A�C�       [  ����    A�CP          $[  ���R    A�CM     D[  ���R    A�CM     d[  ��N    A�CI     �[  1��E    A�C@     �[  V��    A�CW      �[  R��A    A�C|      �[  s��    A�CF                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           E@     ]=@     ��A     ��������        ��������                        Z�A     ��A     ��A      �A     H�A     \�A                                     �A     �A     �A     �A                     6�A     d�A     *�A     ��A     ,�A      �A     v�A     ��A                                     �A     �A     �A     �A     �A     �A                                                    1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `   C     �C     �C     hC     GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             M@           Z@     I       �@     2       �@     -       @            @     "       8@     -      f@     "       �@     �       V@     �       �@     8                       ,    �       @"@     �                       ,           �%@     o                      ,    *       l'@     �                       ,    �       �'@     >                       ,    �       /(@     @                       ,    r       o(@     [                      ,    �       �)@     �                      �   b       O+@     #      r=@             �=@     �       @>@     �      @@            "@@     \       ~@@     �       A@            2A@     6       hA@     Q       �A@            �A@     B       B@            $B@            �B@     �       �C@     #       �C@            �C@     V       6D@     M      �F@     L      �H@           �J@     )       K@            "K@     )       LK@     ,       xK@     )       �K@     h      
O@     �      �S@     #      �U@     +       V@            V@             V@     4       TV@     E       �V@     &       �V@     E       W@     2       8W@     '       `W@     �       (X@     �       �X@     O       4Y@            JY@     I       �Y@     �       �Z@     �       D[@     X       �[@     D      �\@     �       �]@     L        ^@     �       �^@     *       �^@     }       d_@            u_@            �_@            �_@     a      b@            2b@     �      �d@            �d@     j       :e@     (       be@            �e@     7      �f@            �f@     7      h@     a      oj@            �j@     �      m@     d       ~m@     j       �m@     7       o@     7      Xp@     K       �p@     �       uq@     �       r@            *r@            Hr@     1       zr@     �      =x@            Zx@     H       �x@            �x@            �x@     V      8|@            N|@     H       �|@            �|@     1       �|@     �      ��@            Ƃ@     V      �@     W       s�@     1       ��@     �      D�@     �      �@            �@            �@     �      ��@     �      B�@     1       s�@     �      �@     (       D�@     �                       \   �s       ��@           "@@     \       A@            �@           �@     0       �C@     #       �C@            @�@     R       ��@            �J@     )       K@            "K@     )       LK@     ,       V@            V@             V@     4       TV@     E       �V@     &       �^@     *       �p@     �                       |   v�       �@     <	      hA@     Q       �A@            �A@     B       B@            @@            "@@     \       ~@@     �       A@            2A@     6       N�@     *       $B@            �B@     �       �C@     #       �C@            �C@     V       @�@     R       x�@     S       �J@     )       K@            "K@     )       ̨@            ި@            �@     6       LK@     ,       &�@     r       ��@            ��@     >       ֩@     F       �@            .�@     4       b�@     w       ڪ@     �       `�@     !       ��@     %       ��@            ��@            ˫@     O       �@     I       V@            V@             V@     4       TV@     E       c�@     I       �V@     &       ��@     *       �K@     h      ֬@           �^@     *       ٭@           W@     2       8W@     '       `W@     �       (X@     �       �X@     O       4Y@            JY@     I       �Y@     �       
O@     �      �p@     �       D�@     �       ߯@     N       d_@            �]@     L       u_@            �_@            �_@     a      b@            2b@     �      �d@            �d@     j       :e@     (       be@            �e@     7      �f@            �f@     7      �Z@     �       D[@     X       �[@     D      �\@     �        ^@     �       -�@     J       r@            *r@            Hr@     1       zr@     �      =x@            Zx@     H       �x@            �x@            �x@     V      8|@            oj@            N|@     H       �|@            h@     a      �j@     �      m@     d       ~m@     j       �m@     7       o@     7      Xp@     K       w�@     �       s�@     1       ��@     �      D�@     �      �@            �@            ��@            �|@     1       �@     �      ��@     �      �|@     �      Ƃ@     V      �@     U       B�@     1       h�@     �      �@     (                           ��                       �   �       �@     /;      hA@     Q       �A@            �A@     B       B@            @@            "@@     \       ~@@     �       A@            2A@     6       N�@     *       8�@     &       ^�@     H       ��@     e       �@     M       Z�@     &       ��@     <       ��@     g       $�@     c       ��@     6       ��@     Q       �@     S       d�@     O       ��@     .       ��@     	      ��@     L       8�@     S       ��@     O       $B@            �B@     �       �C@     #       �C@            ��@            �C@     V       �U@     +       ��@     *       �@     �      ��@     *       �@     �      �A     +       A     *       0A     �      
O@     �      �J@     )       K@            "K@     )       �@     6       LK@     ,       �A     *       &	A     �      V@            V@            �A            A     1       4A     )       ^A     N       �A     )       �A     N       $A     �      �A     1       .A     )       XA     �      0A     1       bA     )       �A     �      W@     2       8W@     '       JY@     I       �Z@     �       D[@     X       �X@     O       �[@     D      �\@     �       �]@     L       �Y@     �        ^@     �        V@     4       TV@     E       c�@     I       �V@     &       dA     1       �A     )       �A     �      �!A     �       �"A            �"A     ;       �"A     x      V)A     �       0*A     �       +A     �       �+A     �       �,A     �       �-A     �       f.A     �      6A     d       �6A     *       �6A     x      "=A     �       �=A     �       �>A     �       �?A     �       �@A     �       \AA     �       2BA     �      �IA     d       KJA     x      �PA     �       �QA     �       tRA     �       NSA     �       $TA     �       �TA     �       �UA     �      �]A     d       d_@            be@            �f@            h@     a      oj@            �j@     �      �d@            m@     d       4Y@            ~m@     j       :e@     (       u_@            �m@     7      �_@             o@     7      �d@     j       �e@     7      �f@     7      Xp@     K       �^@     *       ٭@           �]A     x      fdA     �       @eA     �       fA     �       �fA     �       �gA     �       �hA     �       viA     �      +qA     d       �qA     J       �qA            �qA     J       4rA     W       @�@     R       ި@            �rA     Y       �rA            �rA     �       �sA     U       �sA     W       CtA     G       �tA     W       �tA     �       �uA     U       �uA     W       ,vA     W       �vA     �       "wA     U       wwA     W       8|@            �|@            �|@     1       �|@     �      ��@            N|@     H       �x@            �x@            Ƃ@     V      r@            b@            Zx@     H       *r@            �x@     V      �p@     �       D�@     �       ߯@     N       �wA     W       %xA     �       �xA     U       yA     W       pyA     �      {A     �      �|A     �      _~A     �      �A     J       Q�A     �      ��A     �      ��A     �      @�A     �      �A     �      ��A     �      8�A     �      ׋A     �      B�@     1       �@     �      ��@     �      �@            �@            =x@            Hr@     1       ��@     �      D�@     �      -�@     J       �A     �      '�A     �      ϐA     �      n�A     �      �@     (       �A     �       w�@     �       ��A     �       �@     U       h�@     �      J�A     �                      ,    ��      ޖA     �                         ��      ��A           hA@     Q       �A@            �A@     B       B@            @@            $B@            �B@     �       ��A            ��A     P       �A            ��A     �       ��A            ��A     *       ʧA     .       ��A     >       6�A           
O@     �      J�A     0       �K@     h      W@     2       8W@     '       JY@     I       �Z@     �       D[@     X       �X@     O       �[@     D      �\@     �       �]@     L       �Y@     �        ^@     �       `W@     �       (X@     �       4Y@            d_@            be@            �f@            h@     a      oj@            �j@     �      �d@            m@     d       ~m@     j       :e@     (       u_@            �m@     7      �_@             o@     7      �d@     j       �e@     7      �f@     7      Xp@     K       �_@     a      b@            2b@     �      8|@            �|@            �|@     1       �|@     �      ��@            N|@     H       �x@            �x@            Ƃ@     V      r@            Zx@     H       *r@            �x@     V      Hr@     1       zr@     �      =x@            B�@     1       �@     �      ��@     �      �@            �@            ��@     �      D�@     �      s�@     1                       ,    t�      z�A     �                       ,   h�      Z�A     @      @@            ��A            ��A     ,       ܫA            �A            ��A     P       H�A            V�A            h�A     %       ��A     {       
�A     $       .�A     7       e�A     
       p�A            ��A     $       ��A                            L   �      ��A     �       ��A     =       ڮA             ��A            
�A            �A     �      ��A     |       "�A     7       Z�A     -       ��A     +       ��A     K       �A     G      H�A           \�A     X      ��A            ԶA            ��A            �A            4�A                            �   9)      T�A     s      @@            "@@     \       ~@@     �       A@            �C@     #       �C@            �C@     V       �J@     )       K@            "K@     )       LK@     ,       ��A     (       V@            V@             V@     4       TV@     E       �V@     &       ��A     C       �^@     *       -�@     J       �p@     �       w�@     �       �@     U       h�@     �      �@     (       D�@     �                       ,    A      4�A     A                       �   �G      u�A           @@            "@@     \       ~@@     �       A@            �C@     #       �C@            �C@     V       ��A     )       ��A            ��A     )       ��A     (       �A     ,       �J@     )       K@            "K@     )       ��A     (       LK@     ,       V@            V@            B�A     4       v�A     E       ��A     C       ��A     &        V@     4       TV@     E       ��A     C       �V@     &       $�A     *       N�A     J       �^@     *       -�@     J       ��A     �       i�A     �       �p@     �       w�@     �       �A     U       �@     U       Z�A     �      h�@     �      �@     (       ��A     �       D�@     �                       �   &d      ��A     B      @@            "@@     \       ~@@     �       A@            2A@     6       �C@     #       �C@            �C@     V       ��A     )       ��A            ��A     )       ��A     )       �A     ,       V@            V@            B�A     4       v�A     E       �A     E       ��A     &       $�A     *       ^�A     }       ��A     �       ��A     �       z�A     W       ��A     �      �@     (       ��A     �                       <   �x      z�A     M      @@            "@@     \       ~@@     �       A@            hA@     Q       �A@            �A@     B       B@            $B@            �B@     �       �C@     #       �C@            �C@     V       ��A     "       ��A     *       �A     �      �J@     )       K@            "K@     )       LK@     ,       �K@     h      ��A     a       �A     �      ��A     )       ��A            ��A     )       �A     ,       �A     +       �U@     +       
O@     �      ��A     3       &�A     #       J�A     (       r�A     2       ��A            �6A     *       ��A     G       �"A            V@            V@            ��A            
�A     0       :�A            L�A             V@     4       TV@     E       �V@     &       W@     2       8W@     '       `W@     �       (X@     �       �X@     O       4Y@            JY@     I       �Y@     �       B�A     4       v�A     E       ��A     &       �Z@     �       D[@     X       �[@     D      �\@     �       �]@     L        ^@     �       f�A     "       ��A     0       CtA     G       ��A     <      ��A            �A            �^@     *       d_@            u_@            �_@            �_@     a      b@            2b@     �      �d@            �d@     j       :e@     (       be@            �e@     7      �f@            �f@     7      $�A     *       h@     a      oj@            �j@     �      m@     d       ~m@     j       �m@     7       o@     7      Xp@     K       �A     J       (�A            �p@     �       r@            *r@            Hr@     1       zr@     �      =x@            Zx@     H       �x@            �x@            �x@     V      8|@            N|@     H       �|@            ��A     �       �|@     1       �|@     �      ��@            Ƃ@     V      �A     �       s�@     1       ��@     �      D�@     �      �@            �@            �@     �      ��@     �      B�@     1       ��A     �       h�@     �      J�A     �      �@     (       D�@     �       6�A     -       d�A     +                       ,    O�      ��A     �                                      �       �  �  �                    5   �  �  H   �  �  [   2N  :  n   -N    	�   �  �  *  �   int �   1    �n   �  u   N  �   �  )   \  <   M  O   Q   b   %   4�   ^  
P  K.  �    `  �   bpp �   �  �   
 ~    ��  �n   	,  �  ^  �  (	�  x 	�    y 		�   K.  	�   `  	�   �  	�   �  	
�   u 		�  x  	

�     
�   V  	  �  '  x 	�    y �    �  	  '  �  r  r �    g �   b �   a �    g  8  "�  �  �  #�     $�   �(  %�   �   &�   
 �  �  n    �  �  '~  ()�  �    *�    K.  +
�   `  ,
�   �   -�   bpp .�   �  /�     0�   �  1
�     2
�   x  3�    �  4�   $ �  5�  �  L  �   
h  
�  |�  /  x �    y �   K.  �   `  �   �  �   Z   /  �  �   l�  �  t  �  (  �    �  ?  n   _   �  !�  @�  �  �      	\  �   #	\      &	\  �  )	\   P  ,	\  (�  -	\  0  2�   8>  5�   < 
�    8"K  @  K�  
�  )  L�  �   M�  (�   Y  �   �    2  �   msg �   �  �   �  �     �   
  �   u  n    �  e  	�C     �  �=�  �  >�   �  ??  pos @'  ��  A�  � oF  fb D
�  	 C     �  EP  	(C     �  F�  	@C     �   %  n    �  H  	hC     Q  I'  	�C        J�  	kC     )  K�  	lC     �   L'  	pC     �  N�  	�C     �  P�  	xC     �  U\  	�C     �  W
�   	�C     �   X
�   	�C       Z�   	�C     �  \
�   	�C     $  ]
�   	�C       kr  	�C     k  l�  	�C     �  n�   	�C     L  H	  [  `   �  �  H	   Z  8  �  �  H	  �    >  !�  �  �  H	      */   �    H	  S	   m  ;�    (  H	  S	   p  L  S	  A  L  H	  [    9  P�  S	  e  p  H	  [    .  Z�  �  �  H	  [   S	   �  d�  �   �  �  H	   �  hM  S	  �  �  H	  [    n  }  S	  �  �  H	   �  ��  S	  	  	  H	   q  ��	   $  ��	  num �[   T S	   
�  H	  
�  G  �	      	�	   �  
�	  obj S	  D  /  �	  �	  �	   T S	   
Y	  �	  �  o�  	�C     �  pS	  	C     �  h  �  E@            ��  
  6
  �  N	     �    !�2  �	    "
  �  Y
  �@     8       ��
  #
  �X$'
  p
  %(
   &'
  �@     )       '(
  �h  (y   @     >       ��
  )>  m�   �l)u  m�   �h *L  �
  V@     �       �4  +�  N	  �X,pos P[   �T-� S�	  �h.�@     8       /i U[   �d  0�  S  �@     �       �~  +�  N	  �H,obj *S	  �@-�2  +�	  �X 1�	  �  �  �  �	   2~  3  �  f@     "       ��  #�  �h 0�  �  8@     -      �b  +�  N	  �H,pos h[   �D-� n�	  �h/obj rS	  �X3^@     	       B  -!Z  jS	  �P .r@     8       /i p[   �d  0(  �  @     "       ��  +�  N	  �h,pos L[   �d *�  �  @            ��  +�  N	  �h �  �  �  �  N	   2�      �@     -       �  #�  �h 4�  ��   �
@     A
      ��  -�  ��  �P-x  ��   �L-[  ��   ��-�  ��  �@-[  ��  ��-�  ��   ��..@     �      5msg @Y  ��~6!Z  _   ��3|@     7         /i ��   �l.�@            /win �S	  ��  3�@     
      �  5i �   �h.�@     �      5win S	  ��.�@     �       6I  Y  ��~6`  �   �d6z  �   �`   3�@     �       �  6I  .Y  ��~6`  0�   �\6z  1�   �X .%@     �       6�  EY  ��~   
�  �    n    7�  ��  @     �      �S  ,win �S	  ��-w  �'  �� 7�  �e   @     �      �(  -�  ��   �L.[@     �      /j �
�   �l.q@     �      -{  ��  �k-�  �?  ��~-�  ��  �X3�@     D         /i ��   �d .
@     �       /win �S	  �P    7  r�  @           ��  -�  s�   �T.S@     �       /i v
�   �l.r@     �       -{  w	�  �k.v@     }       /j x�   �d.�@     e       -�  y?  ��~-�  z�  �X     
?  �  1      �  �   2�  d  3  �@     2       �<  #  �h 7�  _�  M@     �       �n  -e  a�   �h 8�  g  '  Z@     I       ��  ,l 0�  �h,r E�  �` 93   N    k  @"@     0#@     5  src/gfx/sse2.asm NASM 2.14.02 �@"@                 �  i	  �  	  �%@     o      �  �  �  �  G   2N  :  Z   -N  �  �  int 1  M  ;   Q   N   ��  �Z   ,  �  ]	  v   ;	  ��   c	  }    �3  �   8  }   �       Z    �  	   �	  �   
�  !o   ,'@     @       �v  fd !o   �\��  !$�   �PA	  !;v  �Hret "�   �h   
�	  �   �&@     A       ��  fd o   �\�    �   �P�	  ,o   �Xret �   �h 
�	  o   �&@     ?       �8  fd o   �\u %8  �P��  4�   �Hret 	o   �l >  
�	  o   m&@     ?       ��  fd o   �\u �  �P��  -�   �Hret 	o   �l Q	  7&@     6       ��  fd o   �l 
�	  o   �%@     :       �  H	    �X�  *o   �Tfd 	o   �l    �   |  i	  
  	  l'@     �       n  �  �  2N  :  N   -N  �  �  int 1  Q   B   (	�   �   q    2  q   msg q   �  q   �  q     �   }   �	  
�'@     M       �<  	pid 
q   �H	msg 
.�   � 
m q   �h�  q   �`�  q   �X �	  
q   l'@     8       �}  	msg (}  �X
  q   �h �    �    \  i	  N
  	  �'@     >       W  �  �  2N  :  N   -N  �  �  int 1  Q   B   2
  �'@     >       �5
  q   �`:
  &q   �X?
  5q   �PD
  Dq   �Hq
  Sq   �@I
  bq   ��  �    �  i	  v
  	  /(@     @       	    9   �  �  2N  -N  �  �  int 1  �  -   �
  
�   /(@     @       ��   ^  �  &�   �Xptr �   �h 	q   	�    `   K  i	  �
  	  o(@     [      �  �  �  2N  -N  �  �  int 1  �
  �   �(@     �       ��   num ^   �Xstr �   �P.�  %W   �Li W   �lG)@     U       rem &W   �h  	�   �  
�
  o(@     �       �str �   �H��  W   �Dc W   �ld 
�   �`end �   �X!Z  �   �W  �     	  �
  	  �)@     �      �  ��  �9   -N  �
   -   +@     <       ��   s  �   �Xlen !	-   �h#+@     &       i "-   �`  �   �  	�   ��  a  j*@     �       �a  
��  a  �Hsrc 'h  �@
  3-   ��q  t  �X�
  t  �P�*@     4       A  i -   �h �*@     E       i -   �`  a  s  h  �   W�  a  *@     Z       �  
��  c  �Hsrc <n  �@
  H-   ��q  t  �`�
  t  �X0*@     4       i -   �h  ��  a  �)@     F       ��  
��  a  �Xc �  �T
  (-   �Hq  t  �`�)@     )       i -   �h  int  hW   �  c	  
c  	  P          �  ?  5   dint 5   ?�3  M   S   �  S   ?�Q  M   �  k   �  '�  �   2N  �   -N  �   �  �  1  '  ��   'M  ~   �   '%   4�   �   '��  ��   �   '  	  e  @�-  1  �R  5    /rem 5    '�-  	  @�6  e  �R  �    /rem �    '�6  =  @'  �  �R  �   /rem �   ,  ''  q  ffrg h  gg  �	�  On <   pOm <   �P�Z  �   ߰�hmsb �      �P(  �   ���g  A  '  -  �   �!  �W  A  L  �  �    )�R  �n  �   d  j  �   i_st >�   jJa  ?5   �	 AI  �  Q�\   �  6�V  5   ,�  "�6   "�  Rhex  S4D    k0  {#  l�2  |5   0  ~m[      �   B/   .    �  5     �=  �g  8  >  �   �=    S  ^  �  �   �=  4H  s  ~  �  �   �=  �?  �  �  �  �   �=  *�l  �  �  �  �   �=  0]  �  �  �     �=  8�7  �  �  �  5    #�#  = A  
    "  �  �   #fF  Q�1    ;  A     #fF  T�6    Z  `  �   #\?  X�:    y       #�"  \iQ  �  �  �     #�"  `�:  "  �  �  �   #2d  dF  (  �  �  �   ;W  ��  �  �  �   ~  ��   �6  �  T 5    �  4.  2  4.  3�*  >  D  .   )�(  6UB    \  g  .  �   �(  <�   C.  =5   .]  >�  E0  ?  �e  @  �  A  �_  B  rO  C  m3.  BW  �  �  .  5    n4.  �%  �  .  �T      C�  J�  7�0  N�;  W  P   T �   �   �     5   5   5   S    7�  x8  �  P   T �   �   �   5   5   5   S    o6  ��  T �   F   �     �     A~6  

�  Q�  
�  g&  
�  6a  
E ?  �    �      �  �
	|  �  
�2  &  1  �   �    ,�  
?N  E  P  �   �    -�#  
	�*  �   h  s  �   �    �  
Pl  �  �  �   5    )Y4  
"	�c  �   �  �  �   �   R0  
',;  �  �  �   S    R0  
1u?  �  �  �   �   1Ba  
>�    1t 
?Y   1�\  
@
�   �18]  
A  �)�  
	V  �   J  U  T   �      T�5  
	9+  �   p  T �  �   �      )�R  
H $    �  �  �    �0  
MY  �  �  �   �   1�V  
Q   8�    p�-  �   � U   A#  	�  q�i  �   C}C  	�  D!	  V]I      E	  6�-  5   N	  "�6   Rred "�C   �Q  0
  �Q  �+  o	  u	  �   ,�Q  �*  �	  �	  �  �   -�#  �_  �  �	  �	  �  �   �N     �R    �7    \.     >*  !   �R  ")	  ( N	  �R  %W
  7^  '
     9
  T K  �    W�  '�V    T v  �     BD  5�  Xh 8�_  �  }
  �    �N  =j4  �   �
  �    �R  B�i  �   �
  �    �7  E�N  �   �
  �    \.  I�P  �   �
  �    >*  L�  �   �
  �    )  P�,  �       !   9�+  U}O    8  �    9\G  Z�"    S  �    �G  dma  g  m  !   ,�G  g"  �  �  !  !   -�#  i  !  �  �  !  !   )Rr  o_L  �   �  �  !   �(  |�^  �  �  !  �    �e  ��      !  �   �    i  ��=  '  7  !  �   �    �+  ��B  L  W  !  �    $�l  �0  l  w  !  �    %�2  .A  �  �  !  �   �    %Q:  D�  �  �  !  �   �    %�l  xm  �  �  !  �    %�R  ��6  �    !  �    %�  +    &  !  �    $�  �   ;  F  !  �    $�_  #=M  [  f  !  �    3�1  0Z$    �  �  !   3�1  9mI    �  �  !  �   "  !  !   :  �   D �  T v  ;E3  UW  A 
   W
  r�'  ��  &��  &��  &�  &��
  &��
  &��
  FW
   $�b  �@  M  X  .!     $�+  ��m  m  x  .!  �    :�5  �  T v  ;E3  UW  L   A 
   �S  59  Xh 88Y  �  �  �    �N  =�!  �   �  �    �R  BbJ  �     �    �7  E�h  �     �    \.  If  �   5  �    >*  LV/  �   O  �    )  P�[  �   g  m  9!   9�+  U9    �  �    9\G  Z-    �  �    �G  d3<  �  �  9!   ,�G  gn.  �  �  9!  D!   -�#  itF  J!  �  �  9!  D!   )Rr  o�+  �       9!   �(  |�j  2  =  9!  �    �e  �jK  R  b  9!  �   �    i  �A]  w  �  9!  �   �    �+  �6  �  �  9!  �    $�l    �  �  9!  �    %�2  H)  �  �  9!  �   �    %Q:  D�      9!  �   �    %�l  x.8  )  4  9!  �    %�R  �Ld  J  U  9!  �    %�  �  k  v  9!  �    $�  �R  �  �  9!  �    $�_  #	g  �  �  9!  �    3�1  0    �  �  9!   3�1  9�    �  
  9!  �   "  P!  P!   :  �   D >  T K  ;E3  `W  XA 
   �  sX  �&�  &�=  &�b  &��  &�  &�O  F�   $�b  �R%  �  �  V!     $�+  ��  �  �  V!  �    :�5  �  T K  ;E3  `W  XL   A 
    D  V]I      E�  2l  >  tclz �  5   6  �    T �    u%B  �$�  6L3  5   �q  "�6   "�i  "'   L   8  H�	F   8  ��Q  �  �  �   L  �   �    , 8  �&  �  �  �   �    -�#  �
[  �   �  �  �   �    )qe  �ze        �      8  �q   v6  ��   ��  ��   �  ��   v  8  ��	�  Fv   8  �i'  r  �  �   �   �   5    ,8  �E2  �  �  �   �    -�#  ��G  �   �  �  �   �    ��  �<   H�(  ��   L�-  ��   P+  ��  X K  �>  �	z  �>  �Q*  $  *  �    ,�>  �0o  >  I  �   "   -�#  ��>  "  a  l  �   "   �+  ��       �5  �	�  T�R  ��3    �  #!  �   �        �	     �'  �  �  a!   ,+  �	�   �Q  ��   �G  �    '�b  ��  C%  ��Z  !  ,  g!  r!   #N�  �YV    E  P  g!  �    3�&  H
:    j  z  g!    �    %��  z�W  �  �  g!     %Q.  �]  �  �  g!    �    #�:  -	�c  �   �  �  g!   v�\  :�!                         @       G�Z  < �   GkG  = �    =d  D�\  �   D  �      S  �   ^  �    G�&  f<   4�  h�   Oa  k�    �  �    4�e  x�   4�&  {�   w]  ��    H�i  ��U  �   �  �  g!  �    H�i  �C  �   �    g!  5    H'  !�C  �     (  g!  �    $�  3  =  C  g!   $�@  :�5  X  c  g!  �    �=  �
r!   �  ��  '8  ��  +2  �}  �  �	�    Y  ��!  (8�^  �  8D=  �   I�Z  �+N	  IA)  �7>  IA)  �7�  S�Z  x  �c  �l      �!   �c  w  '  7  �!  �  �   �c  =  L  W  �!  �   x�c  !zG  l  w  �!  �!   �c  #�  �  �  �!  �!   �c  (�;  �  �  �!  5    #�#  -4  "  �  �  �!  �   �c  2�n  �  �  �!   a  8p;      �!   #S  >�&    *  0  �!   #+H  BY0    I  T  �!  �   �  G	�   R  H  8D=  �   �  l?  
CI  �  �  T 5   �  �   7�H  �J=  �  F   �    �    7�H  ��(  �  F   �    �    Yb:  2�2    T   F   �8  �    Y�k  2:c  E  T �  F   -9  �    W�Q  
!I  f:  T �   f:  f:    y�  �  *�m  �  *�  �  *lP  �  *H    �  �  �   �  z�   o �  {L  J�  	��A     Z   �  <�  �  �  �  �  <   K5     K�  �  oF      5   5     .  |std  �  �   Jq  4`?  K  T 5   Z�-  [�    �1  J�  4`?  K  T 5   Z�-  [    \@  Nh    \@  NW3     ]�#  Q  ]�?  ~  (N  �  <�  �+  �  �  }J�  	��A     Cde  �  P  [  ~P  
�-  9  ?  �   B�R  �  O  �  �    ^B  +|  �  ^'.  ,�R  �  6�^  5   �  "�6   "�j  "�  "$D  "�7   �  �  /it �   /end �  _fF  Hh    �  �  <    C Z    �7  D  /it H    /end �  _fF  �&    6  <  S    C �   �_  	
  �  j  T �  �  �>   ,R  	
�"  �?  �  T �?  �  �>   I4  	
�e  �@  �  T �@  �  �>   U�     5�  5	  N	  �  
  N	  5�  ^P  �  ^P  �b  	    �   ,^P  �#  #  .  �  �   -�#  PK  �  F  Q  �  �   �c  �!  e  k  �   a  �l    �  �   1je  5     �  �  �  �  �  �-     map �7  �   �  �     �    B�@   H  �     �   �     �  ��  <   �_  �    �f  �     �    �  �   �  <H   �  S   i   �    D|   ��-      Ei   Jn   
        ��>  ��  	 C     �  �     �   |    v  �   F  v  K  �   �  K    �   W
  !  �  W
  �     #!  �  .!  �  9!  9  �  �   >  V!  �  >  g!  �  �   �!  �    x!  *eW  �  *�i    *�    *Gb  ^  `'  l   �`Q5  �   ��:  �     *L  �  �  �!  �    �  �!  x  K�  �  z    5�  5�  �NH  ]=@            ��y   .=@     /       �v"  >  �5   �lu  �5   �h 
�  �"  D�@     �       ��"  �  �   �hs 
'S   �d .}  �@     (       ��"  T 5   a �  �hb #�  �`   s�@     �      �$  P   T �   ��  N�   ��^W  N$�   ��H*  N1  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#S   ��~�  P�  �Xu S$  ��	k T5   �� l�@     E       �#  	i a5   �l  ��@     -       �#  	i d5   �h �@     0       	i f5   �d  S   ($  �    �  B�@     1       �S$  �2  Z�   �h 
U  r$  ��@     �      ��$  �  ?!  ��n �   ��u �   �Xv �   �Pw �   �H 
4  �$  �@     �      �%  �  ?!  ��n ��   ��u ��   �Xv ��   �Pw ��   �H .
  �@            �Q%  T K  �2  '�   �h .9
  �@            ��%  T v  �2  '�   �h 
  �%  D�@     �      ��%  �  !  ��n �   ��u �   �Xv �   �Pw �   �H 
�  &  ��@     �      �O&  �  !  ��n ��   ��u ��   �Xv ��   �Pw ��   �H 8  s�@     1       �z&  �2  Z�   �h W  �@     W       �'  P   T �   ��  x�   �h^W  x!�   �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yS   �P���  {	�     
7  -'  Ƃ@     V      �e'  �  !  �Xn ��   �P�N  ��   �hd4  ��   �` �  ��@            ��'  �  =�   �h 
  �'  �|@     �      ��(  �  ?!  ��n x�   ���N  {�   �Ps ��   �X�R  �)	  �� �}@     �       (  x ��   �H  �~@     z       B(  x ��   �@  w�@     Q       i(  f?  ��   �� Ɓ@     Q       f?  ��   ��  m  �|@     1       ��(  �2  U�   �h 5  �|@            ��(  �  L�   �h 
�  )  N|@     H       �/)  �  ?!  �X�2  #�   �P� $�   �h .�  8|@            �Z)  �  8�   �h 
�  y)  �x@     V      ��)  �  ?!  �Xn ��   �P�N  ��   �hd4  ��   �` 
v  �)  �x@            ��)  �  ?!  �h�2  �   �` 
&  *  �x@            �)*  �  !  �h�2  �   �` 
F  H*  Zx@     H       �u*  �  !  �X�2  #�   �P� $�   �h }
  =x@            ��*  �  =�   �h 
�  �*  zr@     �      ��+  �  !  ��n x�   ���N  {�   �Ps ��   �X�R  �)	  �� Is@     �       .+  x ��   �H  et@     z       R+  x ��   �@  v@     Q       y+  f?  ��   �� Zw@     Q       f?  ��   ��    Hr@     1       ��+  �2  U�   �h �
  *r@            ��+  �  L�   �h .d
  r@            �,  �  8�   �h �  uq@     �       �u,  T �   F   �2  ��   �hfo �/  �`��  �6�   �X 
�  �,  �p@     �       ��,  �  �   �hstr 
1�  �` �  �,  �,  �  �   +�"  �L  +�  �%�   +&8  �6�    (�,  ;R  -  Xp@     K       �0-  �,  �h�,  �d�,  �X�,  �P 
  O-   o@     7      ��-  �  !  �H�N  ��   �@�2  �"�   ��72  ��   �X 
�  �-  �m@     7      ��-  �  !  �H�N  ��   �@�2  �!�   ���l  ��   �X 
�  .  ~m@     j       �.  �  !  �h�2  |�   �` ^  -.  [.  �  �   +�  ��   +&8  �)�   +X[  �65    (.  &Z  ~.  m@     d       ��.  -.  �h6.  �`B.  �XN.  �T 
�  �.  �j@     �      �/  �  ?!  ���2  �   ���   �   ���N  �   �X�R  �   �P�7  �   �H   oj@            �I/  �  I�   �h 
�  h/  h@     a      ��/  �  ?!  ���2  D�   ��f?  D$�   ���l  E�   �X72  F�   �P�N  Z�   �H 
b  �/  �f@     7      �"0  �  ?!  �H�N  ��   �@�2  �"�   ��72  ��   �X   �f@            �M0  �  E�   �h 
=  l0  �e@     7      ��0  �  ?!  �H�N  ��   �@�2  �!�   ���l  ��   �X �  be@            ��0  �  B�   �h 0�  �0  :e@     (       �1  �  )!  �ha �!�   �`b �1�   �X 
  71  �d@     j       �S1  �  ?!  �h�2  |�   �` 0O  r1  �d@            �1  �  ?!  �h 
w  �1  2b@     �      ��1  �  !  ���2  �   ���   �   ���N  �   �X�R  �   �P�7  �   �H �
  b@            �)2  �  I�   �h 
�  H2  �_@     a      ��2  �  !  ���2  D�   ��f?  D$�   ���l  E�   �X72  F�   �P�N  Z�   �H �
  �_@            ��2  �  E�   �h �
  u_@            ��2  �  B�   �h 0�
  3  d_@            �*3  �  !  �h �  �^@     }       �}3  F   �2  � �  ��fo �7  ����  �>�   �� �  �^@     *       ��3  F   �2  � �  �hfo �7  �`��  �>�   �X 
  �3   ^@     �       �)4  �  m!  �H  !=�   �@v6  '�   �Xfra )�   �P 
�  H4  �]@     L       �U4  �  �!  �h 
X  t4  �\@     �       ��4  �  4!  �X�2  ��   �P� ��   �h 
�  �4  �[@     D      �v5  �  m!  ����  95   ��v6  �   �@�  	�   ���H  
	�   �Xslb �   ��Rr  �   �Pk\@     ^       off �   �H�\@     >       �2  �   ��   
�  �5  D[@     X       ��5  �  ?!  �X� p�   �h 
�  �5  �Z@     �       �/6  �  ?!  �H�2  �   �@v  �   �h�\  �   �`�Z@     I       �l  �   �X  
�  N6  �Y@     �       �{6  �  \!  �X�2  ��   �P� ��   �h 0�  �6  JY@     I       ��6  �  �   �Xp �  �P	adr �	�   �h   �6  �6  �  !   2�6  �`  �6  4Y@            �7  �6  �h 
�  &7  �X@     O       �37  �  �!  �h 
W  R7  (X@     �       ��7  �  !  �H�2  �   �@v  �   �h�\  �   �`�X@     I       �l  �   �X  
�  �7  `W@     �       ��7  �  m!  �Xv6  �;�   �P� ��   �h �  8  8  �  �!     <    (�7  �  A8  8W@     '       �J8  8  �h 7  X8  n8  �  �!  +�  �   (J8  dh  �8  W@     2       ��8  X8  �ha8  �`   �  �V@     E       ��8  T   F   �2  2�8  �H��  2!�   �@ 
�  9  �V@     &       �-9  �  �   �ha  
M�  �` �    TV@     E       �}9  T �  F   �2  2-9  �H��  2!�   �@   �9  �9  �  �   +Ca  
�    2}9  �n  �9   V@     4       ��9  �9  �h�9  �`   �9  �9  �  �     <    2�9  =e  :  V@            �":  �9  �h �  0:  ::  �  �   2":  �H  ]:  V@            �f:  0:  �h �   .E  �U@     +       ��:  T �   a f:  �hb #f:  �` 
P  �:  �S@     #      ��;  �  m!  ��W H4  ���=  HD�   ��v6  R�   �X�\  T�  ��fra U�   �P �T@     �       o;  slb [�   �H�  \
�   �@Y  a	  �� U@     �       Y  o	  ��  
,  �;  
O@     �      ��<  �  m!  ��~��  �6�   ��~ JO@     �      }<  ��  �5   �\	bkt �a!  �PsZ  ��  ���2  �   �� �O@     *      I<  slb 	�   �H �P@     �      slb 	�   �@�\  �  ��  �R@     �         6�   ��fra 7�   ���\  9�  ��~  
z  �<  �K@     h      ��=  �  m!  ��~W z0  ��~v6  ��   �X�\  ��  ��fra ��   �Pslb ��   �Hbkt �a!  �@�  �	�   ��sZ  ��  ���-  �  ���2  ��   �� 
+  �=  xK@     )       ��=  T   �  �   �h�2  
  �` 
�  �=  LK@     ,       �>  �  �   �h=�  �  
U  2>  "K@     )       �N>  T �  �  �   �h�2  
�  �` s  \>  o>  �  �      <    2N>  'F  �>  K@            ��>  \>  �h 
�  �>  �J@     )       ��>  �  �   �` M   <�>  D  �H@           ��?  T �  str 	
�  ���  	
#�>  ��Lret 	1�J@     �  �?  	 B     H*  	  ���&  	�  �`	dot 	�  ��	end 	�  ��4  	�  ��	tmp 	�  �XM   	d 	"�  �@  Z   �?  �    �?  ^  j  �F@     L      ��@  T �?  str 	
�  ���  	
#�>  ��Lret 	1�H@     �  �?  	�B     H*  	  �[�&  	�?  �l	dot 	�  �P	end 	�  �H4  	�  �@	tmp 	�  �`M�   	d 	"�?  �\  �  �  6D@     M      �sA  T �@  str 	
�  ���  	
#�>  ��Lret 	1NF@     �  �?  	�B     H*  	  �W�&  	�@  �h	dot 	�  �H	end 	�  �@4  	�  ��	tmp 	�  �`M�   	d 	"�@  �X  �  �A  �A  �  �  +�-  *�   (sA  �b  �A  �C@     V       ��A  �A  �h�A  �` �  �A  �A  �  �     <    (�A   Y  B  �C@            �B  �A  �h #  &B  0B  �  �   (B  �@  SB  �C@     #       �\B  &B  �h !<2  ��@  �<@     3       ��B  �  �*�  �h�  �E�>  �`loc �V�   �X�  �B  	�B      Z   �B  �    �B  !�j  �5   2<@     �       �NC  out �NC  �H�j  �'�   �@  �5�   ��p �  �X�  dC  	�B        Z   dC  �    TC  !�&  ~  \;@     �       ��C  ptr ~  ��~  ~!�   ��~�    �h !�1  u  �:@     �       �D    u�   ��~�  v  �h ���  j�9@     �       �6D  ptr j  ��} D  �B@     �       ��D    S0�   ��	tc U�   �`	e ^�   �X	f _�   �P	ip `�   �H	is a�   �@�B@     :       	i W�   �l  .*  $B@            �5E  idx D6�   ��	tc F�   �h	s K5   �d	ip L�   �X	is M�   �P	f N�   �H !�7  d�   �9@     3       ��E  �  dM   �h�h  d<�  �`�7  dN�   �X�  �B  	�B      !=  L�   L8@     =      ��F  wcs LH   ��mbs L+�  ���V  L7�   ��cc M�F  �hst N   �Py�  O�  �@�W  P�  ���  �B  	�B      �8@     N       �F    S
�   ���8@     H       e T{  �d  9@            e Y
{  �`P9@     7       n ]
�   �X   �  !�  G5   8@     .       �(G  �  GM   �hwc G"�  �d�  8G  	B      Z   8G  �    (G  !�R  >5   �6@     1      ��G  wc > N   ��~mbs >;�  ��~�7  >G�   ��~�  8G  	xB      !h.  /5   �5@           �^H  mbs /�  ���Q  /#�   ��cc 0�F  �Xwc 1
�  �Py�  2�  �@�W  3�  ���  nH  	rB     �6@     Z       e :
{  �T  Z   nH  �    ^H  !F  *	�  �5@     /       ��H  ^W  *�  �h�j  *+�  �`�  nH  	lB      !G  &e  �5@     /       �!I  ^W  &�   �h�j  &�   �`�  1I  	gB      Z   1I  �    !I  �div  1  e5@     &       ��I  ^W   5   �\�j   5   �Xr !1  �h !�-  �  :5@     +       ��I  ^W  �  �h�  nH  	aB      !�-  �   5@     +       �J  ^W  �   �h�  1I  	\B      �abs 5   �4@     *       �_J  ^W  5   �l�  oJ  	XB      Z   oJ  �    _J  N�H  ��3@           ��K  .�  �  ����  ��   ��  �-�   ���0  �	�K  ���3@     �       i  �   �h4@     �       u 	  �P4@     �       j �   �`34@     �       v 
  �H	V  
M   �@;I  	
M   ��w4@     V       k 
�   �X�4@     =       !Z  
S   ��       �5   �K  �  �   �K  �@  �  �2@     �       ��L  key ��  ��.�  �,�  ����  �9�   ��  �G�   ���0  �	�K  ��	i �	�   �h	j �	�   �`�  �?  	PB     (3@     |       	k �
�   �X�^  ��  �P	res �5   �L  Z  �M   �2@     +       ��L  =M   �h�  8G  	BB      dG  �5   �2@     +       �2M  �  ��  �h�  8G  	;B      >�Z  �r2@     *       �sM  o6  �5   �l�  �M  	0B      Z   �M  �   
 sM  >4  �]2@            ��M  o6  �5   �l >�Z  �C2@            ��M  o6  �5   �l �Z  �5   2@     +       �)N  �\  �+N  �h�  AN  	 B      �)N  Z   AN  �    1N  ��  �5   �1@     )       �xN  �\  �+N  �h >�#  ��1@     #       ��N  �  nH  	B      �-  �  v1@     V       ��N  ��  ��   �X  �#�   �P	ptr �  �h �=  �  !1@     U       �YO  m  ��   �X  �.�   �P	ptr �  �`	ret �5   �l N�n  ��0@     Z       ��O  =�   ��~ Nga  ��0@     "       ��O  s ��   �l >3  �5   z0@     +       ��O  =B   �h�  8G  	B      �e4  �5   `0@            �vH  ��  50@     +       �ZP  �  �4�  �hend �N�>  �`.�  �W5   �\ �3  [�   �-@     G      �"Q  �  [.�  ���  [F�>  ��.�  [R5   ���V  ]�   �P	s _"Q  �h	acc `�   ��	c a5   �d3c  b�   �H	neg c5   �`	any c5   �\�3  c5   �D r   �  V�  �-@     +       �xQ  �  V*�  �hend VD�>  �`.�  VM5   �\ \  0�   y,@     J      ��Q  �  0$�  �Xend 0>�>  �P.�  0G5   �L�  8G  	B     H*  ;  �o�&  G�   �` �  -�  @,@     9       �:R  �  -,�  �hend -F�>  �` f[  *�?  ,@     %       �{R  �  *%�  �hend *?�>  �` _[  '�@  �+@     3       ��R  �  '&�  �hend '@�>  �` 	4  $�  �+@     $       ��R  �  $�  �h �  !�   �+@     $       � S  �  !�  �h �  5   |+@     $       �RS  �  �  �h �  �@  O+@     -       ��S  �  �  �h 0k  �S  B@            ��S  �  �  �h 
Q  �S  �A@     B       ��S  �  �  �h�  1I  	�B      .  �A@            �T  x )�   �h [	  &T  0T  �  �   2T  �b  ST  hA@     Q       �\T  &T  �h 
D  {T  2A@     6       ��T  �  4  �`c 63�  �\�  7  �h a�  2�T  �T  �  4     <    (�T    �T  A@            ��T  �T  �h   a�  2U  U  �  4  �T   (�T  �  >U  ~@@     �       �OU  U  �hU  �` *  ]U  gU  �  4   (OU  a  �U  "@@     \       ��U  ]U  �h �F  nH    @@            ��U    #�   �hp /  �` 0L  �U  @>@     �      ��V  �  �  �H��   �V  �P	res 3�   �Xk>@     N      	y -�   �\ k>@     {       �V  	kk #5   �l{>@     e       	y $�   �d  �>@     {       	kk (5   �h�>@     e       	y )�   �`    �   �V  �    �V  0-  �V  �=@     �       �W  �  �  �hs �   �d   W  )W  �  �   (W  j  LW  r=@             �UW  W  �h bv  �  "bK  �  " �   Q  	  t  	  �          B  �r  e6   2N  6   �s  	
N   -N  1  ��  �N   ,  �  L  �  �  �  
6   �  �  int �   M  �   ��  �   	�_  �    	�f  �   	  6    
frg 	u  I  �   �\     �V  �   ,;  �6   �  hex  4D  �  0  {�  �2  |�   0  ~m[  u  {  �   /   .  �  �  �     �=  �g  �  �  �   �=    �  �  �  �    �=  4H  �  �  �  �   �=  �?      �  �   �=  *�l  '  2  �  �   �=  0]  G  R  �  �   �=  8�7  g  r  �  �    �#  = A  �  �  �  �  ;   fF  Q�1  �  �  �  �   fF  T�6  �  �  �  �   \?  X�:  �  �  �  �   �"  \iQ  �      �   �"  `�:  �  +  1  �   2d  dF  �  J  P  �   ;W  ��  d  j  �   	~  �H   	�6  ��  T �    ;  4.  2\  4.  3�*  �  �  �   �(  6UB  �  �  �  �     	�(  <   	C.  =�   	.]  >;  	E0  ?�  	�e  @�  	�  A�  	�_  B�  	rO  C�  3.  BW  P  �  �     �  J�q    q  }r  �  �  �	   q  �q  �  �  �	  �   q  �q  �  �  �	  �  \    �  <s  �  �  �  �	   p  "Yq  �	  	    �	  \      &	�o  \   -  3  �	   �r  *r  �  L  W  �	  d   �r  2�p  �  p  {  �	  d   Mr  6	�o  \   �  �  �	  �  \    jr  >	�s  \   �  �  �	  �   �q  F�s  d  �  �  �	  \   \    	V W�   	��  X	\   �s  �   d  ~6  
  �  #  g&    6a  E ?  U  `  "  �	   �  �	�  �  �2  �  �  -  "   �  ?N  �  �  -  8   �#  	�*  >  �  �  -  8   �  Pl  �  �  -  �    Y4  "	�c  >      -     R0  ',;  $  /  -  �   R0  1u?  C  N  -  �    Ba  >"    t ?D   �\  @
\   � 8]  A�  �!�5  	9+  >  �  T �  -  �    `  �R  H $  `  �  �  "   �0  MY  �  �  "  �    �V  Q�	   �  �	  "�-  N   � #   $�H  ��(  >  F `  �  �  >   %�k  2:c  h  T �  F `  $  >   q  [!d   &
  	@B     '�  �  �  �  'H  �  ';  �  (�   )�   (�  );  (;  oF  �  '�  (�   '�   '�  �  *std  �	  �   J0	  +`?  K�  T �   ,�-  -�    �1  J]	  +`?  K�  T �   ,�-  -�    .@  Nh  �  .@  NW3  �   /�#  	  /�?  =	  (N  'd  �	  '  �	  (�  �+  &(  	AB     0de  �  P  
  1P  
�-  �	  
  �   �R  �  
  �  �    2B  +|  4  2'.  ,�R    �^  �   p
  �6   �j  �  $D  �7   �  �
  3it �   3end �  4fF  Hh  �  �
  �
  �   C �   �r    3it �   3end �  4fF  |o  �  �
     �   C 6    a�  q:  !4s  rbp  ?
  )  �  �	  �    r  #�   5�  t  !4s  0s  ?
  c  �  �  �    6�p  "9q  �  :    '�	  'p
  '6   '=   '�
  '  (:  7  86   �}s   �q  0q  r  ;r  p  q  �s  �r  �p  	Hp  
Xr  �r  ks    9��  '4  "  '`  -  (�  (`  :�  T  ;N    <]	  <o	  =/  }  �p@     �       ��  >�  3  �h?str 1�  �` @  �^@     *       ��  F `  A�2  � �  �h?fo �7�  �`A��  �>>  �X =�    �V@     &       �$  >�  (  �hAa  M�  �` (�  @>  TV@     E       �t  T �  F `  B�2  2$  �HB��  2!>  �@ Cm  �  �  D�  3  ECa  "   Ft  �n  �   V@     4       ��  G�  �hG�  �` C{  �  �  D�  �  D   �    F�  =e    V@            �  G�  �h Ca  '  1  D�  �   F  �H  T  V@            �]  G'  �h =�  |  LK@     ,       ��  >�  3  �hH  �  =�  �  "K@     )       ��  T �  >�  3  �hA�2  �  �` C�  �  �  D�  3  D   �    F�  'F    K@            �   G�  �h =�  ?  �J@     )       �L  >�  (  �` I3  k  ��@            ��  >�  �	  �XA�-  *%d  �@JÞ@     G       Ki -\   �h  C�  �  �  D�  �	  Lcs  �   F�  $p  �  @�@     R       ��  G�  �hG�  �` CR      D�  �  D   �    M�   Y  A  �C@            �J  G  �h C�  X  b  D�  �   MJ  �@  �  �C@     #       ��  GX  �h N'q  #)   ڜ@     *       ��  H)   �lO�  �  	�B      :�  �  ;N    �  N�r  )   ��@     *       �!  H)   �lO�  �  	�B      N�p  �   _�@     Q       ��  Pnc �   �\Qcc �  �hQcp :  �`Js�@     &       Qe 
?
  �d  'F  �  N�r  
�   �@     Q       �  Pnc 
�   �\Qcc �  �hQcp :  �`J"�@     &       Qe 
?
  �d  Ntr  �   ��@     .       �U  H)   �lHB   �`O�  �  	�B      Rvr  �
B   �@     �      ��  ?cs ��  ��|Ks �h  ��} R�p  ��   ϗ@     H       �  ?nc �)   �\Kcc ��  �hKcp �:  �`J�@     %       Ke �
?
  �d  R�r  ��   |�@     S       �m  ?nc �)   �\Kcc ��  �hKcp �:  �`J��@     %       Ke �
?
  �d  R�o  ��   )�@     S       ��  ?nc �)   �\Kcc ��  �hKcp �:  �`J=�@     %       Ke �
?
  �d  R�p  ��   ֖@     S       �E  ?nc �)   �\Kcc ��  �hKcp �:  �`J�@     %       Ke �
?
  �d  RQp  ��   ��@     S       ��  ?nc �)   �\Kcc ��  �hKcp �:  �`J��@     %       Ke �
?
  �d  RDr  ��   0�@     S       �  ?nc �)   �\Kcc ��  �hKcp �:  �`JD�@     %       Ke �
?
  �d  Rbs  ��   ݕ@     S       ��  ?nc �)   �\Kcc ��  �hKcp �:  �`J�@     %       Ke �
?
  �d  R�p  ��   ��@     S       ��  ?nc �)   �\Kcc ��  �hKcp �:  �`J��@     %       Ke �
?
  �d  R�s  ��   7�@     S       �a  ?nc �)   �\Kcc ��  �hKcp �:  �`JK�@     %       Ke �
?
  �d  R|q  ��   �@     S       ��  ?nc �)   �\Kcc ��  �hKcp �:  �`J��@     %       Ke �
?
  �d  R�p  ��   ��@     S       �9  ?nc �)   �\Kcc ��  �hKcp �:  �`J��@     %       Ke �
?
  �d  Rar  x�   >�@     S       ��  ?nc x)   �\Kcc y�  �hKcp z:  �`JR�@     %       Ke {
?
  �d  R s  l�   ��@     J       �  ?nc l�   �\Kcc m�  �hKcp n:  �`J�@     (       Ke o
?
  �d  R�o  d�   ��@     K       �}  ?nc d�   �\Kcc e�  �hKcp f:  �`J��@     (       Ke g
?
  �d  R�p  \�   S�@     V       ��  ?nc \�   �\Kcc ]�  �hKcp ^:  �`Jg�@     (       Ke _
?
  �d  R�s  T�   ��@     V       �U  ?nc T�   �\Kcc U�  �hKcp V:  �`J�@     (       Ke W
?
  �d  Rp  L�   ��@     V       ��  ?nc L�   �\Kcc M�  �hKcp N:  �`J��@     (       Ke O
?
  �d  Rp  D�   Q�@     V       �-  ?nc D�   �\Kcc E�  �hKcp F:  �`Je�@     (       Ke G
?
  �d  R�q  <�   ��@     V       ��  ?nc <�   �\Kcc =�  �hKcp >:  �`J�@     (       Ke ?
?
  �d  R�p  4�   ��@     V       �  ?nc 4�   �\Kcc 5�  �hKcp 6:  �`J��@     (       Ke 7
?
  �d  RZp  ,�   O�@     V       �q  ?nc ,�   �\Kcc -�  �hKcp .:  �`Jc�@     (       Ke /
?
  �d  R�o  $�   ��@     V       ��  ?nc $�   �\Kcc %�  �hKcp &:  �`J�@     (       Ke '
?
  �d  Rts  �   ��@     V       �I  ?nc �   �\Kcc �  �hKcp :  �`J��@     (       Ke 
?
  �d  Rp  �   M�@     V       ��  ?nc �   �\Kcc �  �hKcp :  �`Ja�@     (       Ke 
?
  �d  Rq  �   ��@     V       �!  ?nc �   �\Kcc �  �hKcp :  �`J�@     (       Ke 
?
  �d  St  �@     0       �J  ?c "*:  �l =O  i  �@           �  >�  �  ��?nc 0�  ��?wc 0-�  ��Kuc 1{   �oTy�  7p
  �PT�W  8�
  �@Kst 9�   ��O�    	�B     J��@     .       Ke ;?
  �h  :�    ;N      UC  2(  ;  D�  �  D   �    M    ^  A@            �g  G(  �h C�  u    D�  �   Vg  a  �  "@@     \       �Gu  �h  Q   �  \	  z  	   	          �K  -  5   ]int 5   -�3  M   X   M   �  X   -�Q  M   $��  ��   p   -N  ^1  ,  2N  �   !�  @'  �  M       	p   �   #	p       &	p   �  )	p    P  ,	p   (�  -	p   0  25   8>  55   < $  8"�   -@  K?  '  -)  L?  -�   M?  �  _L  �  i  �  �  �  $  ��   $%   4�  �  `frg �   =#  	�  a�i  �   >}C  	�  ?�  I]I  �     @�  A�-  5     ,�6   Jred ,�C   �Q  0�  �Q  �+  <  B  �    (�Q  �*  V  a  �   �    )�#  �_  �   y  �  �   �    �N  �    �R  �   �7  �   \.   �   >*  !�    �R  "�  (   �R  %$  7^  '
   �     T   L%   K�  '�V  �   T C  5%    BD  5�  Lh 8�_  �   J  5%   �N  =j4  5%  d  5%   �R  B�i  5%  ~  5%   �7  E�N  5%  �  5%   \.  I�P  5%  �  5%   >*  L�  5%  �  5%   %  P�,  5%  �  �  n%   8�+  U}O  �     5%   8\G  Z�"  �      5%   �G  dma  4  :  n%   (�G  g"  N  Y  n%  y%   )�#  i  %  q  |  n%  y%   %Rr  o_L  5%  �  �  n%   �(  |�^  �  �  n%  5%   �e  ��  �  �  n%  5%  5%   i  ��=  �    n%  5%  5%   �+  ��B    $  n%  5%   �l  �0  9  D  n%  5%   �2  .A  Z  j  n%  5%  5%   Q:  D�  �  �  n%  5%  5%   �l  xm  �  �  n%  5%   �R  ��6  �  �  n%  5%   �  +  �  �  n%  5%   �  �       n%  5%   �_  #=M  (  3  n%  5%   2�1  0Z$  �   M  S  n%   2�1  9mI  �   m  �  n%  5%  &"  �%  �%   .  ��    D �  T C  9E3  Q  A �   $  M�'  �t  ��  ��  ��  �d  �~  ��  B$   �b  �@    %  �%  L   �+  ��m  :  E  �%  5%   .�5  �L  T C  9E3  Q  L L  A �   �S  5  Lh 88Y  �   �  L%   �N  =�!  L%  �  L%   �R  BbJ  L%  �  L%   �7  E�h  L%  �  L%   \.  If  L%    L%   >*  LV/  L%    L%   %  P�[  L%  4  :  �%   8�+  U9  �   U  L%   8\G  Z-  �   p  L%   �G  d3<  �  �  �%   (�G  gn.  �  �  �%  �%   )�#  itF  �%  �  �  �%  �%   %Rr  o�+  L%  �  �  �%   �(  |�j  �  
	  �%  L%   �e  �jK  	  /	  �%  L%  L%   i  �A]  D	  T	  �%  L%  L%   �+  �6  i	  t	  �%  L%   �l    �	  �	  �%  L%   �2  H)  �	  �	  �%  L%  L%   Q:  D�  �	  �	  �%  L%  L%   �l  x.8  �	  
  �%  L%   �R  �Ld  
  "
  �%  L%   �  �  8
  C
  �%  L%   �  �R  X
  c
  �%  L%   �_  #	g  x
  �
  �%  L%   2�1  0  �   �
  �
  �%   2�1  9�  �   �
  �
  �%  L%  &"  �%  �%   .  ��    D   T   9E3  Q  XA �   t  bX  ���  �
	  �/	  ��  ��  �  Bt   �b  �R%  f  q  �%  L   �+  ��  �  �  �%  L%   .�5  �L  T   9E3  Q  XL L  A �    ?�  I]I  �     @�  2l    cclz �  5     �    T �    d%B  �$�  AL3  5   �>  ,�6   ,�i  ,'      8  H�	   8  ��Q  d  y  5%    �  p    ( 8  �&  �  �  5%  @%   )�#  �
[  F%  �  �  5%  @%   %qe  �ze  �   �  �  5%  �    8  �>   v6  ��  ��  �|   �  ��   C  8  ��	�  BC   8  �i'  ?  T  L%  �  p   5    (8  �E2  h  s  L%  W%   )�#  ��G  ]%  �  �  L%  W%   ��  �<   H�(  ��   L�-  �c%  P+  ��  X   �>  �	G  �>  �Q*  �  �  c%   (�>  �0o      c%  p&   )�#  ��>  v&  .  9  c%  p&   �+  �c%    �  �5  �	~  N�R  ��3  �   m  �%  @%  @%       �	�    �'  �  �  �%   ,+  �	�    �Q  �L%  �G  ��   $�b  ��  C%  ��Z  �  �  *%  �%   
N�  �YV  �       *%  p    2�&  H
:  �   7  G  *%  �   p    ��  z�W  ]  h  *%  �    Q.  �]  ~  �  *%  �   p    
�:  -	�c  p   �  �  *%   e�\  :�%                         @       C�Z  < �   CkG  = �    =d  D�\  p     �      S  p   +  p    C�&  f<   3�  h|   Oa  k�  �   `  �    3�e  x|   3�&  {|   f]  �|    D�i  ��U  5%  �  �  *%  �   D�i  �C  L%  �  �  *%  5    D'  !�C  5%  �  �  *%  p    �  3  
    *%   �@  :�5  %  0  *%  5%   �=  �
�%   �  ��   $8  ��  +2  �J  �  �	p    Y  �:&  (/�^  {!  /D=  �    =I  �  O�\   �  A�V  5   ,�  ,�6   ,�  Jhex  :4D     g0  {+  h�2  |5   0  ~m[  	    �!   E/   .    �!  5     �=  �g  @  F  �!   �=    [  f  �!  �   �=  4H  {  �  �!  "   �=  �?  �  �  �!  "   �=  *�l  �  �  �!  "   �=  0]  �  �  �!  "   �=  8�7  �    �!  5    
�#  = A  "    *  �!  �   
fF  Q�1  �   C  I   "   
fF  T�6  �   b  h  �!   
\?  X�:  �   �  �   "   
�"  \iQ  "  �  �   "   
�"  `�:  &"  �  �  �!   
2d  dF  ,"  �  �  �!   ;W  ��  �  �  �!   ~  ��   �6  ��   T 5    �  4.  2  4.  3�*  F  L  2"   %�(  6UB  %  d  o  2"  �   �(  <�   C.  =5   .]  >�  E0  ?�   �e  @�   �  A�   �_  B�   rO  C�   i3.  BW  �  �  2"  5    j4.  �%     2"  5O    %  >�  J�  4#�  NE�  _  P   T �   �$  �   �   5   5   5   X    4�}  x=  �  P   T �   �$  �   5   5   5   X    kzx  �U|  T �   F   �   %  �$    :�q  x  q  }r  �  �  N#   q  �q      N#  �!   q  �q  $  4  N#  �!  p    
�  <s  �!  M  S  Y#   
p  "Yq  d#  l  w  Y#  p    
  &	�o  p   �  �  Y#   
�r  *r  �   �  �  Y#  �   
�r  2�p  �   �  �  Y#  �   
Mr  6	�o  p   �    N#  X   p    
jr  >	�s  p      +  N#  X    
�q  F�s  �  D  T  N#  p   p    V W�!   ��  X	p   /�s  X    �  M9{  �  9{  ![w  �  �  q#  |#  p    .t %|#   .  &	p    }  =~6  	
�  O�  	�  g&  	�  6a  	E ?      �$  �#   �  �		�  �  	�2  ;  F  �$  �$   (�  	?N  Z  e  �$  �$   )�#  		�*  �$  }  �  �$  �$   �  	Pl  �  �  �$  5    %Y4  	"	�c  �$  �  �  �$  �   R0  	',;  �  �  �$  X    R0  	1u?  �    �$  �!   0Ba  	>�$   0t 	?�$  0�\  	@
p   �08]  	A�   �%�z  		D{  �$  _  j  T }  �$  }   N�5  		9+  �$  �  T �!  �$  �!      %�R  	H $    �  �  �$   �0  	MY  �  �  �$  �!   0�V  	Q�#   /�  �#  l�-  �   � m   :�~   
�  }w  
�Gt    (  �$  �$   }w  
K~  =  H  �$  �$   }w  
".z  ]  h  �$  �$   M|  
��w  }  �  �$  5    
�#  
)
%�  %  �  �  �$  �   
ux  
�w  %  �  �  �$  %   
ux  
���  %  �  �  �$  %   
%y  
2;}  %      �$  %   
%y  
6�{  %  1  <  �$  %   Fpop 
��x  M   U  [  �$   >  
B6�  p  v  �$   
�  
H�~  �$  �  �  �$   
�  
Lev  %  �  �  %   
  
P	�{  p   �  �  %   
o�  
T��  �   �  �  %   
d 
X�y  �$      �$   
d 
\u�  %  *  0  %   Fend 
`�w  �$  I  O  �$   Fend 
d�  %  h  n  %   
q  
hȁ  %  �  �  �$   
q  
k"x  %  �  �  %   
$  
o�t  %  �  �  �$   
$  
r�u  %  �  �  %   
p  
v�v  %      %  p    
p  
y�|  %  '  2  �$  p    �}  
��t  F  Q  �$  p    G%  
�*%   ,�  
��$    
�	p   �}  
�	p   T M   /�-     �  G�Z  �+  GA)  �7  GA)  �7�  :�Z  P  �c  �l  �  �  S&   �c  w  �    S&  �  u!   �c  =  $  /  S&  u!   n�c  !zG  D  O  S&  ^&   �c  #�  d  o  S&  d&   �c  (�;  �  �  S&  5    
�#  -4  j&  �  �  S&  �   �c  2�n  �  �  S&   a  8p;  �  �  S&   
S  >�&  �       S&   
+H  BY0  �   !  ,  S&  d!   �  G	d!   R  H�   /D=  �    �  l?  
CI  "  {  T 5   "  "   4�H  ���  �  F   �   %  �$   ;�  7�u  �  T �   F   w9  %  �$   ;�H  6y  �  F   }  %  �$   4�H  ��(      F   �!  %  �$   ;~  2܃  J   T }  F   �@  �$   ;�k  2:c  t   T �!  F   NA  �$   $q  [!�   5�  oF  �   5�    �   �    5�  ^P  _!  ^P  �b  �   �   d!   (^P  �#  �   �   d!  o!   )�#  PK  u!  !  !  d!  o!   �c  �!  0!  6!  d!   a  �l  J!  P!  d!   0je  5     �   �   d!  _!  �   �-  �!  omap �7  �  �!  �!  �!  p    E�@   H  �!  �!  �  p     {!  H�  	=B     _   �!  �  �!  �  �!  <   65      6�  �     5   5   %  2"  pstd  3#  �   Ju"  3`?  K�   T 5   P�-  Q"    �1  J�"  3`?  K�   T 5   P�-  Q"    z  �"  $8  M   T %   R@  Nh  �   R@  NW3  �   4�  �z  	#  T M   %  %   $�}  >�"  Kz  !Uu  	#  T %  %    S�#  U"  S�?  �"  (N  �  N#  x  Y#  _   �+  }  q#  �#  qH�  	>B     >de  $  P  �#  rP  
�-  �#  �#  $   E�R  �  �#  $  �!    TB  +|  �  T'.  ,�R  �   �#  ?o$  s)}  w$  U�z  O,$  t    U�z  <H$  t   �!  �    tvw  -u}  ('%  vu�  p   t     @	$  &M   �$  '�     H$  	 C     w�{  �$  	�C     M   �  �$    �$  �    &X   �$  '�    �  �$    �  6�  �  M   S   6M   S   �  %    *%  C  5%    C    L%  �    �  c%  $  n%  �  $  5%  L  �%  �  �%  t  �%    t  L%    �%  ~  {!  &|   �%  '�    �%  7eW  �  7�i  �  7�  �  7Gb  +  V'  9   �VQ5  `   x�:  m     7L  z  &~  J&  '�    y�  �   �  S&  P  6�  �  G  �  5�"  5�"  *U  �@     (       ��&  T 5   a "  �hb #"  �`   h�@     �      ��'  P   T �   ��  N�$  ��^W  N$�   ��H*  N1�   ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�!  �Xu S�'  ��k T5   �� X�@     E       �'  i a5   �l  ��@     -       �'  i d5   �h Բ@     0       i f5   �d  &X   �'  '�    U  B�@     1       �*(  �2  ZL%  �h _  �@     U       ��(  P   T �   ��  x�$  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �TWz�  {	�       �(  Ƃ@     V      �)  �  t%  �Xn �5%  �P�N  �5%  �hd4  �5%  �` �	  2)  �|@     �      �*  �  �%  ��+n xL%  ��	�N  {L%  �Ps �L%  �X	�R  ��  �� �}@     �       �)  x �L%  �H  �~@     z       �)  x �L%  �@  w�@     Q       �)  	f?  �L%  �� Ɓ@     Q       	f?  �L%  ��  "
  /*  ��@     �      �v*  �  �%  ��+n L%  ��u L%  �Xv L%  �Pw L%  �H 
  �*  �@     �      ��*  �  �%  ��+n �L%  ��u �L%  �Xv �L%  �Pw �L%  �H :  �|@     1       �+  �2  UL%  �h �  ��@            �2+  �  =L%  �h *�  �@            �d+  T   �2  'L%  �h *  �@            ��+  T C  �2  '5%  �h �  �+  D�@     �      ��+  �  t%  ��+n 5%  ��u 5%  �Xv 5%  �Pw 5%  �H �  ,  ��@     �      �b,  �  t%  ��+n �5%  ��u �5%  �Xv �5%  �Pw �5%  �H   s�@     1       ��,  �2  Z5%  �h �  w�@     �       ��,  T �   F   �2  ��   �lfo �/%  �`��  �6�$  �X P  �,   -  �  ;%  !�"  �  !�  �%�  !&8  �6p    "�,  ;R  C-  Xp@     K       �d-  �,  �h�,  �d-  �X-  �P �  �-   o@     7      ��-  �  t%  �H�N  �5%  �@�2  �"5%  ��72  �5%  �X �  �-  �m@     7      �.  �  t%  �H�N  �5%  �@�2  �!5%  ���l  �5%  �X �  7.  ~m@     j       �S.  �  t%  �h�2  |5%  �` +  a.  �.  �  R%  !�  ��  !&8  �)p   !X[  �65    "S.  &Z  �.  m@     d       ��.  a.  �hj.  �`v.  �X�.  �T �	  �.  �j@     �      �R/  �  �%  ���2  L%  ���   L%  ��	�N  L%  �X	�R  L%  �P	�7  L%  �H �	  q/  h@     a      ��/  �  �%  ���2  DL%  ��f?  D$L%  ��	�l  EL%  �X	72  FL%  �P	�N  ZL%  �H   �|@            ��/  �  LL%  �h c
  0  N|@     H       �H0  �  �%  �X�2  #L%  �P	� $L%  �h �  oj@            �s0  �  IL%  �h *�  8|@            ��0  �  8L%  �h T	  �0  �x@     V      ��0  �  �%  �Xn �L%  �P�N  �L%  �hd4  �L%  �` C
  1  �x@            �11  �  �%  �h�2  L%  �` �  P1  �x@            �m1  �  t%  �h�2  5%  �`   �1  Zx@     H       ��1  �  t%  �X�2  #5%  �P	� $5%  �h J  =x@            ��1  �  =5%  �h �  2  zr@     �      ��2  �  t%  ��+n x5%  ��	�N  {5%  �Ps �5%  �X	�R  ��  �� Is@     �       r2  x �5%  �H  et@     z       �2  x �5%  �@  v@     Q       �2  	f?  �5%  �� Zw@     Q       	f?  �5%  ��  �  Hr@     1       �3  �2  U5%  �h �  *r@            �73  �  L5%  �h *1  r@            �b3  �  85%  �h {  -�@     J       ��3  F   �2  �!�   �Lfo �8%  �@��  �?�$  �� �  �3   ^@     �       �4  �  0%  �H  !=p   �@	v6  '�  �Xfra )5%  �P %  .4  �\@     �       �[4  �  �%  �X�2  �5%  �P	� �5%  �h �  z4  �[@     D      �05  �  0%  ����  95   ��	v6  �  �@	�  	�   ��	�H  
	p   �Xslb L%  ��	Rr  c%  �Pk\@     ^       off p   �H�\@     >       	�2  c%  ��   �  O5  D[@     X       �k5  �  �%  �X� pL%  �h t	  �5  �Z@     �       ��5  �  �%  �H�2  L%  �@	v  L%  �h	�\  L%  �`�Z@     I       	�l  L%  �X  /	  6  �f@     7      �C6  �  �%  �H�N  �L%  �@�2  �"L%  ��72  �L%  �X �  �f@            �n6  �  EL%  �h 
	  �6  �e@     7      ��6  �  �%  �H�N  �L%  �@�2  �!L%  ���l  �L%  �X �  be@            ��6  �  BL%  �h Y  7  :e@     (       �97  �  �%  �ha �!@%  �`b �1@%  �X �  X7  �d@     j       �t7  �  �%  �h�2  |L%  �`   �7  �d@            ��7  �  �%  �h D  �7  2b@     �      �8  �  t%  ���2  5%  ���   5%  ��	�N  5%  �X	�R  5%  �P	�7  5%  �H �  b@            �J8  �  I5%  �h j  i8  �_@     a      ��8  �  t%  ���2  D5%  ��f?  D$5%  ��	�l  E5%  �X	72  F5%  �P	�N  Z5%  �H ~  �_@            ��8  �  E5%  �h d  u_@            �9  �  B5%  �h �  >9  �]@     L       �K9  �  Y&  �h �  j9  d_@            �w9  �  t%  �h �   �  ߯@     N       ��9  T �   F   �2  7w9  �H+fo 7-%  �@��  74�$  �� �  �9  D�@     �       �:  �  �$  �hs 	'X   �d �  0:  �p@     �       �L:  �  �$  �hstr 	1�!  �` �  k:  
O@     �      �|;  �  0%  ��~��  �6p   ��~ JO@     �      6;  ��  �5   �\bkt ��%  �PsZ  ��  ��	�2  c%  �� �O@     *      ;  slb 	L%  �H �P@     �      slb 	L%  �@	�\  �  ��  �R@     �       	  6�   ��fra 75%  ��	�\  9�  ��~  q  �;  �Y@     �       ��;  �  �%  �X�2  �L%  �P	� �L%  �h �  �;  JY@     I       �<  �  ;%  �Xp ��   �Padr �	�   �h �  <  (<  �  i%   #<  �`  K<  4Y@            �T<  <  �h �  s<  �X@     O       ��<  �  Y&  �h $  �<  (X@     �       ��<  �  t%  �H�2  5%  �@	v  5%  �h	�\  5%  �`�X@     I       	�l  5%  �X  �  =  `W@     �       �J=  �  0%  �Xv6  �;�  �P	� �5%  �h o  X=  k=  �  Y&     <    "J=  �  �=  8W@     '       ��=  X=  �h   �=  �=  �  Y&  !�  u!   "�=  dh  �=  W@     2       ��=  �=  �h�=  �` �  ٭@           ��>  F   �t  '}  ��+fo <%  ����  C�$  ��p �>  �`�@     �      i p   �h�@     �      c 	i  �_   p  �  �^@     *       ��>  F   �2  � �!  �hfo �7%  �`��  �>�$  �X 2  ?  ֬@           ��?  �  �$  ���}  
�4p   ��y  
�	p   �H��  
��$  �@ "�@     ^       f?  i 
�p   �X ��@            i 
�p   �P  G  �?  �K@     h      �Y@  �  0%  ��~W z0�   ��~	v6  ��   �X	�\  ��  ��fra �5%  �Pslb �L%  �Hbkt ��%  �@	�  �	p   ��	sZ  ��  ��	�-  ��   ��	�2  �c%  ��   g@  �@  �  T#  Xs  �!  !��  *p    #Y@  �u  �@  ��@     *       ��@  g@  �hp@  �`z@  �X �  �@  �V@     &       ��@  �  �$  �ha  	M�!  �` �      c�@     I       �NA  T }  F   �2  2�@  �H��  2!�$  �@ �!  J   TV@     E       ��A  T �!  F   �2  2NA  �H��  2!�$  �@ '  �A  �A  �  �$  !Ca  	�$   #�A  �n  �A   V@     4       ��A  �A  �h�A  �`   B  B  �  �!     <    #�A  =e  :B  V@            �CB  B  �h �  QB  [B  �  �!   #CB  �H  ~B  V@            ��B  QB  �h <  �B  �@     I       ��B  �  �$  �X�^  
�M   �h �"  ˫@     O       �C  T M   x %  �Xy %  �P!Z  M   �h *#  ��@            �>C  T %  x *%  �h �  ]C  ��@            �jC  �  %%  �h �  �C  ��@     %       ��C  �  �$  �h   �C  `�@     !       ��C  �  �$  �h��  
yp   �` �  �C  ڪ@     �       �D  �  �$  �H�^  
�#%  �@W 
��$  �X �  :D  b�@     w       �eD  �  �$  �X�^  
�(%  �PW 
��$  �h [  �D  .�@     4       ��D  �  �$  �X6�@            i 
Cp   �h  v  �D  �@            ��D  �  �$  �h h  �D   	E  �  �$     <   W{i 
�p     "�D  �z  ,E  ֩@     F       �bE  �D  �X|�D  CE  }�D   ~�D  �@            �D  �h    pE   �E  �  �$  !H%  
�)�$   #bE  ۂ  �E  ��@     >       ��E  pE  �hyE  �` �  �E  ��@            �F  �  _#  �X�-  *%�  �@Þ@     G       i -p   �h  +  3F  &�@     r       �^F  �  T#  �X �  F&p   �P  F3p   �H �  }F  LK@     ,       ��F  �  �$  �h��  �  @  �F  �@     6       ��F  T }  �  �$  �h�2  	}  �P w  �F  ި@            �G  �  _#  �h 4   G  ̨@            �-G  �  _#  �h j  SG  "K@     )       �oG  T �!  �  �$  �h�2  	�!  �` �  }G  �G  �  �$     <    #oG  'F  �G  K@            ��G  }G  �h �  �G  �J@     )       ��G  �  �$  �` �  H  x�@     S       �OH  �  T#  �Xc 6X   �T�  6#p   �H��@     9       i 7p   �h  �  ]H  rH  �  T#  Xcs  �!   #OH  $p  �H  @�@     R       ��H  ]H  �hfH  �` �  �H  �H  �  �!  !�-  *"   "�H  �b  �H  �C@     V       ��H  �H  �h�H  �` �  I  I  �  �!     <    "�H   Y  BI  �C@            �KI  I  �h +  YI  cI  �  �!   "KI  �@  �I  �C@     #       ��I  YI  �h <�t  �5   �@     >       ��I  �3  ��!  �X <�t  x5   �@     �      �TJ  �3  x�!  ��}`?  x*�!  ��}�~  x55   ��}"q  yt   ��~s z	p   �X�  �M   ��}1�  dJ  	�*B      &_   dJ  '�    TJ  </y  m5   o�@     �       ��J  �  m�!  ��"q  nt   �@s o	p   �X1�  dJ  	�*B      <z  bM   ��@     �       �:K  �3  b�!  ��k c�   �h"q  gt   �@s h	p   �`1�  dJ  	�*B      $  3�@     r      ��K  �3  O)t   �@}w  P%  �X1�  �K  	�*B     k S�   �P &_   �K  '�    �K  ,$  ��@     ?      �$L  �3  <'t   ���  <9�!  ���~  <F�   ��}w  =%  �X1�  4L  	p*B     k @�   �P &_   4L  '�    $L  H$  '�@     �       ��L  }w  .%  �`k�@     P       i 5p   �h  P$  ��@     o       ��L  }w  ).�  	 C        �B@     �       �DM    S0p   ��tc U�   �`e ^�   �Xf _�   �Pip `�   �His a�   �@�B@     :       i W�   �l  *�  $B@            ��M  idx D6�   ��tc F�   �hs K5   �dip L�   �Xis M�   �Pf N�   �H \$  �@     �      �.N  �3  ,t   ��}6�@     o      i p   �X_�@     <      "q  t   ��~s 
p   �P   �  <N  `N  �  w#  Yu !|#  Y  !(p    #.N  ,t  �N  N�@     *       ��N  <N  �hEN  �`RN  �X L  �N  2A@     6       ��N  �  8"  �`c 63�  �\�  7%  �h Z�  2�N  	O  �  8"     <    "�N    ,O  A@            �5O  �N  �h   Z�  2LO  [O  �  8"  5O   ";O  �  ~O  ~@@     �       ��O  LO  �hUO  �` 2  �O  �O  �  8"   "�O  a  �O  "@@     \       ��O  �O  �h �F  nH  �   @@            �P    #p   �hp /�   �` 6!  6P  B@            �CP  �  j!  �h !  bP  �A@     B       ��P  �  j!  �h1�  �P  	g*B      &_   �P  '�    �P  *�  �A@            ��P  x )�   �h (  �P  �P  �  �    #�P  �b  �P  hA@     Q       �Q  �P  �h [C  �  "[  �  " q    �  	  >�  	  )u    4   
       �int �3  Q   	HC     W   �  �Q  Q   	PC      ��   (  r	  g�  	  �          qu  C  5   sint 
5   C�3  M   X   DM   .�  
X   C�Q  M   'ߚ  (|   t�  �   +�   �   /�     .-N  
�   uM�   �   J��   �    J��   �   J!�   �   J̼   �    .2N  
�   v'�  cp   '��  ��   
�   '��    .1  !�  @�  �  M       	�   �   #	�       &	�   �  )	�    P  ,	�   (�  -	�   0  25   8>  55   < '  8"  'E�  9�   
�  C@  K�  �  D�  C)  L�  C�   M�  .�  
�  .�  .�  .�  '�  �  '  ��   '��  /  '%   4  
0  .,  K�r  e�   '��  �  .�  wL  xfrg :,  W#  	
y  y�i  �   X}C  	�  Y�  `]I  F,    Z�  L�-  5   �  $�6   ared $�C   �Q  0�  �Q  �+      P,   >�Q  �*    '  P,  [,   ?�#  �_  a,  ?  J  P,  [,   �N  �    �R  �   �7  �   \.   �   >*  !�    �R  "�  ( 
�  �R  %�  &�  '�V  ?,  �  T 	  �6   [7^  '
   ?,  T �  7    BD  5|  bh 8�_  P,    �6   &�N  =j4  �6  *  �6   &�R  B�i  �6  D  �6   &�7  E�N  �6  ^  �6   &\.  I�P  �6  x  �6   &>*  L�  �6  �  �6   ;  P�,  �6  �  �  47   M�+  U}O  ?,  �  �6   M\G  Z�"  ?,  �  �6   �G  dma  �     47   >�G  g"      47  ?7   ?�#  i  E7  7  B  47  ?7   ;Rr  o_L  �6  Z  `  47   �(  |�^  u  �  47  �6   �e  ��  �  �  47  �6  �6   i  ��=  �  �  47  �6  �6   �+  ��B  �  �  47  �6   0�l  �0  �  
  47  �6   3�2  .A     0  47  �6  �6   3Q:  D�  F  V  47  �6  �6   3�l  xm  l  w  47  �6   3�R  ��6  �  �  47  �6   3�  +  �  �  47  �6   0�  �   �  �  47  �6   0�_  #=M  �  �  47  �6   G�1  0Z$  ?,      47   G�1  9mI  ?,  3  M  47  �6  �-  K7  K7   @  ��    D �  T 	  NE3  ��  A �   
�  <�'  �:  4�`  4��  4��  4�*  4�D  4��  \�   0�b  �@  �  �  \7     0�+  ��m       \7  �6   @�5  �  T 	  NE3  ��  L   A �   �S  5�  bh 88Y  P,  `  7   &�N  =�!  7  z  7   &�R  BbJ  7  �  7   &�7  E�h  7  �  7   &\.  If  7  �  7   &>*  LV/  7  �  7   ;  P�[  7  �   	  g7   M�+  U9  ?,  	  7   M\G  Z-  ?,  6	  7   �G  d3<  J	  P	  g7   >�G  gn.  d	  o	  g7  r7   ?�#  itF  x7  �	  �	  g7  r7   ;Rr  o�+  7  �	  �	  g7   �(  |�j  �	  �	  g7  7   �e  �jK  �	  �	  g7  7  7   i  �A]  

  
  g7  7  7   �+  �6  /
  :
  g7  7   0�l    O
  Z
  g7  7   3�2  H)  p
  �
  g7  7  7   3Q:  D�  �
  �
  g7  7  7   3�l  x.8  �
  �
  g7  7   3�R  �Ld  �
  �
  g7  7   3�  �  �
  	  g7  7   0�  �R    )  g7  7   0�_  #	g  >  I  g7  7   G�1  0  ?,  c  i  g7   G�1  9�  ?,  �  �  g7  7  �-  ~7  ~7   @  ��    D �  T �  NE3  ��  XA �   
:  HX  �4��	  4��	  4��	  4�z  4��  4��  \:   0�b  �R%  ,  7  �7     0�+  ��  L  W  �7  7   @�5  �  T �  NE3  ��  XL   A �    Y�  `]I  F,    Z�  2l  �  zclz �  5   �  �    T �    {%B  �$V  LL3  5   �  $�6   $�i  $'   
�   8  H�	�   8  ��Q  *  ?  �6  �  0  �    > 8  �&  S  ^  �6  7   ?�#  �
[  7  v  �  �6  7   ;qe  �ze  ?,  �  �  �6  �    8  �   v6  �<  ��  �  �  ��%   
	  8  ��	�  \	   8  �i'      7  0  �   5    >8  �E2  .  9  7  7   ?�#  ��G  #7  Q  \  7  7   ��  �<   H�(  ��   L�-  �)7  P+  ��%  X 
�  �>  �	  �>  �Q*  �  �  )7   >�>  �0o  �  �  )7  9   ?�#  ��>  9  �  �  )7  9   �+  �)7    
�  �5  �	D  c�R  ��3  ?,  3  Q7  7  7       �	�    �'  e  k  �7   ,+  �	l,   �Q  �7  �G  ��   '�b  ��%  C%  ��Z  �  �  �7  �7    N�  �YV  �   �  �  �7  �    G�&  H
:  �   �    �7  �   �    3��  z�W  #  .  �7  �    3Q.  �]  D  T  �7  �   �     �:  -	�c  �   m  s  �7   |�\  :�7                         @       ]�Z  < �   ]kG  = �    &=d  D�\  �   �  �    &  S  �   �  �    ]�&  f<   A�  h  &Oa  k�  ?,  &  �    A�e  x  A�&  {  }]  �   ^�i  ��U  �6  h  s  �7  0   ^�i  �C  7  �  �  �7  5    ^'  !�C  �6  �  �  �7  �    0�  3  �  �  �7   0�@  :�5  �  �  �7  �6   �=  �
�7   �  �l,  '8  ��%  +2  �  �  �	�    Y  �8  (�^  4-  D=  l,   WI  
V  d�\   _  L�V  5   ,�  $�6   $�  ahex  O4D    ~0  {�  �2  |5   0  ~m[  �  �  �-   _/   .  �  �-  5     �=  �g      �-   �=    !  ,  �-  V   �=  4H  A  L  �-  �-   �=  �?  a  l  �-  �-   �=  *�l  �  �  �-  �-   �=  0]  �  �  �-  �-   �=  8�7  �  �  �-  5     �#  = A  �-  �  �  �-  �    fF  Q�1  ?,  	    �-    fF  T�6  ?,  (  .  �-    \?  X�:  ?,  G  M  �-    �"  \iQ  �-  f  l  �-    �"  `�:  �-  �  �  �-    2d  dF  �-  �  �  �-   ;W  ��  �  �  �-   ~  ��   �6  �?,  ��  %�  �    U �-  �-  �-   T 5    
�  4.  2�  4.  3�*  3  9  �-   ;�(  6UB    Q  \  �-  p   �(  <p   C.  =5   .]  >�  E0  ??,  �e  @?,  �  A?,  �_  B?,  rO  C?,  3.  BW  �  �  �-  5    �4.  �%  �  �-  ��    
  X�  JS  �  N	�  M  P �#  T 5   =1  5   ?,  5   5   5   X    #�  NE�  �  P �#  T �   =1  �   ?,  5   5   5   X    �}  x=  �  P �#  T �   =1  �   5   5   5   X    ��  x;�  	  P �#  T 5   =1  5   5   5   5   X    zx  �U|  7  T �   F �#  �     =1   �  �ܪ  e  T 5   F �#  5     =1   �  N�  �  P q3  T 0  �=  0  ?,  5   5   5   X    "�  NV�  �  P q3  T �   �=  �   ?,  5   5   5   X    h�  N��  +  P q3  T   �=    ?,  5   5   5   X    �  N��  m  P q3  T �   �=  �   ?,  5   5   5   X    -�  Nh�  �  P �1  T 0  GE  0  ?,  5   5   5   X    ��  N�  �  P �1  T �   GE  �   ?,  5   5   5   X    ǉ  ND�  3  P �1  T   GE    ?,  5   5   5   X    Ǒ  Nέ  u  P �1  T �   GE  �   ?,  5   5   5   X    ĥ  Nt�  �  P �2  T 0  �I  0  ?,  5   5   5   X    I�  N��  �  P �2  T �   �I  �   ?,  5   5   5   X    ��  Nf�  ;  P �2  T   �I    ?,  5   5   5   X    ��  Nݹ  }  P �2  T �   �I  �   ?,  5   5   5   X    9�  N��  �  P C1  T 0  O  0  ?,  5   5   5   X    ��  Nd�    P C1  T �   O  �   ?,  5   5   5   X    D�  Nϧ  C  P C1  T   O    ?,  5   5   5   X    ��  N۸  �  P C1  T �   O  �   ?,  5   5   5   X    V�  xP�  �  P q3  T 0  �=  0  5   5   5   X    1�  x��  �  P q3  T �   �=  �   5   5   5   X    E�  xQ�  <  P q3  T   �=    5   5   5   X    <�  x��  y  P q3  T �   �=  �   5   5   5   X    �  x�  �  P �1  T 0  GE  0  5   5   5   X    �  xJ�  �  P �1  T �   GE  �   5   5   5   X    j�  x�  0  P �1  T   GE    5   5   5   X    �  x�  m  P �1  T �   GE  �   5   5   5   X    ��  x�  �  P �2  T 0  �I  0  5   5   5   X    O�  x�  �  P �2  T �   �I  �   5   5   5   X    ՗  x�  $  P �2  T   �I    5   5   5   X    G�  x*�  a  P �2  T �   �I  �   5   5   5   X    ��  x��  �  P C1  T 0  O  0  5   5   5   X    <�  x`�  �  P C1  T �   O  �   5   5   5   X    f�  x/�    P C1  T   O    5   5   5   X    �h�  x��  P C1  T �   O  �   5   5   5   X     ��  �n  ת  �
�     L�  5   ��  $��   $�  $�  $d�   O�q  J!  q  }r  �  �  0   q  �q  �  �  0  �-   q  �q  �     0  �-  �     �  <s  �-     %   (0    p  "Yq  30  >   I   (0  �       &	�o  �   b   h   (0    �r  *r  ?,  �   �   (0  �    �r  2�p  ?,  �   �   (0  �    Mr  6	�o  �   �   �   0  X   �     jr  >	�s  �   �   �   0  X     �q  F�s  �  !  &!  0  �   �    V W�-   ��  X	�   �s  X    
�  O��   #  q  ��  q!  w!  90   q  ��  �!  �!  90  D0   q  �  �!  �!  90  D0  �     �  �  D0  �!  �!  [0    p  "ؠ  f0  �!  �!  [0  �       &	��  �   "  "  [0    �r  *��  ?,  7"  B"  [0  O!    �r  2��  ?,  ["  f"  [0  O!    Mr  6	�  �   "  �"  90  O0  �     jr  >	Ƅ  �   �"  �"  90  O0    �q  F��  O!  �"  �"  90  �   �    V WD0   ��  X	�   �s  O0   
O!  <9{  W#  09{  ![w  (#  8#  l0  w0  �    @t %w0   @  &	�    
#  W~6  	

\#  d�  	e#  g&  	�%  6a  	E ?  �#  �#  !1  �0   �  �		C%  �  	�2  �#  �#  ,1  !1   >�  	?N  �#  �#  ,1  71   ?�#  		�*  =1  $  $  ,1  71   �  	Pl  $$  /$  ,1  5    ;Y4  	"	�c  =1  G$  R$  ,1  \#   R0  	',;  f$  q$  ,1  X    R0  	1u?  �$  �$  ,1  �-   ,Ba  	>!1   ,t 	?1  ,�\  	@
�   �,8]  	A?,  �;;�  		��  =1  �$  �$  T X   ,1  X    ;�z  		D{  =1  %  %  T #  ,1  #   c�5  		9+  =1  7%  T �-  ,1  �-    
�#  ;�R  	H $  �#  `%  f%  !1   �0  	MY  {%  �%  !1  �-   ,�V  	Q�0   �  �0  ��-  �   � e   ��  K�Z  �+�  KA)  �7�  KA)  �7�  O�Z  m'  �c  �l   &  &  �8   �c  w  &  +&  �8  y  .-   �c  =  @&  K&  �8  .-   ��c  !zG  a&  l&  �8  9   �c  #�  �&  �&  �8  9   �c  (�;  �&  �&  �8  5     �#  -4  9  �&  �&  �8  �%   �c  2�n  �&  �&  �8   a  8p;   '  '  �8    S  >�&  ?,  '  %'  �8    +H  BY0  ?,  >'  I'  �8  -   �  G	-   R  H?,  D=  l,   
�%  &l?  
CI  �-  �'  T 5   �-  �-   �H  ���  �'  F �#  �     =1   �H  ���  �'  F �#  5     =1   (�  7�u  (  T �   F �#  V    =1   (ǟ  2�  ?(  T X   F �#  30  =1   (y�  ���  q(  F q3  �=  X     n  ]5   (I�  p&�  �(  F q3  �=  X     n  ]5   (��  's�  �(  F q3  �=  X     n  ]5   (�H  6y  �(  F �#  #    =1   �H  ��(  $)  F �#  �-    =1   (�  �)�  V)  F �1  GE  X     n  ]5   (��  p��  �)  F �1  GE  X     n  ]5   (ȝ  '.�  �)  F �1  GE  X     n  ]5   (��  ���  �)  F �2  �I  X     n  ]5   (h�  p��  *  F �2  �I  X     n  ]5   (}�  '��  P*  F �2  �I  X     n  ]5   (�  ��  �*  F C1  O  X     n  ]5   (��  p\�  �*  F C1  O  X     n  ]5   (n�  '�  �*  F C1  O  X     n  ]5   �  iK�  +  �-  �-   (~  2܃  ++  T #  F �#  �  =1   (�k  2:c  U+  T �-  F �#  k�  =1   /�  ��  |+  A 8  8  �-  ]5   '�  �Ż  �+  A /6  /6  �-  ]5   &��  	
�  ͛  �+  T �   ͛  ͛   m�  ��  �+  A c5  c5  �-  ]5   �  �z�  ,  A �4  �4  �-  ]5   [�Q  
!I  ͛  T �   ͛  ͛    B�  .oF  
?,  B�  �  
P,  �  �  B�  ^P  -  ^P  �b  �,  �,  -   >^P  �#  �,  �,  -  (-   ?�#  PK  .-  �,  �,  -  (-   �c  �!  �,  �,  -   a  �l  -  	-  -   ,je  5     
l,  l,  
-  -  l,  �-  �-  �map �7  0  Z-  e-  �-  �    _�@   H  u-  �-  0  �     4-  fd  	+B     _   
�-  D�-  �  
�-  �  
�-  <   )5     )�  �    5   5     
�-  �std  0  �   J5.  A`?  KF,  T 5   P�-  Q�-    �1  Jb.  A`?  KF,  T 5   P�-  Q�-    �  �.  '8  5   T �-   ��  J�.  A`?  KF,  T 5   P�-  Q�-    ��  J�.  A`?  KF,  T 5   P�-  Q�-    ��  �.  '8  ?,  T 3c   R@  Nh  F,  R@  NW3  F,  R@  N�  F,  R@  N��  F,  ��  
��  h/  T ?,  3c  3c   '�}  >�.  &��  
!�  h/  �/  T 3c  3c   A�  
>�  �/  T 5   �-  �-   &��  
ۈ  �-  �/  T �-  �   '�}  >o.  [��  
!X�  �/  T �-  �-    S�#  .  S�?  B.  .(N  �  
0  J!  
(0  _   O!  
90  V0  DD0  .�+  
O0   #  
[0  V0  #  
l0  }0  �fj#  	+B     Xde  1  P  �0  �P  
�-  �0  �0  1   _�R  �  �0  1  �-    gB  +|  v#  g'.  ,�R  �%  e$  �0  �0  +X   !1  /�    v#  
!1  �#  
,1  C%  �#  R�  D�1  R�  EI�  d1  o1  �1  �   R0  H��  �1  �1  �1  X    R0  M��  �1  �1  �1  �-   R0  R�  �1  �1  �1  �-  �    4�  W�   ��  X	�    C1  
�1  P�  [�2  P�  \b�  2  #2  �2  M    R0  _�  72  B2  �2  X    R0  d�  V2  a2  �2  �-   R0  l��  u2  �2  �2  �-  �    u tM    ��  u	�    �1  
�2  ��  xf3  ��  y'�  �2  �2  f3  M   �    R0  |�  �2  �2  f3  X    R0  �ζ  3  3  f3  �-   R0  �2�  .3  >3  f3  �-  �    u �M    �Q  �	�   ��  �	�    �2  
f3  ��  �<4  ��  ���  �3  �3  <4   ��  �4�  �3  �3  <4   R0  �ϫ  �3  �3  <4  X    R0  �W�  �3  �3  <4  �-   R0  ��  4  4  <4  �-  �    u �M    �Q  �	�   ��  �	�    q3  
<4  Y�4  ��   �
$��   $L�  $u�  $L�  $��  $�  $L�  $�    Z�G4  y�  R5  ��  ��  �4  �4  R5  �1  ]5   �R  �  �4  �4  R5  X    �R  ��  �4  5  R5  �-  �    �R  G�  5  .5  R5  X     n   ,��  @�1   ,��  A]5  F C1   �4  
R5  S  ��  $6  ��  ��  �5  �5  $6  f3  ]5   �R  E�  �5  �5  $6  X    �R  ��  �5  �5  $6  �-  �    �R  )�  �5   6  $6  X     n   ,��  @f3   ,��  A]5  F �2   c5  
$6  ��  �6  ��  N�  P6  `6  �6  �2  ]5   �R  �  t6  6  �6  X    �R  �  �6  �6  �6  �-  �    �R  ��  �6  �6  �6  X     n   ,��  @�2   ,��  A]5  F �1   /6  
�6  	  
�6  �  	  �  
7  �  �  �  
)7  �  
47  |  �  �6    
Q7  �  
\7  :  
g7  �  :  7  �  
�7  D  �  
�7  4-  +  �7  /�    
�7  IeW  s  I�i  �  I�  �  IGb  �  h'  �   �hQ5  &   ��:  3     IL  @  +D  8  /�    6�  �8  ��  ��  =8  M8  �8  <4  ]5   �R  ׯ  a8  l8  �8  X    �R  ��  �8  �8  �8  �-  �    �R  �  �8  �8  �8  X     n   ,��  @<4   ,��  A]5  F q3   8  
�8  S(�  �.  S��  �.  �%  
�8  m'  )�%  �%    �  B�.  B/  B"/  B4/    J�A     �      �e:  P �#  T 5   ��  N=1  ��^W  N$5   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ��/�A     E       ":  i a5   �l ~�A     -       E:  i d5   �h ��A     0       i f5   �d  +X   u:  /�    M  h�@     �      ��;  P �#  T �   ��  N=1  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ��X�@     E       ^;  i a5   �l ��@     -       �;  i d5   �h Բ@     0       i f5   �d  �  �@     U       �3<  P �#  T �   ��  x=1  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �T12�  {	�     �  ��A     �       ��<  P �#  T 5   ��  x=1  �X^W  x!5   �T�b  x-5   �PK.  x85   �L.]  y5   �H]  yX   �DהA     ;       �  {	�   �l  	  w�@     �       �/=  T �   F �#  �2  ��   �lfo �/  �`��  �6=1  �X 7  �A     �       ��=  T 5   F �#  �2  �5   �lfo �/  �`��  �6=1  �X 5r'  �@     (       ��=  T 5   a �-  �hb #�-  �` q3  e  n�A     �      ��>  P q3  T 0  ��  N�=  ��^W  N$0  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��g�A     E       �>  i a5   �l ��A     -       �>  i d5   �h �A     0       i f5   �d  �  ϐA     �      �!@  P q3  T �   ��  N�=  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ����A     E       �?  i a5   �l �A     -       @  i d5   �h ;�A     0       i f5   �d  �  '�A     �      �MA  P q3  T   ��  N�=  ��^W  N$  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   �� �A     E       
A  i a5   �l o�A     -       -A  i d5   �h ��A     0       i f5   �d  +  �A     �      �yB  P q3  T �   ��  N�=  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��x�A     E       6B  i a5   �l ǎA     -       YB  i d5   �h �A     0       i f5   �d  �'  -�@     J       ��B  F �#  �2  �!�   �Lfo �8  �@��  �?=1  �� �  �B  D�@     �      �0C  	�  :7  ��n �6  ��u �6  �Xv �6  �Pw �6  �H w  OC  ��@     �      ��C  	�  :7  ��n ��6  ��u ��6  �Xv ��6  �Pw ��6  �H �  Hr@     1       ��C  �2  U�6  �h   =x@            ��C  �  =�6  �h 5�  �@            �D  T 	  �2  '�6  �h 5�  �@            �PD  T �  �2  '7  �h �
  oD  ��@     �      ��D  	�  m7  ��n 7  ��u 7  �Xv 7  �Pw 7  �H �
  �D  �@     �      �E  	�  m7  ��n �7  ��u �7  �Xv �7  �Pw �7  �H 	  B�@     1       �GE  �2  Z7  �h �1  m  ׋A     �      �yF  P �1  T 0  ��  NGE  ��^W  N$0  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��ЌA     E       6F  i a5   �l �A     -       YF  i d5   �h L�A     0       i f5   �d  �  8�A     �      ��G  P �1  T �   ��  NGE  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ��(�A     E       bG  i a5   �l w�A     -       �G  i d5   �h ��A     0       i f5   �d  �  ��A     �      ��H  P �1  T   ��  NGE  ��^W  N$  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ����A     E       �H  i a5   �l ؉A     -       �H  i d5   �h �A     0       i f5   �d  3  �A     �      ��I  P �1  T �   ��  NGE  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ���A     E       �I  i a5   �l 0�A     -       �I  i d5   �h ]�A     0       i f5   �d  �2  u  @�A     �      �/K  P �2  T 0  ��  N�I  ��^W  N$0  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��9�A     E       �J  i a5   �l ��A     -       K  i d5   �h ��A     0       i f5   �d  �  ��A     �      �[L  P �2  T �   ��  N�I  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ����A     E       L  i a5   �l ��A     -       ;L  i d5   �h �A     0       i f5   �d  �  ��A     �      ��M  P �2  T   ��  N�I  ��^W  N$  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ���A     E       DM  i a5   �l A�A     -       gM  i d5   �h n�A     0       i f5   �d  ;  Q�A     �      ��N  P �2  T �   ��  N�I  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��J�A     E       pN  i a5   �l ��A     -       �N  i d5   �h ƁA     0       i f5   �d  �'  �A     J       �O  F �#  �2  �5   �Lfo �/  �@��  �6=1  �� C1  }  _~A     �      �6P  P C1  T 0  ��  NO  ��^W  N$0  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��XA     E       �O  i a5   �l �A     -       P  i d5   �h �A     0       i f5   �d  �  �|A     �      �bQ  P C1  T �   ��  NO  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ���  P�-  �Xu Se:  ��k T5   ���}A     E       Q  i a5   �l �}A     -       BQ  i d5   �h ,~A     0       i f5   �d    {A     �      ��R  P C1  T   ��  NO  ��^W  N$  ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��|A     E       KR  i a5   �l `|A     -       nR  i d5   �h �|A     0       i f5   �d  C  pyA     �      ��S  P C1  T �   ��  NO  ��^W  N$�   ��H*  N1?,  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#X   ��~�  P�-  �Xu Se:  ��k T5   ��izA     E       wS  i a5   �l �zA     -       �S  i d5   �h �zA     0       i f5   �d  �  yA     W       �LT  P q3  T 0  ��  x�=  �h^W  x!0  �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	0    �  �xA     U       ��T  P q3  T �   ��  x�=  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �T12�  {	�     �  %xA     �       ��U  P q3  T   ��  x�=  �X^W  x!  �P�b  x-5   �LK.  x85   �H.]  y5   �D]  yX   �@LxA     ?       �  {	�   �h  <  �wA     W       �V  P q3  T �   ��  x�=  �h^W  x!�   �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	�     �   �'  ߯@     N       �vV  T �   F �#  �2  7V  �Hfo 7-  �@��  74=1  �� R$  �V  D�@     �       ��V  	�  21  �hs 	'X   �d q$  �V  �p@     �       ��V  	�  21  �hstr 	1�-  �` 
  	W  �x@     V      �AW  	�  m7  �Xn �7  �P�N  �7  �hd4  �7  �` x  *r@            �lW  �  L�6  �h �  �W  Zx@     H       ��W  	�  :7  �X�2  #�6  �P� $�6  �h ^  b@            ��W  �  I�6  �h 5�  r@            �X  �  8�6  �h �  -X  Ƃ@     V      �eX  	�  :7  �Xn ��6  �P�N  ��6  �hd4  ��6  �` �  �X  �x@            ��X  	�  :7  �h�2  �6  �` 	  �X  �x@            ��X  	�  m7  �h�2  7  �` )  �X  N|@     H       �)Y  	�  m7  �X�2  #7  �P� $7  �h `  ��@            �TY  �  =7  �h �
  sY  �|@     �      �QZ  	�  m7  ��n x7  ���N  {7  �Ps �7  �X�R  ��  ���}@     �       �Y  x �7  �H �~@     z       Z  x �7  �@ w�@     Q       -Z  f?  �7  �� Ɓ@     Q       f?  �7  ��   	  �|@     1       �|Z  �2  U7  �h �  �|@            ��Z  �  L7  �h 5G  8|@            ��Z  �  87  �h y  wwA     W       �d[  P �1  T 0  ��  xGE  �h^W  x!0  �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	0    �  "wA     U       ��[  P �1  T �   ��  xGE  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �T12�  {	�     �  �vA     �       ��\  P �1  T   ��  xGE  �X^W  x!  �P�b  x-5   �LK.  x85   �H.]  y5   �D]  yX   �@�vA     ?       �  {	�   �h  0  ,vA     W       �-]  P �1  T �   ��  xGE  �h^W  x!�   �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	�     m  �uA     W       ��]  P �2  T 0  ��  x�I  �h^W  x!0  �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	0    �  �uA     U       �Q^  P �2  T �   ��  x�I  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �T12�  {	�     �  �tA     �       ��^  P �2  T   ��  x�I  �X^W  x!  �P�b  x-5   �LK.  x85   �H.]  y5   �D]  yX   �@uA     ?       �  {	�   �h  $  �tA     W       ��_  P �2  T �   ��  x�I  �h^W  x!�   �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	�     (  CtA     G       ��_  T X   F �#  �2  230  �H��  2!=1  �@ a  �sA     W       �d`  P C1  T 0  ��  xO  �h^W  x!0  �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	0    �  �sA     U       ��`  P C1  T �   ��  xO  �h^W  x!�   �d�b  x-5   �`K.  x85   �\.]  y5   �X]  yX   �T12�  {	�     �  �rA     �       ��a  P C1  T   ��  xO  �X^W  x!  �P�b  x-5   �LK.  x85   �H.]  y5   �D]  yX   �@sA     ?       �  {	�   �h  6�!  �a  �rA            ��a  	�  a0  �h !w!  �a  �a  �  ?0  Ecs  D0   *�a  ��  b  �rA     Y       �b  �a  �h�a  �` 6I   =b  ި@            �Jb  	�  .0  �h !�  Xb  mb  �  #0  Ecs  �-   *Jb  $p  �b  @�@     R       ��b  Xb  �hab  �`   4rA     W       �3c  P C1  T �   ��  xO  �h^W  x!�   �`�b  x-5   �\K.  x85   �X.]  y5   �T]  yX   �P12�  {	�     ?,  F/  �qA     J       ��c  T ?,  x 
3c  �Xy 
3c  �P!Z  
?,  �o 5t/  �qA            ��c  T 3c  x 
*3c  �h �/  �qA     J       �d  T 5   x 
�-  �Xy 
�-  �P!Z  
5   �l ?(  +qA     d       �sd  F q3  ��  ��=  �ht �*X   �d��  �<  �Xà  �n  �`vsp �%]5  �P q(  viA     �      ��i  F q3  ��  p�=  ��t p(X   ����  p:  ��à  qn  ��vsp q%]5  ���iA           e  ^W  w  �X "   )e  3�  �)e  �@ <;�  ��f  b�  c�  He  _e  Me  )e  Xe  ))e   b�  <�  pe  �e  Me  ze  �e  
)e   7b�  ��  �e  �e  Me   a�  �  �e  �e  Me  5    #��  ��i   #��  ��=  8E�  Q�  
f  @eA     �       �Hf  g�  �   g�  �   	�  f  �X
j  ^W  ��   �T��  �i  �X��  �=  �X# 9��  �  yf  fdA     �       �g�  �   g�  �   	�  f  �X^W  ��   �P��  �i  �X��  �=  �X#  "0  �f  3�  ��f  �� <��  �Xh  b�  \�  �f  g  �f  �f  �f  )�f   b�  �  g  +g  �f  g  %g  
�f   7b�  �  <g  Bg  �f   a�  '�  Sg  ^g  �f  5    #��  ��i   #��  ��=  8E�  ��  �g  �fA     �       ��g  ��  �   ��  �   	�  �g  �X
j  ^W  ��   �T��  �i  �X��  �=  �X# 9��  ��  h  fA     �       ���  �   ��  �   	�  �g  �X^W  ��   �P��  �i  �X��  �=  �X#  "`  sh  3�  �sh  �� H�  �b�  ��  �h  �h  �h  sh  �h  )sh   b�  p�  �h  �h  �h  �h  �h  
sh   7b�  ��  �h  �h  �h   a�  ֮  �h  �h  �h  5    #��  ��i   #��  ��=  8E�  0�  Pi  �hA     �       ��i  ��  �   ��  �   	�  \i  �X
 j  ^W  ��   �T��  �i  �X��  �=  �X# 9��  j�  �i  �gA     �       ���  �   ��  �   	�  \i  �X^W  ��   �P��  �i  �X��  �=  �X#     �h  %g  �e  �(  �]A     x      �l  F q3  ��  '�=  ��t ')X   ����  ';  ��~à  (n  ��vsp (%]5  ��~�`A     �      Hk  s @	�-  �h��  D5   �dkaA     J       �j  i I5   �` �aA     -       k  i K5   �\ �aA     )       'k  i N5   �X bA     R       i P5   �T  ]bA     �      s U	D0  �H��  Y5   �DCcA     V       �k  i ^5   �@ �cA     -       �k  i `5   �� �cA     )       �k  i c5   �� �cA     V       i e5   ��   �(  ٭@           ��l  F �#  �t  '#  ��fo <  ����  C=1  ��p �l  �`�@     �      i �   �h�@     �      c 	�  �_   �  �(  �^@     *       �m  F �#  �2  � �-  �hfo �7  �`��  �>=1  �X !  m  >m  �  7  %�"  ��  %�  �%0  %&8  �6�    :m  ;R  am  Xp@     K       ��m  m  �hm  �d%m  �X1m  �P �	  �m  �f@     7      ��m  	�  m7  �H�N  �7  �@�2  �"7  ��72  �7  �X �	  �m  �e@     7      �6n  	�  m7  �H�N  �7  �@�2  �!7  ���l  �7  �X �	  Un  �d@     j       �qn  	�  m7  �h�2  |7  �` �  �n   o@     7      ��n  	�  :7  �H�N  ��6  �@�2  �"�6  ��72  ��6  �X D  �_@            ��n  �  E�6  �h �  o  �m@     7      �Po  	�  :7  �H�N  ��6  �@�2  �!�6  ���l  ��6  �X *  u_@            �{o  �  B�6  �h 6  �o  :e@     (       ��o  	�  W7  �ha �!7  �`b �17  �X `  �o  ~m@     j       ��o  	�  :7  �h�2  |�6  �` !�  
p  p  �  /7   *�o  �`  7p  4Y@            �@p  
p  �h !�  Np  |p  �  7  %�  �0  %&8  �)�   %X[  �65    :@p  &Z  �p  m@     d       ��p  Np  �hWp  �`cp  �Xop  �T 6�  �p  �d@            ��p  	�  m7  �h Z
  q  �j@     �      �kq  	�  m7  ���2  7  ���   7  ���N  7  �X�R  7  �P�7  7  �H �  oj@            ��q  �  I7  �h �
  �q  h@     a      �r  	�  m7  ���2  D7  ��f?  D$7  ���l  E7  �X72  F7  �P�N  Z7  �H �  �f@            �@r  �  E7  �h z  be@            �kr  �  B7  �h 6�  �r  d_@            ��r  	�  :7  �h $)  �]A     d       �	s  F �1  ��  �GE  �ht �*X   �d��  �<  �Xà  �n  �`vsp �%]5  �P V)  �UA     �      ��x  F �1  ��  pGE  ��t p(X   ����  p:  ��à  qn  ��vsp q%]5  ��#VA           �s  ^W  w  �X "p  �s  3�  ��s  �@ <;�  �Iu  b�  W�  �s  �s  �s  �s  �s  )�s   b�  Z�  t  t  �s  t  t  
�s   7b�  ��  -t  3t  �s   a�  �  Dt  Ot  �s  5    #��  ��i   #��  �GE  8E�  v�  �t  �QA     �       ��t  g�  �   g�  �   	�  �t  �X
�x  ^W  ��   �T��  �i  �X��  GE  �X# 9��  3�  u  �PA     �       �g�  �   g�  �   	�  �t  �X^W  ��   �P��  �i  �X��  GE  �X#  "�  du  3�  �du  �� <��  ��v  b�  g�  �u  �u  �u  du  �u  )du   b�  ]�  �u  �u  �u  �u  �u  
du   7b�  6�  �u  �u  �u   a�  ��  �u  �u  �u  5    #��  ��i   #��  �GE  8E�  ��  Ev  NSA     �       ��v  ��  �   ��  �   	�  Qv  �X
�x  ^W  ��   �T��  �i  �X��  GE  �X# 9��  ��  �v  tRA     �       ���  �   ��  �   	�  Qv  �X^W  ��   �P��  �i  �X��  GE  �X#  "�  	w  3�  �	w  �� H�  �b�  �  $w  ;w  )w  	w  4w  )	w   b�  ��  Lw  bw  )w  Vw  \w  
	w   7b�  ��  sw  yw  )w   a�  }�  �w  �w  )w  5    #��  ��i   #��  �GE  8E�  d�  �w  �TA     �       �$x  ��  �   ��  �   	�  �w  �X
�x  ^W  ��   �T��  �i  �X��  GE  �X# 9��  �  Ux  $TA     �       ���  �   ��  �   	�  �w  �X^W  ��   �P��  �i  �X��  GE  �X#   \w  �u  t  �)  KJA     x      ��z  F �1  ��  'GE  ��t ')X   ����  ';  ��~à  (n  ��vsp (%]5  ��~MA     �      �y  s @	�-  �h��  D5   �d�MA     J       oy  i I5   �` NA     -       �y  i K5   �\ @NA     )       �y  i N5   �X iNA     R       i P5   �T  �NA     �      s U	D0  �H��  Y5   �D�OA     V       +z  i ^5   �@ �OA     -       Pz  i `5   �� $PA     )       uz  i c5   �� MPA     V       i e5   ��   �)  �IA     d       �
{  F �2  ��  ��I  �ht �*X   �d��  �<  �Xà  �n  �`vsp �%]5  �P �)  2BA     �      ���  F �2  ��  p�I  ��t p(X   ����  p:  ��à  qn  ��vsp q%]5  ���BA           �{  ^W  w  �X "�  �{  3�  ��{  �@ <;�  �J}  b�  �  �{  �{  �{  �{  �{  )�{   b�  �  |  |  �{  |  |  
�{   7b�  ^�  .|  4|  �{   a�  )�  E|  P|  �{  5    #��  ��i   #��  ��I  8E�  k�  �|  �=A     �       ��|  g�  �   g�  �   	�  �|  �X
��  ^W  ��   �T��  �i  �X��  �I  �X# 9��  m�  }  "=A     �       �g�  �   g�  �   	�  �|  �X^W  ��   �P��  �i  �X��  �I  �X#  "  e}  3�  �e}  �� <��  ��~  b�  M�  �}  �}  �}  e}  �}  )e}   b�  ��  �}  �}  �}  �}  �}  
e}   7b�  ��  �}  �}  �}   a�  М  �}  �}  �}  5    #��  ��i   #��  ��I  8E�  0�  F~  �?A     �       ��~  ��  �   ��  �   	�  R~  �X
��  ^W  ��   �T��  �i  �X��  �I  �X# 9��  X�  �~  �>A     �       ���  �   ��  �   	�  R~  �X^W  ��   �P��  �i  �X��  �I  �X#  "@  
  3�  �
  �� H�  �b�  .�  %  <  *  
  5  )
   b�  L�  M  c  *  W  ]  

   7b�  ��  t  z  *   a�  ��  �  �  *  5    #��  ��i   #��  ��I  8E�  ��  �  \AA     �       �%�  ��  �   ��  �   	�  �  �X
��  ^W  ��   �T��  �i  �X��  �I  �X# 9��  ��  V�  �@A     �       ���  �   ��  �   	�  �  �X^W  ��   �P��  �i  �X��  �I  �X#   ]  �}  |  *  �6A     x      ���  F �2  ��  '�I  ��t ')X   ����  ';  ��~à  (n  ��vsp (%]5  ��~f9A     �      ف  s @	�-  �h��  D5   �d(:A     J       p�  i I5   �` r:A     -       ��  i K5   �\ �:A     )       ��  i N5   �X �:A     R       i P5   �T  ;A     �      s U	D0  �H��  Y5   �D <A     V       ,�  i ^5   �@ V<A     -       Q�  i `5   �� �<A     )       v�  i c5   �� �<A     V       i e5   ��   �$  ��  �6A     *       �ۂ  T X   	�  21  �h�2  	X   �d P*  6A     d       �M�  F C1  ��  �O  �ht �*X   �d��  �<  �Xà  �n  �`vsp �%]5  �P �*  f.A     �      �Ԉ  F C1  ��  pO  ��t p(X   ����  p:  ��à  qn  ��vsp q%]5  ���.A           �  ^W  w  �X "P  �  3�  ��  �@ <;�  ���  b�  l�  "�  9�  '�  �  2�  )�   b�  ��  J�  `�  '�  T�  Z�  
�   7b�  3�  q�  w�  '�   a�  k�  ��  ��  '�  5    #��  ��i   #��  �O  8E�   �  �  0*A     �       �"�  g�  �   g�  �   	�  ��  �X
��  ^W  ��   �T��  �i  �X��  O  �X# 9��  ��  S�  V)A     �       �g�  �   g�  �   	�  ��  �X^W  ��   �P��  �i  �X��  O  �X#  "�  ��  3�  ���  �� <��  �2�  b�  E�  ǅ  ޅ  ̅  ��  ׅ  )��   b�  M�  �  �  ̅  ��  ��  
��   7b�  ��  �  �  ̅   a�  �  -�  8�  ̅  5    #��  ��i   #��  �O  8E�  ��  ��  �+A     �       �ǆ  ��  �   ��  �   	�  ��  �X
ڈ  ^W  ��   �T��  �i  �X��  O  �X# 9��  3�  ��  +A     �       ���  �   ��  �   	�  ��  �X^W  ��   �P��  �i  �X��  O  �X#  "�  M�  3�  �M�  �� H�  �b�  ��  h�  �  m�  M�  x�  )M�   b�  �  ��  ��  m�  ��  ��  
M�   7b�  k�  ��  ��  m�   a�  ��  ·  ه  m�  5    #��  ��i   #��  �O  8E�  ��  *�  �-A     �       �h�  ��  �   ��  �   	�  6�  �X
Ԉ  ^W  ��   �T��  �i  �X��  O  �X# 9��  ��  ��  �,A     �       ���  �   ��  �   	�  6�  �X^W  ��   �P��  �i  �X��  O  �X#   ��  ��  Z�  �*  �"A     x      �܊  F C1  ��  'O  ��t ')X   ����  ';  ��~à  (n  ��vsp (%]5  ��~�%A     �      �  s @	�-  �h��  D5   �d[&A     J       ��  i I5   �` �&A     -       ׉  i K5   �\ �&A     )       ��  i N5   �X �&A     R       i P5   �T  M'A     �      s U	D0  �H��  Y5   �D3(A     V       o�  i ^5   �@ �(A     -       ��  i `5   �� �(A     )       ��  i c5   �� �(A     V       i e5   ��   l  ��  �"A     ;       ��  	�  �-  �h �/  5�/  �"A            �>�  T �-  x 
.�  �h �*  �!A     �       ���  Rr  i�-  �H �  i.�-  �@�!A     0       ��  tmp o5   �\ @"A     0       tmp s5   �X  �8  ݋  �A     �      �L�  	�  �8  ��}t X   ��}��  /  ��}à  Jn  ��}�  \�  	8TB     � A     |       p 4	�-  �X  +_   \�  /�   
 
L�  M8  ��  �A     )       ���  	�  �8  �hc X   �d l8  ��  dA     1       ���  	�  �8  �hc �-  �`n )�   �X f%  ��  �V@     &       ��  	�  '1  �ha  	M�-  �` W#  +  c�@     I       �k�  T #  F �#  �2  2�  �H��  2!=1  �@ �-  ++  TV@     E       ���  T �-  F �#  �2  2k�  �H��  2!=1  �@ !�#  ɍ  ߍ  �  21  %Ca  	!1   *��  �n  �   V@     4       ��  ɍ  �hҍ  �` �  2�   ^@     �       �o�  	�  �7  �H  !=�   �@v6  '0  �Xfra )�6  �P 7  ��  �Y@     �       ���  	�  �7  �X�2  �7  �P� �7  �h �&  ڎ  �]@     L       ��  	�  9  �h �  �  �\@     �       �3�  	�  b7  �X�2  ��6  �P� ��6  �h s  R�  �[@     D      ��  	�  �7  ����  95   ��v6  0  �@�  	�   ���H  
	�   �Xslb 7  ��Rr  )7  �Pk\@     ^       off �   �H�\@     >       �2  )7  ��   �&  '�  �X@     O       �4�  	�  9  �h �	  S�  D[@     X       �o�  	�  m7  �X� p7  �h :
  ��  �Z@     �       ��  	�  m7  �H�2  7  �@v  7  �h�\  7  �`�Z@     I       �l  7  �X  6�  �  JY@     I       �5�  	�  7  �Xp ��   �Padr �	�   �h !�&  C�  V�  �  9     <    :5�  �  y�  8W@     '       ���  C�  �h !+&  ��  ��  �  9  %�  .-   :��  dh  ɑ  W@     2       �ڑ  ��  �h��  �` �6  ��  �A     �      �h�  	�  �6  ��}t X   ��}��  /  ��}à  Jn  ��}�  \�  	SB     TA     |       p 4	�-  �X  `6  ��  bA     )       ���  	�  �6  �hc X   �d 6  ��  0A     1       ��  	�  �6  �hc �-  �`n )�   �X �5  �  XA     �      �u�  	�  *6  ��}t X   ��}��  /  ��}à  Jn  ��}�  \�  	�RB      A     |       p 4	�-  �X  �5  ��  .A     )       ���  	�  *6  �hc X   �d �5  ͓  �A     1       ���  	�  *6  �hc �-  �`n )�   �X 5  �  $A     �      ���  	�  X5  ��}t X   ��}��  /  ��}à  Jn  ��}�  \�  	�RB     �A     |       p 4	�-  �X  !�  ��  ��  U �-  �  �-  %`?  %�-   :��  |�  ה  �A     N       ��  U �-  ��  �X��  �P �  �  �A     )       �$�  	�  �-  �h�-  = �  �` !L  2�  H�  �  �-  %�2  �-   :$�  `�  k�  ^A     N       �|�  2�  �X;�  �P �4  ��  4A     )       ���  	�  X5  �hc X   �d �4  ԕ  A     1       ���  	�  X5  �hc �-  �`n )�   �X 5�/  �A            �+�  T �-  x 
*�-  �h !�  9�  L�  �  �-     <    *+�  =e  o�  V@            �x�  9�  �h !�  ��  ��  �  �-   *x�  �H  ��  V@            ���  ��  �h U+  &	A     �      ���  A 8  ��  �8  ��~s �)�-  ��~vsp �7]5  ��~h	A     �      ��  �  ��à  n  �`v	A     c       `�  n ��   �h eA     ~       ��  w �5   �d �A     �       `?  	5   ��   !)8  ��  ؗ  �  �8  %��  <4  Evsp ,]5   *��  ۢ  ��  �A     *       ��  ��  �h��  �`˗  �X /$  3�  LK@     ,       �H�  	�  21  �h\#  �  �$  n�  �@     6       ���  T #  	�  21  �h�2  	#  �P %  ��  "K@     )       �̘  T �-  	�  21  �h�2  	�-  �` !$  ژ  �  �  21     <    *̘  'F  �  K@            ��  ژ  �h H%  8�  �J@     )       �E�  	�  '1  �` �  d�  
O@     �      �u�  	�  �7  ��~��  �6�   ��~JO@     �      /�  ��  �5   �\bkt ��7  �PsZ  ��%  ���2  )7  ���O@     *      ��  slb 	7  �H �P@     �      slb 	7  �@�\  �%  ��  �R@     �         6�   ��fra 7�6  ���\  9�%  ��~  |+  0A     �      �a�  A /6  ��  �/6  ��~s �)�-  ��~vsp �7]5  ��~rA     �      ��  �  ��à  n  �`�A     c       �  n ��   �h oA     ~       <�  w �5   �d �A     �       `?  	5   ��   !<6  o�  ��  �  �6  %��  �2  Evsp ,]5   *a�  �  ��  A     *       �͛  o�  �hx�  �`��  �X �   5�+  �A     +       ��  T �   a 	͛  �hb 	#͛  �` �+  �@     �      ���  A c5  ��  �c5  ��~s �)�-  ��~vsp �7]5  ��~P�@     �      ��  �  ��à  n  �`^�@     c       ��  n ��   �h M�@     ~       ל  w �5   �d ��@     �       `?  	5   ��   !p5  
�  ,�  �  *6  %��  f3  Evsp ,]5   *��  )�  O�  ��@     *       �h�  
�  �h�  �`�  �X i��  %5   x�@     �      ��  H ��  �  %��  ��y��  fmt %-�-  ��yת  %A�  ��y��  &	5   �l��@     t      ��  8�   �`K.  B5   �\8  [�   �X.�  \�   �T"�  E�  c 3X   ��~ "   m�  res �$0  �Hc �X   �G "0  ��  res �$0  ��c �X   �� "`  ��  res �$0  ��c �X   �� "�  ��  ��  �M   ��~c �X   ����  �5   �� "�  7�  ��  	M   ��~c 
X   ����  5   �� "�  ��  ��  5   ����  �  ��z��  5M   ��~��  65   ��c 7X   ��l�@     F       c /#X   ��  ��@     @      ��  res F$0  ��c GX   ��~��  _-�  ��~ F   ��  d�-  ��~   �   +X   -�  ��     �   �+  �@     �      ��  A �4  ��  ��4  ��~s �)�-  ��~vsp �7]5  ��~Z�@     �      ��  �  ��à  n  �`h�@     c       נ  n ��   �h W�@     ~       ��  w �5   �d ��@     �       `?  	5   ��   !�4  -�  O�  �  X5  %��  �1  Evsp ,]5   *�  ��  r�  ��@     *       ���  -�  �h6�  �`B�  �X i��  %5   ��@     �      �8�  H �  �  %ơ  ��y�  fmt %-�-  ��yת  %A�  ��y��  &	5   �l��@     t      ��  8�   �`K.  B5   �\8  [�   �X.�  \�   �T"P  h�  c 3X   ��~ "�  ��  res �$0  �Hc �X   �G "�  ��  res �$0  ��c �X   �� "�  �  res �$0  ��c �X   �� "  �  ��  �M   ��~c �X   ����  �5   �� "@  Z�  ��  	M   ��~c 
X   ����  5   �� "p  أ  ��  5   ����  �  ��z��  5M   ��~��  65   ��c 7X   ����@     F       c /#X   ��  ��@     @      �  res F$0  ��c GX   ��~��  _-�  ��~ F�  ��  d�-  ��~   5,  �U@     +       �u�  T �   a ͛  �hb #͛  �` !l  ��  ��  �  �-  %�-  *�-   :u�  �b  ��  �C@     V       �ͤ  ��  �h��  �` 6  �  ��@            ���  	�  �-  �h !�  �  �  �  �-     <    :��   Y  =�  �C@            �F�  �  �h !�  T�  ^�  �  �-   :F�  �@  ��  �C@     #       ���  T�  �h �  aM   ��@     2       �٥  M   �h5   �d�  �X�  �  	PTB      +_   �  /�    
٥  R�  ,�   L�@     ;      ���  u ,$w0  ��|  ,3�   ��|��  ,@�   ��|)�  ,M�  ��|� -1  �P��@     �       ��  �_  4
�   �hF�  ?�  6�   ��}  �@     �       i G�   �`��@     �       �_  H�   �XF   ?�  J�   ��}    ��  ��   �@     ;      �
�  u ��   ��|  �,�   ��|��  �9�   ��|)�  �F�  ��|� �1  �P��@     �       ��  �_  �
�   �hF�  ?�  �   ��}  D�@     �       i �   �`]�@     �       �_  �   �XF�  ?�  �   ��}    ��  �5   ��@     D       �L�  4�  ��  �Xd ��  �o T{�  �5   ��@            ���  )�  ��  �h T��  �5   ��@            ���  )�  ��  �h j�  ���@            ��  )�  ��  �h ?�  �5   4�@     [       ��  �  ��~ k>�  ���@     [       �:�  �  ��~ k&�  �~�@     [       �c�  �  ��~ V�  �5   ��@     �       �ة  out �ة  ����  �'�-  ��ת  �>�  ��vs �S  �@p �q3  �� M   W�  �5   /�@     �       �G�  out �ة  ��~��  �&�-  ��~-ת  �
�   ��~�&  �5   ��~ ڼ  �		  ��@     6       ���  
% �ة  �hn �'��  �`ݼ  �.5   �\)�  �;�  �P�  Ҫ  	(TB      �   +_   Ҫ  /�    
ª  ��  �		  :�@     �      �Z�  
% �ة  ��~n �&��  ��~)�  �/�  ��}u �M   �X�}  �	�   �Pk �	�   �H �  �B@     �       ��    S0�   ��tc U�   �`e ^�   �Xf _�   �Pip `�   �His a�   �@�B@     :       i W�   �l  5�  $B@            �Y�  idx D6�   ��tc F�   �hs K5   �dip L�   �Xis M�   �Pf N�   �H �  �5   ��@     �       ���  �  ��-  �X�^  �5   �l Tp�  �5   ��@            �Ѭ  )�  ��  �h T
�  �5   ��@            ��  )�  ��  �h j��  �y�@            �5�  )�  ��  �h ƶ  ~5   J�@     /       ���  4�  ~�  �ht�  ~)��  �`�  ��  	TB      �  +_   ��  /�    
��  ��  y5   �@     /       ���  4�  y�  �ht�  y9�  �`�  ��  	TB      �  D��  q�  u�   ��@     2       �m�  u uw0  �h  u*�   �`��  u8�   �X)�  uE�  �P Y�  q�   ��@     2       �Ѯ  u q�   �h  q#�   �`��  q0�   �X)�  q=�  �P ��  oH  ��@     .       ��  H  �l�  �`�  ��  	TB      �  nH  _�@     *       �W�  O0  �l�  Ҫ  	�SB      !�  mH  1�@     .       ���  O0  �l�  �`�  ��  	�SB      +_   ��  /�    
��  S�  lH  �@     #       ��  �  Ҫ  	�SB      M�  kH  ��@     +       �)�  �  �h�  ��  	�SB      ��  j5   ��@     .       �p�  �  �h5   �d�  ��  	�SB      4�  i5   ��@     /       ���  J0  �h�  �`�  ǰ  	�SB      +_   ǰ  /�    
��   �  hH  X�@     .       ��  O0  �l�  �`�  ǰ  	�SB      ��  g
b�  &�@     2       �b�  h�  �h5   �d�  �X�  ǰ  	�SB      O0  Db�  L�  fH  ��@     +       ���  �  �h�  ǰ  	�SB      $�  M5   �@     �       �C�  �  M�-  ��� N1  �`�_  P	�   �hlen Q	�   �X۩  ^	�   �Pt�@     O       ?�  S
�   �H  ��  I5   �@            �u�  c I5   �l ��  F5   ��@     $       ���  c F5   �l ��  B5   ��@     "       ��  c B5   �l4�  B�  �` m�  <5   x�@     I       �9�  c <5   �\4�  < �  �Pd =X   �o lx�  85   `�@            �l>�  45   H�@            ��  05   .�@            ���  4�  0�  �h ��  ,5   �@            �߳  4�  ,�  �h #�  (5   ��@     %       �#�  �  ("�-  �h4�  (;�  �` ɠ  #5   ��@     P       �g�  �  #+�-  �h4�  #D�  �` ��  5   }�@     "       ���  c 5   �l4�  �  �` l�  5   2�@     K       ���  c 5   �\4�  !�  �Pd X   �o s�  �M   ]�@     �       ���  u �S   �X�7  �-�   �P4�  �H�  �H�  ��  	�SB     ��@     �       i ��   �h��@     �       c �5   �d   �  �5   �@     D       ��  4�  ��  �Xc �X   �gܓ  ��   �h _�  �5   ��@     /       �9�  J0  �h�  �`�  ��  	�SB      8�  �5   ��@     /       ���  J0  �h�  �`�  Ҫ  	�SB      ɜ  �5   C�@     x       ���  J0  ��~-�  ǰ  	�SB      y�  �5   ��@     x       ��  J0  ��~-�  ��  	�SB      �  �5   ��@     7       �Y�  h�  �h�   �`J0  �X�  �P�  Ҫ  	�SB      R�  �5   ]�@     7       ���  h�  �h�   �`J0  �X�  �P�  ��  	pSB      +_   ��  /�   	 
��  �  �5   �@     x       ��  h�  ��~�   ��~J0  ��~-�  ��  	hSB      S�  �5   m�@     x       �k�  h�  ��~�   ��~J0  ��~-�  Ҫ  	XSB      ǜ  �5   :�@     3       ���  �  �hJ0  �`�  �X�  Ҫ  	HSB      w�  �5   �@     3       �	�  �  �hJ0  �`�  �X�  ��  	8SB      Ȝ  �5   ��@     x       �S�  �  ��~J0  ��~-�  ��  	0SB      x�  �5   �@     x       ���  �  ��~J0  ��~-�  Ҫ  	 SB      A�  �5   �@     3       ��  u �$�-  �h��  �C�-  �`ת  �Z�  �X�  ��  	SB      y�  �5   Y�@     �       �y�  u �S   ����  �>�-  ��ת  �U�  ��vs �S  �@p ��1  �� �  �5   w�@     �       � �  u � S   ��~�7  �/�   ��~��  ��-  ��~ת  �1�  ��~vs �S  ��p ��2  �� �  �5   H�@     /       �W�  ��  �#�-  �hת  �:�  �`�  ǰ  	�RB      �  �5   �@     /       ���  ��  �$�-  �hת  �;�  �` ^�  �5   ��@     `       �S�  4�  ��  �H��  �=�-  �@ת  �T�  ��� �1  �h��	B�  U��  �  (�  �  ��  5    U��  5�  F�  �  ?�  )��   U��  S�  i�  �  ]�  c�  
��   U��  v�  |�  �   m��  �X   ��  ��@     b       �μ  	�  �  �Xc �	X   �o�  ��   �` m?�  �X   ��  ^�@     [       �%�  	�  �  �X
�  c �	X   �o�  ��   �` #� �1   #!�  �5    �  ���  �P ��  �5   ~�@     }       �Ƚ  4�  ��  ����  �>�-  ��ת  �U�  ��vs �S  �@p �C1  �� B�  �5   ��@     �       �Q�  u �#�-  ��}��  �B�-  ��}-���  V��  '�  8�  ,�  �  5    V��  F�  W�  ,�  P�  )�   V��  e�  {�  ,�  o�  u�  
�   V��  ��  ��  ,�   n��  �X   ��  b�@            �ľ  	�  ��  �h n?�  �X   �  v�@     0       ���  	�  ��  �h
,�   @u ��-   @!�  �5    �  ��  ��~ת  ��   ��~�&  �	5   ��~ X�  z5   ��@     �       ���  u zS   ��~��  z=�-  ��~-ת  {
�   ��~�&  }5   ��~ �  s5   ��@     �       �4�  u sS   ��~�7  s.�   ��~��  sO�-  ��~-ת  t
�   ��~�&  v5   ��~ `�  o5   ~�@     x       �}�  ��  o"�-  ��~-�  ��  	�RB      ���  Զ@     �       ���  ��  �   �h  0�   �di I0  �X =��  �5   �@     �       � �  ��  �#�-  ��~-ת  �
�   ��~�&  �5   ��~ =_�  �5   i�@     �       ���  4�  ��  ��~��  �<�-  ��~-ת  �
�   ��~�&  �5   ��~ =��  �5   ��@     �       ���  4�  ��  ��~��  �=�-  ��~-ת  �
�   ��~�&  �5   ��~ ��  ���@     2       �9�  4�  ��  �hu �7S   �`�  ǰ  	�RB      =1�  ��  P�@     3       ���  H	  �&�-  �h  �G�-  �`4�  �^�  �X�  ��  	�RB      =P�  �M   %�@     +       ���  u �M   �h�  ǰ  	�RB      =��  ��  �@     #       ��  �  ��  	�RB      =^�  �5   ͳ@     5       ���   �  �5   �lw�  �(�-  �`��  �65   �h5�  �L�-  �X�  Ҫ  	�RB      =�  �5   3�@     �       ���  {�  ��-  �X5�  �*�-  �P�  ǰ  	�RB     ��@     ;       e �	5   �l  =�l  �5   �@     +       �A�  H	  ��-  �h�  ǰ  	�RB      �3  `�  ��@     O       ���  	�  B4  �Xstr ��-  �Pn �&�   �H��@     8       i ��   �h  �3  ��  8�@     S       ��  	�  B4  �Xstr ��-  �PH�@     @       i ��   �h  �3  !�  ��@     L       �;�  	�  B4  �hc �X   �d �3  Z�  ��@     	      ���  	�  B4  �H�  ǰ  	CTB     �@     �       ��  �	�   �h��  �	M   �P  !~3  ��  ��  �  B4   *��  ��  ��  ��@     .       ���  ��  �h 3  �  d�@     O       �U�  	�  l3  �Xstr ��-  �Pn �&�   �Hx�@     8       i ��   �h  �2  t�  �@     S       ���  	�  l3  �Xstr ��-  �P �@     @       i ��   �h  6�2  ��  ��@     Q       ���  	�  l3  �hc |X   �d !�2  ��  �  �  l3  %u yM   %�Q  y&�    *��  �  ;�  ��@     6       �T�  ��  �h��  �`�  �X 6a2  s�  $�@     c       ���  	�  �2  �Xstr l�-  �Pn l&�   �H4�@     P       i n�   �h  6B2  ��  ��@     g       ��  	�  �2  �Xstr d�-  �P��@     X       i f�   �h  6#2  4�  ��@     <       �N�  	�  �2  �hc _X   �d !2  \�  r�  �  �2  %u \M    *N�  ��  ��  Z�@     &       ���  \�  �he�  �` �1  ��  �@     M       ���  	�  �1  �hstr R�-  �`n R&�   �X �1  �  ��@     e       �)�  	�  �1  �Xstr M�-  �P o1  H�  ^�@     H       �b�  	�  �1  �hc HX   �d !P1  p�  ��  �  �1  %4�  E�   *b�  	�  ��  8�@     &       ���  p�  �hy�  �` !#  ��  ��  �  r0  ou !w0  o  !(�    *��  ,t  �  N�@     *       �(�  ��  �h��  �`��  �X 9  G�  2A@     6       �q�  	�  �-  �`c 63p  �\�  7  �h p�  2��  ��  �  �-     <    :q�    ��  A@            ���  ��  �h �  p�  2��  ��  �  �-  ��   :��  �  
�  ~@@     �       ��  ��  �h��  �` !  )�  3�  �  �-   :�  a  V�  "@@     \       �_�  )�  �h �F  nH  �   @@            ���    #�   �hp /�   �` 6�,  ��  B@            ���  	�  #-  �h �,  ��  �A@     B       ��  	�  #-  �h�  �  	 TB      +_   �  /�    
�  5�  �A@            �L�  x )�   �h !�  Z�  d�  �  V,   *L�  �b  ��  hA@     Q       ���  Z�  �h q	  �%  "q�  �%  " �   �(  	  1�  	  ޖA     �      ��  ��  �9   -N    L   int �3  _   j   _   �  j   �Q  _   2N  	�  
��  _   H�A     H       ��   ��  e   �Xsrc <�   �Pn 9   �h q   �   
s�  �   �A     7       �C  ��  �   �hsrc 'C  �`len 3-   �X I  
��  L   ��A     ]       ��  e L   �\u _   �P��  ,-   �Hs _   �h (�  �_   t�A     @      ��  e �L   �\s ��   �h ��  �
5  B�A     2       �5  5  �h@  �d-   �X�  \  	(^B      @  5  �+  @  q   \  9    L  ��  �-   �A     +       ��  �  �h�  �  	^B      G  �  q   �  9    �  �  �
5  ��A     f       �9  s �!�  �Xc �,@  �T  �6-   �H��  ��  �`ȢA     H       i �-   �h  ��  �
5  ~�A     3       ��  ;  �h�  �`�  �X�  �  	^B      5  �  ��  �
5  O�A     /       ��  �  �h�  �`�  �  	^B      *�  �-    �A     /       �  �  �h�  �`�  �  	^B      ��  �
5  �A     .       �d  �  �h@  �d�  \  	 ^B      d�  �
5  áA     /       ��  �  �h�  �`�  \  	�]B      ��  �-   ��A     /       ��  �  �h�  �`�  \  	�]B      l�  �
5  f�A     .       �6  �  �h@  �d�  �  	�]B      ��  �L   3�A     3       ��  �  �h�  �`-   �X�  \  	�]B      F�  �L    �A     3       ��  ;  �h�  �`-   �X�  \  	�]B      {�  �L   ͠A     3       �   �  �h�  �`-   �X�  \  	�]B      �  �L   ��A     /       �f  �  �h�  �`�  \  	�]B      ��  �L   o�A     /       ��  �  �h�  �`�  �  	�]B      ��  �
5  <�A     3       ��  ;  �h�  �`-   �X�  \  	�]B      ��  �
5  �A     /       �@  ;  �h�  �`�  �  	�]B      ��  �
5  ڟA     3       ��  5  �h�  �`-   �X�  �  	�]B      q   �  9    �  V�  �
5  ��A     3       ��  ;  �h�  �`-   �X�  \  	�]B      ��  �
5  t�A     3       �?  ;  �h�  �`-   �X�  \  	�]B      ��  �
5  E�A     /       ��  ;  �h�  �`�  �  	�]B      �  ��  �A     2       ��  �  �h�  �`L   �\�  �  	�]B      (N  ��  �9   �A     2       �(	  �  �h�  �`L   �\�  \  	�]B       �  �v	  ��A     2       �v	  �  �h�  �`L   �\�  \  	x]B      ,  �  ��	  }�A     2       ��	  �  �h�  �`L   �\�  �  	p]B      1  �  �
  N�A     /       �
  �  �h�  �`�  \  	h]B      �  ��  �e
  �A     /       �e
  �  �h�  �`�  �  	^]B      ^  ��  ��
  �A     /       ��
  �  �h�  �`�  �  	W]B      �  ��  �_   ��A     \       �  s ��   �Xc �$L   �Ti �	-   �h ��  �_   e�A     /       �U  s �e   �hZ�  �9�   �`�  �  	P]B      ?�  �_   ��A     �       ��  s ��   �H��  �)�   �@��A     �       i �-   �hܜA     x       $�  ��  �g��A     a       j �-   �X    oF  �  �-   E�A     m       �F  s ��   �X�  �*�   �Pn �	-   �h N�  �_   ՛A     p       ��  s ��   �Xc �"L   �T��  �	-   �`��A     J       i �-   �h  f�  �_   g�A     n       ��  s ��   �X�  �*�   �Pn �	-   �h ��  }-   ��A     m       �I  s }�   �X�  }+�   �Pn ~	-   �h ��  r_   ��A     i       ��  s r�   �Xc r!L   �Ti s	-   �h �  k�   8�A     Y       �  s kC  �Xc k!L   �T  k+-   �H��  l  �`O�A     ;       i m-   �h    �    �  f-   �A     3       ��  ��  f!e   �hsrc f>�   �`�7  fJ-   �X�  \  	H]B      ^�  UL   ~�A     �       �  a U�   �Xb U(�   �P�7  U2-   �Hi V	-   �h��A     k       ��  Z  �g��  [  �f  ��  PL   Y�A     %       �H  a P�   �hb P(�   �` 8�  @L   �A     r       ��  a @�   �Xb @'�   �Pi A	-   �h��A     Z       ��  C  �g��  D  �f  ��  5L   u�A     r       �]  a 5C  �Xb 5'C  �P  51-   �H��A     [       i 6-   �h��A     B       ��  7  �g��  8  �f   ��  (_   �A     �       ��  ��  ( e   �Hsrc (=�   �@�7  (I-   ��q  )_   �h�
  *�   �`i ,	-   �X 1�  $_   ��A     ;       �  ��  $e   �hsrc $<�   �` ��  _   1�A     �       ��  ��   e   �Hsrc 2�   �@�7  >-   ��q  _   �h�
  �   �`i 	-   �X ��  _   ޖA     S       ���  e   �Xsrc 1�   �Pq  _   �h�
  _   �`  �5   @*  	  ��  	  P$          0�  ��  
�:   )   -N  1  ,  �  L  �  �  2N  i   �  �  int �     �:   %   4�   �   frg 	�  #  		�   	�i  	�    
}C  	�
  �   ]I  �    �   �-  �      �6   red �C   �Q  0�  �Q  �+  A  G  �   �Q  �*  [  f  �  �   �#  �_  �  ~  �  �  �   �N  �   �R  �  �7  �  \.   �  >*  !�   �R  "�   (    �R  %)  �  '�V  �    T H  �   7^  '
   �  T   �    BD  5�  h 8�_  �  O  �   �N  =j4  �  i  �   �R  B�i  �  �  �   �7  E�N  �  �  �   \.  I�P  �  �  �   >*  L�  �  �  �     P�,  �  �  �     �+  U}O  �  
  �   \G  Z�"  �  %  �   �G  dma  9  ?     �G  g"  S  ^    #   �#  i  )  v  �    #   Rr  o_L  �  �  �     �(  |�^  �  �    �   �e  ��  �  �    �  �   i  ��=  �  	    �  �   �+  ��B    )    �   �l  �0  >  I    �    �2  .A  _  o    �  �    Q:  D�  �  �    �  �    �l  xm  �  �    �    �R  ��6  �  �    �    �  +  �  �    �   �  �         �   �_  #=M  -  8    �   !�1  0Z$  �  R  X     !�1  9mI  �  r  �    �  /  5  5   "  ��   D �  T H  #E3  �5  A �   )  $�'  �y  %��  %��  %��  %�i  %��  %��  &)   �b  �@    *  F  Q   �+  ��m  ?  J  F  �   "�5  �Q  T H  #E3  �5  L Q  A �   �S  5
  h 88Y  �  �  �   �N  =�!  �  �  �   �R  BbJ  �  �  �   �7  E�h  �  �  �   \.  If  �    �   >*  LV/  �  !  �     P�[  �  9  ?  Q   �+  U9  �  Z  �   \G  Z-  �  u  �   �G  d3<  �  �  Q   �G  gn.  �  �  Q  \   �#  itF  b  �  �  Q  \   Rr  o�+  �  �  �  Q   �(  |�j      Q  �   �e  �jK  $  4  Q  �  �   i  �A]  I  Y  Q  �  �   �+  �6  n  y  Q  �   �l    �  �  Q  �    �2  H)  �  �  Q  �  �    Q:  D�  �  �  Q  �  �    �l  x.8  �  	  Q  �    �R  �Ld  	  '	  Q  �    �  �  =	  H	  Q  �   �  �R  ]	  h	  Q  �   �_  #	g  }	  �	  Q  �   !�1  0  �  �	  �	  Q   !�1  9�  �  �	  �	  Q  �  /  h  h   "  ��   D 
  T   #E3  �5  XA �   y  'X  �%��  %�  %�4  %��  %��  %�!  &y   �b  �R%  k
  v
  n  Q   �+  ��  �
  �
  n  �   "�5  �Q  T   #E3  �5  XL Q  A �    �
  ]I  �    �
  2l    (clz �  �     :    T :    )%B  �$�  L3  �   �C  �6   �i  '      8  H�	   8  ��Q  i  ~  �    �   )     8  �&  �  �  �  �   �#  �
[  �  �  �  �  �   qe  �ze  �  �  �  �  �   8  �C   v6  ��   ��  �5   �  ��   H  8  ��	�  &H   8  �i'  D  Y  �  �   )   �    8  �E2  m  x  �     �#  ��G    �  �  �     ��  ��   H�(  �i   L�-  �  P+  ��  X   �>  �	L  �>  �Q*  �  �     �>  �0o        �   �#  ��>  �  3  >    �   �+  �    �  �5  �	�  *�R  ��3  �  r  ;  �  �       �	�    �'  �  �  y   ,+  �	�   �Q  ��  �G  ��   �b  ��  C%  ��Z  �  �  �     +N�  �YV  �    "  �  )    !�&  H
:  �  <  L  �  �  )     ��  z�W  b  m  �  �    Q.  �]  �  �  �  �  )    +�:  -	�c  )   �  �  �   ,�\  :�                         @       -�Z  < p   -kG  = p    =d  D�\  )     i      S  )   0  )    -�&  f�   .�  h5   Oa  k�  �  e  i    .�e  x5   .�&  {5   /]  �5    0�i  ��U  �  �  �  �  �    0�i  �C  �  �  �  �  �    0'  !�C  �  �  �  �  )    �  3      �   �@  :�5  *  5  �  �   �=  �
   �  ��  8  �  +2  �O  �  �	)    Y  ��  (1�^  �  1D=  �   2�   0  }w  �)�  �  �  V  a   }w  ��  �  �  V  g   }w  "��  �    V  m   M|  �s�    "  V  �    +�#  )
n�  s  ;  F  V  �   +ux  �]�  y  _  j  V     +ux  ���  y  �  �  V  �   +%y  2��  y  �  �  V     +%y  6�  y  �  �  V  �   3pop ���  �  �  �  V   >  B��  
    V   +�  H��  �  )  /  V   +�  LC�  �  H  N  �   +  P	?�  )   g  m  �   +o�  T��  �  �  �  �   +d X��  �  �  �  V   +d \��  �  �  �  �   3end ``�  �  �  �  V   3end d��  �      �   +q  h��  y  !  '  V   +q  k��    @  F  �   +$  oJ�  y  _  e  V   +$  r��    ~  �  �   +p  v�    �  �  �  )    +p  y3�  y  �  �  V  )    �}  ��  �  �  V  )    G%  ��   ,�  ��    �	)   �}  �	)   T �  1�-     �  4��     ��  ��  W  ]  �   u �   #  :    #{�  :    5��   �  3get  �  s  �  �  �   6��  %)5   ��  N�  �  �  7�-  �  8a   �  a   T �   9�Z  �+   9A)  �7
  9A)  �7�  2�Z  	�  �c  	�l  :  @  �   �c  	w  U  e  �  �   �   �c  	=  z  �  �  �   :�c  	!zG  �  �  �  �   �c  	#�  �  �  �  �   �c  	(�;  �  �  �  �    +�#  	-4  �  �  	  �     �c  	2�n    $  �   a  	8p;  9  ?  �   +S  	>�&  �  X  ^  �   ++H  	BY0  �  w  �  �  �   �  	G	�   R  	H�  1D=  �      ;�   oF  �  ;�   <   �  =�  =   >;�
  ^P  �  ^P  �b      �   ^P  �#    &  �  �   �#  PK  �  >  I  �  �   �c  �!  ]  c  �   a  �l  w  }  �   ?je  �     �  <�  �  =�  =�  �-  �  @map �7  �   �  �  �  )    A�@   H  �  �  �   )     <�  ��  4  ��  D   ��  �  S�  �   �  BD  �   <9  ��  <�  <�  V  =  =0  C�  =�  =�  =4  C�  <�  <4  <0  �  <  �  <5  �  D�  �  E:    �  �  <  �  <H  �  =  =H  <  �  =�  =  <�    <)    =�  =)  =�   =�  <Q  ;  <�  F  <y  Q  =
  =y  =�  <
  n  <�  =�  D5   �  E:    �  FeW  �  F�i  �  F�  �  FGb  0  G'  >   �GQ5  e   H�:  r     FL    D�  �  E:    Istd  �  ��  &  8    T a   ��  G  8  �  T y   �}  >3  V�  !��  G  t  T y  y   ��  �  a  �  T a  E2   �}  >   <  �  =�  C  =  =L  =�  J
  s�@     1       ��  K�2  Z�  �h L�    D�@     �      �\  M�    ��Nn �  ��Ou �  �XOv �  �POw �  �H L�  {  ��@     �      ��  M�    ��Nn ��  ��Ou ��  �XOv ��  �POw ��  �H P�  �@            ��  T H  K�2  '�  �h P  �@            �&  T   K�2  '�  �h L'	  E  ��@     �      ��  M�  W  ��Nn �  ��Ou �  �XOv �  �POw �  �H L	  �  �@     �      ��  M�  W  ��Nn ��  ��Ou ��  �XOv ��  �POw ��  �H JZ  B�@     1       �  K�2  Z�  �h JO  =x@            �H  K�  =�  �h L�  g  zr@     �      �E  M�    ��Nn x�  ��Q�N  {�  �POs ��  �XQ�R  ��   ��RIs@     �       �  Ox ��  �H Ret@     z       �  Ox ��  �@ Rv@     Q       !  Qf?  ��  �� SZw@     Q       Qf?  ��  ��  J�  Hr@     1       �p  K�2  U�  �h LY  �  �x@     V      ��  M�  W  �XTn ��  �PU�N  ��  �hUd4  ��  �` J�  *r@            ��  K�  L�  �h L    Zx@     H       �>  M�    �XV�2  #�  �PQ� $�  �h P6  r@            �i  K�  8�  �h L	  �  Ƃ@     V      ��  M�    �XTn ��  �PU�N  ��  �hUd4  ��  �` L�  �  �x@            ��  M�    �hV�2  �  �` LH	     �x@            �8   M�  W  �hV�2  �  �` Lh	  W   N|@     H       ��   M�  W  �XV�2  #�  �PQ� $�  �h J�  ��@            ��   K�  =�  �h L�  �   �|@     �      ��!  M�  W  ��Nn x�  ��Q�N  {�  �POs ��  �XQ�R  ��   ��R�}@     �       =!  Ox ��  �H R�~@     z       a!  Ox ��  �@ Rw�@     Q       �!  Qf?  ��  �� SƁ@     Q       Qf?  ��  ��  J?  �|@     1       ��!  K�2  U�  �h J  �|@            �"  K�  L�  �h P�  8|@            �-"  K�  8�  �h LI  L"  2b@     �      ��"  M�    ��V�2  �  ��V�   �  ��Q�N  �  �XQ�R  �  �PQ�7  �  �H J�  b@            ��"  K�  I�  �h Lo  �"  �_@     a      �V#  M�    ��V�2  D�  ��Vf?  D$�  ��Q�l  E�  �XQ72  F�  �PQ�N  Z�  �H WU  d#  �#  X�  �  Y�"  �  Y�  �%�   Y&8  �6)    ZV#  ;R  �#  Xp@     K       ��#  [d#  �h[m#  �d[y#  �X[�#  �P L4  �#  �f@     7      �0$  M�  W  �HK�N  ��  �@K�2  �"�  ��U72  ��  �X L  O$  �e@     7      ��$  M�  W  �HK�N  ��  �@K�2  �!�  ��U�l  ��  �X L�  �$  �d@     j       ��$  M�  W  �hK�2  |�  �` L�  �$   o@     7      �%  M�    �HK�N  ��  �@K�2  �"�  ��U72  ��  �X J�  �_@            �J%  K�  E�  �h L�  i%  �m@     7      ��%  M�    �HK�N  ��  �@K�2  �!�  ��U�l  ��  �X Ji  u_@            ��%  K�  B�  �h \^  �%  :e@     (       �&  M�  A  �hTa �!�  �`Tb �1�  �X L�  4&  ~m@     j       �P&  M�    �hK�2  |�  �` W0  ^&  �&  X�  �  Y�  ��   Y&8  �))   YX[  �6�    ZP&  &Z  �&  m@     d       ��&  [^&  �h[g&  �`[s&  �X[&  �T \!  �&  �d@            ��&  M�  W  �h L�  '  �j@     �      �{'  M�  W  ��V�2  �  ��V�   �  ��Q�N  �  �XQ�R  �  �PQ�7  �  �H J�  oj@            ��'  K�  I�  �h L�  �'  h@     a      �%(  M�  W  ��V�2  D�  ��Vf?  D$�  ��Q�l  E�  �XQ72  F�  �PQ�N  Z�  �H J�  �f@            �P(  K�  E�  �h J�  be@            �{(  K�  B�  �h \�  �(  d_@            ��(  M�    �h W�  �(  �(  X�     ]�(  �`  �(  4Y@            ��(  [�(  �h L)  
)  (X@     �       �i)  M�    �HV�2  �  �@Qv  �  �hQ�\  �  �`S�X@     I       Q�l  �  �X  L�  �)  `W@     �       ��)  M�  �  �XVv6  �;�   �PQ� ��  �h L�  �)   ^@     �       �*  M�  �  �HV  !=)   �@Qv6  '�   �XOfra )�  �P Lv
  0*  �Y@     �       �]*  M�  t  �XV�2  ��  �PQ� ��  �h L	  |*  �]@     L       ��*  M�  �  �h L*  �*  �\@     �       ��*  M�  L  �XV�2  ��  �PQ� ��  �h L�  �*  �[@     D      ��+  M�  �  ��V��  9�   ��Qv6  �   �@Q�  	:   ��Q�H  
	)   �XOslb �  ��QRr    �PSk\@     ^       Ooff )   �HS�\@     >       Q�2    ��   L$  �+  �X@     O       ��+  M�  �  �h L�  �+  D[@     X       �,  M�  W  �XU� p�  �h Ly  0,  �Z@     �       ��,  M�  W  �HV�2  �  �@Qv  �  �hQ�\  �  �`S�Z@     I       Q�l  �  �X  \�  �,  JY@     I       ��,  M�  �  �XTp ��  �P^adr �	:   �h W�  �,  �,  X�  �  X   �    Z�,  �  -  8W@     '       �$-  [�,  �h We  2-  H-  X�  �  Y�  	�   Z$-  dh  k-  W@     2       �|-  [2-  �h[;-  �` LL  �-  �K@     h      �O.  M�  �  ��~VW z0�  ��~Qv6  �:   �XQ�\  �  ��Ofra ��  �POslb ��  �HObkt �y  �@Q�  �	)   ��QsZ  �  ��Q�-  ��  ��Q�2  �  �� PS  J�A     0       �.  T y  Tx *y  �` L�  �.  
O@     �      ��/  M�  �  ��~K��  �6)   ��~RJO@     �      i/  U��  ��   �\^bkt �y  �PUsZ  �  ��Q�2    ��R�O@     *      5/  Oslb 	�  �H S�P@     �      Oslb 	�  �@Q�\    ��  S�R@     �       Q  6:   ��Ofra 7�  ��Q�\  9  ��~  L�  �/  6�A           �J0  M�  \  �HK�}  �4)   �@Uy  �	)   �XU��  ��  �PR��A     l       *0  ^i �)   �h S��A            ^i �)   �`  W�  X0   n0  X�  \  YH%  �)a   ]J0  y�  �0  ��A     >       ��0  [X0  �h[a0  �` WC  �0  �0  X�  �   ]�0  ��  �0  ʧA     .       ��0  [�0  �h \�  1  ��A     *       �!1  M�  \  �hK��  y)   �` \N  @1  ��A            �M1  M�  �  �h LF  l1  ��A     �       ��1  M�  \  �XK�^  �(  �PUW ��  �h \�  �1  �A            ��1  M�  �  �h W�  �1  �1  7�-  �1  8a   X�  �  _a    Z�1  ��  &2  ��A     P       �E2  7�-  &2  8a   [�1  �X`<2  a�1   [�1  �P =�  Pt  ��A            �{2  T a  Tx .E2  �h b��  #��  1�A     a       ��2  ^eq $�2  �`SB�A     M       ^i %)   �hSY�A     /       U�  &�  �X   =J  c��  �   �A     J       �R3  K��  $D  �HK��  =�  �@K�  M�  ��U�  �  �P d~�  i�  �2  ��A     W       ��3  U��  !  	`C      J  �B@     �       �4  K  S0)   ��^tc U:   �`^e ^:   �X^f _:   �P^ip `:   �H^is a:   �@S�B@     :       ^i Wi   �l  P�  $B@            ��4  Tidx D6i   ��^tc F:   �h^s K�   �d^ip L:   �X^is M:   �P^f N:   �H eF  nH  �  @@            ��4  K  #)   �hTp /�  �` \c  �4  B@            ��4  M�  �  �h LI  5  �A@     B       �<5  M�  �  �hf�  L5  	OoB      D�  L5  E:    <5  P�
  �A@            �z5  Tx ):   �h W-  �5  �5  X�  �   ]z5  �b  �5  hA@     Q       ��5  [�5  �h gH  �  "g  �  " �   1  	  ��  	  z�A     �       � �  �  2N  -N  �  �  int 1    �B   %   4e   ��  �B   ,  �  L  de    t�  �  ��  W�  W   �   	  	}    E�  
��  W   �   	}   	X   
<�  '�  	W     �   D�A            ��   1�A            �X  W   �h  *}   �`   �   ��A     �       ��    
}   �hW 
,X  �`�  �  	�oB      �  �  B    �  �  �  �   z�A     3       �o6  W   �l  �   "2  	  ��  	  P)          � ��  �:   )   -N  1  ,  �  L  �  �  2N  i   �  �  int �     	�:   %   
4�   �   frg 	<  #  	�   	�i  �    
}C  	�
  �   ]I  H    �   �-  �      �6   red �C   �Q  0�  �Q  �+  A  G  R   �Q  �*  [  f  R  X   �#  �_  ^  ~  �  R  X   �N  d   �R  d  �7  d  \.   d  >*  !d   �R  "�   (    �R  %BD  5x  h 8�_  R    �   �N  =j4  �  &  �   �R  B�i  �  @  �   �7  E�N  �  Z  �   \.  I�P  �  t  �   >*  L�  �  �  �     P�,  �  �  �     �+  U}O  A  �  �   \G  Z�"  A  �  �   �G  dma  �  �     �G  g"           �#  i    3  >       Rr  o_L  �  V  \     �(  |�^  q  |    �   �e  ��  �  �    �  �   i  ��=  �  �    �  �   �+  ��B  �  �    �   �l  �0  �      �   �2  .A    ,    �  �   Q:  D�  B  R    �  �   �l  xm  h  s    �   �R  ��6  �  �    �   �  +  �  �    �   �  �   �  �    �   �_  #=M  �  �    �   �1  0Z$  A         �1  9mI  A  /  I    �    "  "      �d   !D }  !T �
  "E3  }  !A �   �  #�'  �6  $�\  $�|  $��  $�&  $�@  $��  %�   �b  �@  �  �  .  h   �+  ��m  �    .  �    �5  �h  !T �
  "E3  }  !L h  !A �   �S  5�	  h 88Y  R  \  �   �N  =�!  �  v  �   �R  BbJ  �  �  �   �7  E�h  �  �  �   \.  If  �  �  �   >*  LV/  �  �  �     P�[  �  �  �  9   �+  U9  A    �   \G  Z-  A  2  �   �G  d3<  F  L  9   �G  gn.  `  k  9  D   �#  itF  J  �  �  9  D   Rr  o�+  �  �  �  9   �(  |�j  �  �  9  �   �e  �jK  �  �  9  �  �   i  �A]      9  �  �   �+  �6  +  6  9  �   �l    K  V  9  �   �2  H)  l  |  9  �  �   Q:  D�  �  �  9  �  �   �l  x.8  �  �  9  �   �R  �Ld  �  �  9  �   �  �  �  	  9  �   �  �R  	  %	  9  �   �_  #	g  :	  E	  9  �   �1  0  A  _	  e	  9   �1  9�  A  	  �	  9  �    P  P      �d   !D �	  !T �  "E3  �  X!A �   6  &X  �$��  $��  $��  $�v  $��  $��  %6   �b  �R%  (
  3
  V  h   �+  ��  H
  S
  V  �    �5  �h  !T �  "E3  �  X!L h  !A �    �
  ]I  H    �
  '%B  �$�  L3  �   ��
  �6   �i  '   �
   8  H�	�   8  ��Q  �
    �  �
  �   )     8  �&     +  �  �   �#  �
[  �  C  N  �  �   qe  �ze  A  f  q  �  d   8  ��
   v6  ��   ��  �5   �  �Y   �
  8  ��	^  %�
   8  �i'  �  �  �  �   )   �    8  �E2  �    �  �   �#  ��G  �    )  �  �   ��  ��   H�(  �i   L�-  ��  P+  �Y  X �  (�>  �5  �	�  )�R  ��3  A  �  (  �  �       �	�    �'  �  �  a   ,+  �	k   �Q  ��  �G  ��   �b  �f  C%  ��Z  
    l  �   *N�  �YV  d  .  9  l  )    �&  H
:  d  S  c  l  d  )    ��  z�W  y  �  l  d   Q.  �]  �  �  l  d  )    *�:  -	�c  )   �  �  l   +�\  :�                         @       ,�Z  < p   ,kG  = p    =d  D�\  )   -  i      S  )   G  )    ,�&  f�   -�  h5   Oa  k�  A  |  i    -�e  x5   -�&  {5   .]  �5    /�i  ��U  �  �  �  l  �    /�i  �C  �  �  �  l  �    /'  !�C  �      l  )    �  3  &  ,  l   �@  :�5  A  L  l  �   �=  �
�   �  �k  8  �s  +2  �f  �  �	)    Y  ��  (0�^  3  0D=  k   1��  �  ��  ��  �  �  �   u �   "  :   "{�  :    2F�  Y  3get  \�  �    #  �   4��  %)�   ��  ��  K  Q  5�-  �   !T 3   6�Z  �+   6A)  �7�	  6A)  �7}  7p�  ��  ��  ��  �  �  �   u �   8  :   �"{�  :    9`�  �3get  �     �  �     4��  %)�   ��  �  (  3  :�-  (  ;�     �   !T �
    <�   oF  A  <�   =   >�  >   ?<�
  ^P    ^P  �b  �  �     ^P  �#  �  �    '   �#  PK  -  �  �    '   �c  �!  �  �     a  �l         @je  �     k  =k    >  >k  �-  �  Amap �7  �   X  c  �  )    B�@   H  s  �  �   )     =3  �  ��  #>�
  �  �  Cde  -=�  �  D�  �  E:     >3  =�  �  =�
  >�  >�
  =�  >^  >�  =c  =�    >x  >�  >�   >�  =h  =}  .  =6  9  >�	  >6  >�  =�	  V  =�  a  =�
  l  D5   �  E:    w  FeW  �  F�i  �  F�    FGb  G  F'  U  FQ5  |  F�:  �  FL  �  D�  �  E:    =�  �  D�     G:   � >�
  =�    Hstd  �  ��  =  8  3  !T �   ��  ^  8  h  !T �   �}  >J  ��  !!�  ^  �  !T �  �   U�  m�  �  �  !T �  �   �}  >)   I2  �  �  J�  ?   K�  ��  �  ��A            ��  L�  �h I
    "  J�  \  M�5  �h   N�  �  E  ��A     $       �V  L  �hL  �  I�  d  n  J�     KV  G�  �  p�A            ��  Ld  �h >h  Oj  e�A     
       ��  !T �  Px *�  �h I�  �  �  J�  g   N�  ��    .�A     7       �  L�  �h I�  "  9  J�  4  M�5  �h   N  ��  \  
�A     $       �m  L"  �hL+  �  I�  {   �  J�  r  Q�=  �7�   Nm  ��  �  ��A     {       ��  L{  �XL�  �P I�  �  �  J�  �   K�  �     h�A     %       �	  L�  �h I�    !  J�  �   K	  ��  D  V�A            �M  L  �h R�  l  H�A            �y  S�    �h I  �  �  :�-  �  ;�   J�    T�    Ny  �  �  ��A     P       ��  :�-  �  ;�   L�  �XU�  V�   L�  �P >�  O�  �A            �1  !T �  Px .�  �h R  P  ܫA            �]  S�  �  �h I1  p  ~  5�-  J�  �  W N]  �  �  ��A     ,       ��  5�-  Lp  �hW Xc  �  H�A     R       �  S�  �  �hYv6  (�   �`Y��  8)   �XZ�  #  	KpB      D�  #  E:      X@  J  ��A     Q       ��  S�  �  �XY��  ()   �P[ptr d  �hZ�  �  	GpB      D�  �  E:    �  \��  ��  �  Z�A     �       ��  ]��  (�  	�C     ]��  '�  	�C      >�  Ix      J�  "   K�  ��  1  ��A            �:  L  �h ^F  nH  d  @@            �}  Y  #)   �hPp /d  �` _�
  Y  "_�  Y  " 9   @8  	  I�  	  �*          8 ��  �5   -N  �  �  �  V   2N  V   �  �  int p   1  M  J   frg 8  I  �   �\   �   	4D    
0  {  �2  |p   0  ~m[  �   �   �   /   .    �  p     �=  �g  &  ,  �   �=    A  L  �  �    �=  4H  a  l  �  �   �=  �?  �  �  �  �   �=  *�l  �  �  �  �   �=  0]  �  �  �  �   �=  8�7  �  �  �  p    �#  = A  �      �  �    fF  Q�1  �  )  /  �   fF  T�6  �  H  N  �   \?  X�:  �  g  m  �   �"  \iQ  �  �  �  �   �"  `�:  �  �  �  �   2d  dF  �  �  �  �   ;W  ��  �  �  �   ~  ��    �6  ��  T p    �   �  J~6  
  �    g&      E  �  >  ,  �  L  �   	`pB     ��  �  �_  i    �f  i     V    �   �   w   p     �   �   oF  �    p   p   std  u  �   	J#  `?  	K�  T p   �-   �    �1  	JP  `?  	K�  T p   �-   �    !@  	Nh  �  !@  	NW3  �   "�#    "�?  0  (N  �  �+  �  !  	apB     #de  
c  $B  
+|  -  $'.  
,�R  2  %�^  p     &�6   &�j  &�  &$D  &�7   �  Z  'it 8   'end 8  (fF  Hh  �  L  R  c   C E   �r  �  'it n   'end t  (fF  |o  �  �  �  z   C V    �7  �  'it �   'end �  (fF  �&  �  �  �  �   C �   a�  q$  )4s  rbp  �    �  �  �    r  #�   M�  	/  ��  	�  ��  m�  ^  d  �   *�_  ,�  �  |  �  �   *  ��  �  �  �  �   *�R  �  �  �  �  �  �   +�_  5p    +  6$   ��  9	  )�R  <�  �    �  �  �    ,��  
�  ,��  �    [�  {  'it �   'end 8  (fF  R�  �  m  s  �   C >   o�  �  'it t   'end t  (fF  ��  �  �  �  �   C ]    :�    'it �   'end �  (fF  ��  �      �   C �   -��  Q~	  y	  .~	   /��  �  ;  F       /��  ��  W  b    "   ��  R��  v  |     0��  U��  �    �  �    �  (  .   0;�  qR�  �    �  �    �  4  .   0��  �A�  �    	  	    �  :  .   0��  �~�  �    ;	  P	    �  @  .   1��  ��    f	  q	    p    G 0     -�  ,~	  =  /�  �  �	  �	  F  Q   2��  b   3+�  ,��  ~	  �	  �	  F  p    *4s  0s  �  �	  
  F  >  �   *8�  D��  �  
  *
  F  >  r   �  W��  >
  N
  F  �  �   0��  ZQ�  �  ~	  n
  �
  F  �  (  .   0;�  ]��  �  ~	  �
  �
  F  �  4  .   0��  `i�  �  ~	  �
  �
  F  �  :  .   0��  c��  �  ~	    "  F  �  @  .   ��  g�  ��  j�  	 ~	  4��  ���  �  4�  ���  F     c  V   ]   Z  z  �  �  �  �  �  $  =  �  ��    �  �  /  {  5
�    5j�     {  >  /  �  �  �  6�  �        y	  Z  l  �  )   �  ~	  F  =  7p   b  8 h  9t�  W  �  :P  :b  ;�  �  4�A            ��  <�    �h ;U  �  �A            ��  <�  �  �h ;�  �  ��A            �  <�  �  �h ;�  %  ԶA            �2  <�  �  �h ;4  Q  ��A            �^  <�  i  �h =	  }  \�A     X      �-  <�    ��>y�  �3�  ��>�W  �R@  ��?st �.  ��@�  =  	pqB     AF�  �/  �PBes ��  �OC�A     �       Bcp �$  �HBcps �{  ��Dp*  Be ��  �l   EE  =  F5    -  =�  a  H�A           ��  <�    ��>y�  �@�  ��?n �N:  ��?st �.  ��@�  �  	�qB     Ar�  �  �PBds �=  �HCŴA     !       Be ��  �l  EE  �  F5    �  =�     �A     G      ��  <�    ��>y�  q9�  ��>�W  qR4  ��?st r.  ��@�  =  	�qB     Ar�  u  �PBds v=  �HC��A     $       Be z�  �l  =|  �  ��A     K      �W  <�    ��>y�  U.�  ��>�W  UI(  ��?st V.  ��@�  g  	�qB     Ar�  Y  �@Bds Z=  ��CK�A     $       Be ^�  �\  EE  g  F5    W  GP	  Q}  �  H�    H   w    Il  o�  �  ��A     +       ��  J}  �h Il  ��  �  Z�A     -       ��  J}  �h Kb  �     H�     I�  (�  #  "�A     7       �,  J�  �h LB  ��A            �^  AZ�  ��  	�C      M�  ��  p�A            ��  <�  �  �h?nc �/�  �d?wc �>�  �X NR  	�A     g       ��  A��  �5  	�C      K�	  �   �  H�  L  H   w    I�  K�    ޭA     +       �(  J�  �h O�  ��  K  ��A            �T  J�  �h =�  s  ��A     |       ��  <�  �  �X>y�  <.�  �P>�W  <O�  �HBwc =	V   �l@�  �  	�qB      EE  �  F5   
 �  =�  �  �A     �      �0  <�  �  �X?seq 4�  �PBuc 	<   �o@�  �  	�qB      P�  V   S  
�A            �`  <�  �  �h Pd  p   �  ��A            ��  <�  �  �h KJ  �  �  H�  �   O�  �  �  ڮA             ��  J�  �h K*
  �    H�  L  Q^�  W�  QK�  W8�   R�  ]�  #  ��A     =       �J�  �hJ�  �dJ�  �`  �   G=  	  �  	  �+          �$ 1  ��  �<   -N  ,  �  L  �  �  �  p   2N  p   �  �  int �   M  	d   frg 	�  	I  �   
�\   �   �V  �   ,�   �6   �  hex  4D  @  0  {K  �2  |�   0  ~m[  )  /  �   /   .  ?  �  �     �=  �g  `  f     �=    {  �    �    �=  4H  �  �       �=  �?  �  �       �=  *�l  �  �       �=  0]  �      !   �=  8�7    &    �    �#  = A  '  ?  J    �    fF  Q�1  -  c  i  9   fF  T�6  -  �  �     \?  X�:  -  �  �  9   �"  \iQ    �  �  9   �"  `�:  ?  �  �     2d  dF  E  �       ;W  ��         ~  ��    �6  �-  T �    �   4.  2,  4.  3�*  f  l  K   �(  6UB  E  �  �  K  �    �(  <�    C.  =�   .]  >�   E0  ?-  �e  @-  �  A-  �_  B-  rO  C-  3.  BW      K  �    4.  �%     K      E  �  J�  #�  NE�    P -  T p   �  p   -  �   �   �   �   �}  x=  �  P -  T p   �  p   �   �   �   �   zx  �U|  T p   F -  p   E  �    	~6  
�  
�  �  g&  	  6a  E ?  "  -  �  	   �  �	�  �  �2  N  Y  �  �    �  ?N  m  x  �  �   !�#  	�*  �  �  �  �  �   �  Pl  �  �  �  �    Y4  "	�c  �  �  �  �  �   R0  ',;  �  �  �  �   R0  1u?      �  �   "Ba  >�   "t ?�  "�\  @
0   �"8]  A-  �D�  	�  �  r  }  T p   �  p    #�5  	9+  �  �  T �  �  �    -  �R  H $  -  �  �  �   �0  MY  �  �  �  �   "�V  Q	   $�  	  %�-  <   � &   'l?  
CI    4  T �        �H  ���  [  F -  p   E  �   �H  ��(  �  F -  �  E  �   (�  2X�  �  T p   F -  Q  �   )�k  2:c  T �  F -  �  �    *�   	�qB     +�  �  �  �  +�   �  +�     ,�   -�   ,@  -�   ,�   oF  -  +@  ,�   +�   +E  K  .std  �  �   
J�  /`?  
K4  T �   0�-  1    �1  
J�  /`?  
K4  T �   0�-  1!    2@  
Nh  4  2@  
NW3  4   3�#  n  3�?  �  (N  �+  *�  	�qB     de  �  P  a	  4P  
�-  ?	  E	  �   �R  �  U	  �  �    5B  +|    5'.  ,�R  	  r  #�   ��  |  ��  ��  -  �	  �	  �    �  ��  -  �	  �	  �  �	   )�  ��  -  �	  �	  �  �	   9�  ��  -  
  !
  �  �	   O�  2�  -  9
  D
  �  �	   ��  �  -  \
  g
  �  �	   ��  n�  -  
  �
  �  �	   ��  E�  -  �
  �
  �  �	   ��  ��  -  �
  �
  �  �	   0�  b�  -  �
  �
  �  �	   '�  ��  -      �  �	   �  ��  -  .  9  �  �	   ��  
�  �	  Q  \  �  �	   #;�  �  �	  p  �  �	    6^�  �
(�  �   +	  +�	  �  +  �  +-  �  ,�  ,-  7�  �  8<    9�  9�  :�  �  D�@     �       �  ;�  �  �h<s '�  �d =  �@     (       �P  T �   <a   �h<b #  �` >=  h�@     �      �|  P -  T p   ?��  N�  ��?^W  N$p   ��?H*  N1-  ��?�b  N?�   ��?K.  O�   ��?.]  O�   ��?]  O#�  ��@�  P�  �X@u S|  ��Ak T�   ��BX�@     E       9  Ai a�   �l B��@     -       \  Ai d�   �h CԲ@     0       Ai f�   �d  7�  �  8<    >  �@     U       �  P -  T p   ?��  x�  �h?^W  x!p   �d?�b  x-�   �`?K.  x8�   �\?.]  y�   �X?]  y�  �TDE�  {	p     >�  w�@     �       �u  T p   F -  ?�2  �p   �l<fo �/E  �`?��  �6�  �X :�  �  �p@     �       ��  ;�  �  �h<str 1�  �` >4  -�@     J       �  F -  ?�2  �!p   �L<fo �8E  �@?��  �?�  �� >[  �^@     *       �Q  F -  ?�2  � �  �h<fo �7E  �`?��  �>�  �X ,w   >�  ��A     C       ��  T p   F -  F�2  2Q  �HF��  2!�  �@ :�  �  �V@     &       ��  ;�  �  �h?a  M�  �` ,�  >�  TV@     E       �,  T �  F -  F�2  2�  �HF��  2!�  �@ G:  :  P  H�  �  ICa  �   J,  �n  s   V@     4       ��  K:  �hKC  �` G/  �  �  H�  �  H   �    J�  =e  �  V@            ��  K�  �h G  �  �  H�  �   J�  �H    V@            �  K�  �h :S  ;  ��A     (       �W  T p   ;�  �  �h?�2  p   �d :�  v  LK@     ,       ��  ;�  �  �hL�  �  :}  �  "K@     )       ��  T �  ;�  �  �h?�2  �  �` G�  �  �  H�  �  H   �    J�  'F    K@            �  K�  �h :�  9  �J@     )       �F  ;�  �  �` G�  T  j  H�  
  I�-  *   MF  �b  �  �C@     V       ��  KT  �hK]  �` G  �  �  H�  
  H   �    M�   Y  �  �C@            ��  K�  �h GK  �    H�  
   M�  �@  &  �C@     #       �/  K�  �h =|  ��A            �a  @��  ��	  	�C      N\  ��  �A     �       ��  ;�  �  ��~<c �'�	  ��~ N9  v�  J�A     �       ��  ;�  �  ��~<c v'�	  ��~ N  m�  ��A     �       �  ;�  �  ��~<c m"�	  ��~ N�
  d=  ֿA     �       �Y  ;�  �  ��~<c d"�	  ��~ N�
  [{  �A     �       ��  ;�  �  ��~<c ["�	  ��~ N�
  R�  >�A     �       ��  ;�  �  ��~<c R"�	  ��~ N�
  I�  p�A     �       �  ;�  �  ��~<c I"�	  ��~ Ng
  @5  ��A     �       �Q  ;�  �  ��~<c @"�	  ��~ ND
  1s  ��A           ��  ;�  �  ��~<c 1"�	  ��~ N!
  (�  ȹA     �       ��  ;�  �  ��~<c ("�	  ��~ N�	  �  �A     �       �  ;�  �  ��~<c #�	  ��~ N�	  -  0�A     �       �I  ;�  �  ��~<c "�	  ��~ N�	  k  d�A     �       ��  ;�  �  ��~<c "�	  ��~ O�	  �  T�A            ��  ;�  �  �h P�  2�  �  H�  Q  H   �    M�    �  A@            �  K�  �h ,,  P  2  ,  H�  Q     M  �  O  ~@@     �       �`  K  �hK&  �` GR  n  x  H�  Q   M`  a  �  "@@     \       ��  Kn  �h QF  nH  �   @@            �?  #0   �h<p /�   �`  �   RB  	  8�  	  4�A     A       b1 1  -N  ,  �  L  2N  �  �  �  �  int q   frg 	:  I  �   �\   �   	4D  �  
0  {�   �2  |q   0  ~m[  �   �   [   /   .  �   [  q     �=  �g      a   �=    /  :  a  �    �=  4H  O  Z  a  g   �=  �?  o  z  a  m   �=  *�l  �  �  a  s   �=  0]  �  �  a  y   �=  8�7  �  �  a  q    �#  = A    �  �  a  �    fF  Q�1  �      �   fF  T�6  �  6  <  a   \?  X�:  �  U  [  �   �"  \iQ  g  t  z  �   �"  `�:  �  �  �  a   2d  dF  �  �  �  a   ;W  ��  �  �  a   ~  ��    �6  ��  T q    �   �  J~6  
  �  
  g&  �  6a  E ?  <  G  )  j   �  �R  H $  G  d  j  )   �0  MY    �  )  I   �V  Qj   �  j  �-  4   �    6a  E��  �  �  A  �   �  �R  H��  �  �  �  A   �0  MC�      A  I   �V  Q�   �  �  �-  4   �  �   	jwB     V  �  O  �   �   x   q   �  �   �   oF  �  �  q   q    std  -  �   J�  !`?  K�  T q   "�-  #s    �1  J  !`?  K�  T q   "�-  #y    $@  Nh  �  $@  NW3  �   %�#  �  %�?  �  (N  �+    	kwB     &de    P  �  'P  
�-  �  �     �R  �  �    I    ��  �  '��  �  �  �     �R  �  �    I    (B  +|    ('.  ,�R  �   j    �      )�  $	�C     �  )  	%	�C     *  *  +�  �  T�A     !       ��  ,�  $  �h-a  )I  �` .�  �  4�A            �,�    �h-a  (I  �`  )   E  	  ��  	  �-          �2 1  ��  	�<   -N  ,  �  L  2N  V   �  �  �  �  int �   frg 	  	I  �   
�\   �   �V  �   ,�   �6   �  hex  4D  (  0  {3  �2  |�   0  ~m[      3   /   .  '  3  �     �=  �g  H  N  >   �=    c  n  >  �    �=  4H  �  �  >  I   �=  �?  �  �  >  O   �=  *�l  �  �  >  U   �=  0]  �  �  >  [   �=  8�7      >  �    �#  = A  a  '  2  >  �    fF  Q�1  g  K  Q  s   fF  T�6  g  j  p  >   \?  X�:  g  �  �  s   �"  \iQ  I  �  �  s   �"  `�:  y  �  �  >   2d  dF    �  �  >   ;W  ��       >   ~  ��    �6  �g  T �    �   4.  2  4.  3�*  N  T  �   �(  6UB  -  l  w  �  �    �(  <�    C.  =�   .]  >�   E0  ?g  �e  @g  �  Ag  �_  Bg  rO  Cg  3.  BW  �  �  �  �    4.  �%    �  O    -  �  J|  #�  NE�  g  P �  T V   Z  V   g  �   �   �   '   �  Nf�  �  P �  T V   (  V   g  �   �   �   '   �}  x=  �  P �  T V   Z  V   �   �   �   '   @  x��  #  P �  T V   (  V   �   �   �   '   zx  �U|  Q  T V   F �  V   -  Z   ��  ��  T V   F �  V   -  (    	~6  
|  
�  �  g&  �  6a  E ?  �  �  >  W   �  �	9  �  �2  �  �  I  >    �  ?N      I  T   !�#  	�*  Z  %  0  I  T   �  Pl  D  O  I  �    Y4  "	�c  Z  g  r  I  |   R0  ',;  �  �  I  '   R0  1u?  �  �  I     "Ba  >>   "t ?.  "�\  @
0   �"8]  Ag  �D�  	�  Z      T V   I  V    #�5  	9+  Z  -  T   I      �  �R  H $  �  V  \  >   �0  MY  q  |  >     "�V  QW   $�  W  %�-  <   �    �	  6a  E��  �  �    �   �  �	A	  �  �  �  �        �  ��  
      "   !�#  	��  (  -  8    "   �  �  L  W    �    Y4  "	��  (  o  z    |   R0  'G�  �  �    '   R0  1��  �  �       "Ba  >   "t ?.  "�\  @
0   �"8]  Ag  �D�  	� (  	  	  T V     V    #�5  	��  (  5	  T         �  �R  H��  �  ^	  d	     �0  MC�  y	  �	       "�V  Q�   $�  �  %�-  <   � &l?  
CI  I  �	  T �   I  I   �H  ���  �	  F �  V   -  Z   �H  ��(  
  F �    -  Z   ^�  �d A
  F �  V   -  (   ^�  �"�  h
  F �    -  (   '�  2X�  �
  T V   F �  F  Z   '�k  2:c  �
  T   F �  �  Z   '��  2 �
  T V   F �  F  (   (��  2U�  T   F �  �  (    )�   	pwB     *.    �  '  *�   3  *�   >  +�   ,�   +(  ,�   +�   oF  g  *(  +�   *�   *-  �  -std 
   �   J�  .`?  Kn  T �   /�-  0U    �1  J�  .`?  Kn  T �   /�-  0[    1@  Nh  n  1@  NW3  n   2�#  �  2�?  �  (N  �+  )�  	qwB     de     P  �  3P  
�-  y        �R  �  �         ��  �  3��  �  �  �     �R  �  �        4B  +|  �  4'.  ,�R  �   *W  *�  *�    *�    +A	  +�  5'  >  6<    *�  >  *�  I  +9  +�  7�  7  8r  �  D�@     �       ��  9�  O  �h:s ''  �d 8z  �  ��A     �       ��  9�    �h:s ''  �d ;�	  �@     (       �  T �   :a I  �h:b #I  �` <%  h�@     �      �E  P �  T V   =��  NZ  ��=^W  N$V   ��=H*  N1g  ��=�b  N?�   ��=K.  O�   ��=.]  O�   ��=]  O#'  ��>�  P  �X>u SE  ��?k T�   ��@X�@     E         ?i a�   �l @��@     -       %  ?i d�   �h AԲ@     0       ?i f�   �d  5'  U  6<    <g  Z�A     �      ��  P �  T V   =��  N(  ��=^W  N$V   ��=H*  N1g  ��=�b  N?�   ��=K.  O�   ��=.]  O�   ��=]  O#'  ��>�  P  �X>u SE  ��?k T�   ��@J�A     E       >  ?i a�   �l @��A     -       a  ?i d�   �h A��A     0       ?i f�   �d  <�  �@     U       �  P �  T V   =��  xZ  �h=^W  x!V   �d=�b  x-�   �`=K.  x8�   �\=.]  y�   �X=]  y'  �TBC�  {	V     <�  �A     U       ��  P �  T V   =��  x(  �h=^W  x!V   �d=�b  x-�   �`=K.  x8�   �\=.]  y�   �X=]  y'  �TBC�  {	V     <#  w�@     �       ��  T V   F �  =�2  �V   �l:fo �/-  �`=��  �6Z  �X 8�    �p@     �       �7  9�  O  �h:str 1  �` <Q  i�A     �       ��  T V   F �  =�2  �V   �l:fo �/-  �`=��  �6(  �X 8�  �  ��A     �       ��  9�    �h:str 1  �` <�	  -�@     J       �  F �  =�2  �!V   �L:fo �8-  �@=��  �?Z  �� <�	  �^@     *       �j  F �  =�2  �   �h:fo �7-  �`=��  �>Z  �X <
  N�A     J       ��  F �  =�2  �!V   �L:fo �8-  �@=��  �?(  �� <A
  $�A     *       �  F �  =�2  �   �h:fo �7-  �`=��  �>(  �X 8\  *  �V@     &       �F  9�  D  �h=a  M  �` +]   <h
  ��A     C       ��  T V   F �  D�2  2F  �HD��  2!Z  �@ +"  <�
  TV@     E       ��  T   F �  D�2  2�  �HD��  2!Z  �@ E�  �  
  F�  O  GCa  >   H�  �n  -   V@     4       �>  I�  �hI�  �` 8d	  ]  ��A     &       �y  9�    �h=a  M  �` <�
  ��A     C       ��  T V   F �  D�2  2F  �HD��  2!(  �@ <�
  v�A     E       �  T   F �  D�2  2�  �HD��  2!(  �@ E�    1  F�    GCa     H  ��  T  B�A     4       �e  I  �hI$  �` E  s  �  F�  9  F   �    He  =e  �  V@            ��  Is  �h E�   �  �  F�  9   H�  �H  �  V@            ��  I�  �h 8O    LK@     ,       �*  9�  O  �hJ|  �  8�  P  ��A     (       �l  T V   9�  O  �h=�2  V   �d 8  �  "K@     )       ��  T   9�  O  �h=�2    �` E0  �  �  F�  O  F   �    H�  'F  �  K@            ��  I�  �h 8>    �J@     )       �'  9�  D  �` 8W  F  �A     ,       �[  9�    �hJ|  �  8�  �  ��A     (       ��  T V   9�    �h=�2  V   �d 8	  �  ��A     )       ��  T   9�    �h=�2    �` E8  �     F�    F   �    H�  m�  #  ��A            �,  I�  �h 8F	  K  ��A     )       �X  9�    �` E�  f  |  F�  D  G�-  *U   KX  �b  �  �C@     V       ��  If  �hIo  �` E�  �  �  F�  D  F   �    K�   Y  �  �C@            ��  I�  �h E3      F�  D   K�  �@  8  �C@     #       �A  I  �h L_�  ��A           ��  =    ��~=� 7  ��~=
% JV   ��~=��    ��~ L� u�A           ��  =    ��~=� 7  ��~=
% JV   ��~=��    ��~ M�  2  #  F�  �  F   �    K�    F  A@            �O  I  �h +  M�  2f  u  F�  �  O   KU  �  �  ~@@     �       ��  If  �hIo  �` E:  �  �  F�  �   K�  a  �  "@@     \       ��  I�  �h NF  nH  b   @@            �=  #0   �h:p /b   �`  y   �I  	  � 	  `0          h< 1  ��  �<   -N  ,  �  L    b   �  �  �  |   2N  �  �  *  �   int �   � )     �<   N  	�   �   R   	�   �  	V   M  	p   %   	4�     frg 	8  	I    
�\     �V  �   ,T  �6   �  hex  4D  �  0  {�  �2  |�   0  ~m[  �  �  ^   /   .  �  ^  �     �=  �g  �  �  i   �=    �  �  i     �=  4H       i  t   �=  �?     +  i  z   �=  *�l  @  K  i  �   �=  0]  `  k  i  �   �=  8�7  �  �  i  �    �#  = A  �  �  �  i  T   fF  Q�1  �  �  �  �   fF  T�6  �  �  �  i   \?  X�:  �      �   �"  \iQ  t  %  +  �   �"  `�:  �  D  J  i   2d  dF  �  c  i  i   ;W  ��  }  �  i   ~  �a   �6  ��  T �    T  4.  2�  4.  3�*  �  �  �   �(  6UB  �  �  �  �  /   �(  </   C.  =�   .]  >T  E0  ?�  �e  @�  �  A�  �_  B�  rO  C�  3.  BW  m  x  �  �    4.  �%  �  �  �    �  �  JL   Np �  P �  T <   �
  <   �  �   �   �   R   � x+ !  P �  T <   �
  <   �   �   �   R   	 �� T <   F �  <   �  �
    	~6  
L  
�  U   g&     s  6a  E��  �  �  �
  �	   �  �	  �  �  �  �  �
  �
   !�  ��  �  �  �
  �
   "�#  	��  �
  �    �
  �
   �  �    $  �
  �    Y4  "	��  �
  <  G  �
  L   R0  'G�  [  f  �
  R   R0  1��  z  �  �
  G   #Ba  >�
   #t ?�	  #�\  @
0   �#8]  A�  ��  	X �
  �  �  T   �
     $�5  	��  �
    T G  �
  G    �  �R  H��  �  +  1  �
   �0  MC�  F  Q  �
  G   #�V  Q�	   %�  �	  &�-  <   � 'l?  
CI  t  �  T �   t  t   ^�  �J �  F �  g	  �  �
   ^�  �"�  �  F �  G  �  �
   (� 2�   T   F �  `  �
   )��  2U�  T G  F �  �  �
    *#  	�yB     +Y  G  �  R  +a  ^  +T  i  ,�   -�   ,�  -T  ,T  oF  �  +�  ,�   +�   +�  �  .std  E	  �   
J�  /`?  
K�  T �   0�-  1�    �1  
J 	  /`?  
K�  T �   0�-  1�    2@  
Nh  �  2@  
NW3  �   3�#  �  3�?   	  (N  �+  +m	  4*Z  	�yB     de  �	  ��  �	  5��  �  �	  �	  �	   �R  �  �	  �	  G    6B  +|  f  6'.  ,�R  k   +�	  7R  
  8<    9h
  :% ;V  �   <�c  0
  6
  u
   <a  F
  L
  u
   A !
�    �  $�     =	
  >
  +	
  u
  +k  �
  +�  �
  ,  ,�  > 	  >2	  ?G  �
  ��A     �       ��
  @�  �
  �hAs 'R  �d Bs  �@     (       �"  T �   Aa t  �hAb #t  �` C�  ��A     �      �N  P �  T <   D��  N�
  ��D^W  N$<   ��DH*  N1�  ��D�b  N?�   ��DK.  O�   ��D.]  O�   ��D]  O#R  ��~E�  PG  �XEu SN  ��Fk T�   ��G��A     E         Fi a�   �l G�A     -       .  Fi d�   �h HF�A     0       Fi f�   �d  7R  ^  8<    C�  z�A     W       ��  P �  T <   D��  x�
  �hD^W  x!<   �`D�b  x-�   �\DK.  x8�   �XD.]  y�   �TD]  yR  �PIJ�  {	<     C!  ��A     �       �G  T <   F �  D�2  �<   �hAfo �/�  �`D��  �6�
  �X ?f  f  ��A     �       ��  @�  �
  �hAstr 1G  �` C�  ^�A     }       ��  F �  D�2  � g	  ��Afo �7�  ��D��  �>�
  �� C�  $�A     *       �%  F �  D�2  � G  �hAfo �7�  �`D��  �>�
  �X ?1  D  ��A     &       �`  @�  �
  �hDa  MG  �` ,  C�  �A     E       ��  T   F �  K�2  2`  �HK��  2!�
  �@ ,M  C  v�A     E       �   T G  F �  K�2  2�  �HK��  2!�
  �@ L�    $  M�  �
  NCa  �
   O   ��  G  B�A     4       �X  P  �hP  �` L�  f  y  M�  d  M   �    OX  =e  �  V@            ��  Pf  �h Lz  �  �  M�  d   O�  �H  �  V@            ��  P�  �h ?$    �A     ,       �  @�  �
  �hQL  �  ?�  C  ��A     )       �_  T   @�  �
  �hD�2    �` ?�  �  ��A     )       ��  T G  @�  �
  �hD�2  G  �` L  �  �  M�  �
  M   �    O�  m�  �  ��A            ��  P�  �h ?    ��A     )       �  @�  �
  �` L+  (  >  M�  o  N�-  *�   R  �b  a  �C@     V       �r  P(  �hP1  �` Lk  �  �  M�  o  M   �    Rr   Y  �  �C@            ��  P�  �h L�  �  �  M�  o   R�  �@  �  �C@     #       �  P�  �h S� <1��A     .       �@  Aptr <N@  �XE ]  =u
  �h +�   T� 00�   x�A     J       ��  Aptr 0M@  �XE ]  1u
  �h U] +1�A     f       �V6
  �  ��A            ��  @�  {
  �h ? 
  �  ��A     J       �  @�  {
  �XFv �   �l ?�  %  2A@     6       �O  @�  �  �`Ac 63/  �\E�  7�  �h W\  2`  s  M�  �  M   �    RO    �  A@            ��  P`  �h ,�  Wx  2�  �  M�  �  �   R�  �  �  ~@@     �       ��  P�  �hP�  �` L�      M�  �   R�  a  4  "@@     \       �=  P  �h XF  nH    @@            �D  #0   �hAp /  �`  �p   YO  v	  �% 	  02          sC 5  5   wint 5   5�3  M   S   "�  S   5�Q  M   ��  �|   k   "-N  |   x"1  ",  "�  "�  "2N  �   "�  "�    �|   %   4�   �   ��  �   !�  @l  �  M       	k   �   #	k       &	k   �  )	k    P  ,	k   (�  -	k   0  25   8>  55   <   8"�   5@  K�  l  5)  L�  5�   M�  ]	  �   "�  yL  zfrg 	�"  AI  �  [�\   �  :�V  5   ,  !�6   !�  \hex  ]4D  V  {0  {a  |�2  |5   0  ~m[  ?  E  �"   B/   .  U  �"  5     �=  �g  v  |  #   �=    �  �  #  �   �=  4H  �  �  #  #   �=  �?  �  �  #  #   �=  *�l  �  �  #  #   �=  0]      #  %#   �=  8�7  1  <  #  5    '�#  = A  +#  U  `  #     'fF  Q�1  1#  y    =#   'fF  T�6  1#  �  �  #   '\?  X�:  1#  �  �  =#   '�"  \iQ  #  �  �  =#   '�"  `�:  C#  �  �  #   '2d  dF  I#      #   ;W  ��  .  4  #   ~  �   �6  �1#  T 5      4.  2B  4.  3�*  |  �  O#   �(  6UB  [  �  �  O#  �   �(  <�   C.  =5   .]  >  E0  ?1#  �e  @1#  �  A1#  �_  B1#  rO  C1#  }3.  BW    )  O#  5    ~4.  �%  6  O#  �o    [  C�  J?  3�  N	�  �  P �  T 5   �.  5   1#  5   5   5   S    3#�  NE�  �  P �  T �   �.  �   1#  5   5   5   S    3��  x;�    P �  T 5   �.  5   5   5   5   S    �  �ܪ  T 5   F �  5   [  �.    A~6  	
?  [�  	H  g&  	a  6a  	E ?  z  �  q.  �%   �  �		�  �  	�2  �  �  |.  q.   -�  	?N  �  �  |.  �.   .�#  		�*  �.  �  �  |.  �.   �  	Pl      |.  5    Y4  	"	�c  �.  *  5  |.  ?   R0  	',;  I  T  |.  S    R0  	1u?  h  s  |.  �"   Ba  	>q.   t 	?�-  �\  	@
k   �8]  	A1#  �;�  		��  �.  �  �  T S   |.  S    K�5  		9+  �.  �  T �"  |.  �"    �  �R  	H $  �      q.   �0  	MY  4  ?  q.  �"   �V  	Q�%   �  �%  ^�-  |   �    	?
  6a  	E��  �  �  �/  �%   �  �		�	  �  	�  �  �  �/  �/   -�  	��  �  �  �/  �/   .�#  		��  �/  �  �  �/  �/   �  	�  	  	  �/  5    Y4  	"	��  �/  2	  =	  �/  ?   R0  	'G�  Q	  \	  �/  S    R0  	1��  p	  {	  �/  �"   Ba  	>�/   t 	?�-  �\  	@
k   �8]  	A1#  �K�5  		��  �/  �	  T �"  �/  �"    �  �R  	H��  �  �	  �	  �/   �0  	MC�  
  
  �/  �"   �V  	Q�%   �  �%  ^�-  |   � A#  	?
  ��i  H
   C}C  	N  D{
  L]I  8#    Mh
  :�-  5   �
  !�6   \red !�C   �Q  0`  �Q  �+  �
  �
  �,   -�Q  �*  �
  �
  �,  �,   .�#  �_  �,      �,  �,   �N  �    �R  �   �7  �   \.   �   >*  !�    �R  "�
  ( �
  �R  %�  7^  '
   1#  �  T �  �.   _�  '�V  1#  T �  �.    BD  5C  `h 8�_  �,  �  �.   �N  =j4  �.  �  �.   �R  B�i  �.    �.   �7  E�N  �.  %  �.   \.  I�P  �.  ?  �.   >*  L�  �.  Y  �.     P�,  �.  q  w  �.   E�+  U}O  1#  �  �.   E\G  Z�"  1#  �  �.   �G  dma  �  �  �.   -�G  g"  �  �  �.  �.   .�#  i  �.  �  	  �.  �.   Rr  o_L  �.  !  '  �.   �(  |�^  <  G  �.  �.   �e  ��  \  l  �.  �.  �.   i  ��=  �  �  �.  �.  �.   �+  ��B  �  �  �.  �.   #�l  �0  �  �  �.  �.   $�2  .A  �  �  �.  �.  �.   $Q:  D�      �.  �.  �.   $�l  xm  3  >  �.  �.   $�R  ��6  T  _  �.  �.   $�  +  u  �  �.  �.   #�  �   �  �  �.  �.   #�_  #=M  �  �  �.  �.   1�1  0Z$  1#  �  �  �.   1�1  9mI  1#  �    �.  �.  C#  �.  �.   F  ��    D H  T �  ;E3  �p  A e   �  N�'  �  (�'  (�G  (�l  (��  (�  (�Y  <�   #�b  �@  �  �  �.  �   #�+  ��m  �  �  �.  �.   F�5  ��  T �  ;E3  �p  L �  A e   �S  5�  `h 88Y  �,  '  �.   �N  =�!  �.  A  �.   �R  BbJ  �.  [  �.   �7  E�h  �.  u  �.   \.  If  �.  �  �.   >*  LV/  �.  �  �.     P�[  �.  �  �  �.   E�+  U9  1#  �  �.   E\G  Z-  1#  �  �.   �G  d3<      �.   -�G  gn.  +  6  �.  
/   .�#  itF  /  N  Y  �.  
/   Rr  o�+  �.  q  w  �.   �(  |�j  �  �  �.  �.   �e  �jK  �  �  �.  �.  �.   i  �A]  �  �  �.  �.  �.   �+  �6  �    �.  �.   #�l      !  �.  �.   $�2  H)  7  G  �.  �.  �.   $Q:  D�  ]  m  �.  �.  �.   $�l  x.8  �  �  �.  �.   $�R  �Ld  �  �  �.  �.   $�  �  �  �  �.  �.   #�  �R  �  �  �.  �.   #�_  #	g      �.  �.   1�1  0  1#  *  0  �.   1�1  9�  1#  J  d  �.  �.  C#  /  /   F  ��    D �  T �  ;E3  �p  XA e     aX  �(�w  (��  (��  (�A  (�[  (��  <   #�b  �R%  �  �  /  �   #�+  ��      /  �.   F�5  ��  T �  ;E3  �p  XL �  A e    Da  L]I  8#    MN  2l  �  bclz �  5   �  |    T |    �%B  �$   :L3  5   ��  !�6   !�i  !'   �   8  H�	�   8  ��Q  �    �.  �  �   k    - 8  �&    &  �.  �.   .�#  �
[  �.  >  I  �.  �.   qe  �ze  1#  a  l  �.  �    8  ��   v6  ��   ��  �w   �  ��   �  8  ��	Y  <�   8  �i'  �  �  �.  �   k   5    -8  �E2  �    �.  �.   .�#  ��G  �.    $  �.  �.   ��  �<   H�(  ��   L�-  ��.  P+  ��  X �  �>  �	�  �>  �Q*    �  �.   -�>  �0o  �  �  �.  �0   .�#  ��>  �0  �  �  �.  �0   �+  ��.    ^  �5  �	  K�R  ��3  1#  �  �.  �.  �.       �	[    �'  -  3  '/   ,+  �	�,   �Q  ��.  �G  �[   �b  ��  C%  ��Z  |  �  -/  8/   'N�  �YV  �   �  �  -/  k    1�&  H
:  �   �  �  -/  �   k    $��  z�W  �  �  -/  �    $Q.  �]      -/  �   k    '�:  -	�c  k   5  ;  -/   ��\  :N/                         @       O�Z  < �   OkG  = �    =d  D�\  k   �  �      S  k   �  k    O�&  f<   =�  hw   Oa  k�  1#  �  �    =�e  xw   =�&  {w   �]  �w    P�i  ��U  �.  2  =  -/  �    P�i  �C  �.  V  a  -/  5    P'  !�C  �.  z  �  -/  k    #�  3  �  �  -/   #�@  :�5  �  �  -/  �.   �=  �
8/   �  ��,  8  ��  +2  ��  �  �	k    Y  ��/  (�^  �-  D=  �,   C�    A7! � �  � �# V  \  �-   Q $�-      \   w &�-  ; u  & 1#   �-  � �-   �+$ QQ   R�Z   E�#  ch %z ).  �  �  /.  �   Rw "6u  D *	  QQ   ch -	}& ).  &  1  O.  �   D 2 E  P  O.  �   �"  5Y �  h  n  Z.   �r  9� 1#  �  �  Z.  e.   �r  <` 1#  �  �  Z.  e.   �" @i k.  �  �  O.   �" D� �  �  �  O.  5    � K�    �  x' N �  !  ,  /.  �   � S� @  F  /.   � VP �  ^  i  /.  i   RQ !4\  %y  gd �  �  �  /.  i   �+  x� �  �  �  /.  �  i   o�  �} 1#  �  �  /.   q  ��! �  �  �  /.   $  �0 �      /.   /" ��' i  3  9  /.   }# �$ i  Q  W  /.   �$ �~ i  o  z  /.  �   !! � �  �  /.  �  :.   d �� �  �  �  /.   dend �� �  �  �  /.   p  �i   #  ��  T �&  �     b	 Q  �R  ' .  -  8  .  .   T �&  H 5  ;E3  �p  X c 
�  Q   bget 
�" .    #.   Tag ,  T    ] �  �! 	 �-  �  �-   T �&   �-  � �-   S�Z  �+�
  SA)  �7�  SA)  �7H  ]�Z  �   �c  �l       �0   �c  w  5  E  �0  ?
  ~-   �c  =  Z  e  �0  ~-   ��c  !zG  {  �  �0  �0   �c  #�  �  �  �0  �0   �c  (�;  �  �  �0  5    '�#  -4  �0  �  �  �0  �   �c  2�n  �     �0   a  8p;         �0   'S  >�&  1#  9   ?   �0   '+H  BY0  1#  X   c   �0  m-   �  G	m-   R  H1#  D=  �,   �  � �5  l?  

CI  #  �   T 5   #  #   3�H  ���  �   F �  5   [  �.   3^�  �"�  !  F �  �"  [  �/   3�H  ��(  3!  F �  �"  [  �.   % 
� .  ]!  Tag ,  T   #.   Tǟ  2�  �!  T S   F �  m%  �.   T��  2U�  �!  T �"  F �  <J  �/   T�k  2:c  �!  T �"  F �  <J  �.   G	
 1  %"  T �*  �-  �  H�-  "  /C#  /r]   �O  C#  "  6r]   G� 1  o"  T �*  �-  �  H�-  Y"  /C#  /�^   �O  C#  h"  6�^   3� �  �"  T �&  �-  �  �O  �-   �Q  

!I  ,T  �"  T |   ,T  ,T   _��  
	
�  ,T  T |   ,T  ,T    4�  	|B     Z   �"    �"    #  <   65   V  6    "oF  1#  V  5   5   [  O#  �std  R%  �   J�#  =`?  K8#  T 5   e�-  /#    �1  J�#  =`?  K8#  T 5   e�-  /%#    fR !f! 3�# �#  8  5  T .   �}  >�#  �  $  8  5   T C#   y" ?$  8  �-  T �N   \ `$  8  �^  T �^   B! �$  8  r]  T r]   g@  Nh  8#  g@  NW3  8#  �}  >+$  }  ! �$  �$  T �N  �N   G "  �$  T r]  QP   �}  >m$  ��  ۈ  C#  %  T C#  Q   �}  >
$  G�
 h"  E%  T �^  OQ   �}  >L$   h�#  s#  h�?  �#  "(N  Z   "�+  4M  	|B     Cde  �,  P  �%  iP  
�-  �%  �%  �,   B�R  �  �%  �,  �"    ��  &  i��  �  �%  &  �,   B�R  �  &  �,  �"    jB  +|  Y  j'.  ,�R  a  :� 5   
b&  !  !: !�	  :�" 5   �&  !  !�$ !p !�  k$ p�&  c*  <�   � i1   $ 0� �&  �&  �-  21   -$ X" �&  �&  �-  z1   .�#  � .  '  '  �-  z1   �� @ �&  *'  5'  �-  5    [# L� I'  O'  �-   �W	  #| 5   �&  p'  v'  �-   �	  VM 5   �'  �'  �-  M   k   P1   �	  �� 5   �'  �'  �-  �"  k   P1   � �. �'  �'  �-  S    h �� 5   (  (  �-  b&   G � &(  ,(  �-   �' �� 5   D(  J(  �-   � �4& 5   b(  m(  �-  V1   �	  �  5   �(  �(  �-  �  5    >(! 2' 5   �&  �(  �(  �-  D1   > 3' 5   �&  �(  �(  �-  J1   >I 4� 5   �&  )  #)  �-  M   k   P1   >� 5M 5   �&  D)  Y)  �-  �"  k   P1   >� 6� 5   �&  z)  �)  �-  �  5   V1   1Y 2 5   �)  �)  �-   1� "J 5   �)  �)  �-   1� ,j 5   �)  �)  �-   1;W  N�
 5   	*  *  �-   $� _� %*  +*  �-   8  A=&  H Bb&  LW# C%21  P� G(�   X �&  D�*  L� $8#   V !�  �O 'z*   Mh*  k� xJ�&  �,  <�&   l�  �*  �*  1  &1   l� c# �*  �*  1  ,1   #� l�  +  +  1  5   21   �fd o 5   )+  /+  1   �W	  s� 5   �*  Q+  W+  1   ?(! | 5   �*  y+  �+  1  D1   ? �� 5   �*  �+  �+  1  J1   ?I ��% 5   �*  �+  �+  1  M   k   P1   ?� �V' 5   �*  
,  ,  1  �"  k   P1   ?� �9" 5   �*  A,  V,  1  �  5   V1   �_fd [5   p�� R �*  x,  1  5     �*   �%  �%  7M
  7m
  �
  �,  `  �
  7S  ^P  h-  ^P  �b  �,  �,  m-   -^P  �#  �,  -  m-  x-   .�#  PK  ~-  -  %-  m-  x-   �c  �!  9-  ?-  m-   a  �l  S-  Y-  m-   je  5     �,  �,  m-  h-  �,  �-  �-  dmap �7  �   �-  �-  �-  k    B�@   H  �-  �-  �   k     �-  �&  �-  5  �-  %S   .  &|    7m*  5    .  �&    Q  �  �  /.  �  4�*  	�C     �  O.    Z.    �  Y  q.  �  |.  �  �  �  �.  �  �  �  �.  Y  �  ^  �.  �  �.  C  �  �.  �  �.  H  �.    �.  �    �.  �  /    �  -/  �-  %w   N/  &|    >/  @eW  ;  @�i  j  @�  x  @Gb  �  m'  �   �mQ5  �   ��:  �     @L  	  %  �/  &|    a  �/  �  �/  �	  �  DP0  Ir& ��*  I�
 ��*  I ��*  N�% �	B0  ��% �"0  (0  �0   �'& �60  �0  5     I�% �0   ���/  4�/  	�C     4�/  	`C     4�/  	�C     0  �0  4B0  	XC     Ux  �	�C     U�  �	�C     U�  �	�C     �  �0  �   6�  �  �  ^  �^  �^  r]  �]  �*  1  6�*  �,  81  �D1  �-   =&  b&  k   �  �5   i1  � o1  �t�  \1  c*  ��  �   7�$  7�$  �_ ��A            ��y   ��A     �       ��1  	>  _5   �l	u  _5   �h Ve,  J�1  2  �  !1     <    �1  & 02  d�A     +       �92  �1  �h �1   \2  6�A     -       �e2  �1  �h 5  �2  D�@     �       ��2  �  �.  �hs 	'S   �d  �   �@     (       ��2  T 5   a 
#  �hb 
##  �` S  J�A     �      �4  P �  T 5   ��  N�.  ��^W  N$5   ��H*  N11#  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#S   ���  P�"  �Xu S4  ��k T5   ��/�A     E       �3  i a5   �l ~�A     -       �3  i d5   �h ��A     0       i f5   �d  %S   4  &|    �  h�@     �      �C5  P �  T �   ��  N�.  ��^W  N$�   ��H*  N11#  ���b  N?5   ��K.  O5   ��.]  O5   ��]  O#S   ���  P�"  �Xu S4  ��k T5   ��X�@     E        5  i a5   �l ��@     -       #5  i d5   �h Բ@     0       i f5   �d  �  ��A     �       ��5  P �  T 5   ��  x�.  �X^W  x!5   �T�b  x-5   �PK.  x85   �L.]  y5   �H]  yS   �DהA     ;       �  {	�   �l  �  B�@     1       �6  �2  Z�.  �h �  26  ��@     �      �y6  �  /  ��2n �.  ��
u �.  �X
v �.  �P
w �.  �H �  �6  �@     �      ��6  �  /  ��2n ��.  ��
u ��.  �X
v ��.  �P
w ��.  �H  r  �@            �7  T �  �2  '�.  �h  �  �@            �C7  T �  �2  '�.  �h _  b7  D�@     �      ��7  �  �.  ��2n �.  ��
u �.  �X
v �.  �P
w �.  �H >  �7  ��@     �      �8  �  �.  ��2n ��.  ��
u ��.  �X
v ��.  �P
w ��.  �H �  s�@     1       �:8  �2  Z�.  �h   �A     �       ��8  T 5   F �  �2  �5   �lfo �/[  �`��  �6�.  �X �  �8  Ƃ@     V      ��8  �  �.  �Xn ��.  �P�N  ��.  �hd4  ��.  �` '  ��@            �9  �  =�.  �h m  29  �|@     �      �:  �  /  ��2n x�.  ���N  {�.  �P
s ��.  �X�R  ��
  ���}@     �       �9  
x ��.  �H �~@     z       �9  
x ��.  �@ w�@     Q       �9  f?  ��.  �� Ɓ@     Q       f?  ��.  ��  �  �|@     1       �;:  �2  U�.  �h \	  Z:  ��A     �       �v:  �  �/  �hstr 	1�"  �` �  �|@            ��:  �  L�.  �h �  �:  N|@     H       ��:  �  /  �X	�2  #�.  �P� $�.  �h    8|@            �;  �  8�.  �h �  7;  �x@     V      �o;  �  /  �Xn ��.  �P�N  ��.  �hd4  ��.  �` �  �;  �x@            ��;  �  /  �h	�2  �.  �` �  �;  �x@            ��;  �  �.  �h	�2  �.  �` �  <  Zx@     H       �3<  �  �.  �X	�2  #�.  �P� $�.  �h �  =x@            �^<  �  =�.  �h   }<  zr@     �      �[=  �  �.  ��2n x�.  ���N  {�.  �P
s ��.  �X�R  ��
  ��Is@     �       �<  
x ��.  �H et@     z       =  
x ��.  �@ v@     Q       7=  f?  ��.  �� Zw@     Q       f?  ��.  ��  w  Hr@     1       ��=  �2  U�.  �h ?  *r@            ��=  �  L�.  �h  �  r@            ��=  �  8�.  �h T  �=  �p@     �       �>  �  �.  �hstr 	1�"  �`  e  (�A            �@>  p 
%#.  �h �   �A     J       ��>  F �  �2  �5   �Lfo �/[  �@��  �6�.  �� �  �>  �>  �  �.  )�"  ��  )�  �%�   )&8  �6k    �>  ;R  �>  Xp@     K       �?  �>  �h�>  �d�>  �X�>  �P l  0?   o@     7      �k?  �  �.  �H�N  ��.  �@�2  �"�.  ��72  ��.  �X G  �?  �m@     7      ��?  �  �.  �H�N  ��.  �@�2  �!�.  ���l  ��.  �X '  �?  ~m@     j       � @  �  �.  �h�2  |�.  �` �  @  <@  �  �.  )�  ��   )&8  �)k   )X[  �65     @  &Z  _@  m@     d       ��@  @  �h@  �`#@  �X/@  �T !  �@  �j@     �      ��@  �  /  ��	�2  �.  ��	�   �.  ���N  �.  �X�R  �.  �P�7  �.  �H u  oj@            �*A  �  I�.  �h G  IA  h@     a      ��A  �  /  ��	�2  D�.  ��	f?  D$�.  ���l  E�.  �X72  F�.  �P�N  Z�.  �H �   $�A     *       ��A  F �  �2  � �"  �hfo �7[  �`��  �>�/  �X �  B  �f@     7      �SB  �  /  �H�N  ��.  �@�2  �"�.  ��72  ��.  �X [  �f@            �~B  �  E�.  �h �  �B  �e@     7      ��B  �  /  �H�N  ��.  �@�2  �!�.  ���l  ��.  �X A  be@            �C  �  B�.  �h 0�  "C  :e@     (       �IC  �  �.  �ha �!�.  �`b �1�.  �X w  hC  �d@     j       ��C  �  /  �h�2  |�.  �` 0�  �C  �d@            ��C  �  /  �h �  �C  2b@     �      �/D  �  �.  ��	�2  �.  ��	�   �.  ���N  �.  �X�R  �.  �P�7  �.  �H %  b@            �ZD  �  I�.  �h �  yD  �_@     a      ��D  �  �.  ��	�2  D�.  ��	f?  D$�.  ���l  E�.  �X72  F�.  �P�N  Z�.  �H   �_@            �E  �  E�.  �h �  u_@            �/E  �  B�.  �h 0Y  NE  d_@            �[E  �  �.  �h !  �^@     *       ��E  F �  �2  � �"  �hfo �7[  �`��  �>�.  �X 0  �E  �A            ��E  �  .  �hx .  �` 3!  ��A            �F  Tag ,  T   p 
#.  �h �  <F  ��A     <      ��F  �  3/  ��	W �6�   ��	  �Fk   ��v6  �|   �X
slb ��.  �P
bkt �'/  �H�  �	k   �@sZ  ��  ���-  �1#  ���2  ��.  �� ]!  CtA     G       �)G  T S   F �  	�2  2m%  �H	��  2!�.  �@   HG  ��A     0       �dG  �  U.  �hptr -�  �` 0n  �G  f�A     "       ��G  �  `.  �h�-  9$e.  �` a  �G   ^@     �       ��G  �  3/  �H	  !=k   �@v6  '�   �X
fra )�.  �P �  H  �]@     L       �'H  �  �0  �h �  FH  �\@     �       �sH  �  �.  �X	�2  ��.  �P� ��.  �h =  �H  �[@     D      �HI  �  3/  ��	��  95   ��v6  �   �@�  	|   ���H  
	k   �X
slb �.  ��Rr  �.  �Pk\@     ^       
off k   �H�\@     >       �2  �.  ��   Y  gI  D[@     X       ��I  �  /  �X� p�.  �h   �I  �Z@     �       �J  �  /  �H	�2  �.  �@v  �.  �h�\  �.  �`�Z@     I       �l  �.  �X  �	   J  ��A     &       �<J  �  �/  �ha  	M�"  �` �"  �!  v�A     E       ��J  T �"  F �  	�2  2<J  �H	��  2!�/  �@ �  �J  �J  �  �/  )Ca  	�/   +�J  ��  �J  B�A     4       ��J  �J  �h�J  �` �  K  �Y@     �       �0K  �  "/  �X	�2  ��.  �P� ��.  �h 0I  OK  JY@     I       �xK  �  �.  �Xp ��   �Padr �	|   �h k  �K  �K  �  �.   +xK  �`  �K  4Y@            ��K  �K  �h    �K  �X@     O       ��K  �  �0  �h �  L  (X@     �       �fL  �  �.  �H	�2  �.  �@v  �.  �h�\  �.  �`�X@     I       �l  �.  �X    �L  `W@     �       ��L  �  3/  �X	v6  �;�   �P� ��.  �h �  �L  �L  �  �0     <    �L  �  �L  8W@     '       ��L  �L  �h E  M  #M  �  �0  )�  ~-   �L  dh  FM  W@     2       �WM  M  �hM  �`   vM  �V@     &       ��M  �  w.  �ha  	M�"  �` �!  TV@     E       ��M  T �"  F �  	�2  2<J  �H	��  2!�.  �@ �  �M   N  �  �.  )Ca  	q.   +�M  �n  #N   V@     4       �4N  �M  �h�M  �` 1  BN  XN  �  U.  )� 2�   +4N  � {N  L�A            ��N  BN  �hKN  �` �-   �$  :�A            ��N  T �N  x *�N  �h �  �N  
�A     0       ��N  �  5.  �hptr %�  �`  �  ��A            �(O  � �-  �h E  6O  IO  �  #     <    +(O  =e  lO  V@            �uO  6O  �h +  �O  �O  �  #   +uO  �H  �O  V@            ��O  �O  �h �  �!  ;�A     �       �QP  T �*  �-  �  H�-  �O  /C#  /r]   H%  �O  ��n+!P  C#  "   W �   �H�! +C#  ���  +"  �� �$   �$  -�A            ��P  T r]  x .QP  �h %"  ��A     �       �Q  T �*  �-  �  H�-  �P  /C#  /�^   H%  �O  ��n+�P  C#  h"   W �   �H�! +C#  ���  +h"  �� %   �$  �"A            �OQ  T C#  x .Q  �h E%   (%  ��A            ��Q  T �^  x .OQ  �h o"  ��A     G       ��Q  T �&  �-  �  H%  �O  �hW (�-  �` �  �Q  �6A     *       �R  T S   �  �.  �h�2  	S   �d 0P  0R  ��A            �=R  �  `.  �h �  \R  r�A     2       �iR  �  U.  �h �  �R  J�A     (       ��R  �  `.  �h�-  <$e.  �` �  �R  &�A     #       ��R  �  5.  �X �  �R  ��A     3       ��R  �  5.  �X �  S  
O@     �      �,T  �  3/  ��~��  �6k   ��~JO@     �      �S  ��  �5   �\bkt �'/  �PsZ  ��  ���2  �.  ���O@     *      �S  
slb 	�.  �H �P@     �      
slb 	�.  �@�\  �  ��  �R@     �         6|   ��
fra 7�.  ���\  9�  ��~  �    �"  �U@     +       �oT  T |   a 
,T  �hb 
#,T  �`  �"  �A     +       ��T  T |   a 
	,T  �hb 
	#,T  �` 	  �T  �A     ,       ��T  �  �/  �hJ?  �  �	  U  ��A     )       �"U  T �"  �  �/  �h�2  	�"  �` �  0U  CU  �  �/     <    +"U  m�  fU  ��A            �oU  0U  �h �	  �U  ��A     )       ��U  �  �/  �` W  �U  �A     �      �V  �  5.  ��it ��  ��    �i  �H; ��  �P
 �i  �X 	  #V  ��A     a       �?V  �  5.  �Xptr N&�  �P �  ^V  �K@     h      �W  �  3/  ��~	W z0�   ��~v6  �|   �X�\  ��  ��
fra ��.  �P
slb ��.  �H
bkt �'/  �@�  �	k   ��sZ  ��  ���-  �1#  ���2  ��.  ��   1W  LK@     ,       �FW  �  �.  �hJ?  �  �  lW  "K@     )       ��W  T �"  �  �.  �h�2  	�"  �` �  �W  �W  �  �.     <    +�W  'F  �W  K@            ��W  �W  �h   �W  �J@     )       �X  �  w.  �` v   X  �A     �      �KX  �  5.  �H�^  g#i  �@� i�  �X B  YX  cX  �  �-   +KX   �X  ��A     *       ��X  YX  �h ,  �X  �X  �  5.   +�X  � �X  ��A     "       ��X  �X  �h �  �X  �X  �  #  )�-  *#   �X  �b  Y  �C@     V       �+Y  �X  �h�X  �`   9Y  LY  �  #     <    +Y   Y  oY  �C@            �xY  9Y  �h a  �Y  �Y  �  #   xY  �@  �Y  �C@     #       ��Y  �Y  �h oD \f�A     5       ��Y  	)�  \�  �X� ]�-  �h ,�$ V5   $�A     B       �NZ  2c V5   �\	)�  V�  �P� W�-  �h o  P��A     R       ��Z  	)�  P�  �X� Q�-  �h ,A 65   ��A           �l[  	)�  6�  �H	u 6$M   �@	  605   ��	  6=k   ��� 8�-  �h��A     @       '[  
e :
5   �d 6�A     9       K[  
e ?
5   �` u�A     9       
e D
5   �\  ,�' 25   ��A            ��[  	)�  2�  �h ,�' ,5   V�A     I       ��[  	)�  ,�  �X� -�-  �h ,� "�   ��A     i       �X\  	)�  "�  �H� #�-  �hq $�  �X�A     =       
e %	5   �d  ,� 5   {�A     r       ��\  	)�  �  �X	�   !�   �P	�	  -5   �L� �-  �h��A     >       
e 	5   �d  ,� 5   ��A     �       �.]  	)�  �  �X� �-  �`
e 5   �l , �  ]�A     �       �,^  2fd 5   ��~	  "�"  ��~a< pa�  �]  �]  1  5    q�R  �]  �A     *       ��]  r]  � ^  �h	t �-  �` rT  21  �]  L�A            �
^  �  ^  �h1   s�' ,�A            �J�-  �h   ,�  ��  ��A     Q      �_  	{�  ��"  ��}	  �+�"  ��}�  �5   �l �1#  �k
fd �5   ��}N< ^_  pa�  �^  �^  1  5    q�R  �^  V�A     *       �_  �^  � 7_  �h	t �-  �` rT  21  +_  ��A            �=_  �  7_  �h	1   s�' ��A            �J�-  �h  ��A     C       
e �	5   �d  ,� �5   ;�A            ��_  	)�  ��  �h ,� �5   �A     4       ��_  	)�  ��  �X� �1  �h (0  `  N`  �  �0     <   Wtit ��-  X :.  X^ �  X� �  Wte �5      ��_  n`  �A     �       ��`  `  ��~u`  �`  8`  8$`  8-`  86`  �?`  8@`    Y`  0�A     �       9`  �`9$`  �h9-`  ��~96`  ��~Y?`  ��A     [       9@`  �\   0  a  a  �  �0   ��`  0a  �A            �9a  a  �h ,  Xa  ��A     E       ��a  �  !1  �X	�   ��  �P	�	  �(5   �L	e �7V1  �@��A     '       
e �	5   �l  �+  �a  v�A     U       �?b  �  !1  �X	u �#�"  �P	�7  �2k   �H	�  �DP1  �@
s �
�   �`��A     (       
e �	5   �l  �+  ^b   �A     U       ��b  �  !1  �X	u �M   �P	�7  �+k   �H	�  �=P1  �@
s �
�   �`8�A     (       
e �	5   �l  �+  �b  ,�A     �       �:c  �  !1  ��~	  �-J1  ��~*�  Jc  	��B     ��A     �       
e �	5   �l  %Z   Jc  &|    :c  W+  nc  ��A     h       ��c  �  !1  �X	8  |*D1  �P�   }�  �`
e ~5   �l /+  �c  *�A     �       ��c  �  !1  ��~��A            
e w	5   �l  0+  d  �A            �"d  �  !1  �h �*  0d   Ud  �  !1  �fd l5   �X# l!21   "d  �' xd  ��A     E       ��d  0d  �h9d  �dFd  �X *  �d  \�A     u       ��d  �  �-  �X*�  �d  	��B     
ptr d�   �h %Z   �d  &|    �d  �)  e  ��A     �       �Te  �  �-  �X*�  de  	|�B     ��A            
e O	5   �l  %Z   de  &|    Te  �)  �e  ��A     �      �Tf  �  �-  �H*�  df  	p�B     ��A            �e  
e -	5   �l ��A     Z       f  e 6	�  �X��A     J       
e 7
5   �h  ��A     �       v A
k   �P��A     i       
e B
5   �d   %Z   df  &|    Tf  �)  �f  �A     �       ��f  �  �-  �h*�  �f  	`�B      %Z   �f  &|    �f  �)  �f  ��A            �g  �  �-  �X*�  ,g  	P�B     ��A     0       
e 	5   �l  %Z   ,g  &|   
 g  m(  Pg  ��A           �(h  �  �-  �H�   ��  �@�	  �+5   ��e �  �P*�  8h  	G�B     ��A            �g  e �	5   �l ��A     e       h  M �   �`��A     D       
e 
5   �\  J�A     @       
e 
5   �X  %Z   8h  &|    (h  J(  \h  �A     n       ��h  �  �-  �Xq � V1  �PM ��  �`&�A     3       e �	5   �l  ,(  �h  ��A            ��h  �  �-  �h 0(  �h  ��A     ?       ��h  �  �-  �h �'  i  h�A     T       �Li  �  �-  �h  �/b&  �d*�  \i  	8�B      %Z   \i  &|    Li  �'  �i  ��A     m       ��i  �  �-  �hc � S   �d*�  �i  	2�B      %Z   �i  &|    �i  �'  �i  2�A     �      ��j  �  �-  ��~u �&�"  ��~�7  �5k   ��}�  �GP1  ��}*�  �i  	,�B     ?�  �|   ��~% �1#  �o��A     �       �j  v �
k   ��~��A     Y       e �
5   �h  ��A             �j  e �
5   �d ��A             �j  e �
5   �` ��A     @       nl �M   �X  v'  k  ��A     �      �Gl  �  �-  ��~u VM   ��~�7  V.k   ��~�  V@P1  ��~*�  8h  	'�B     ?�  �|   �X�A     �       �k  v \
k   ��~�A     Y       e ]
5   �l  G�A           v x
k   ��~G�A             l  e q
5   �h g�A             &l  e s
5   �d ��A     a       e y
5   �`   5'  fl  f�A     /       �sl  �  �-  �h '  �l   �l  �  �-     <   W�it H�    sl  5 �l  :�A     +       ��l  �l  �h sl  U& �l  N�A     �       �)m  �l  ��~u�l  	m  8�l   Y�l  u�A     �       9�l  ��~  �  �B@     �       ��m    S0k   ��tc U|   �`e ^|   �Xf _|   �Pip `|   �His a|   �@�B@     :       i W�   �l   �  $B@            �(n  idx D6�   ��tc F|   �hs K5   �dip L|   �Xis M|   �Pf N|   �H �&  6n   Ln  �  �-  )X# 0%21   (n  � on  z�A     �       ��n  6n  �h?n  �` 0?-  �n  B@            ��n  �  s-  �h %-  �n  �A@     B       ��n  �  s-  �h*�  8h  	"�B       v  �A@            �o  x )|   �h �
  "o  ,o  �  �,   +o  �b  Oo  hA@     Q       �Xo  "o  �h V  2io  |o  �  U#     <    Xo    �o  A@            ��o  io  �h B  V)  2�o  �o  �  U#  �o   �o  �  �o  ~@@     �       �p  �o  �h�o  �` h  p  p  �  U#   p  a  =p  "@@     \       �Fp  p  �h �F  nH  �   @@            ��p    #k   �hp /�   �` Z�&  �   "Z�  �  "Z�  �  " �    Z  	  �( 	  ��A     �      Rx 1  ��  �@   -N  ,  �  L  ��  -   ]	  -   int 2N  �  �  �  �  �  �   de  �  �( D�( �   	�   
e( ;�( r   �   	�  	r    
p( 5B) r     	r    
) *�( r   '  	�  	r   	<   
X) a) r   P  	r   	f   	r   	�   
z( �) r   y  	r   	  	4   	   	) &) r   	r   	�  	4   	    �   �   #�A            ��  �  �h �   ��A     A       �  H	  ;�  �X  ;+r   �Tret <r   �l �   ��A            �<  fd 5r   �l r     ��A     E       ��  H	  *�  �X�  *)r   �Tfd *5<  �H_fd +r   �l f   '  3�A     N       �  fd r   �\�   f   �P�	  )r   �Xe 8�  �Hoff 	f   �h) r    Z   P  ��A     R       ��  fd r   �\buf   �P��  )4   �Hܓ  9  �@ret Z   �h) r    �  y  ��A     R       �fd r   �\u $�  �P��  34   �H{) C  �@z) Z   �h  %U   :;9I  $ >  $ >  & I  :;9   :;9I8   :;9I8  	   
 I  :;9n  I  ! I/  ;   .?n4<d   I4  4 :;9I?<  4 :;9I?  4 :;9I?  :;9  .?:;9n2<d   I  .?:;9nI2<d   :;9I82   :;9I82  / I  .?n42<d  4 I?4<  . 4@�B  .Gd    I4     !4 :;9I  ".1nd@�B  # 1  $1  %4 1  &1  '4 1  (.4@�B  ) :;9I  *.Gd@�B  + I4  , :;9I  -4 :;9I  .  /4 :;9I  0.Gd@�B  1.G:;9d   2.1nd@�B  3  4.?:;9I@�B  54 :;9I  64 :;9I  7.?:;9n@�B  8.?:;9nI@�B  9 I   %  . @   %  $ >   :;9I  $ >  :;9   :;9I8  I  ! I/  	& I  
.?:;9'I@�B   :;9I   :;9I  4 :;9I   I  &      .?:;9'@�B   %  $ >   :;9I  $ >  :;9   :;9I8   :;9I8  .?:;9'@�B  	 :;9I  
4 :;9I  4 :;9I  .?:;9'I@�B   I   %  $ >   :;9I  $ >  .?:;9'@�B   :;9I   %   :;9I  $ >  $ >  .?:;9'I@�B   <   :;9I  4 :;9I  	 I   %  $ >  $ >  .?:;9'I@�B   :;9I   :;9I  4 :;9I    	 I  
.?:;9'@�B  4 :;9I   %   :;9I  $ >  .?:;9I@�B   :;9I  4 :;9I     I  	& I  
 :;9I  4 :;9I       7 I  &   $ >    I   I4   :;9I  4 :;9I  / I  & I   I4   :;9I  	4 :;9I  
.Gd@�B  4 :;9I   :;9I8   I   :;9I   I  4 :;9I   1    .G@�B  .?:;9n2<d  4 I4   I4  :;9  .?:;9n<d  .?:;9I@�B  .?:;9nI<   :;9I  $ >  I  .Gd   ! I/     !.?:;9I@�B  "(   #.?:;9nI2<d  $.?:;9n<d  %.?:;9n2<d  & :;9  ' :;9I  (.1nd@�B  ).?:;9nI<d  *4 nG  + :;9I  ,.?:;9n<�d  -.?:;9nI<�d  ..G@�B  / :;9I8  0.Gd@�B  1 :;9I82  2.1nd@�B  3.?:;9nI2<d  4 :;9I?<l   54 G  6m>I:;9  7.?:;9n<  8/ I  9.?:;9nI2<  : :;9I82  ;0 I  <7 I  = I  >.?:;9�@�B  ?4 :;9I?<  @:;9n  A :;9  B.?:;9n<d  C9:;9  D9  E: :;9  F I8  G :;9I?<l   H.?:;9nI<d  I :;9I  J4 G  KB I  L
 :;9  MU  N.?:;9@�B  O :;9I?<l   P :;9I?<l   Q4 :;9I<l  R(   S:;9  T.?:;9nI<d  U <  V4 :;9I<l  W.?:;9nI<  X.?:;9nI2<  Y.?:;9n<  Z��  [/ I  \4 :;9nI?<l   ]4 nG  ^4 :;9nI?<  _.?:;9nI<cd  `4 nG  a.G:;9d   b IJ  c%U  d$ >  e   f9:;9  g:;9  h :;9I?<l   i :;9I82  j :;9I82  k:;9  l :;9I  m.?n4<d  n.?n4<d  o.?:;9n<  p0 I  q4 :;9I<
l  r:;9  s:;9  t.?:;9nI<  u:;9  v :;9I?<
l   w :;9I?<l   x.?:;9n2<�d  y4 Gn  z! I/  {;   |9:;  }&   ~.?:;9n<�d  .?:;9nI<d  �4 :;9I<  �4 :;9I?  �4 nG  �. 4@�B  �.4@�B  �  �4 :;9I  �.?:;9@�B  �.?:;9I@�B  �.?:;9I@�B  �I  �   �. ?:;9I@�B  �.?:;9nI@�B  �4 :;9Il   %U   :;9I  $ >  & I   :;9I  ;   $ >  :;9  	 :;9I8  
9:;9   :;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d  / I  .?:;9nI<d  .?n4<d  9 :;9  / I  .?:;9n<�d  .?:;9nI<�d    :;9I82  !.?:;9nI<d  "0 I  # <  $.?:;9n<  %.?:;9n<  &4 G  ' I  ( I  )B I  *9:;  + :;9I?<l   ,��  -/ I  .4 :;9nI?<l   /4 nG  09:;9  1.?:;9n<�d  24 :;9nI?<  3 :;9I8  4.?:;9nI<cd  5<  6.?:;9nI<  79  8>I:;9  9: :;9  :I  ;! I/  <4 G  =.Gd@�B  > I4  ? :;9I  @.G@�B  A :;9I  B :;9I  C.Gd   D I4  E :;9I  F.1nd@�B  G 1  H I  I.Gd@�B  J  K4 :;9I  L :;9I  M.1nd@�B  N.?:;9I@�B  O4 I4  P :;9I  Q4 :;9I  R.?:;9I@�B  S.G@�B  T4 :;9I  U.G:;9d   V.1nd@�B    I   I4   :;9I  / I   I4  & I   :;9I8  .Gd@�B  	4 :;9I  
.?:;9nI2<d   1   I   I  .?:;9n2<d  4 :;9I  .G@�B  4 :;9I  4 :;9I   :;9I   I4  :;9   :;9I  .?:;9n<d    .Gd   .?:;9nI<  .Gd@�B  $ >  .?:;9n<d  .?:;9n2<d   :;9     ! :;9I  ".1nd@�B  #.1nd@�B  $ :;9I  %.?:;9nI<d  &I  '! I/  (.?:;9n<�d  ).?:;9nI<�d  *.G@�B  + :;9I  ,(   -4 :;9I?<  . :;9I82  // I  0 :;9I82  14 I4  2.?:;9nI2<d  3 :;9I?<l   4.?:;9n<  54 G  6B I  74 nG  8.?:;9nI2<  90 I  ::;9  ;.?:;9n<  <.?:;9I@�B  = :;9  >9:;9  ?9  @: :;9  Am>I:;9  B I8  C :;9I?<l   D.?:;9nI<d  E.?:;9n<d  F.?:;9nI2<d  G :;9I  H4 G  I4 :;9I<l  J(   K.?:;9nI<  L.?:;9nI2<  M:;9  N.?:;9nI<d  O4 :;9I<l  P��  Q/ I  R4 :;9nI?<l   S4 nG  T4 :;9nI?<  U.:;9<  V4 nG  W  X :;9I  Y :;9I  Z.G:;9d   [ IJ  \%U  ]$ >  ^   _;   `9:;9  a4 :;9I<
l  b:;9  c.?:;9nI<  d:;9  e :;9I?<
l   f :;9I?<l   g:;9  h :;9I  i.?n4<d  j.?n4<d  k.?:;9n<  l0 I  m <  n.?:;9n2<�d  o.?:;9nI<d  p9:;  q&   r.?:;9n<�d  s4 :;9I<  t. :;9<  u. :;9I<  v.:;9I<  w4 :;9I?  x4 nG  y4 I?4<  z4 :;9I  {4 :;9I  |1  }4 1  ~1  4 1  � I  �.?:;9nI@�B   %  4 :;9I?  $ >   I  $ >    I   :;9I  / I   I4   :;9I  4 :;9I  4 :;9I  4 :;9I  	 I4  
& I  4 I4    .G@�B   I     :;9I  4 :;9I  .Gd@�B  .?:;9I@�B   :;9I8   1   I  / I   I  .?:;9n<d  .?:;9n<   :;9I  .?n4<d   I4  :;9  .?:;9n2<d   .?:;9nI2<d  !.Gd   "U  # :;9I8  $(   % :;9I  &.?:;9nI<  ' :;9I  (.?:;9n<  )B I  *.1nd@�B  +I  , :;9I82  -   .$ >  /! I/  0.?:;9n<d  1  24 :;9I  3.?:;9n2<d  4 :;9  5.G@�B  6.Gd@�B  7.?n4<�d  8.?n4d@�B  9.?n4d@�B  :.1nd@�B  ;.?:;9nI<d  <:;9  =.?:;9I@�B  >.?:;9n<�d  ?.?:;9nI<�d  @ :;9I82  A :;9I?<l   B4 G  C4 :;9I?<  D7 I  E :;9I  FU  G.?:;9nI2<d  H:;9  I4 nG  J :;I8  K :;9I  Lm>I:;9  M.?:;9nI2<  N0 I  O:;9  P��  Q/ I  R4 :;9nI?<l   S4 nG  T.?:;9I@�B  U.4<d  V.42<d  W :;9  X9:;9  Y9  Z: :;9  [.?:;9nI<  \ I8  ] :;9I?<l   ^.?:;9nI<d  _.?:;9n<d  `4 :;9I<l  a(   b.?:;9nI2<  c.?:;9nI<d  d4 :;9I<l  e <  f4 G  g4 :;9nI?<  h4 nG  i.:;9I@�B  j.?:;9@�B  k.?:;9@�B  l. ?:;9I@�B  m.:;9Id@�B  n.:;9I2d@�B  o :;9I  p.G:;9d   q IJ  r%U  s$ >  t I  u:;  v   w;   x9:;9  y4 :;9I<
l  z.?:;9nI<  {:;9  | :;9I?<
l   } :;9I?<l   ~:;9   :;9I  �.?n4<d  �.?:;9n<  �0 I  �9 :;9  �.?:;9n2<�d  �.?:;9nI<d  �9:;  �&   �.?:;9n<�d  �>I:;9  �4 nG  �! I/  �:;9  �:;9  �.:;9@�B  �.?:;9@�B  �.?:;9nI@�B   %   :;9I  $ >  4 :;9I?<  $ >   I  7 I  & I  	   
.?:;9I@�B   :;9I   :;9I  4 :;9I  &   .?:;9I@�B   :;9I  4 :;9I  .?:;9I@�B   I  4 I4  I  ! I/   :;9I  4 :;9I    .?:;9I@�B   %U   :;9I  & I  $ >  ;   $ >  9:;9   :;9  	4 :;9I<
l  
9:;9  9  4 :;9I<l  : :;9  m>I:;9  (   (   :;9  .?:;9n<d   I4  .?:;9n<�d   I  .?:;9nI<�d   :;9I8  .?:;9nI<  / I  .?:;9nI<  .?:;9nI2<  .?:;9nI<d  .?:;9nI2<  .?:;9n2<d  .?:;9n<d   .?:;9n2<d  !.?:;9nI2<d  " :;9I82  #0 I  $:;9  % :;9  & I8  ':;9  (.?:;9nI<  ):;9  *.?:;9nI<d  +.?:;9nI2<d  , :;9I?<
l   - :;9I?<l   . :;9I?<l   / :;9I?<l   0.?:;9nI<d  1/ I  2:;9  3.?:;9nI2<d  4�:;9  5�:;9  6 :;9I�8  7��  8/ I  9 :;9I  :.?:;9n2<�d  ;4 G  < I  = I  >   ? :;9I82  @.?:;9nI<d  A.?:;9n<d  B  CB I  DI  E! I/  F4 nG  G4 nG  H4 nG  I9:;  J.G@�B  K :;9I  L.Gd@�B  M I4  N :;9I  O4 :;9I  P.G@�B  Q4 :;9I  R  S  T :;9I  U4 :;9I  V :;9I  W.Gd   X I4  Y :;9I  Z.1nd@�B  [ 1  \.Gd@�B  ].1nd@�B  ^4 :;9I  _��:;9  `��:;9  a 1  b.?:;9n@�B  c.?:;9I@�B  d.?:;9nI@�B  e.?:;9nI@�B  f4 I4  g IJ   %  $ >  $ >   :;9I  ;   9:;9  . ?:;9n<  .?:;9nI<  	 I  
.?:;9n<  . G@�B     .G@�B   :;9I   I  .G@�B  4 I4  I  ! I/  & I  .G@�B   %U   :;9I  & I  $ >  ;   $ >  9:;9   :;9  	4 :;9I<
l  
9:;9  9  4 :;9I<l  : :;9  m>I:;9  (   (   :;9  .?:;9n<d   I4  .?:;9n<�d   I  .?:;9nI<�d   :;9I8  .?:;9nI2<  .?:;9nI<  .?:;9nI<d  .?:;9nI2<  .?:;9n2<d  .?:;9n<d  .?:;9n2<d  .?:;9nI2<d    :;9I82  !/ I  "0 I  #:;9  $ :;9  % I8  &:;9  ':;9  ( <  ).?:;9nI<d  *.?:;9nI2<d  + :;9I?<
l   , :;9I?<l   - :;9I?<l   . :;9I?<l   /.?:;9nI<d  0/ I  1�:;9  2�:;9  3.?:;9nI2<d  4 :;9I�8  5��   6 :;9I  7�:;9  80 I  9�:;9  :��  ;/ I  <4 G  = I  > I  ?   @ :;9I82  A.?:;9nI<d  B.?:;9n<d  C9 :;9  DI  E! I/  F4 nG  G! I/  H9:;  I.Gd   J I4  K.1nd@�B  L 1  M :;9I  N.1nd@�B  O.G@�B  P :;9I  Q :;9I  R.Gd@�B  S I4  T��:;9  U��:;9  V 1  W�� :;9  X.G:;9d@�B  Y :;9I  Z4 I4  [4 :;9I  \.?:;9nI@�B  ]4 :;9I  ^.?:;9nI@�B  _ IJ   %U   :;9I  $ >  & I  $ >  9:;9   :;9  4 :;9I<l  	:;9  
:;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  9 :;9   <   I  ;   4 G  :;9      I  B I  9:;   :;9I?<l   ��   / I  !4 :;9nI?<l   "4 nG  #9:;9  $4 :;9nI?<  %m>I:;9  &(   ' :;9I8  (.?:;9nI<cd  ).?:;9nI<d  *.?:;9nI<d  + :;9I82  , :;9I?<l   -:;9  . I8  /.?n4<d  0.?:;9nILM<d  1.?nL4<d  2 I84  3.?:;9nL<�d  4. ?:;9nI<  54 nG  64 I?4<  7I  8   9 I  :4 G  ;.Gd@�B  < I4  =.Gd@�B  > :;9I  ? :;9I  @4 I4  A4 :;9I  B4 :;9I  C  DU  EI  F! I/  G.G:;9d   H I4  I.1nd@�B  J 1  K.Gd   L.G@�B  M.G:;9d@�B  N.G@�B  O.1nd@�B  P.GId@�B  Q :;9I  R.1nd@�B   %U  $ >   :;9I  ;   & I  $ >     9:;9  	 :;9  
4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  :;9  .?:;9nI<d  .?n4<d  .?n4<d  9:;9  .?:;9n<  .?:;9n<   .?:;9n<�d  !.?:;9nI<�d  " :;9I82  #.?:;9nI<d  $/ I  %0 I  & <  '.?:;9nI<  (.?:;9n<  ).?:;9n<  *4 G  + I  , I  -B I  .9:;  / :;9I?<l   0��  1/ I  24 :;9nI?<l   34 nG  4.?:;9n<�d  54 :;9nI?<  6. ?:;9nI<  7I  8! I/  94 G  :.Gd@�B  ; I4  < :;9I  =.G@�B  >.G@�B  ? :;9I  @4 :;9I  A4 :;9I  B  C  D  E4 :;9I  F :;9I  G.Gd   H I4  I :;9I  J.1nd@�B  K 1  L I  M.1nd@�B  N.G:;9d@�B  O.G:;9d@�B  P.G:;9d   Q.?:;9nI@�B   %  $ >  ;   $ >  & I  9:;9   :;9  4 :;9I<l  	:;9  
:;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  9 :;9  :;9   <  .?:;9nI<d   :;9I82  / I  0 I  :;9  4 G   I   I  B I   9:;  ! :;9I?<l   "��  #/ I  $4 :;9nI?<l   %4 nG  &9:;9  '.?:;9n<�d  (4 :;9nI?<  )4 G:;9  *4 G  +.G:;9d@�B  , I4  - :;9I  ..G:;9d@�B   %U  $ >   :;9I  ;   & I     $ >  9:;9  	 :;9  
4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  :;9  .?:;9nI<d  .?n4<d  .?n4<d  9:;9  .?:;9n<  .?:;9n<   .?:;9n<�d  !.?:;9nI<�d  " :;9I82  #.?:;9nI<d  $/ I  %0 I  &.?:;9nI<  '.?:;9n<  (.?:;9n<  )4 G  * I  + I  ,B I  -9:;  . :;9I?<l   /��  0/ I  14 :;9nI?<l   24 nG  3.?:;9n<�d  44 :;9nI?<  5I  6! I/  74 G  8.Gd@�B  9 I4  : :;9I  ;.G@�B  <.G@�B  = :;9I  >4 :;9I  ?4 :;9I  @  A  B  C4 :;9I  D :;9I  E.Gd   F I4  G :;9I  H.1nd@�B  I 1  J I  K.1nd@�B  L.?:;9@�B  M.G:;9d   N.?:;9nI@�B   %U  $ >   :;9I  ;   $ >  & I     9:;9  	 :;9  
4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  :;9  .?:;9nI<d  .?n4<d  .?n4<d  9:;9  .?:;9n<  .?:;9n<    <  !.?:;9n<�d  ".?:;9nI<�d  # :;9I82  $.?:;9nI<d  %/ I  &0 I  '.?:;9nI<  (.?:;9n<  ).?:;9n<  *4 G  + I  , I  -B I  .9:;  / :;9I?<l   0��  1/ I  24 :;9nI?<l   34 nG  4&   5.?:;9n<�d  64 :;9nI?<  7I  8! I/  99  ::;9  ; :;9I<l   <.:;9<d  =: :;9  >4 G  ?.Gd@�B  @ I4  A :;9I  B.G@�B  C.G@�B  D :;9I  E4 :;9I  F4 :;9I  G  H  I  J4 :;9I  K :;9I  L.Gd   M I4  N :;9I  O.1nd@�B  P 1  Q I  R.1nd@�B  S.?:;9@�B  T.?:;9I@�B  U. ?:;9@�B  V.Gd@�B  W.G:;9d   X.?:;9nI@�B    I   I4  / I   I4   :;9I  .Gd@�B  4 :;9I  & I  	 :;9I  
4 :;9I   :;9I8   I   I   1   I4  .?:;9nI<d     :;9I  :;9  .?:;9n<d  4 :;9I  .G@�B  4 :;9I  .?:;9n2<d    .Gd    :;9I  .?:;9nI<   :;9I82  / I  .1nd@�B   .G@�B  !(   "$ >  #.?:;9n<d  $.?:;9n2<d  %I  &! I/  '.?:;9nI2<d  ( :;9  ) :;9I  *4 I4  +.1nd@�B  ,.?:;9I@�B  -.?:;9n<�d  ..?:;9nI<�d  // I  0.Gd@�B  1.?:;9nI2<d  2 :;9I  3.?:;9n<  44 G  54 :;9I?<  6B I  74 G  84 1  94 1  :m>I:;9  ;0 I  < I8  = :;9I?<l   >.?:;9nILM2<d  ?.?:;9nILM2<d  @4 nG  A :;9  B.?:;9n<d  C9:;9  D9  E.?:;9nI2<  F :;9I82  G.:;9I<  H��  I4 :;9I<  J I  K.?:;9nI<d  L4 :;9I<l  M: :;9  N:;9  O :;9I?<l   P.?:;9nI<d  Q I82  R :;9I2  S :;9I  T.?:;9n<  U4 G:;9  V.G:;9d   W  X4 I4  Y1  Z IJ  [4 :;9I<l  \(   ]:;9  ^0 I  _.?:;9nI<  `.?:;9nI2<  a:;9  b.?:;9nI<  c.?:;9nI2<d  d.?:;9nI<d  e��  f9 :;9  g4 :;9nI?<l   h4 nG  i.?:;9n<�d  j4 :;9nI?<  k:;9  l.?n4<�d  m4 nG  n��:;9  o.?:;9@�B  p.4<d  q.4d@�B  r.I4d@�B  s.4@�B  t4 :;9I  u1  v%U  w$ >  x   y;   z9:;9  {:;9  | :;9I  }.?n4<d  ~.?n4<d  .?:;9n<  �4 :;9I<
l  �:;9  � :;9I?<
l   � :;9I?<l   �:;9  �.?:;9n2<�d  �9:;  � I84  �.?:;9nL<d  �.?:;9nILM<d  �4 :;9I<  �.?:;9nI<d  �.?:;9nILM<d  � :;9I82  �.?nL4<d  �4 nG  �.:;9<d  �.:;9<d  �: :;9  �  �I  �   � I  �4 I?4<  �. 4@�B  �.4@�B  �.1d@�B  �1  �.1d@�B  � :;9I  � :;9I  �4 :;9I  �.?:;9nI@�B   %  $ >   :;9I  ;   $ >  & I  9:;9  .?:;9n<  	 I  
.?:;9nI<  .?:;9nI<   I  .G@�B   I  .G@�B   :;9I  4 :;9I   :;9I  4 :;9I     &   .G@�B  4 :;9I   1     �      /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx/window /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/bits /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/lemon /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include  graphics.h   main.cpp    window.h   list.h   types.h   stdint.h   fb.h   stddef.h   surface.h   types.h   stdio.h   ipc.h    G 	Z@     
�ff!.  tt!.�  	M@     � 	�2(K�d�tu�'t��g���
<	�'
�' t �	�K t��+��<tKxfftK� ot�>	�'
� t�K
�+�( t ���<tKK +mt%����'��= jt�>Zt<ZK
�H<
t&$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�.K�k�<60B�4�B �8R:�<(.*�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9 %)!D<K/>/�LT���.��u\,	tD.	J�(!@![�, t � / �kv>f��f���u,fftJg,fftJg�& J( t��& J( t�tf � ��"u%�* f�/f�, �9 fG �; �  .Y �f fM �t �� f� �� �h .���u�<f5 J; t& <K+f �7.Df9�J�trX�t<K'f�J='f�JZ'f�)J<='f�)J<">4<;tf6K�K- g.�� J	�w  �" t f�	u*ut �* f �8 �H fY �J �, .k �{ f_ �� �� f� �� �} .�!u�<f: J@ �( <���<K)f�J=)f�JZ)f�+J<=)f�+J<! >3 <: t f8 K � K0���t � t�tJ" X' t <Y$�)t/<�h$�(t�.L�K00tg\+tgZy.mh X0�4C4RfIfY<<4.t��*[� f�~���<J  	�@     �*  	�@     ����  	@     � 
�u  	@     � �  	8@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K  	f@     �  	�@     )�#���tY��Y����  	V@     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	�@     �	 � t J / �    '   �       src/gfx/sse2.asm      	@"@     !>==ALLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""�� �   D  �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../sysdeps/lemon/include/lemon  filesystem.c   types.h   stdint.h   stddef.h   off_t.h   filesystem.h    0 	�%@     �&=0�(3>0'=:00'=30")KB00'K �    �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include ../sysdeps/lemon/include/lemon  ipc.c   types.h   stdint.h   ipc.h    , 	l'@     �	&K20����& �    �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include  syscall.c   types.h   stdint.h    g 	�'@     �� �    �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include  fb.c   types.h   stdint.h    - 	/(@     ��&K 1   6   �      ../sysdeps/lemon/generic  itoa.c     	o(@     ���t
 /! W J f[t 0 � t g �
 Y yX J �	X?/v��t=
�=� =% f f1 J f . � t / f�{	�>	K �   �   �      ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  essential.cpp   stddef.h    . 	�)@     �� � � � W	vKN0�� � � � � < -	vK90��� � � � � < -w �. �5 � � �5 � < -	wK0	�� � ! W	vK v/   �  �      ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  random.hpp   new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   stdlib-stubs.cpp   optional.hpp   strtofp.hpp   logging.hpp   utility.hpp   mutex.hpp   errno.h   types.h   stdint.h   stddef.h   locale_t.h 	  stdlib.h   type_traits   debug.hpp   charcode.hpp   mbstate.h   <built-in>      	r=@     �  	�=@     
�� � �# u( �+ <4 �9 �< <> �- < .H f �F � . � �"  	@>@     ���� t � �, t/ f1 � X Y �  � X0 .3 f& f J �k t � �, t/ f1 � X Y �& �! X6 .9 f, f J �k�,t.fXY!�X1.4f'f.	�����f=fX=fX=f
>= 2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	2A@     5//
�!  	hA@     �F  	�A@     ��  	�A@     �6J7tXK�  	B@     �Ju ! 	O+@     �X�/�Y/�Y%/�YE/�+t�D/�/K/$�0��M/2	tKt�X	LU0$ ��KtK	K[g f�#X\�	tKt J tK<$�X	xzX	.u� f t .J!S/0YX00��	w�<g��1g	u�<	�g�<g f  fgt  J t
K�gYvg f t X&=	f&/$f	 =�u�XKg�X�� J t X?�# f J4 f, J> f��u! r�<g]>	 g	�gtKu f � JuK]/0Y2-L<�Y0���=>�?X��4>��	u
g	v L)/�K
uu	�K3K ��	YY'/���Y���� ����/�	��
��
�<uA���gg	
g�%�i �	�Y/0v �*�&�	tK �+�'�
tK<X
N�� � �
 � g � � < / � co  ��>���#��"��	t=�	=K&/�2��-�#6�,�6�,K)�,�L�A;�#�&g�J KQu��AX�� �� �� �� ���t<	/Y&/�A�#=�//�3�)�3.L;v+�Jg
�2i#�Jg�J
�K	�.
g LX0=�"!�f��� ���Y5�?����!>!%�Z!�fK����	�K'0�$��!�fK��  +��	�K;0KJ
g��t
Yu7�".!
uw <�	�Y[v=�� f�}���<J  	$B@     � v
�<g�ut�t!J�u �&�)J�  	�B@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/ 	 	6D@     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	ZY 	 	�F@     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	LY 	 	�H@     	�t�t J tKZt J! � <1 J6 �( <K�Z K&�J� t � J K��X�!�
�f�S6����<# J( � <8 J= �/ <K��YX"L)����	s.<
z<'u�g	�= 
 	�J@     � �/ 
 	K@     � 
	 	"K@     
�/K 
	 	LK@     !�t��K 
	 	xK@     
�/K  	�K@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	
O@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	�S@     �Nu�u
/� ���g�u � .
�f�*�$t��	�gu	�g
0� � � .� � � .��g	hgu%u	�/
0_J #� 
 	�U@     �� X J . K  	V@     � �  	V@     � � 
 	 V@     -�1%  	TV@     ��2 
 	�V@     � �/  	�V@     ��2  	W@     $�/�  	8W@     '��K�  	`W@     ��=��'g !3�(�	<(g" � � � .�	jY  	(X@     ����uf	u.u
fy.�"k  	�X@     7� � � .���  	4Y@     ���  	JY@     �	���# f- �+ � < f t Y  	�Y@     ���fK/[���fKg0#�fKg0t�X  	�Z@     ����uf	u.u
fy.�"k  	D[@     � ��uu���
0K  	�[@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�\@     ���fK/[���fKg0#�fKg0t�X  	�]@     1� � � .���  	 ^@     � � � .�t�J/	PK  	�^@     �=/  	�^@     �=/S  	d_@     �  �u  	u_@     � �(�K  	�_@     � �)�K  	�_@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	b@     � �/�K  	2b@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�d@     �  �u  	�d@     � � � � .��/1  	:e@     ����  	be@     � �(�K  	�e@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�f@     � �)�K  	�f@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	h@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	oj@     � �/�K  	�j@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	m@     �6h:J  	~m@     � � � � .��/1  	�m@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	 o@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	Xp@     �3g71 
 	�p@     0��  � .��gt��������y�	X  	uq@     �	=fY&* � � � .�&  	r@     7��  	*r@     � �-�K  	Hr@     � �uu�(<g  	zr@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	=x@     <�*�=  	Zx@     ���u�<L�0#  	�x@     ���  	�x@     ���  	�x@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	8|@     7��  	N|@     ���u�<L�0#  	�|@     � �-�K  	�|@     � �uu�(<g  	�|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��@     <�*�=  	Ƃ@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�@     � �4  	s�@     � �uu�(<g  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	D�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	�@     &
�Y  	�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	B�@     � �uu�(<g  	s�@     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K 
 	D�@     &  � .��gt���J����� g	   
  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/ansi/include ../options/internal/include/bits ../options/internal/include ../subprojects/cxxshim/stage2/include  formatting.hpp   charcode.hpp   charset.hpp   ctype-stubs.cpp   optional.hpp   string.hpp   logging.hpp   stddef.h   wctype.h   types.h   stdint.h   mbstate.h   type_traits   debug.hpp   <built-in>      	"@@     2&�*M  	A@     1�  	�@     /KJ	=J J �K�)�&�)�(K%�(�K$0�JgZ �� �� Y - 	�@     !1u" f1 f? f1 � t 
Y  	��@     #���
g+u.J =0#���
g+u.J =0#���
g,u/J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g"u%� =0#���
gu� =4)��t
g+u.J =0)��t
g+u.J =0)��t
g,u/J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g"u%� =!.!�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 Ju�/�5 T��	� Y 0��#���
g+Y K0#���
g+Y K4���  	�C@     �<  	�C@     7�  	@�@     �h��K;0  	��@     )��JYu � �gt�$J�K r
wY  	�J@     � �/  	K@     � 	 	"K@     
�/K 	 	LK@     !�t��K  	V@     � �  	V@     � �  	 V@     -�1%  	TV@     ��2  	�V@     � �/  	�^@     �=/  	�p@     0��  � .��gt��������y�	X �)   O  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   environment.cpp   optional.hpp   string.hpp   logging.hpp   vector.hpp   utility   mutex.hpp   utility.hpp   errno.h   stdio.h   stddef.h   types.h   stdint.h   type_traits   debug.hpp   <built-in>      	hA@     �F  	�A@     ��  	�A@     �6J7tXK�  	B@     �Ju 2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	2A@     5//
�!  	N�@     ��#f 2 	�@     % �"�#JK� � �" �1  	 7: � ���K vf
�u4�CK �B JC X	8u0������ � � � � �v�
�w�
 Q0)� #�gu�J.[ ��J�=�
��/��� #�g t � .�   < t X J)��4��w
�� ��*
u!�"J!� t%�,�/� = 0�/�u�Y	5Y@v"����!�0 57��	�K� 2� ��Y	D Y ��Y	&Y  	$B@     � v
�<g�ut�t!J�u �&�)J�  	�B@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/  	@�@     �h��K;0 	 	x�@     5" �  �gt�Y dxu 	 	�J@     � �/ 	 	K@     � 		 	"K@     
�/K  	̨@     
�u 	 	ި@     %
�� 		 	�@     
�/K 		 	LK@     !�t��K  	&�@     � = t � .�1t#  	��@     )��JYu � �gt�$J�K r
wY 
 	��@     �D�H/ 
 	֩@     �� � � fvt�� 
 	�@     � 
�� 
 	.�@     � � � � fv� 
 	b�@     ���/��J<��
=K 
 	ڪ@     ��2/���J<�u
=K 
 	`�@     � 
���= 
 	��@     � 
����= 
	 	��@     � 
�� ! 	��@     0�u  	˫@     ��
K�
u�u 
 	�@     ��="�!�t	�K  	V@     � �  	V@     � � 	 	 V@     -�1%  	TV@     ��2  	c�@     ��6 	 	�V@     � �/  	��@     �#f  	�K@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�   
 	֬@     ��	��tg � �# g, �" � � � ew � � fvt���t�   	�^@     �=/  	٭@     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	W@     $�/�  	8W@     '��K�  	`W@     ��=��'g !3�(�	<(g" � � � .�	jY  	(X@     ����uf	u.u
fy.�"k  	�X@     7� � � .���  	4Y@     ���  	JY@     �	���# f- �+ � < f t Y  	�Y@     ���fK/[���fKg0#�fKg0t�X  	
O@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
 	 	�p@     0��  � .��gt��������y�	X 	 	D�@     &  � .��gt���J�����  	߯@     �=7  	d_@     �  �u  	�]@     1� � � .���  	u_@     � �(�K  	�_@     � �)�K  	�_@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	b@     � �/�K  	2b@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�d@     �  �u  	�d@     � � � � .��/1  	:e@     ����  	be@     � �(�K  	�e@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�f@     � �)�K  	�f@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	�Z@     ����uf	u.u
fy.�"k  	D[@     � ��uu���
0K  	�[@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�\@     ���fK/[���fKg0#�fKg0t�X  	 ^@     � � � .�t�J/	PK  	-�@     �/4  	r@     7��  	*r@     � �-�K  	Hr@     � �uu�(<g  	zr@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	=x@     <�*�=  	Zx@     ���u�<L�0#  	�x@     ���  	�x@     ���  	�x@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	8|@     7��  	oj@     � �/�K  	N|@     ���u�<L�0#  	�|@     � �-�K  	h@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	�j@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	m@     �6h:J  	~m@     � � � � .��/1  	�m@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	 o@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	Xp@     �3g71  	w�@     �	/fY%* � � � .�%  	s�@     � �uu�(<g  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	D�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	�@     &
�Y  	��@     <�*�=  	�|@     � �uu�(<g  	�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	Ƃ@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�@     � �3  	B�@     � �uu�(<g  	h�@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K D    >   �      ../options/ansi/generic  errno-stubs.cpp    l~   �  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   stdio-stubs.cpp   optional.hpp   utility.hpp   logging.hpp   utility   mutex.hpp   string.hpp   errno.h   <built-in>    stdarg.h   stddef.h   ssize_t.h   stdio.h   types.h   stdint.h 	  type_traits   debug.hpp   list.hpp     	hA@     �F  	�A@     ��  	�A@     �6J7tXK�  	B@     �Ju 2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	2A@     5//
�!  	N�@     ��#f  	8�@     � �f  	^�@     � 	���  	��@     � 	*	�/  	�@     � 	=�g  	Z�@     � �f  	��@     � �
t�<g��  	��@     � � � ! � t � < < /	 � �x  	$�@     � � � � � t � < < /	 � �x  	��@     � )�-#  	��@     � ���Yt�<g��  	�@     �� � !
 � �v  	d�@     �> � �
 � �v  	��@     �&�*#  	��@     ����)�"� �3t5�@�K �
��
t	�t�
�� J�  	��@     �	�
t�<g��  	8�@     �� � !
 � �v  	��@     �= � �
 � �v " 	�@     ��4���	�KvX	ug	vYV/Y�K��f�=?���J?Y-	&gI/Y-	&g00Y-	)gL.�-�0�0�0� 0� 0�0�2�"/�<Y\�Y-	*gJ/Y-	&g2�	�0�t�t	�Ov.YX�-&g[/>�02KA�tuJYt � fY0�tuJYt� � fYZl.= t � X J � �' f !@/��@/�7�"
u�'��5J)�f*<,<= K[�>�02JJ<=K`/=@�Y?�YL�<K�<�YJ�YW�tV�t-�Y,�Y9��8��ؼ�
u	u uP0= t���g�=i�
fu�=iw�[g�=`f"XY)0�g�t
K	u Y /�L0�/'t
K	uYC/�/!0��0��0K!0K!(0�g�t
K	u =/�0�g/��08�� X � X	 L ��'WLu	JYww�.�X
K	w Y0�=�. ��9����׺�J��׬ ��H�uuP0uuC0�3�� ���>�$t=0�$t= 0�= t t
K	"+:B� �	�K�	���
Y��2u<X��fK�
��=�=�E�O1�����F�g3�Y-	&gD0>��
2�JJ<=JuK2!�NX��>!�PX��>!�QX��)>��$>�$t=&0�$t="0
��t
K	uJ =Q0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��&�-�t�WM�Y��/t]s�
X&� mf
�vX0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��-�4�t�WM�Y��/t]s�
X&� mf
�v+0/�y�	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=�}.	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=  	$B@     � v
�<g�ut�t!J�u �&�)J�  	�B@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	�C@     �<  	�C@     7�  	��@     � 
��  	�C@     )���u�K&<f/ 
 	�U@     �� X J . K  	��@     #�'f  	�@     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	��@     #�'f  	�@     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X 
 	�A     �� X J . K  	A     #�'f  	0A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	
O@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
 	 	�J@     � �/ 	 	K@     � 		 	"K@     
�/K 		 	�@     
�/K 		 	LK@     !�t��K  	�A     #�'f  	&	A     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	V@     � �  	V@     � � 
! 	�A     0�g  	A     =�  	4A     K  	^A     "=�/  	�A     <�/K  	�A     $(=�K  	$A     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	�A     =�  	.A     K  	XA     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	0A     =�  	bA     K  	�A     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	W@     $�/�  	8W@     '��K�  	JY@     �	���# f- �+ � < f t Y  	�Z@     ����uf	u.u
fy.�"k  	D[@     � ��uu���
0K  	�X@     7� � � .���  	�[@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�\@     ���fK/[���fKg0#�fKg0t�X  	�]@     1� � � .���  	�Y@     ���fK/[���fKg0#�fKg0t�X  	 ^@     � � � .�t�J/	PK 	 	 V@     -�1%  	TV@     ��2  	c�@     ��6 	 	�V@     � �/  	dA     =�  	�A     K  	�A     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	�!A     � �  J �*KJJ�	�' J � < KJ�*>�0./�	<' J �!KJ�)>� 1��� 
 	�"A     �K  	�"A     � � � � .�K  	�"A     ��� � � .� � � .� � � .� � � .�0/.%Z � � .� � � .� � � .� � � .� f � .� < � .�-Z � � .� � � .��	J.u$��= <) � . X t XK�Z�K t � = �h" f t � �i" f t Y �h t � u �j f � .�	J.u3��= <) � . X t XK�Z�� t � � 'h" f t � �i" f t Y �h t � � 'l � . �*$   	V)A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	0*A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	+A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�+A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�,A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�-A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	f.A     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	6A     ��_/0 � .� 		 	�6A     
/K  	�6A     ��� � � .� � � .� � � .� � � .�0/.%Z � � .� � � .� � � .� � � .� f � .� < � .�-Z � � .� � � .��	J.u$��= <) � . X t XK�Z�K t � = �h" f t � �i" f t Y �h t � u �j f � .�	J.u3��= <) � . X t XK�Z�� t � � 'h" f t � �i" f t Y �h t � � 'l � . �*$   	"=A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�=A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�>A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�?A     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�@A     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	\AA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	2BA     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	�IA     ��_/0 � .�  	KJA     ��� � � .� � � .� � � .� � � .�0/.%Z � � .� � � .� � � .� � � .� f � .� < � .�-Z � � .� � � .��	J.u$��= <) � . X t XK�Z�K t � = �h" f t � �i" f t Y �h t � u �j f � .�	J.u3��= <) � . X t XK�Z�� t � � 'h" f t � �i" f t Y �h t � � 'l � . �*$   	�PA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�QA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	tRA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	NSA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	$TA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�TA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	�UA     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	�]A     ��_/0 � .�  	d_@     �  �u  	be@     � �(�K  	�f@     � �)�K  	h@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	oj@     � �/�K  	�j@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�d@     �  �u  	m@     �6h:J  	4Y@     ���  	~m@     � � � � .��/1  	:e@     ����  	u_@     � �(�K  	�m@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�_@     � �)�K  	 o@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	�d@     � � � � .��/1  	�e@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�f@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	Xp@     �3g71  	�^@     �=/  	٭@     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	�]A     ��� � � .� � � .� � � .� � � .�0/.%Z � � .� � � .� � � .� � � .� f � .� < � .�-Z � � .� � � .��	J.u$��= <) � . X t XK�Z�K t � = �h" f t � �i" f t Y �h t � u �j f � .�	J.u3��= <) � . X t XK�Z�� t � � 'h" f t � �i" f t Y �h t � � 'l � . �*$   	fdA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	@eA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	fA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�fA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�gA     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�hA     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	viA     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	+qA     ��_/0 � .� 
 	�qA     ��
=�
g�g 
! 	�qA     0�u 
 	�qA     ��
=�
g�g  	4rA     � �4  	@�@     �h��K;0 	 	ި@     %
��  	�rA     �h�K;0 	 	�rA     %
��  	�rA     � �Fu	Ju4,4  	�sA     � �3  	�sA     � �4  	CtA     ��4  	�tA     � �4  	�tA     � �Fu	Ju4,4  	�uA     � �3  	�uA     � �4  	,vA     � �4  	�vA     � �Fu	Ju4,4  	"wA     � �3  	wwA     � �4  	8|@     7��  	�|@     � �-�K  	�|@     � �uu�(<g  	�|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��@     <�*�=  	N|@     ���u�<L�0#  	�x@     ���  	�x@     ���  	Ƃ@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	r@     7��  	b@     � �/�K  	Zx@     ���u�<L�0#  	*r@     � �-�K  	�x@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/  	 	�p@     0��  � .��gt��������y�	X 	 	D�@     &  � .��gt���J�����  	߯@     �=7  	�wA     � �4  	%xA     � �Fu	Ju4,4  	�xA     � �3  	yA     � �4  	pyA     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	{A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�|A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	_~A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     �/4  	Q�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	@�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	8�A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	׋A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	B�@     � �uu�(<g  	�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	�@     &
�Y  	=x@     <�*�=  	Hr@     � �uu�(<g  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	D�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	-�@     �/4  	�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	'�A     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	ϐA     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	n�A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K  	�A     �	/fY%* � � � .�%  	w�@     �	/fY%* � � � .�%  	��A     � �Fg	<Y3,3  	�@     � �3  	h�@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	J�A     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h K   �   �      ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  string-stubs.cpp   errno.h   stddef.h    6 	ޖA     ���	t K�<�-0	uKH/�	��t J ��<�/V
2��=V	2KA0��	YKS/=���	K�t J ��<�/V2	uK70� �8��8g�g�u� zt	|Y*/	���=�= fgv�u�uY/+0�/<0	���u�=�= fgv�u�uY/T/=1��� ���<2K �	wY$/	��	!#Y�U3"g	�Y1/	�
�� J �  X t XKgV 20/	��!�f#K�U	3Y%/�� ����*Y.� �	xY0/	�
��  J �  X t XKgV 22/� �YK �!� J �+ � �
MK+|#g u�	�YD/�'�	��	!#Y�U!3�@0�?��F��C�.I�.M�.S�.A��J�<�<7�<A��J�<.��/��7�<E�<7�<+��2��4��,��1��3��W�<<��� ��J)Y,� �	wY 0�.�.�v35�Y.�Y2�Y3�Y0�Y4�Y0�Y&�Y5�/9�/-�/D�/9�/7�/*�/1�/7�0�K33/	�h�t
K	uY80=*�uA0���� �   �  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/lsb/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   dso_exit.cpp   utility   eternal.hpp   vector.hpp   mutex.hpp   stddef.h   types.h   stdint.h   type_traits   <built-in>      	hA@     �F  	�A@     ��  	�A@     �6J7tXK�  	B@     �Ju 2 	@@     	�K  	$B@     � v
�<g�ut�t!J�u �&�)J�  	�B@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	��A     9M �8 J9 X��U0>����	�Y0�� � u � t �x  	��A     �K  	��A     '���  	�A     *�K  	��A     ���/���<��
=K 	 	��A     � 
��  	��A     � 
��=  	ʧA     �#  	��A     �D�H/  	6�A     ���	��t� � � g <# f, �" < �w � � fvt���t�   	
O@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
 ! 	J�A     0��  	�K@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�   	 	W@     $�/� 	 	8W@     '��K�  	JY@     �	���# f- �+ � < f t Y  	�Z@     ����uf	u.u
fy.�"k  	D[@     � ��uu���
0K 	 	�X@     7� � � .���  	�[@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�\@     ���fK/[���fKg0#�fKg0t�X 	 	�]@     1� � � .���  	�Y@     ���fK/[���fKg0#�fKg0t�X  	 ^@     � � � .�t�J/	PK  	`W@     ��=��'g !3�(�	<(g" � � � .�	jY  	(X@     ����uf	u.u
fy.�"k  	4Y@     ���  	d_@     �  �u  	be@     � �(�K  	�f@     � �)�K  	h@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	oj@     � �/�K  	�j@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�d@     �  �u  	m@     �6h:J  	~m@     � � � � .��/1  	:e@     ����  	u_@     � �(�K  	�m@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�_@     � �)�K  	 o@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	�d@     � � � � .��/1  	�e@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�f@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	Xp@     �3g71  	�_@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	b@     � �/�K  	2b@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	8|@     7��  	�|@     � �-�K  	�|@     � �uu�(<g  	�|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��@     <�*�=  	N|@     ���u�<L�0#  	�x@     ���  	�x@     ���  	Ƃ@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	r@     7��  	Zx@     ���u�<L�0#  	*r@     � �-�K  	�x@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	Hr@     � �uu�(<g  	zr@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	=x@     <�*�=  	B�@     � �uu�(<g  	�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	�@     &
�Y  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	D�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	s�@     � �uu�(<g ?   �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  lemon.cpp   types.h   stdint.h   stddef.h     	z�A     
�%5>� �
�	-tY
uY00
�Y0K� g 6   �  �      ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/internal/generic ../subprojects/frigg/include/frg /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  new   allocator.hpp   allocator.cpp   eternal.hpp   utility   slab.hpp   rbtree.hpp   stddef.h   types.h   stdint.h   mutex.hpp   type_traits   sysdeps.hpp   <built-in>     2 	@@     	�K  	��A     �� ! 	Z�A     (M � JGu � J'�0B� ��K@>= ��  	��A     ��  	ܫA     *�K  	�A     �K  	��A     '���  	H�A     *�K  	V�A     �t  	h�A     ��  	��A     �/ G X  
  	
�A     ����  	.�A     ��( ! 	e�A     �  	p�A     � ��  	��A     ����  	��A     � �� �   �  �      ../options/internal/include/mlibc ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include  charcode.hpp   charcode.cpp   stddef.h   types.h   stdint.h   optional.hpp   logging.hpp   mbstate.h   type_traits   debug.hpp   hash.hpp   formatting.hpp   <built-in>      	��A     � S!W(  	ڮA     � J  	��A     �'f  	
�A     �#t  	�A     .�)t	<=f�JL��u�u��u�u��u�u� � ��x ��t$Xt.uf
�t�Y  	��A     ;=	tY f
�tYt�t�Y  	��A     +�X�*��5K � J
5uB0��Y)0
Lu  	"�A     � E�I(  	Z�A     � �!  	��A     � �  	��A     � � ��/� � � t X�Xg�LJuKut�/tt�XKu Y  	 �A     � v ��/� � � t X�Xg�KJvKu�t/tt�XKu Y  	H�A     �v ��/���XgZKJvKuv XKu Y  	\�A     �v ��1 � � t X�tY<K�+��K�
hgZ ��t�Jx�y XJtYu Y  	��A     
�t�  	ԶA     
�t�  	��A     
�t�  	�A     
�t�  	4�A     
�t� �   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   charset.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   debug.hpp   charcode.hpp   charset.hpp   <built-in>     2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1� # 	T�A     	�Y%>u# � � J t X!K �! �. �! �9 X! .9 X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y&0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X)�z� �+ �7 �C �� � �* �6 �B �� � �� � �) �5 �A ��� � �* �6 �B � � � �) � �1 X) 	.1 	X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��)�3��	�Y%>u# � � J t XGK �  �- �: �G 
� �O XG .O X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y*0u# � � J t XK �����-X�	�g*0u# � � J t XK �����-X�	�g0
Lu  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/  	�J@     � �/  	K@     � 	 	"K@     
�/K 	 	LK@     !�t��K 	 	��A     
�/K  	V@     � �  	V@     � �  	 V@     -�1%  	TV@     ��2  	�V@     � �/  	��A     ��0  	�^@     �=/  	-�@     �/4  	�p@     0��  � .��gt��������y�	X  	w�@     �	/fY%* � � � .�%  	�@     � �3  	h�@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K  	D�@     &  � .��gt���J����� *      �      ../options/internal/generic ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc  debug.cpp   optional.hpp   logging.hpp   type_traits   debug.hpp   formatting.hpp   <built-in>     1 	4�A     
��2L�� �	   m  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic ../options/internal/include/mlibc /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  new   formatting.hpp   ensure.cpp   optional.hpp   logging.hpp   utility.hpp   type_traits   debug.hpp   stddef.h   <built-in>     2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	u�A     &�,�!  # +�� # 6���?&�+�!  # +�� # 6���  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/  	��A     � �/  	��A     � 	 	��A     
�/K 	 	��A     
�/K 	 	�A     !�t��K  	�J@     � �/  	K@     � 	 	"K@     
�/K 	 	��A     
�/K 	 	LK@     !�t��K  	V@     � �  	V@     � �  	B�A     -�1%  	v�A     ��2  	��A     ��0  	��A     � �/  	 V@     -�1%  	TV@     ��2  	��A     ��0  	�V@     � �/  	$�A     �=/  	N�A     �/4  	�^@     �=/  	-�@     �/4  	��A     0��  � .��gt��������y�	X  	i�A     �	/fY%* � � � .�%  	�p@     0��  � .��gt��������y�	X  	w�@     �	/fY%* � � � .�%  	�A     � �3  	�@     � �3  	Z�A     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	h�@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K  	��A     &  � .��gt���J�����  	D�@     &  � .��gt���J�����    �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/gcc /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   guard-abi.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   debug.hpp   <built-in>     2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	2A@     5//
�!  	��A     �"u!��N�+$0��uF<��)�3���R>���J8<XK
�vZS/��Ju�  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/  	��A     � �/  	��A     � 	 	��A     
�/K 	 	��A     
�/K 	 	�A     !�t��K  	V@     � �  	V@     � �  	B�A     -�1%  	v�A     ��2  	�A     ��2  	��A     � �/  	$�A     �=/  	^�A     �=/S  	��A     0��  � .��gt��������y�	X  	��A     �	=fY&* � � � .�&  	z�A     � �4  	��A     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	�@     �� J J . K  	��A     &  � .��gt���J����� �4   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include/mlibc ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/posix/include/bits/posix  new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   file-io.cpp   optional.hpp   list.hpp   logging.hpp   utility.hpp   allocation.hpp   utility   intrusive.hpp   mutex.hpp   file-io.hpp   errno.h   stddef.h   types.h   stdint.h 	  ssize_t.h 
  stdio.h   off_t.h 
  type_traits   debug.hpp   <built-in>     2 	@@     	�K  	"@@     2&�*M  	~@@     1��  	A@     1�  	hA@     �F  	�A@     ��  	�A@     �6J7tXK�  	B@     �Ju  	z�A     /V�D��������!�/> K��Y�Y���Y��-��Yv<
����Z��"MB' ���XK!��0��g��tY�
�� J �Y�Y������ g� g�;�)g��tY���!$ ��/�-�fBJ� ��JY�	� YT>' ���XK!��� �1��g�� ��
���Y g� g�� J �Y�Y��� ��(�&�:�X:<wK�,Y�u�
tuM ���	t��<"��+Y�3��<'�0��7��<�����-��$�:��<��g�XKw	 Y#> ��
����<g5L� J�	�Y0������M��00.���
g)Z#�;<3� <t	u Y30/�
g�&g �8<0�<6��<�/[ f f1��<g/^	� Y!>�t
K"v�f
gY �	�Y$>�t
K v�!<XKu �	�Y">��
g���
Y�tVZ��3<��g��� �� J���V�3�A��f&�$�J.g/Z ��gxf	XY>��
g�tY J� J���	�Y*0� ���[$�g�$B$/(/L	�u>!��Y�Y��<
g	YY0>�"	g
�u	�
�v >30��	�
��<	g
�u	�
�v�&X��ZJ>v�
gY	� YQ>v�
gY	� YC>g�
g	YY
<�L" 1 � / �g�Y� � �]&D� t � X K �0��&-<E�7�S�&<S�&<S�1U��"<��K
g���K
g�	v��6�7�?�K����	���K�	�K�	�
Ku��7�? K���v�X�	u
g5v'�TY X f Y&6E�7�S�&<S�&<S�(z�u�Y��5�'�TY X fY0� t � X K u � XKu��XKu	�=50/ t � X K �	ug	vY0� t � X L X	ug	� K&0� t � X K � X
K	uY/��C0h t � X K"g<
�g�"g<
ugv"g<
ug	�K	wY0� t � X K Y /$>� t � X K	 = = 0� t � X K ��{<�Kv.�*K3�*<	�3�	J3�=��Kv.�*K3�*<	�3�	J3�=��� ��{���X�X�X��&<J  	$B@     � v
�<g�ut�t!J�u �&�)J�  	�B@     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	�C@     �<  	�C@     7�  	�C@     )���u�K&<f/  	��A     � "�&f  	��A     3�7�  	�A     �  � � .(�� � � .� � � .� � � .��Y���.K�f>�.Kg 	 	�J@     � �/ 	 	K@     � 		 	"K@     
�/K 		 	LK@     !�t��K  	�K@     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	��A     � � � � .�g  	�A     � � � .� � � .1�!.�,K.�JY  � .�� 0 � .�J�Nu � � .�J�� / � .#�. ��.? � � .�.u.�.
LK 	 	��A     � �/ 	 	��A     � 		 	��A     
�/K 		 	�A     !�t��K 

 	�A     �� X J . K 

 	�U@     �� X J . K  	
O@     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	��A     �(�%  	&�A     ��K  	J�A     ;�.=  	r�A     ?��uK  	��A     4�u 		 	�6A     
/K  	��A     �v/�#  	�"A     �K  	V@     � �  	V@     � �  	��A     
�K  	
�A     $��� ! 	:�A     0�u  	L�A     1�� 	 	 V@     -�1%  	TV@     ��2 	 	�V@     � �/  	W@     $�/�  	8W@     '��K�  	`W@     ��=��'g !3�(�	<(g" � � � .�	jY  	(X@     ����uf	u.u
fy.�"k  	�X@     7� � � .���  	4Y@     ���  	JY@     �	���# f- �+ � < f t Y  	�Y@     ���fK/[���fKg0#�fKg0t�X 	 	B�A     -�1%  	v�A     ��2 	 	��A     � �/  	�Z@     ����uf	u.u
fy.�"k  	D[@     � ��uu���
0K  	�[@     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�\@     ���fK/[���fKg0#�fKg0t�X  	�]@     1� � � .���  	 ^@     � � � .�t�J/	PK  	f�A     8�t� 	 	��A     ,� ��  	CtA     ��4  	��A     �K��/[4��K � � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY s�k�$  
 	��A     !��  	�A     ��  	�^@     �=/  	d_@     �  �u  	u_@     � �(�K  	�_@     � �)�K  	�_@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	b@     � �/�K  	2b@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�d@     �  �u  	�d@     � � � � .��/1  	:e@     ����  	be@     � �(�K  	�e@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	�f@     � �)�K  	�f@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	$�A     �=/  	h@     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	oj@     � �/�K  	�j@     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	m@     �6h:J  	~m@     � � � � .��/1  	�m@     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	 o@     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	Xp@     �3g71  	�A     �/4 
 	(�A     �K 	 	�p@     0��  � .��gt��������y�	X  	r@     7��  	*r@     � �-�K  	Hr@     � �uu�(<g  	zr@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	=x@     <�*�=  	Zx@     ���u�<L�0#  	�x@     ���  	�x@     ���  	�x@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	8|@     7��  	N|@     ���u�<L�0#  	�|@     � �-�K 	 	��A     0��  � .��gt��������y�	X  	�|@     � �uu�(<g  	�|@     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��@     <�*�=  	Ƃ@     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	�A     �	/fY%* � � � .�%  	s�@     � �uu�(<g  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	D�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�@     &
�Y  	�@     &
�Y  	�@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��@     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	B�@     � �uu�(<g  	��A     � �Fg	<Y3,3  	h�@     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	J�A     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 

 	�@     �� J J . K 	 	D�@     &  � .��gt���J�����  	6�A     � �!  	d�A     � � j   �   �      ../sysdeps/lemon/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  filesystem.cpp   stddef.h   ssize_t.h   off_t.h    K 	��A     !g3Jhuv
�YE0jJhuv
�YD0\vuv
�Y81/>uv
�Y1�
�Y01�>g�uY 0�         __io_offset mouseDown __in_chrg next uintptr_t _ZN4ListIP8Window_sE8add_backES1_ uint64_t title _ZN4ListIP8Window_sEC4Ev __static_initialization_and_destruction_0 dragOffset __offset handle_t lastUptimeMilliseconds 13ipc_message_t stdout colourPlanes senderPID __mlibc_uintptr RemoveDestroyedWindows long long int __mlibc_uint64 mouseEventMessage closeInfoHeader closeButtonSurface fb_info_t redrawWindowDecorations __buffer_ptr _ZN4ListIP8Window_sE10get_lengthEv mouseDevice Vector2i lastUptimeSeconds active remove_at _ZN4ListIP8Window_sE9get_frontEv stdin _ZN8ListNodeIP8Window_sEC4Ev List<Window_s*> uint16_t _Z13AddNewWindowsv linePadding _ZN10win_info_tC4Ev this closeButtonBuffer _windowCount long double compression _Z15UpdateFrameRatev currentUptimeSeconds GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions __initialize_p _ZN4ListIP8Window_sE9remove_atEj get_front colourNum RGBAColour _Z10DrawWindowP8Window_s 20bitmap_file_header_t data short unsigned int AddNewWindows UpdateFrameRate depth _ZN4ListIP8Window_sE8get_backEv _ZN4ListIP8Window_sEC2Ev recieverPID __status_bits decltype(nullptr) FBInfo difference operator[] windowFound __mlibc_uint16 vector2i_t fbInfo windowInfo 20bitmap_info_header_t pitch /home/computerfido/Desktop/Lemon/Applications/Init frameRate __mlibc_int8 _ZN4ListIP8Window_sEixEj _ZN8ListNodeIP8Window_sEC2Ev __dirty_begin float _ZN10win_info_tC2Ev closeButtonFd operator+ _ZN4ListIP8Window_sE6get_atEj importantColours unsigned char _ZN4ListIP8Window_sED2Ev short int magic main.cpp 10win_info_t __mlibc_uint8 vres FILE currentUptimeMilliseconds clear ListNode uint32_t surface_t mouseX _ZplRK8Vector2iS1_ mouseY __mlibc_uint32 get_length info __dirty_end data2 _ZN4ListIP8Window_sE9add_frontES1_ _ZN4ListIP8Window_sE10replace_atEjS1_ _ZN4ListIP8Window_sE5clearEv hdrSize add_back drag replace_at get_at stderr ListNode<Window_s*> closeButtonLength add_front renderPos _Z22RemoveDestroyedWindowsv prev lastKey fbSurface uint8_t DrawWindow windows renderBuffer flags windowHandle __valid_limit hres backgroundColor __io_mode __buffer_size __mlibc_int32 _ZN4ListIP8Window_sED4Ev mousePos ~List height rgba_colour_t __priority main mouseData __dso_handle get_back ownerPID frameCounter keyMsg _GLOBAL__sub_I_keymap_us lemon_readdir ../sysdeps/lemon/generic/filesystem.c /home/computerfido/Desktop/Lemon/LibC/build lemon_dirent filename lemon_close off_t inode GNU C17 8.2.0 -mtune=generic -march=x86-64 -g -fno-builtin -fPIC lemon_open whence lemon_dirent_t lemon_write lemon_read lemon_seek ReceiveMessage SendMessage queue_size ../sysdeps/lemon/generic/ipc.c syscall arg0 arg1 arg2 arg4 ../sysdeps/lemon/generic/syscall.c arg3 ../sysdeps/lemon/generic/fb.c lemon_map_fb itoa reverse ../sysdeps/lemon/generic/itoa.c strlen src_bytes ../options/internal/generic/essential.cpp GNU C++17 8.2.0 -mtune=generic -march=x86-64 -g -std=c++17 -fno-builtin -fno-rtti -fno-exceptions -fPIC dest_bytes _ZN5mlibc10infoLoggerE mb_chr _ZN3frg11unique_lockI13AllocatorLockEC4EOS2_ aggregate<frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame> size_to_bucket _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14size_to_bucketEm _ZN3frg7mt19937C2Ev _stor _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE6bucketC4Ev alignment _ZN3frg11unique_lockI13AllocatorLockEC4ENS_11dont_lock_tERS1_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ replacement _ZN3frg7mt199371nE _ZN3frg8optionalIiE6_resetEv mag01 item_size code_seq<char const> _ZN3frg14format_optionsD2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4ERKSB_ stack_buffer_logger<mlibc::PanicSink, 128> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN3frg8optionalIiEC4ENS_13null_opt_typeE mbstowcs lldiv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE12huge_paddingE __func__ _tree_mutex digits strtold nptr strtoll plus_becomes_space print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> lsbs _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ get_root dont_lock_t ~storage_union __mlibc_rand_engine _is_locked _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg10bitop_implImE3clzEm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ operator<< <void*> absv _verify_integrity max_bucket_size _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ _ZN3frg11unique_lockI13AllocatorLockED2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EaSERKSB_ atof rotateRight _fmt_basics locale_t __cpoint _ZN5mlibc7strtofpIeEET_PKcPPc _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic endptr _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ _ZN3frg14format_optionsC2ERKS0_ aggregate_node _usedPages _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ atoi atol illegal_input endlog decimal mb_string address_ frame_hook _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ ~item _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE23test_bucket_calculationEj InfoSink _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ _ZN5mlibc8InfoSinkclEPKc wctomb _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14small_step_expE _ZN3frg7mt199378matrix_aE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE17_verify_integrityEv message insert_right left_ptr __mlibc_errno copy _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ area_size _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEv _ZN3frg9_redblack15null_aggregator9aggregateINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ is_constructible<int, const frg::optional<int>&> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ seed _ZN13AllocatorLock4lockEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ operator* _ZN5mlibc7strtofpIfEET_PKcPPc type_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ abort _ZN13AllocatorLockC4ERKS_ operator= _ZNSt16is_constructibleIiJRKN3frg8optionalIiEEEE5valueE _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEv slab_allocator _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ _ZN3frg14format_optionsC4ERKS0_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameC4ERKS4_ stack_buffer_logger<mlibc::InfoSink, 128> _ZN5mlibc8code_seqIwEcvbEv _ZN3frg11unique_lockI13AllocatorLockE9is_lockedEv realloc result num_buckets slabsize _construct_large 7lldiv_t _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE15max_bucket_sizeE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameC4Emmi tree_struct<frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> num_reserved with_conversion insert_root _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ rbtree _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ successor negative _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistC4Ev _ZN3frg14format_optionsC4Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemaSERKS4_ _ZN3frg9_redblack11hook_structC4ERKS1_ partial_hook bucket_mutex _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ isRed wchar_t link fix_insert _ZN3frg9_redblack11hook_structC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv _ZN5mlibc8InfoSinkC4Ev llabs other color_type mblen_state calloc 5div_t Limit Args VirtualAllocator was_unavailable _ZN3frg8optionalIiE13storage_unionD4Ev panicLogger ~format_options minimum_width deallocate predecessor mblen _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4ERKSB_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ left_justify append _ZN3frg11unique_lockI13AllocatorLockE8protectsEPS1_ _emit print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> compare _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ malloc _ZNK3frg8optionalIiEcvbEv check_invariant is_constructible<int, frg::optional<int>&&> _frame_tree succ strtod_l _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameC4ERKS4_ object _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ replace_node _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4EPS3_ rand_r Member frame_type _ZSt18is_constructible_vIiJON3frg8optionalIiEEEE program_invocation_name strtoul cutlim _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ atoll _Exit dot_end _ZN3frg11unique_lockI13AllocatorLockEaSES2_ strtofp<double> operator<< grand _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE9page_sizeE operator<< <char const*> frame_less _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE23_verify_frame_integrityEPNS3_5frameE format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> status address endlog_t 6ldiv_t _non_null _ZN3frg8optionalIiEcvbEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ _ZN3frg8optionalIiED4Ev output_overflow code_seq<wchar_t> wcstombs max_size get_right _ZN16VirtualAllocator3mapEm frame_tree_type slab_frame length_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE7reallocEPvm remove_half_leaf format<void*, frg::stack_buffer_logger<mlibc::InfoSink>::item> numUsedPages _ZNK3frg8optionalIiE9has_valueEv _ZN3frg8optionalIiEdeEv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8slabsizeE _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc _ZN3frg11unique_lockI13AllocatorLockE6unlockEv _ZN3frg11unique_lockI13AllocatorLockED4Ev _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4Ev _ZN3frg11unique_lockI13AllocatorLockEC4ERS1_ Mutex _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ aligned_alloc ~optional _plcy new_length _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ freelist _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistaSERKS4_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEC4ES2_ has_value child max<int> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZNSt16is_constructibleIiJON3frg8optionalIiEEEE5valueE _ZN3frg8optionalIiEC4EOi is_constructible_v _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ _ZN3frg8optionalIiEC2Ev unmap _verify_frame_integrity bsearch _ZN3frg8optionalIiEaSES1_ _ZN3frg7mt19937C4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ infoLogger slab_allocator<VirtualAllocator, AllocatorLock> _ZN3frg14format_options15with_conversionENS_17format_conversionE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ _redblack _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE16_construct_largeEm _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE15_construct_slabEi input_underflow optional<int> tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::_redblack::null_aggregator> operator new _ZN3frg8optionalIiEptEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev operator bool _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EaSERKSB_ isBlack system small_step_exp _ZN3frg11unique_lockI13AllocatorLockEC4ERKS2_ partial_tree tree_crtp_struct _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameaSERKS4_ _ZN3frg7mt199374lsbsE protects _ZN3frg8optionalIiEC4ERKi _GLOBAL__sub_I_stdlib_stubs.cpp _ZnwmPv strtoull _ZN16VirtualAllocator5unmapEmm format_object<frg::stack_buffer_logger<mlibc::InfoSink>::item> qsort overhead _ZN3frg8optionalIiE13storage_unionC2Ev null_opt_type _ZN3frg3maxImEERKT_S3_S3_ v_bytes _ZN3frg3maxIiEERKT_S3_S3_ enable_checking _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ _ZN13AllocatorLockaSERKS_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5firstEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ long long unsigned int _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4ERKS4_ get_parent _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ fill_zeros _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ AllocatorLock _ZN3frg7mt199373msbE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _ZNK3frg8optionalIiEdeEv mb_limit max<long unsigned int> program_invocation_short_name hook_struct head_slb _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameC4ENS3_10frame_typeEmm strtofp<float> _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm mbtowc get_left rotateLeft null_aggregator operator() _ZN5mlibc11panicLoggerE quot parent_color _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::_redblack::null_aggregator> _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE11_find_frameEm u_bytes _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm wc_limit format_conversion ULONG_MAX _sink _ZN3frg9_redblack15null_aggregator9aggregateINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ _reset _ZN3frg14format_optionsD4Ev number _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10tiny_sizesE _ZN3frg7mt199374seedEj wseq _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv tree_struct<frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> _bkts new_pointer _ZN3frg8optionalIiED2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ mktemp _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi bucket_guard unique_lock<AllocatorLock> matrix_a rbtree_hook at_quick_exit small_base_exp _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC4ERS1_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameaSERKS4_ index_ strtod strtof _ZN3frg8optionalIiE13storage_unionC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv strtol tiny_sizes null_opt right_ptr _off func _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj tree_guard huge_padding _ZN3frg8optionalIiEC4EOS1_ precision _emitted _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ aggregate<frg::slab_allocator<VirtualAllocator, AllocatorLock>::slab_frame> charcode_error element Policy _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ alt_conversion aggregate_path _ZN3frg9_redblack11hook_structaSERKS1_ __progress strtofp<long double> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistC2Ev unlock _ZN3frg14format_optionsC2Ev stack_buffer_logger _ctr test_bucket_calculation srand _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE11num_bucketsE partial_tree_type _ZN13AllocatorLockC4Ev tree_struct _ZN3frg8optionalIiEC2ERKS1_ radix _ZN3frg9_redblack11hook_structC2Ev ../options/ansi/generic/stdlib-stubs.cpp cutoff _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ ~unique_lock _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE12numUsedPagesEv operator-> bucket_to_size _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ _ZN3frg8optionalIiE13storage_unionD2Ev mlibc _futex contains _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frame8containsEPv always_sign insert_left page_size _ZN5mlibc7strtofpIdEET_PKcPPc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ __shift mt19937 _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ _ZN3frg8optionalIiEC4Ev _ZSt18is_constructible_vIiJRKN3frg8optionalIiEEEE _ZN5mlibc8code_seqIKcEcvbEv _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ wc_string _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14small_base_expE _find_frame dont_lock _construct_slab _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ dirty denom posix_memalign _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ format<char const*, frg::stack_buffer_logger<mlibc::InfoSink>::item> bitop_impl<long unsigned int> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD4Ev pred _ZN3frg8optionalIiEC4ERKS1_ _ZN13AllocatorLock6unlockEv fix_remove _ZN3frg11unique_lockI13AllocatorLockEC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ _ZN3frg7mt199371mE _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN3frg7mt19937clEv srandom _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistC4ERKS4_ _ZN5mlibc8code_seqIjEcvbEv iswlower iscntrl isalnum _ZN3frg17basic_string_viewIcE10find_firstEcm _ZNK3frg17basic_string_viewIcE4sizeEv isprint isdigit isspace ct_digit _ZN3frg17basic_string_viewIcEC2EPKc ct_space iswspace ispunct _ZN5mlibc13wide_charcode7promoteEwRj _ZNK3frg17basic_string_viewIcEneES1_ isupper ct_punct iswcntrl toupper generic_is_control iswdigit iswpunct isgraph iswprint ct_graph isalpha basic_string_view towupper ct_alpha _ZN5mlibc18generic_is_controlEj _ZNK3frg17basic_string_viewIcEixEm iswxdigit _ZN3frg17basic_string_viewIcEC4EPKc basic_string_view<char> _ZN3frg17basic_string_viewIcEC4EPKcm ct_alnum isblank sub_string ct_blank codepoint _ZNK3frg17basic_string_viewIcEeqES1_ ct_cntrl iswblank find_first ct_upper iswalpha find_last iswctype _ZN3frg17basic_string_viewIcEC4Ev iswupper tolower operator== ct_print operator!= ct_xdigit code_seq<unsigned int> wint_t towlower isascii _ZN5mlibc20polymorphic_charcode7promoteEcRj promote _ZNK3frg17basic_string_viewIcE4dataEv iswgraph ct_count isxdigit ct_null _ZN3frg17basic_string_viewIcE9find_lastEc iswalnum islower Char _ZN3frg17basic_string_viewIcE10sub_stringEmm wctype_t ct_lower ../options/ansi/generic/ctype-stubs.cpp _ZN3frg10escape_fmtC2EPKvm _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERS5_ unsetenv self _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ _ZN3frg17basic_string_viewIcEC2EPKcm _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ _ZN3frg10escape_fmtC4EPKvm update_vector _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED4Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv push format_integer<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv new_capacity push_back putenv _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv move<char*&> getenv remove_reference<char*&> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4EOS6_ ../options/ansi/generic/environment.cpp _ZSt4swapIPcEvRT_S2_ unassign_variable operator<< <frg::escape_fmt> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev escape_fmt _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv environ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backEOS1_ ~vector _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm get_vector empty_environment _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backERKS1_ print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> _ensure_capacity remove_reference_t format<frg::escape_fmt, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERKS6_ overwrite vector<char*, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic swap<char*> _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv format<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic new_array _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> empty _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv start_from _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEaSES6_ find_environ_index _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5emptyEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ERS5_ _elements _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ ../options/ansi/generic/errno-stubs.cpp print_int<StreamPrinter, long int> _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic _ZN3frg17basic_string_viewIwE9find_lastEw do_printf_ints<StreamPrinter> fgetc printf_format<PrintfAgent<StreamPrinter> > chunk print_int<ResizePrinter, long int> print_int<StreamPrinter, long unsigned int> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev format_integer<int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic vfprintf _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN11PrintfAgentI14LimitedPrinterEclEc fputc_unlocked ferror_unlocked _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_digits<BufferPrinter, long int> vswscanf fread_unlocked print_digits<ResizePrinter, long unsigned int> _ZN13ResizePrinter6expandEv BufferPrinter renameat _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev vasprintf _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _vsp putchar __mlibc_intmax remove_reference<int&> print_digits<BufferPrinter, long long unsigned int> ~<lambda> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev print_int<ResizePrinter, long long unsigned int> fgetpos new_buffer ssize_t clearerr _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic _ZN13StreamPrinter6appendEPKcm SCANF_TYPE_INT _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic ftrylockfile SCANF_TYPE_SIZE_T vfscanf _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN13StreamPrinter6appendEPKc print_digits<BufferPrinter, long unsigned int> do_scanf<sscanf(char const*, char const*, ...)::<unnamed class> > vwprintf swap<int> _ZN3frg4swapERNS_8optionalIiEES2_ printf_format<PrintfAgent<LimitedPrinter> > _ZNK3frg17basic_string_viewIwEneES1_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ print_digits<LimitedPrinter, long int> bytes_read print_int<BufferPrinter, unsigned int> _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ vscanf _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ print_digits<ResizePrinter, long long unsigned int> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN3frg17basic_string_viewIwEC2EPKw PrintfAgent _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ <lambda(auto:1)> fgetwc getwchar _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_int<LimitedPrinter, long int> fgetws _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ do_printf_chars<LimitedPrinter> feof_unlocked _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE native_size _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ __builtin_va_list do_scanf<vfscanf(FILE*, char const*, __va_list_tag*)::<unnamed struct> > _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ do_printf_floats<LimitedPrinter> __gnuc_va_list handler _ZNK3frg17basic_string_viewIwE4sizeEv clearerr_unlocked _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZN13BufferPrinterC2EPc _ZN11PrintfAgentI13StreamPrinterEC4EPS0_PN3frg9va_structE move<bool&> print_int<BufferPrinter, long unsigned int> _ZN14LimitedPrinter6appendEPKcm fwrite_unlocked _ZN13BufferPrinterC4EPc _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE vfwscanf _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE print_digits<StreamPrinter, long unsigned int> do_printf_chars<BufferPrinter> actual_size do_printf_floats<BufferPrinter> _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic ungetwc fp_offset ptrdiff_t new_limit _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg8optionalIiEC4IRivEEOT_ stream operator<< <char> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ format<char, frg::stack_buffer_logger<mlibc::InfoSink>::item> vsnprintf _ZN11PrintfAgentI13BufferPrinterEclEc new_path _ZSt4swapIiEvRT_S1_ vswprintf _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE szmod fputs_unlocked _ZNK3frg17basic_string_viewIwEixEm fwide _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic funlockfile _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _ZSt18is_constructible_vIiJRiEE putchar_unlocked _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ print_int<StreamPrinter, unsigned int> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE putwchar SCANF_TYPE_PTRDIFF print_int<ResizePrinter, unsigned int> _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ remove_reference<bool&> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN3frg17basic_string_viewIwE10find_firstEwm print_digits<StreamPrinter, long int> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ rename _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ print_digits<ResizePrinter, long int> <lambda(auto:2)> format do_printf_ints<BufferPrinter> print_digits<LimitedPrinter, long long unsigned int> _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ ferror vfwprintf move<int&> _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic _ZN3frg17basic_string_viewIwEC4EPKwm _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic print_int<StreamPrinter, long long unsigned int> unused _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ args _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN13ResizePrinter6appendEc _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic _ZNSt16is_constructibleIiJOiEE5valueE _ZN11PrintfAgentI13BufferPrinterEC4EPS0_PN3frg9va_structE _ZN3frg17basic_string_viewIwEC4Ev _ZN11PrintfAgentI13ResizePrinterEC4EPS0_PN3frg9va_structE _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE PrintfAgent<ResizePrinter> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic printf_size_mod second printf_format<PrintfAgent<BufferPrinter> > StreamPrinter _ZN3frg8optionalIiEC2EOi PrintfAgent<StreamPrinter> _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev SCANF_TYPE_SHORT _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN11PrintfAgentI13ResizePrinterEclEc gp_offset _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic print_digits<LimitedPrinter, unsigned int> _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE vprintf flockfile _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> _ZN11PrintfAgentI13BufferPrinterEclEPKcm perror do_printf_floats<StreamPrinter> consume print_int<LimitedPrinter, long unsigned int> position _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN14LimitedPrinter6appendEc _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN11PrintfAgentI13StreamPrinterEclEc _ZN3frg3minImEERKT_S3_S3_ _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE agent _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN13ResizePrinter6appendEPKcm overflow_arg_area _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev operator()<long unsigned int> fsetpos _ZN14LimitedPrinter6appendEPKc _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ <lambda(auto:3)> SCANF_TYPE_LL setbuf feof _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE print_int<BufferPrinter, long int> intmax_t LimitedPrinter expand __opts _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic olddirfd _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg8optionalIiEC2IRivEEOT_ swap<bool> va_struct _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic swap _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN13ResizePrinterC4Ev _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE fgets_unlocked num_consumed _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13ResizePrinterEclEPKcm default_size reg_save_area getdelim _ZN14LimitedPrinterC2EPcm _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE invert _ZN13StreamPrinter6appendEc _ZN11PrintfAgentI14LimitedPrinterEC4EPS0_PN3frg9va_structE _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ getchar_unlocked print_int<LimitedPrinter, unsigned int> old_path print_digits<BufferPrinter, unsigned int> _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic match_count ~<constructor> _ZNSt16is_constructibleIiJRiEE5valueE print_int<BufferPrinter, long long unsigned int> _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic __formatter _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev longlong_size _ZN14LimitedPrinterC4EPcm vsscanf do_printf_ints<ResizePrinter> ../options/ansi/generic/stdio-stubs.cpp fputc SCANF_TYPE_CHAR _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ fputs _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev getline _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN13BufferPrinter6appendEPKc print_int<ResizePrinter, long unsigned int> do_printf_ints<LimitedPrinter> _ZNK3frg17basic_string_viewIwEeqES1_ _ZN3frg17basic_string_viewIwE10sub_stringEmm print_int<LimitedPrinter, long long unsigned int> _ZNK3frg17basic_string_viewIwE4dataEv freopen print_digits<StreamPrinter, long long unsigned int> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ min<long unsigned int> _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE tmpnam _ZN13ResizePrinter6appendEPKc SCANF_TYPE_INTMAX scanset newdirfd look_ahead optional<int&> _ZSt4swapIbEvRT_S1_ tmpfile print_digits<StreamPrinter, unsigned int> auto:2 auto:3 _ZN13BufferPrinter6appendEc print_digits<ResizePrinter, unsigned int> SCANF_TYPE_L fread vwscanf auto:1 do_printf_chars<StreamPrinter> print_digits<LimitedPrinter, long unsigned int> _ZN13BufferPrinter6appendEPKcm _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE fpos_t _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ PrintfAgent<LimitedPrinter> fgetc_unlocked _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev basic_string_view<wchar_t> _ZN3frg17basic_string_viewIwEC4EPKw fputwc _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZSt18is_constructible_vIiJOiEE fputws _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic typed_dest store_int is_constructible<int, int&> is_constructible<int, int&&> PrintfAgent<BufferPrinter> _ZN13StreamPrinterC2EP17__mlibc_file_base _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ printf_format<PrintfAgent<ResizePrinter> > _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev vsprintf _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev ResizePrinter print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> _ZN13StreamPrinterC4EP17__mlibc_file_base fgets do_printf_floats<ResizePrinter> forward<int&> do_printf_chars<ResizePrinter> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ operator()<unsigned int> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ typedef __va_list_tag __va_list_tag fwrite getchar _ZN13ResizePrinterC2Ev wcsrchr strchrnul pattern wmemmove wmemcmp wcsncat bufsz wmemset wcstod wcscpy wcstof wcsncpy stpcpy wcstok wcstold wcstoull wcstol chrs wcstoll strerror ../options/ansi/generic/string-stubs.cpp delimiter wcspbrk wcschr mempcpy wcsncmp wcsstr b_byte strtok wcscspn wcscat wcslen s_bytes strchr strncat strcspn wcstoul wcscmp strncpy strerror_r strcoll strcpy a_byte strxfrm wmemchr strspn wcscoll found wcsspn strcat strcmp strstr wcsxfrm strrchr wmemcpy strncmp strpbrk _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEaSES6_ _Z19__mlibc_do_finalizev _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv forward<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> remove_reference<ExitHandler&> _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv move<ExitHandler&> _Z12getExitQueuev Align _ZSt4moveIR11ExitHandlerENSt16remove_referenceIT_E4typeEOS3_ aligned_storage ../options/lsb/generic/dso_exit.cpp _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4EOS6_ _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEEC4IJRS6_EEEDpOT_ eternal<frg::vector<ExitHandler, frg::slab_allocator<VirtualAllocator, AllocatorLock> > > _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm argument __cxa_atexit ExitHandler _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEEC2IJRS6_EEEDpOT_ _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED4Ev _ZN3frg15aligned_storageILm32ELm8EEC4Ev _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ dsoHandle _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backEOS1_ getExitQueue _ZN3frg15aligned_storageILm32ELm8EEC2Ev _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERKS6_ _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEE3getEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ERS5_ _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm __mlibc_do_finalize _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv remove_reference<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv aligned_storage<32, 8> _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5emptyEv vector<ExitHandler, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZSt7forwardIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE function _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv eternal<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERS5_ singleton _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backERKS1_ _ZN5mlibc14sys_libc_panicEv _ZN5mlibc8sys_exitEi sys_exit sys_anon_allocate _ZN5mlibc13sys_anon_freeEPvm sys_libc_panic _ZN5mlibc17sys_anon_allocateEmPPv ../sysdeps/lemon/generic/lemon.cpp sys_anon_free move<frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less&> _ZN3frg15aligned_storageILm456ELm8EEC2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ _ZN3frg15aligned_storageILm1ELm1EEC2Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE6bucketC2Ev _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ _ZN3frg7eternalI16VirtualAllocatorE3getEv eternal<> eternal<VirtualAllocator&> _Z12getAllocatorv _ZN3frg7eternalI16VirtualAllocatorEC4IJEEEDpOT_ _ZN3frg15aligned_storageILm456ELm8EEC4Ev _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ eternal<VirtualAllocator> eternal<frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev MemoryAllocator virtualAllocator getAllocator _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ forward<VirtualAllocator&> aligned_storage<456, 8> remove_reference<frg::slab_allocator<VirtualAllocator, AllocatorLock>::frame_less&> _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2ERS1_ _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE aligned_storage<1, 1> _ZN13AllocatorLockC2Ev _ZN3frg15aligned_storageILm1ELm1EEC4Ev _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ ../options/internal/generic/allocator.cpp remove_reference<VirtualAllocator&> _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4IJRS2_EEEDpOT_ global_wide_charcode code_seq<unsigned int const> _ZN5mlibc16current_charcodeEv _ZN5mlibc8code_seqIKwEcvbEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate promote_wtranscode has_shift_states_ _ZN5mlibc20polymorphic_charcodeC2Ebb platform_wide_charcode _ZN5mlibc20polymorphic_charcodeD4Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED4Ev preserves_7bit_units _ZN5mlibc20polymorphic_charcodeC4ERKS0_ decode_wtranscode utf8_charcode code_seq<char> _ZN5mlibc13utf8_charcode16has_shift_statesE _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4Ev decode_wtranscode_length _ZN5mlibc20polymorphic_charcode17decode_wtranscodeERNS_8code_seqIKcEERNS1_IwEER15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode6decodeERNS_8code_seqIKcEERNS1_IjEER15__mlibc_mbstate _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4ERKS2_ auto has_shift_states _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE encode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate decode polymorphic_charcode_adapter<mlibc::utf8_charcode> _ZN5mlibc13utf8_charcode20preserves_7bit_unitsE code_seq<wchar_t const> _ZN5mlibc8code_seqIcEcvbEv _ZN5mlibc13utf8_charcode12decode_stateC4Ev global_charcode _ZN5mlibc20polymorphic_charcodeD2Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE ../options/internal/generic/charcode.cpp decode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _vptr.polymorphic_charcode current_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN5mlibc20polymorphic_charcode24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode17encode_wtranscodeERNS_8code_seqIcEERNS1_IKwEER15__mlibc_mbstate ~polymorphic_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13utf8_charcode12decode_state6cpointEv encode_wtranscode _ZN5mlibc13utf8_charcode12decode_stateC2Ev _ZN5mlibc13utf8_charcode12decode_state8progressEv preserves_7bit_units_ __vtbl_ptr_type ~polymorphic_charcode_adapter _ZN5mlibc8code_seqIKjEcvbEv _ZN5mlibc22platform_wide_charcodeEv _ZN5mlibc20polymorphic_charcodeC4Ebb _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4EOS2_ _ZN5mlibc20polymorphic_charcodeD0Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev encode_state _ZN5mlibc20polymorphic_charcode18promote_wtranscodeEcRw decode_state _ZN5mlibc7charset8is_punctEj is_upper _ZN5mlibc15current_charsetEv _ZN5mlibc7charset8is_blankEj _ZN5mlibc7charset8is_printEj _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZN5mlibc7charset8is_alphaEj is_graph _ZN5mlibc7charset17is_ascii_supersetEv ../options/internal/generic/charset.cpp to_upper operator<< <unsigned int> current_charset _ZN5mlibc7charset8is_graphEj _ZN5mlibc7charset8is_upperEj _ZN5mlibc7charset8is_digitEj to_lower global_charset _ZN5mlibc7charset8is_spaceEj is_space _ZN5mlibc7charset8to_upperEj is_alpha is_digit _ZN5mlibc7charset8is_alnumEj is_alnum _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ is_blank _ZN5mlibc7charset8is_lowerEj is_punct _ZN5mlibc7charset9is_xdigitEj is_ascii_superset _ZN5mlibc7charset8to_lowerEj is_lower is_print is_xdigit _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEC4ES2_ PanicSink _ZN5mlibc9PanicSinkC4Ev _ZN5mlibc9PanicSinkclEPKc ../options/internal/generic/debug.cpp format_object<frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc format<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> format_integer<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ format<char const*, frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemaSERKS4_ print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4ERKS4_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD4Ev _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ ../options/internal/generic/ensure.cpp _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4EPS3_ __ensure_warn _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ assertion _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ __ensure_fail _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ Guard _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic __mlibc_int64 ../options/internal/gcc/guard-abi.cpp _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ complete _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ __cxa_guard_acquire __cxa_guard_release format<void*, frg::stack_buffer_logger<mlibc::PanicSink>::item> format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> __cxa_pure_virtual _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE4backEv default_list_hook _ZN5mlibc13abstract_file7io_readEPcmPm _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ owner intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*> fclose _init_bufmode _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC4Ev _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> pipe_like erased construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > stdout_file _ZN5mlibc13abstract_file6_resetEv forward<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > __for_range rewind _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ ~fd_file fileno _write_back destruct<mlibc::abstract_file, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN5mlibc7fd_fileD2Ev _ZN5mlibc13abstract_file14determine_typeEPNS_11stream_typeE composition<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8pop_backEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN5mlibc13abstract_file8io_writeEPKcmPm io_size _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE _vptr.abstract_file _ZN5mlibc13abstract_file10_init_typeEv _init_type _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ fileno_unlocked unknown _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN5mlibc13abstract_file13_init_bufmodeEv abstract _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5emptyEv OwnerPointer _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE _void_impl intrusive_traits<mlibc::abstract_file, mlibc::abstract_file*, mlibc::abstract_file*> borrow _ZN5mlibc13abstract_fileC4EPFvPS0_E __closure stream_type _ZN5mlibc13abstract_file7disposeEv fdopen _ZN5mlibc13abstract_fileD4Ev file_like iterator seek_offset _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv _ZN5mlibc7fd_fileC4EiPFvPNS_13abstract_fileEE _ZN5mlibc13abstract_file4seekEli setvbuf io_read owner_pointer _GLOBAL__sub_I_file_io.cpp _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ determine_bufmode _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ new_offset line_buffer _ZN5mlibc13abstract_file5closeEv intrusive_list Locate _ZN5mlibc13abstract_fileaSERKS0_ _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE10push_frontES6_ unget _ensure_allocation has_plus _ZN5mlibc13abstract_file5purgeEv _ZN5mlibc13abstract_file5ungetEc global_file_list _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _current _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6spliceENS9_8iteratorERS9_ _ZN5mlibc13abstract_file18_ensure_allocationEv io_write _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE _ZN5mlibc7fd_file2fdEv _ZN5mlibc13abstract_fileD0Ev _ZN5mlibc7fd_fileD4Ev update_bufmode borrow_pointer _ZN5mlibc13abstract_file7io_seekEliPl push_front BorrowPointer fseek ftell _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEi _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv _ZN5mlibc7fd_fileC4EOS0_ forward<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > __for_begin _ZN5mlibc13abstract_file11_write_backEv _ZN5mlibc7fd_file5closeEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev previous __fpurge _ZN5mlibc13abstract_file4readEPcmPm current_offset ~abstract_file globallyDisableBuffering _ZN5mlibc13abstract_file5flushEv _ZN5mlibc13abstract_fileC2EPFvPS0_E intrusive_list_hook stderr_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC4ES6_ _ZN5mlibc13abstract_file5writeEPKcmPm io_seek __for_end _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE full_buffer _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv _ZN5mlibc7fd_fileD0Ev <lambda(mlibc::abstract_file*)> remove_reference<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6insertENS9_8iteratorES6_ operator void (*)(mlibc::abstract_file*) move<mlibc::abstract_file*&> args#1 fopen _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ _result_of_impl splice determine_type locate_tag remove_reference<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > args#0 decay _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5frontEv pop_front _ZN5mlibc7fd_file7io_seekEliPl _ZN5mlibc13abstract_fileC4ERKS0_ remove_reference<mlibc::abstract_file*&> operator++ buffer_mode _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ _do_dispose _ZN5mlibc7fd_fileC4ERKS0_ pop_back _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC4Ev remove_reference<frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>&> intrusive_list<mlibc::abstract_file, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > ungetc erase no_buffer flush_line get<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > global_stdio_guard ../options/ansi/generic/file-io.cpp _ZN5mlibc7fd_file7io_readEPcmPm in_list ~stdio_guard _ZN5mlibc13abstract_file4tellEPl _ZN5mlibc13abstract_fileD2Ev stdin_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ _ZN5mlibc13abstract_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc7fd_file8io_writeEPKcmPm iterator_to _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE fflush _FUN fflush_unlocked _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9pop_frontEv sys_access sys_close sys_read _ZN5mlibc8sys_openEPKciPi sys_libc_log _ZN5mlibc12sys_libc_logEPKc _ZN5mlibc10sys_accessEPKci ../sysdeps/lemon/generic/filesystem.cpp sys_write sys_open sys_errno _ZN5mlibc9sys_writeEiPKvmPl _ZN5mlibc9sys_closeEi sys_seek _ZN5mlibc8sys_seekEiliPl _written _ZN5mlibc8sys_readEiPvmPl                 M@     Z@     Z@     �@     �@     �@     �@     @     @     @     @     8@     8@     e@     f@     �@     �@     V@     V@     �@     �@     @                     �E@     GF@     MF@     NF@                     �G@     �H@     �H@     �H@                     
J@     �J@     �J@     �J@                     O+@     r=@     r=@     �=@     �=@     ?>@     @>@     @@     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     2A@     hA@     hA@     �A@     �A@     �A@     �A@     B@     B@     $B@     $B@     �B@     �B@     �C@     �C@     �C@     �C@     �C@     �C@     6D@     6D@     �F@     �F@     �H@     �H@     �J@     �J@     K@     K@     !K@     "K@     KK@     LK@     xK@     xK@     �K@     �K@     
O@     
O@     �S@     �S@     �U@     �U@     V@     V@     V@     V@     V@      V@     TV@     TV@     �V@     �V@     �V@     �V@     W@     W@     8W@     8W@     _W@     `W@     (X@     (X@     �X@     �X@     3Y@     4Y@     JY@     JY@     �Y@     �Y@     �Z@     �Z@     D[@     D[@     �[@     �[@     �\@     �\@     �]@     �]@      ^@      ^@     �^@     �^@     �^@     �^@     c_@     d_@     u_@     u_@     �_@     �_@     �_@     �_@     b@     b@     1b@     2b@     �d@     �d@     �d@     �d@     :e@     :e@     be@     be@     �e@     �e@     �f@     �f@     �f@     �f@     h@     h@     oj@     oj@     �j@     �j@     m@     m@     ~m@     ~m@     �m@     �m@     o@      o@     Wp@     Xp@     �p@     �p@     uq@     uq@     r@     r@     *r@     *r@     Hr@     Hr@     yr@     zr@     =x@     =x@     Zx@     Zx@     �x@     �x@     �x@     �x@     �x@     �x@     8|@     8|@     N|@     N|@     �|@     �|@     �|@     �|@     �|@     �|@     ��@     ��@     Ƃ@     Ƃ@     �@     �@     s�@     s�@     ��@     ��@     D�@     D�@     �@     �@     �@     �@     �@     �@     ��@     ��@     B�@     B�@     s�@     s�@     �@     �@     C�@     D�@     ��@                     ��@     �@     "@@     ~@@     A@     1A@     �@     �@     �@     @�@     �C@     �C@     �C@     �C@     @�@     ��@     ��@     �@     �J@     K@     K@     !K@     "K@     KK@     LK@     xK@     V@     V@     V@     V@      V@     TV@     TV@     �V@     �V@     �V@     �^@     �^@     �p@     uq@                     �@     M�@     hA@     �A@     �A@     �A@     �A@     B@     B@     $B@     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     2A@     hA@     N�@     x�@     $B@     �B@     �B@     �C@     �C@     �C@     �C@     �C@     �C@     6D@     @�@     ��@     x�@     ˨@     �J@     K@     K@     !K@     "K@     KK@     ̨@     ݨ@     ި@     �@     �@     &�@     LK@     xK@     &�@     ��@     ��@     �@     ��@     ֩@     ֩@     �@     �@     .�@     .�@     b�@     b�@     ٪@     ڪ@     _�@     `�@     ��@     ��@     ��@     ��@     ��@     ��@     ˫@     ˫@     �@     �@     c�@     V@     V@     V@     V@      V@     TV@     TV@     �V@     c�@     ��@     �V@     �V@     ��@     ֬@     �K@     
O@     ֬@     ٭@     �^@     �^@     ٭@     ߯@     W@     8W@     8W@     _W@     `W@     (X@     (X@     �X@     �X@     3Y@     4Y@     JY@     JY@     �Y@     �Y@     �Z@     
O@     �S@     �p@     uq@     D�@     ��@     ߯@     -�@     d_@     u_@     �]@      ^@     u_@     �_@     �_@     �_@     �_@     b@     b@     1b@     2b@     �d@     �d@     �d@     �d@     :e@     :e@     be@     be@     �e@     �e@     �f@     �f@     �f@     �f@     h@     �Z@     D[@     D[@     �[@     �[@     �\@     �\@     �]@      ^@     �^@     -�@     w�@     r@     *r@     *r@     Hr@     Hr@     yr@     zr@     =x@     =x@     Zx@     Zx@     �x@     �x@     �x@     �x@     �x@     �x@     8|@     8|@     N|@     oj@     �j@     N|@     �|@     �|@     �|@     h@     oj@     �j@     m@     m@     ~m@     ~m@     �m@     �m@     o@      o@     Wp@     Xp@     �p@     w�@     �@     s�@     ��@     ��@     D�@     D�@     �@     �@     �@     �@     �@     ��@     Ƃ@     �|@     �|@     �@     ��@     ��@     B�@     �|@     ��@     Ƃ@     �@     �@     h�@     B�@     s�@     h�@     �@     �@     C�@                     ��@     5�@     :�@     ;�@                     v�@      �@     %�@     &�@                     ��@     p�@     u�@     v�@                     ��@     [�@     `�@     a�@                     ��@     ��@     b�@     e�@                     |�@     ��@     B�@     E�@                     ��@     0�@     E�@     H�@                     0�@     z�@     H�@     K�@                     z�@     3�@     K�@     N�@                     3�@     ��@     N�@     Q�@                     ��@     ��@     Q�@     R�@                     �@     B�@     e�@     f�@                     P�@     ��@     !�@     $�@                     ;�@     ]�@     �@     �@                     ]�@     ��@     �@     �@                     ��@     9�@     �@     
�@                     9�@     ��@     
�@     �@                     ��@     ��@     �@     �@                     ��@     ��@     �@     �@                     ��@     �@     $�@     %�@                     �0A     Q1A     V1A     �1A                     �1A     U2A     Z2A     �2A                     �2A     Y3A     ^3A     �3A                     �DA     EA     "EA     }EA                     �EA     !FA     &FA     �FA                     �FA     %GA     *GA     eGA                     )XA     �XA     �XA     YA                     $YA     �YA     �YA     #ZA                     (ZA     �ZA     �ZA     [A                     �kA     alA     flA     �lA                     �lA     emA     jmA     �mA                     �mA     inA     nnA     �nA                     �@     7�@     hA@     �A@     �A@     �A@     �A@     B@     B@     $B@     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     2A@     hA@     N�@     x�@     8�@     ^�@     ^�@     ��@     ��@     �@     �@     Y�@     Z�@     ��@     ��@     ��@     ��@     #�@     $�@     ��@     ��@     ��@     ��@     �@     �@     c�@     d�@     ��@     ��@     ��@     ��@     ��@     ��@     8�@     8�@     ��@     ��@     ��@     $B@     �B@     �B@     �C@     �C@     �C@     �C@     �C@     ��@     ��@     �C@     6D@     �U@     V@     ��@     �@     �@     ��@     ��@     �@     �@     �A     �A     A     A     0A     0A     �A     
O@     �S@     �J@     K@     K@     !K@     "K@     KK@     �@     &�@     LK@     xK@     �A     &	A     &	A     �A     V@     V@     V@     V@     �A     A     A     3A     4A     ]A     ^A     �A     �A     �A     �A     $A     $A     �A     �A     -A     .A     WA     XA     /A     0A     aA     bA     �A     �A     cA     W@     8W@     8W@     _W@     JY@     �Y@     �Z@     D[@     D[@     �[@     �X@     3Y@     �[@     �\@     �\@     �]@     �]@      ^@     �Y@     �Z@      ^@     �^@      V@     TV@     TV@     �V@     c�@     ��@     �V@     �V@     dA     �A     �A     �A     �A     �!A     �!A     �"A     �"A     �"A     �"A     �"A     �"A     U)A     V)A     /*A     0*A     +A     +A     �+A     �+A     �,A     �,A     �-A     �-A     f.A     f.A     6A     6A     6A     �6A     �6A     �6A     "=A     "=A     �=A     �=A     �>A     �>A     �?A     �?A     �@A     �@A     [AA     \AA     2BA     2BA     �IA     �IA     KJA     KJA     �PA     �PA     �QA     �QA     tRA     tRA     MSA     NSA     $TA     $TA     �TA     �TA     �UA     �UA     �]A     �]A     �]A     d_@     u_@     be@     �e@     �f@     �f@     h@     oj@     oj@     �j@     �j@     m@     �d@     �d@     m@     ~m@     4Y@     JY@     ~m@     �m@     :e@     be@     u_@     �_@     �m@     o@     �_@     �_@      o@     Wp@     �d@     :e@     �e@     �f@     �f@     h@     Xp@     �p@     �^@     �^@     ٭@     ߯@     �]A     edA     fdA     ?eA     @eA     fA     fA     �fA     �fA     �gA     �gA     �hA     �hA     viA     viA     +qA     +qA     �qA     �qA     �qA     �qA     �qA     �qA     4rA     4rA     �rA     @�@     ��@     ި@     �@     �rA     �rA     �rA     �rA     �rA     �sA     �sA     �sA     �sA     CtA     CtA     �tA     �tA     �tA     �tA     �uA     �uA     �uA     �uA     ,vA     ,vA     �vA     �vA     "wA     "wA     wwA     wwA     �wA     8|@     N|@     �|@     �|@     �|@     �|@     �|@     ��@     ��@     Ƃ@     N|@     �|@     �x@     �x@     �x@     �x@     Ƃ@     �@     r@     *r@     b@     1b@     Zx@     �x@     *r@     Hr@     �x@     8|@     �p@     uq@     D�@     ��@     ߯@     -�@     �wA     %xA     %xA     �xA     �xA     yA     yA     pyA     pyA     {A     {A     �|A     �|A     _~A     _~A     �A     �A     Q�A     Q�A     ��A     ��A     ��A     ��A     @�A     @�A     �A     �A     ��A     ��A     8�A     8�A     ׋A     ׋A     �A     B�@     s�@     �@     ��@     ��@     B�@     �@     �@     �@     �@     =x@     Zx@     Hr@     yr@     ��@     D�@     D�@     �@     -�@     w�@     �A     '�A     '�A     ϐA     ϐA     n�A     n�A     �A     �@     C�@     �A     ��A     w�@     �@     ��A     J�A     �@     h�@     h�@     �@     J�A     ޖA                     ��A     ��A     hA@     �A@     �A@     �A@     �A@     B@     B@     $B@     @@     !@@     $B@     �B@     �B@     �C@     ��A     ��A     ��A     �A     �A     ��A     ��A     ��A     ��A     ��A     ��A     ʧA     ʧA     ��A     ��A     6�A     6�A     J�A     
O@     �S@     J�A     z�A     �K@     
O@     W@     8W@     8W@     _W@     JY@     �Y@     �Z@     D[@     D[@     �[@     �X@     3Y@     �[@     �\@     �\@     �]@     �]@      ^@     �Y@     �Z@      ^@     �^@     `W@     (X@     (X@     �X@     4Y@     JY@     d_@     u_@     be@     �e@     �f@     �f@     h@     oj@     oj@     �j@     �j@     m@     �d@     �d@     m@     ~m@     ~m@     �m@     :e@     be@     u_@     �_@     �m@     o@     �_@     �_@      o@     Wp@     �d@     :e@     �e@     �f@     �f@     h@     Xp@     �p@     �_@     b@     b@     1b@     2b@     �d@     8|@     N|@     �|@     �|@     �|@     �|@     �|@     ��@     ��@     Ƃ@     N|@     �|@     �x@     �x@     �x@     �x@     Ƃ@     �@     r@     *r@     Zx@     �x@     *r@     Hr@     �x@     8|@     Hr@     yr@     zr@     =x@     =x@     Zx@     B�@     s�@     �@     ��@     ��@     B�@     �@     �@     �@     �@     ��@     D�@     D�@     �@     s�@     ��@                     Z�A     ��A     @@     !@@     ��A     ��A     ��A     ܫA     ܫA     �A     �A     ��A     ��A     H�A     H�A     V�A     V�A     h�A     h�A     ��A     ��A     	�A     
�A     .�A     .�A     e�A     e�A     o�A     p�A     ��A     ��A     ��A     ��A     ��A                     �A     B�A     ��A     ��A                     ��A     ��A     ��A     ٮA     ڮA     ��A     ��A     
�A     
�A     �A     �A     ��A     ��A     "�A     "�A     Y�A     Z�A     ��A     ��A     ��A     ��A     ��A      �A     G�A     H�A     \�A     \�A     ��A     ��A     ӶA     ԶA     �A     ��A     �A     �A     3�A     4�A     S�A                     T�A     ��A     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     �C@     �C@     �C@     �C@     �C@     6D@     �J@     K@     K@     !K@     "K@     KK@     LK@     xK@     ��A     ��A     V@     V@     V@     V@      V@     TV@     TV@     �V@     �V@     �V@     ��A     3�A     �^@     �^@     -�@     w�@     �p@     uq@     w�@     �@     �@     h�@     h�@     �@     �@     C�@     D�@     ��@                     u�A     ��A     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     �C@     �C@     �C@     �C@     �C@     6D@     ��A     ��A     ��A     ��A     ��A     ��A     ��A     �A     �A     B�A     �J@     K@     K@     !K@     "K@     KK@     ��A     ��A     LK@     xK@     V@     V@     V@     V@     B�A     v�A     v�A     ��A     ��A     ��A     ��A     $�A      V@     TV@     TV@     �V@     ��A     3�A     �V@     �V@     $�A     N�A     N�A     ��A     �^@     �^@     -�@     w�@     ��A     i�A     i�A     �A     �p@     uq@     w�@     �@     �A     Z�A     �@     h�@     Z�A     ��A     h�@     �@     �@     C�@     ��A     ��A     D�@     ��@                     ��A     ��A     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     2A@     hA@     �C@     �C@     �C@     �C@     �C@     6D@     ��A     ��A     ��A     ��A     ��A     ��A     ��A     �A     �A     B�A     V@     V@     V@     V@     B�A     v�A     v�A     ��A     �A     ^�A     ��A     $�A     $�A     N�A     ^�A     ��A     ��A     i�A     ��A     z�A     z�A     ��A     ��A     y�A     �@     C�@     ��A     ��A                     z�A     ��A     @@     !@@     "@@     ~@@     ~@@     A@     A@     1A@     hA@     �A@     �A@     �A@     �A@     B@     B@     $B@     $B@     �B@     �B@     �C@     �C@     �C@     �C@     �C@     �C@     6D@     ��A     ��A     ��A     �A     �A     ��A     �J@     K@     K@     !K@     "K@     KK@     LK@     xK@     �K@     
O@     ��A     �A     �A     ��A     ��A     ��A     ��A     ��A     ��A     ��A     �A     B�A     �A     A     �U@     V@     
O@     �S@     ��A     %�A     &�A     I�A     J�A     r�A     r�A     ��A     ��A     ��A     �6A     �6A     ��A     ��A     �"A     �"A     V@     V@     V@     V@     ��A     
�A     
�A     :�A     :�A     K�A     L�A     f�A      V@     TV@     TV@     �V@     �V@     �V@     W@     8W@     8W@     _W@     `W@     (X@     (X@     �X@     �X@     3Y@     4Y@     JY@     JY@     �Y@     �Y@     �Z@     B�A     v�A     v�A     ��A     ��A     $�A     �Z@     D[@     D[@     �[@     �[@     �\@     �\@     �]@     �]@      ^@      ^@     �^@     f�A     ��A     ��A     ��A     CtA     �tA     ��A     ��A     ��A     �A     �A     (�A     �^@     �^@     d_@     u_@     u_@     �_@     �_@     �_@     �_@     b@     b@     1b@     2b@     �d@     �d@     �d@     �d@     :e@     :e@     be@     be@     �e@     �e@     �f@     �f@     �f@     �f@     h@     $�A     N�A     h@     oj@     oj@     �j@     �j@     m@     m@     ~m@     ~m@     �m@     �m@     o@      o@     Wp@     Xp@     �p@     �A     Q�A     (�A     6�A     �p@     uq@     r@     *r@     *r@     Hr@     Hr@     yr@     zr@     =x@     =x@     Zx@     Zx@     �x@     �x@     �x@     �x@     �x@     �x@     8|@     8|@     N|@     N|@     �|@     �|@     �|@     ��A     i�A     �|@     �|@     �|@     ��@     ��@     Ƃ@     Ƃ@     �@     �A     ��A     s�@     ��@     ��@     D�@     D�@     �@     �@     �@     �@     �@     �@     ��@     ��@     B�@     B�@     s�@     ��A     J�A     h�@     �@     J�A     ޖA     �@     C�@     D�@     ��@     6�A     c�A     d�A     ��A                                                          � @                    @                   q�A                   ��A                   șB                     C                     C                    C                  	 ( C                  
 8 C                   `C                   �C                                                                                                                                                                                                                                             ��                      C                 	 ( C             (     șB             ;      @             =     P@             P     �@             f     �C            u     �C            �      @             �     �C     0           ��                �       C             �     ��B             �     0�A             �    ��                �    ��                     @                ��                #    @     >       S    E@            l   ��                x   ��                �     M"@             �     q"@             �     �"@             �     �"@             �     #@             �     #@             �     #@               ��                   ��                   ��                &   ��                ,   ��                6   ��                ;   ��                B   ��                P   ��                a    ��A            t    ��A            �    ��A            �    ��A            �    ��A            �    �B                               :    B            O    B            d    B            x     B            �    0B            �    ;B            �    BB            �    PB            �    XB                \B                aB            (    gB            ;    lB            O    rB            c    xB            x    B            �    �B     	       �    �B     	       �    �B            �    �B     	       �    �B                �B            B     B            #    .=@     /       k    ]=@            �   ��                a    @B            t    AB            �    �B            �    �B     	       �    �B     	            �B     	          ��                �    �B            �    �B            �    �B            �    g*B            a    =B            t    >B            '     C            M    �@     �      �     C             �    @C            �    ��@     o           '�@     �       '    ��@     ?      k    p*B            �    3�@     r      �    �*B            I    �*B            ^    �*B            s    �*B            �   ��                �   ��                �    �*B            �    �*B            �    �*B            �     TB            a    +B            t    +B            �    CTB            �    �RB            �    �RB            �    �RB     	       	    �RB            &	    �RB            ;	    �RB            Q	    �RB            f	    Զ@     �       x	    �RB            �	    b�@            �	    v�@     0       �	    ��@     �      �	    ��@     b       
    ^�@     [       /
    x�@     �      a
    �RB            v
    SB            �
     SB     	       �
    0SB            �
    8SB     
       �
    HSB     	       �
    XSB     	       �
    hSB                pSB     
       -    �SB     	       D    �SB            Z    �SB            o    �SB     	       �    �SB            �    �SB            �    �SB            �    �SB            �    �SB            �    �SB                �SB                �SB            ,    �SB     	       C    �SB            W    �SB     	       n    TB            �    TB            �    TB            �    (TB     	       �    PTB            �    �RB            B    �RB            �    SB            �    8TB            Z   ��                k    H]B            �    P]B            �    W]B            �    ^]B            �    h]B            �    p]B            �    x]B                �]B                �]B     	       .    �]B            C    �]B            Y    �]B            o    �]B     	       �    �]B            �    �]B            �    �]B            �    �]B            �    �]B            �    �]B                �]B                �]B            3    �]B            I    �]B            _     ^B            u    ^B            �    ^B            �    ^B            �    ^B            �    (^B            �   ��                �    0^B            �    1^B            �    2^B            �    OoB            �    `C             
    �C            *   ��                4    �oB            a   ��                �    �oB            �    �oB            �    �oB            o    �C            �    �C            �    �C     �      �    �C            �    GpB            "    KpB            L   ��                a    `pB            t    apB            Y    �qB            �    �qB            �    �C            !    �C            T    �C            �    �qB                �qB            �    �qB                pqB            �   ��                a    �qB            t    �qB            �    �C            �   ��                a    jwB            t    kwB            �   ��                a    pwB            t    qwB            �   ��                a    �yB            t    �yB                �yB            &    ��A     J       E    ��A            f   ��                a    |B            t    |B            �    |B            �    |B            �    |B            �    "�B            r    m|B            �    �C            �    '�B                 ,�B            1    2�B            ]    8�B            �    G�B            �    P�B                `�B            6    p�B            i    |�B            �    ��B            �    ��B                �C     x       2    `C     x       R    �C     x       r    �A            �    �A            �    �A     �       �    �A     �       �    XC            %    V�A     *       T    ��A            �    ��A            �    ��A     �       G    �A     *       w    ,�A            �    L�A            �    ;�A     �       m    ��A            �    -�A            #    ��A     �           ��A            7   ��                F    �@     #       O  "  -�@     J       �  "  �PA     �       6    H�A     H       =    �@            E  "  oj@            7  "  �6A     x      �  "  A     *       �    �A     �       �    ޖA     S       �     @                "  ��A            �     �@     o      (!  "  "@@     \       D!  "  .�A     7       �!  "  �?A     �       	"  "  �x@            �"    �A     n       #    �@     >       #  "  �C@     V       :#  "  �IA     d       �#    ȹA     �       �#  "  r�A     2       Y$  "  �UA     �      �$  "  ��A     �       %  "  B�A     4       J%  "  �A     N       i%  "  �A     U       �%  "  ��@     >        &  "  K@            _&    �@     #       g&    �C            p&    d�A     �       �&  "  �A     )       �&  "  ��A     >       '    H�@     /       
'  "  Z�@     &       "'  "  ��A     P       �'  ! 
 x C     @       �'    ~�A     3       �'    @ @     (       �'    @C     (       ��    �@     �       (    �C            	(    Y�@     �       (  "  �C@     #       *(    �A     /       1(  "  �x@     V      ")  "  �gA     �       �)  "  @�@     R       �)    ]�@     7       �)    ��A     �      �)  "  ��@            $*  "  B�A     4       ��    x�@     I       g*  "  ��A     "       �*  "  0A     1       +  "  ��A            :+  "  
O@     �      �+    $�A     B       �+  "  u_@            k,  "  ��A     P       �,  "  x�@     S       -  "  �Y@     �       �-    t�A     @      �-    ��A     A       �-  "  �^@     *       M.  "  A     1       v.  "  b@            ^/  "  uq@     �       �/  "  Xp@     K       00  "  �,A     �       �0  "  8�@     &       �0  "  �@            O1  "  �>A     �       ��    j*@     �       �1  "  D�@     �      �2    h�A     T       �2  "  ��A     <      <3  "  �tA     �       M    ��@     �       z3    �'@     >       �3  "  ��A     =       �3  "  NSA     �       %4   ��A     E       ?4  "  ٭@           �4    o(@     �       �4    �A     4       �4    �C            �4  "  f.A     �      D5  "  CtA     G       �5  "  �U@     +       �5    �A     2       �5  "  6�A     -       �5    �+@     $       �5    ��A            �5  "  b�@     w       G6    �C            ^6    l'@     8       m6  "  �J@     )       �    �@            �6  "  ��@            �6    p�A            7  "  V)A     �       �7  "  Xp@     K       �7  "  V@            8    ��@     �        8  "  p�A            �8  "  �K@     h      =9    �A     +       D9    ϗ@     H       M9  "  ��@     <       i9  "  ��A     P       �9    ��@     S       �9  "  �!@            �9    m&@     ?       �9    @,@     9       �9    ��@     V       6�    5@     +       �9    ��A     2       �9    >�@     S       �9    0�@     S       :    �2@     �       :    `@     o      ::  "  �\@     �       �:  "  ~@@     �       ;  "  wwA     W       A;  "  d_@            "<  "  xK@     )       j<  "  �uA     U       �<    �@     3       �<  "  ��A     )       �<  "  _~A     �      <=  "  6D@     M      Z=    �3@           `=  "  ڮA             �=  "  8|@            r>    �A     .       z>  "  ��A     )       �    i�@     �       �>    ]�@     �       �>  "  $�A     *       6?    ��@     /       ??     @     �      R?    �@     S       \?  "  $TA     �       �?  "  \AA     �       Y@  "  "=A     �       �@  "  �A     N       �@    �A     �        A  "  �A     �      T�    .�@            bA    N�A     �       A  "  ��A     +       �A  "  �fA     �       >B  "  �xA     U       {B  "  �f@            jC  "  f@     "       X    *@     Z       �C    T�A     !       �C  "  Z@     I       �C    ��A           �C   �C             �C  ! 
 8 C     @       D  "  &�A     #       �D    ͳ@     5       �D    ��@     �       �D    �'@     M       �D  "  �A@            �D  "  ��A            E  	 0 C             #E    T�A            JE  "  �wA     W       �E  "  LK@     ,       �E  "  �V@     &       F  "  f�A     "       �    �@     �       �F  "  �rA     Y       �F    pC            �F    �%@     :       �F   3�A     N       G    ��@     V       
G    ��A            .G    f�A     5       7G    �@     Q       ?G  "  �_@     a      /H    ޭA     +       SH  "  L�A            �H  "  XA     �      @I    )�@     S       II  "  %xA     �       �I    �2@     +       �I  "  ��A            &J    ��@            +J    &�@     2       2J    áA     /       :J  "  �F@     L      XJ    }�A     2       _J    N�A     �       |J  "  8�A     �      �J  "  +qA     d       'K    �:@     �       .K    �@     +       �|    r2@     *       5K    ��@     S       >K  "  &	A     �      �K  "  ��A            �K  "  �@     �      �L  !   B             �L  "  n�A     �      M    w�@     �       'M    �-@     +       /M    \�A     u       ^M  "  ��A     *       �M  "  �QA     �       N  "  ��@     O       >N    �A            UN    ͠A     3       ]N  "  �6A     *       �N  "  m@     d       �N    �-@     G      �N   `C             O    �(@     �       O  "  ��@            $O  "  Z�A     -       eO    O�A     /       ~�    C�@     x       lO  "  J�A     (       	P  "  4�A            %P  "  Z�@     &       =P  "  �"A     x      �P    �2@     +       �P    ��A     ?       �P    O�@     V       �P  "  �A     1       �P  "  ��A     *       CQ                  QQ  "  ��A     =       vQ    8@     .       }Q   #�A            �Q  "  ^�@     H       �Q    �C            �Q    �9@     3       �Q  "  :e@     (       2R  "  f@     "       OR  "  �C@     V       kR  "  ��A            �R  "  �d@     j       �S  "  h�@     �      T  "  �@     �       )T  "  �A     �      �T    ��@            �T    Q�@     V       �T    ��@     /       �T    f�A     /       U  "  �@     W       sU    �A     7       {U    ��A            �U  "  :�A            �U  "  B@            �U  ! 
 � C     P       �U    /(@     @       V  "  (�A            �V  "  �@     S       �V  "  �@     �      W    0�A     �       0W  "  �X@     O       _W    L8@     =      hW    ��A            �W  "  �vA     �       �W    o�@     �       �W  "  ֩@     F       X    ��A     3       &X  "  �A     �      xX  "   "@            X  "  �@     M       �X  "  ��A     �       Y    ��@     7       #Y    ]2@            )Y  "  �A     �      �Y    ��A     m       �Y    lC            �Y  "  �@            9Z    �C            IZ    �1@     #       OZ  "  @     "       hZ  "  ^A     N       V     C            �Z  "  v�A     E       �Z    ��A     /       �Z  "  4Y@            '[  "   o@     7      \    4�@     [        \    ��@     V       )\    � @             /\  "  ��@     >       �\    Z�A     �       �\    y,@     J      �\  "  �rA     �       �\  "  ��A     "       e]    J�@     /       m]     C     �	      �]    �A     /       �]    �5@           �]    ֖@     S       �]  "  �p@     �       �]    ��A     �       b    �C            �]  "  0*A     �       |^    xC            �^    C            �^  "  A     *       �^  "  6A     d       ._  "  ��A     {       p_  "  �A            �_    3�@     �       �_  "  �@     2       �_     @     k       �_  "  ̨@            `  "  ��A     �      U`    @           q`  "  "�A     7       �`  "  �|A     �      �`    ՛A     p       �`  "  H�A            Ka    E�A     /       Ra  "  �Z@     �       >b    v1@     V       Eb    d"@             [b    �C            eb    hC            ob    �+@     3       vb  "  h�A     %       �b  "  @>@     �      �b  "  2b@     �      �c  "  �qA     J       �c  "  dA     1       �c  "  r=@             �c    ��A     f       �c  "  N|@     H       �d    O+@     -       �d  "  �x@            �e    �C            �e  "  be@            ��    ��@     �       �f    ��@     P       �f    ݕ@     S       �f  "  $�@     c       g  "  ��@     *       9g    ��A     Q       Ug    `@     k       og  "  L�A            	h    ��A     ;       h    ��A           {�    1�@     .       h  "  ��@     .       5h    �A     �       Rh  "  ��A     �       �h    z0@     +       �h  "  ��A     )       �h    �@     /       �h    �C     (       �h  "  �A            i  "  fA     �       �i   D�A            �i  "  '�A     �      �i  "  �A     �      �)    m�@     x       'j  "  ��@     L       Cj    *�A     �       ]j    �"@             kj  "  �A     �      �j  "  ��@     *       �j    {�A     r       �j  "  ^A     N       k  "  ��A     K      �k  "  ֩@     F       �k  "  ��A     ,       l  "  �j@     �      �l  "  �"A            2m  "  V@            Ym    �&@     ?       em    ��@     6       nm     �A     U       �m    ��A           �m  ! 
 C     P       �m    N�A     /       �c    8�A     Y       �m    0#@     R      �m  "  ��A            .n  "  .�A     7       tn    �C            zn  "  ��@     g       �n  "  �@     2       �n  "  zr@     �      �o    4�A            �o  "  ��A     �      �o    >�A     �       p  "  
�A     $       �p    �C            �p  "  ԶA            u�     @            �p    ��A            q  "  ܫA            0q    ��@            7q    ��A     �       >q  "  �A            �q  "  ��A     �      ��    `0@            r   �A     f       %r  "  *r@            
s  "  6�A           ss  "  ߯@     N       �s  "  ֬@           8t  "  ��@     *       rt  "  �tA     W       �t  "  J�A     �      u    ��@     .       #u  "  s�@     �      �u    Y�A     %       �u    ��A     h       �u    S�@     V       �u  "  �A     *       v  "  �|@     �      �v    ~�A     �       w  "  V@     �       #w  "   ^@     �       rw  "  �H@           �w    B�A     2       �w  "  m@     d       �w  "  "@            �w    �@     �       x    1�A     �       #    �@     �      x  "  V�A            7x    PC            Ux  "  �sA     W       �x    ��A     E       �x  "  4rA     W       �x  "  �rA     Y       y    ��@     [       y  "  8�@     S       <y  "  �A     *       vy    ��@     J       ~y  "  �!A     �       �y    \;@     �       �y  "  W@     2       �y    �C            �y    ڜ@     *       �y  "  6�A     -        z  "  �sA     U       =z    ��A     �       Zz    �A     J       gz  "  ި@            �z    �@             �z  "  fdA     �       /{  "  �|@            |  "  ��@     e       <|  "  �@            �|    e�A     /       �|    2@     +       �    u�A     r       �|  "  �C@            �|    kC            �|  "  {A     �      &}    ]�A     �       -}  "  r=@             �<    ��@     �       A}    @     I      d}    0@     �       �}    ��@     V       �}  "  ڮA             �}    ��A     /       �}  "  �[@     D      	~    �A     2       ~  "  r@            �~    �A     �       �~  "  ��A     0       �  "  �e@     7      ��    f�A     .       ��  "  ��A     3       �  "  N�@     *       :�    �%@     m       Y�  "  �@     -       r�    ��@     2       x�  "  �A     +       ��  "  �C@            ��  "  �@     �      ��  "  $A     �      I�    ��A     E       w�  "  Ƃ@     V      }�    ��@     x       ^�  "  �A     �      ��    �C            ��  "  �A     E       �    50@     +       �  "  N�A     J       {�  "  ^�A     }       �  "  2BA     �      P�  "  ��@     6       j�    ��A     Q      p�    �C             |�    <�A     3       ��    �@            ��  "  `�@     !       ��    _�@     *       �w    �)@     F       �  "  �uA     W       ?�  "  �f@     7      5�    �
@     A
      :�     �A     /       A�  "  ��@     *       |�    ��A     i       ��    ֿA     �       ��    �0@     "       ��    �A     3       ��  "  ��A            ɇ    �@     3       Ӈ    �C            ��    @            �  "  �A@     B       u    �@     �      �    y�@            �  "  ʧA     .       5�  "  ��A     *       ��    v�A     U       ��  "   "@            ��  "  @@            ��  "  V�A            �    ��A     �       �  "  �A     �       h�    `�@            p�  "  
�A     0       �  "  ��A     $       ��  "  ��@            ��  "  .�@     4       ��    �C            �    ��@     V       �    t�A     3       �  "  ��A     ,       G�    �@     /       O�    ��@     V       W�  "  �C@     #       o�  "  �B@     �       ��    %�@     +       ʇ    �@     x       Ì    ��@     V       ˌ  "  �@     8       �  "  �@     8       ��  "  h@     a      I�    ��@     "       ��    	�A     g       �  "  �rA            ;�  "  A@            W�    �@     ;      f�  "  ��A     &       ��  "  ��A     �       �    �A     r       �  "  &�@     r       ;�  "  �-A     �       ��    �A     �       ׏  "  V@            ��  "  ��A     |       C�  "  ��@     Q       `�    �"@             n�  "  "wA     U       ��    q�A             ��  "  ׋A     �      �  "  ��A            
�  "  �V@     E       ^�  "  ʧA     .       ��  "  KJA     x      �  "  ��A     �       S�    �@     D       ��    ��@     �       ��    /�@     �       Y�    ��A     ]       d�  "  �S@     #      ��    ��A     �      Ӓ    ,@     %       ڒ    �<@     3       `z    �1@     )       �   ��A     .       ��    ��A     m       ��  "  @�@     R       #�  "  ��A     C       w�  "  ��A     a       �  "  Hr@     1       ��  "  ��@     	      �  "  �@     U       u�    ~�@     [       �  "  �A            ��  "  4Y@            ?�    ��@     S       H�  "  @            k�  "  �_@            P�  "  `W@     �       ��  "  bA     )       �    ~�@     x       ��    �C            Ǘ  "  0A     �      �  "  �=A     �       ��    M@     �       ��  "  $B@            ��    �C            �  "  
�A     $       ��    �0@     Z       ��  "  ��A     C       �  "  "�A     7       L�    H�A     R       k�  "   V@     4       ��  "  ��A            �  "  �A            K�  "  pyA     �      ��  "  d�@     O       ��  "  +A     �       +�  "  �d@            �    ��@     $       H�    �5@     /       '�  "  �]A     d       v�    ��@     +       ��  "  �hA     �       �  "  hA@     Q       1�  "  ��@     .       H�    }�@     "       N�  "  ��@     6       h�  "  D[@     X       P�  "  �!@            V�    ��@            d�  "  ��A     {       ��  "  ��@     %       ��    �@     3       �  "  @eA     �       ��    H�@            ��  "  .A     )       Ҡ    ��@     .       ؠ    |�@     S       �    u�A           �  "  e�A     
       d�  "  (X@     �       F�    ��A            g�    V�A     I       w�  "  ~@@     �       ��  "  c�@     I       ��  "  ϐA     �      ;�    ��@     /       B�  "  "@@     \       ^�  "  �]@     L       ��  "   �A     G      	�    L�@     ;      �    3�A     3       !�  "  4A     )       G�    �5@     /       M�  "  W@     2       z�    ��A     W       ��    ڟA     3       ��  "  �TA     �       �    z�A     �       7�    M�@     V       ?�   1�A            \�    ��@     2       c�    �C             j�  "  s�@     1       M�  "  w�@     �       Ȧ    1�A     a       �    `C             �  "  \�A     X      d�   ��A            z�  "  �@     -       ��    �C            ��  "  Q�A     �      �    ��@     `       ��  "  ��A     >       R�  "  2A@     6       ��    ��A     R       ��  "  hA@     Q       ��    P�@     3       Ũ  "  yA     W       �    ��@     D       �  "  A@            -�  "  ~m@     j       �    ��@     .       �    �&@     A       (�  "  i�A     �       ��  "  ��A            N�  "  �@A     �       �|    C2@            ͫ  "  �=@     �       �    ,�A     �       �    z�A     �       @�    ��A            d�  "  ��A     �      ��  "  �]A     x      �    ��@     *       �    ��A     �       5�    :5@     +       ;�  "  TV@     E       ��   ��A     R       ��    ��@     2       ��  "  �@           ߭    7�@     S       Y    �@     x       �    o�A     /       �  "  ��A     G       Y�  "  Z�A     -       ��  "  ��A     $       F�    |+@     $       K�  "  �A     )       q�    ��@     K       y�  "  �|@     1       d�    @     �      }�  "  8W@     '       ��    ��@            ��    :�A     +       ԰  "  �A     J       >�  "  tRA     �       ��    ;�A            ñ  "  �A     ,       �    ��@     2       �    :�@     �      &�    p @     �       J�  "  
�A            z�  "  "K@     )       ò  "  �qA            ��    �A     /       ��  "  h�A     %       $�  "  Zx@     H       �    E�A     m       �  "  Z�A     �      ��  "  D�@     �       Ŵ    +@     <       ̴  "   V@     4       �  "  ��A     (       U�  "  �+A     �       ӵ    HC            �  "  N�@     *       �    _�@     Q       ˇ    ��@     x       �    7&@     6       �  "  ��A            L�    �+@     $       R�    ��A           o�  "  �"A     ;       ��  "  ,vA     W       Ķ  "  ��@     �      ��  "  K@            ��  "  J�A     0       2�     �A     3       :�  "  ��A     P       ��  "  8@     -      I�    e5@     &       7�    �4@     *       ��  "  viA     �      �    ��A     i       "�   z�A     3       7�  "  ��A            �    ��@     %       !�  "  ˫@     O       6�   ��A     �       X�  "  �@     (       r�    �C            {�  "  �^@     }       �   ��A     R       �  "  JY@     I       N�  "  V@            u�    ��@     +       |�    :�@     3       ��  "  �qA     J       ��    ��@     �       ��    (C            ��    2�@     K       ��    ��A     \       û  "  8W@     '       �  "  ڪ@     �       A�  "  �@     I       ��  "  =x@            x�  "  z�A     W       ޽  "  ��@     *       �  "  0"@             �    ,'@     @       .�    p�A     �       K�    @"@             W�    J�A     �       t�  "  �m@     7      _�    !1@     U       m�  "  B�@     1       Z�   x�A     J       n�    2<@     �       }�  "  ��@            ��  "  d�A     +       ��    �C            ��  "  8�@     &       ��    ��A     E       �    �6@     1      �  "  �@     6       u�  "  @�A     �      ��    ~�@     }       ��    g�A     n       ��     !@     �       ��  "  ��@     *       �  "  ��A            z�    X�@     .       ��  "  H�A           ��    2�A     �      %�  "  ��A     (       m�    �9@     �       r�  "  p�A            L�  "  ��@     �      3�  "  �@     0        crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.5415 dtor_idx.5417 frame_dummy object.5427 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux graphics.cpp /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_keymap_us runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp filesystem.c ipc.c syscall.c fb.c itoa.c essential.cpp stdlib-stubs.cpp _ZN3frgL8null_optE _ZN3frgL6endlogE _ZN3frgL9dont_lockE _ZN3frg9_redblack12_GLOBAL__N_1L15enable_checkingE _ZN3frg12_GLOBAL__N_1L15enable_checkingE _ZZN13AllocatorLock4lockEvE8__func__ _ZN12_GLOBAL__N_111mblen_stateE _ZZ6strtolE8__func__ _ZZ6rand_rE8__func__ _ZZ5abortE8__func__ _ZZ13at_quick_exitE8__func__ _ZZ10quick_exitE8__func__ _ZZ6systemE8__func__ _ZZ6mktempE8__func__ _ZZ7bsearchE8__func__ _ZZ3absE8__func__ _ZZ4labsE8__func__ _ZZ5llabsE8__func__ _ZZ4ldivE8__func__ _ZZ5lldivE8__func__ _ZZ5mblenE8__func__ _ZZ6mbtowcE8__func__ _ZZ6wctombE8__func__ _ZZ8mbstowcsE8__func__ _ZZ8wcstombsE8__func__ _ZZ14posix_memalignE8__func__ _ZZ8strtod_lE8__func__ _ZZN5mlibc7strtofpIdEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIfEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIeEET_PKcPPcE8__func__ _GLOBAL__sub_I_stdlib_stubs.cpp ctype-stubs.cpp _ZZN5mlibc20polymorphic_charcode7promoteEcRjE8__func__ _ZZ8iswctypeE8__func__ _ZZ8towlowerE8__func__ _ZZ8towupperE8__func__ environment.cpp _ZN12_GLOBAL__N_117empty_environmentE _ZN12_GLOBAL__N_118find_environ_indexEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_110get_vectorEvE6vector _ZGVZN12_GLOBAL__N_110get_vectorEvE6vector _ZN12_GLOBAL__N_110get_vectorEv _ZN12_GLOBAL__N_113update_vectorEv _ZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcb _ZZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcbE8__func__ _ZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEEE8__func__ _ZZ6getenvE8__func__ _ZZ6putenvE8__func__ _ZZ6setenvE8__func__ errno-stubs.cpp stdio-stubs.cpp _ZZN13ResizePrinter6expandEvE8__func__ _ZZ6removeE8__func__ _ZZ6renameE8__func__ _ZZ8renameatE8__func__ _ZZ7tmpfileE8__func__ _ZZ6tmpnamE8__func__ _ZZ7freopenE8__func__ _ZZ6setbufE8__func__ _ZL9store_intPvjy _ZZ5scanfE8__func__ _ZZ6sscanfENUt_10look_aheadEv _ZZ6sscanfENUt_7consumeEv _Z8do_scanfIZ6sscanfEUt_EiRT_PKcP13__va_list_tag _ZZ7vfscanfENUt_10look_aheadEv _ZZ7vfscanfENUt_7consumeEv _Z8do_scanfIZ7vfscanfEUt_EiRT_PKcP13__va_list_tag _ZZ6vscanfE8__func__ _ZZ7vsscanfE8__func__ _ZZ8fwprintfE8__func__ _ZZ7fwscanfE8__func__ _ZZ9vfwprintfE8__func__ _ZZ8vfwscanfE8__func__ _ZZ8swprintfE8__func__ _ZZ7swscanfE8__func__ _ZZ9vswprintfE8__func__ _ZZ8vswscanfE8__func__ _ZZ7wprintfE8__func__ _ZZ6wscanfE8__func__ _ZZ8vwprintfE8__func__ _ZZ7vwscanfE8__func__ _ZZ5fgetsE8__func__ _ZZ6fgetwcE8__func__ _ZZ6fgetwsE8__func__ _ZZ6fputwcE8__func__ _ZZ6fputwsE8__func__ _ZZ5fwideE8__func__ _ZZ5getwcE8__func__ _ZZ8getwcharE8__func__ _ZZ5putwcE8__func__ _ZZ8putwcharE8__func__ _ZZ7ungetwcE8__func__ _ZZ7fgetposE8__func__ _ZZ7fsetposE8__func__ _ZZ8getdelimE8__func__ _ZZ14fgets_unlockedE8__func__ _ZZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ string-stubs.cpp _ZZ7strxfrmE8__func__ _ZZ6strtokE8__func__ _ZZ6wcstodE8__func__ _ZZ6wcstofE8__func__ _ZZ7wcstoldE8__func__ _ZZ6wcstolE8__func__ _ZZ7wcstollE8__func__ _ZZ7wcstoulE8__func__ _ZZ8wcstoullE8__func__ _ZZ6wcscpyE8__func__ _ZZ7wcsncpyE8__func__ _ZZ7wmemcpyE8__func__ _ZZ8wmemmoveE8__func__ _ZZ6wcscatE8__func__ _ZZ7wcsncatE8__func__ _ZZ6wcscmpE8__func__ _ZZ7wcscollE8__func__ _ZZ7wcsncmpE8__func__ _ZZ7wcsxfrmE8__func__ _ZZ7wmemcmpE8__func__ _ZZ6wcschrE8__func__ _ZZ7wcscspnE8__func__ _ZZ7wcspbrkE8__func__ _ZZ7wcsrchrE8__func__ _ZZ6wcsspnE8__func__ _ZZ6wcsstrE8__func__ _ZZ6wcstokE8__func__ _ZZ6wcslenE8__func__ _ZZ7wmemsetE8__func__ dso_exit.cpp _ZZ12getExitQueuevE9singleton _ZGVZ12getExitQueuevE9singleton lemon.cpp _ZZN5mlibc17sys_anon_allocateEmPPvE8__func__ allocator.cpp _ZZ12getAllocatorvE16virtualAllocator _ZGVZ12getAllocatorvE16virtualAllocator _ZZ12getAllocatorvE9singleton _ZGVZ12getAllocatorvE9singleton _ZZN16VirtualAllocator3mapEmE8__func__ _ZZN16VirtualAllocator5unmapEmmE8__func__ charcode.cpp _ZZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEEE8__func__ _ZZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEEE8__func__ _ZZN5mlibc16current_charcodeEvE15global_charcode _ZGVZN5mlibc16current_charcodeEvE15global_charcode _ZZN5mlibc22platform_wide_charcodeEvE20global_wide_charcode _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstateE8__func__ charset.cpp _ZZN5mlibc15current_charsetEvE14global_charset debug.cpp ensure.cpp guard-abi.cpp _ZN12_GLOBAL__N_15Guard6lockedE _ZN12_GLOBAL__N_15Guard4lockEv _ZN12_GLOBAL__N_15Guard6unlockEv file-io.cpp _ZN5mlibc12_GLOBAL__N_1L24globallyDisableBufferingE _ZN5mlibc12_GLOBAL__N_116global_file_listE _ZZN5mlibc13abstract_file4readEPcmPmE8__func__ _ZZN5mlibc13abstract_file5writeEPKcmPmE8__func__ _ZZN5mlibc13abstract_file5ungetEcE8__func__ _ZZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeEE8__func__ _ZZN5mlibc13abstract_file4seekEliE8__func__ _ZZN5mlibc13abstract_file10_init_typeEvE8__func__ _ZZN5mlibc13abstract_file13_init_bufmodeEvE8__func__ _ZZN5mlibc13abstract_file11_write_backEvE8__func__ _ZZN5mlibc13abstract_file6_resetEvE8__func__ _ZZN5mlibc13abstract_file18_ensure_allocationEvE8__func__ _ZZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeEE8__func__ _ZN12_GLOBAL__N_110stdin_fileE _ZN12_GLOBAL__N_111stdout_fileE _ZN12_GLOBAL__N_111stderr_fileE _ZN12_GLOBAL__N_111stdio_guardC2Ev _ZN12_GLOBAL__N_111stdio_guardC1Ev _ZN12_GLOBAL__N_111stdio_guardD2Ev _ZN12_GLOBAL__N_111stdio_guardD1Ev _ZN12_GLOBAL__N_118global_stdio_guardE _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ5fopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ5fopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ6fdopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ6fdopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZSt7forwardIZ5fopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _ZSt7forwardIZ6fdopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _GLOBAL__sub_I_file_io.cpp filesystem.cpp getwchar _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ stpcpy putchar _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13BufferPrinterEC1EPS0_PN3frg9va_structE _ZN5mlibc7charset8to_upperEj strcpy _Z12GetVideoModev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC1Ev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN3frg14format_optionsC2Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE6bucketC1Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ _ZN5mlibc13abstract_file4tellEPl unsetenv _ZN3frg8optionalIiEC2ERKS1_ _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN5mlibc7charset8is_alnumEj _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ _ZN3frg8optionalIiEC2IRivEEOT_ _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1ERS5_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev tmpfile mousePos _ZN5mlibc7charset8is_alphaEj _ZN3frg8optionalIiEaSES1_ _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ERS5_ vscanf _ZN13BufferPrinterC1EPc _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEEC2IJRS6_EEEDpOT_ _ZTVN5mlibc20polymorphic_charcodeE wcstok _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer stdout vsprintf _ZN3frg8optionalIiEC2Ev wcstof _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg17basic_string_viewIcEC2EPKc vswprintf _ZN5mlibc13abstract_file4readEPcmPm _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC1EPS3_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev _ZN11PrintfAgentI13BufferPrinterEclEPKcm _ZN5mlibc8code_seqIwEcvbEv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm ungetc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEEC1IJRS6_EEEDpOT_ _ZN3frg17basic_string_viewIcE10find_firstEcm _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ strerror _ZN5mlibc10sys_accessEPKci _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN13StreamPrinterC1EP17__mlibc_file_base _ZN3frg9_redblack15null_aggregator9aggregateINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic syscall _ZN5mlibc20polymorphic_charcodeC1Ebb _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN5mlibc8sys_openEPKciPi _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ reverse fileno_unlocked frameCounter _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg3maxImEERKT_S3_S3_ wcstoull _ZN5mlibc7fd_fileD1Ev atol _ZN5mlibc15current_charsetEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ lastUptimeMilliseconds ReceiveMessage _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv _ZN5mlibc13wide_charcode7promoteEwRj _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameC1ENS3_10frame_typeEmm _ZN3frg8optionalIiE13storage_unionC2Ev getenv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC1Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv wcslen iswcntrl _ZN13BufferPrinter6appendEc _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ iswpunct _Znwm lemon_read strtold isblank wcstoll iswalpha iswblank bsearch _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg14format_optionsC1ERKS0_ _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic vsscanf _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZN5mlibc7strtofpIdEET_PKcPPc qsort _ZN5mlibc13utf8_charcode12decode_stateC2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ wcsrchr _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ fgets _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ vwprintf _Z13AddNewWindowsv iswxdigit _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg8optionalIiEC1IRivEEOT_ _ZN5mlibc13abstract_file13_init_bufmodeEv _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic _ZN5mlibc13abstract_fileD2Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ _ZN8ListNodeIP8Window_sEC2Ev _ZN5mlibc9PanicSinkclEPKc _ZplRK8Vector2iS1_ setvbuf __TMC_END__ _ZTVN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEE _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv renameat perror SendMessage _ZN3frg10bitop_implImE3clzEm _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ __DTOR_END__ _ZN5mlibc7charset17is_ascii_supersetEv _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ _ZN3frg17basic_string_viewIwEC2EPKw dragOffset lemon_open _ZN5mlibc8sys_seekEiliPl islower _ZN5mlibc20polymorphic_charcodeD1Ev __fpurge tolower _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ _ZN5mlibc20polymorphic_charcodeD0Ev _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE iswlower _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic system _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv feof fgetws wcspbrk _ZN5mlibc7strtofpIfEET_PKcPPc wcstol _ZN5mlibc13abstract_fileD1Ev _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE malloc remove iswspace _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE _ZN13AllocatorLockC2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10tiny_sizesE _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic vsnprintf strtoll _ZN5mlibc13abstract_file18_ensure_allocationEv _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN13ResizePrinter6appendEPKcm _ZN5mlibc7fd_file2fdEv wcsncmp _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameC1Emmi strtoul __dso_handle itoa _ZN3frg8optionalIiEcvbEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED1Ev wcsstr _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _ZN5mlibc8code_seqIKwEcvbEv _ZN13BufferPrinterC2EPc _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE mktemp _ZN5mlibc13abstract_file5purgeEv ispunct _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC1Ev __mlibc_errno _ZN5mlibc20polymorphic_charcodeC2Ebb wctomb _ZN5mlibc12sys_libc_logEPKc _ZN13StreamPrinter6appendEc currentUptimeMilliseconds wcstombs _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ _ZN8ListNodeIP8Window_sEC1Ev _ZN3frg8optionalIiEC1ERKS1_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic _ZN4ListIP8Window_sE8add_backES1_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE clearerr_unlocked isspace vwscanf _ZN5mlibc13abstract_file7disposeEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic mempcpy fflush _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ _ZN13AllocatorLock6unlockEv _ZTVN5mlibc7fd_fileE lemon_map_fb _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ _ZN14LimitedPrinter6appendEPKc _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE _ZN5mlibc7charset8is_digitEj _ZN3frg11unique_lockI13AllocatorLockE6unlockEv mbstowcs _ZN5mlibc22platform_wide_charcodeEv _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic putenv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED1Ev wmemcpy _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZdlPv _ZN13StreamPrinter6appendEPKcm _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ vswscanf _Exit _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ _ZN5mlibc13abstract_file5ungetEc drag _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv backgroundColor abort _ZN4ListIP8Window_sEixEj _ZN3frg8optionalIiEC2EOi _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ wcscoll _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistC1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ ftrylockfile isxdigit _init _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ERS5_ _Z12getAllocatorv strtol _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC1Ev fsetpos __mlibc_rand_engine wcstod mblen iswprint _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZN5mlibc13abstract_file6_resetEv _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ lastKey active _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2ERS1_ _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE rename _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm _ZNK3frg17basic_string_viewIcE4dataEv _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _Z22RemoveDestroyedWindowsv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic strrchr _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv wcscpy _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ calloc memcpy_sse2_unaligned frameRate mouseData strtod _ZN3frg15aligned_storageILm456ELm8EEC1Ev _ZN3frg7mt19937clEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ _ZSt4swapIbEvRT_S1_ _ZN11PrintfAgentI13ResizePrinterEclEPKcm _ZN3frg7mt19937C2Ev wmemchr _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ atof _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ environ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ fputs_unlocked iswgraph _ZN13BufferPrinter6appendEPKcm _ZN3frg17basic_string_viewIcEC1EPKcm _ZN16VirtualAllocator3mapEm _Z16memcpy_optimizedPvS_m _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC1ES6_ strcat __ensure_warn _ZN13ResizePrinterC1Ev _ZN5mlibc7charset8is_printEj _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc rand_r _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv vprintf closeButtonSurface _ZN5mlibc8code_seqIcEcvbEv _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN5mlibc14sys_libc_panicEv _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE _ZN13ResizePrinter6appendEc _ZN5mlibc7fd_file5closeEv memset32_sse2 _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE fseek _ZN3frg8optionalIiEC1EOi _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev _ZN3frg7eternalI16VirtualAllocatorEC1IJEEEDpOT_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg8optionalIiE13storage_unionD2Ev lemon_write getdelim _ZN5mlibc7fd_file7io_readEPcmPm _ZN5mlibc13abstract_file4seekEli _ZTVN5mlibc13abstract_fileE wcstold _Z8DrawCharciihhhP7Surface _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE6bucketC2Ev stdin _ZN13BufferPrinter6appendEPKc _ZN10win_info_tC1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ _ZN5mlibc8InfoSinkclEPKc _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic _ZN5mlibc7charset8is_spaceEj _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ currentUptimeSeconds _ZN5mlibc8code_seqIjEcvbEv _ZN5mlibc13abstract_file10_init_typeEv _ZN3frg7eternalI16VirtualAllocatorE3getEv ferror strstr _ZN3frg7eternalINS_6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEE3getEv _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic __cxa_pure_virtual _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZN11PrintfAgentI13StreamPrinterEC1EPS0_PN3frg9va_structE _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic iswctype _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic strcoll _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE isupper _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ strncmp _ZN4ListIP8Window_sE6get_atEj _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE16_construct_largeEm _ZN5mlibc7strtofpIeEET_PKcPPc wmemset _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi _ZdlPvm _Z18memset64_optimizedPvmm strncpy _ZN3frg15aligned_storageILm1ELm1EEC2Ev program_invocation_short_name _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic _ZN5mlibc7fd_file7io_seekEliPl _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic _ZN3frg17basic_string_viewIwEC1EPKw funlockfile _ZN13ResizePrinter6appendEPKc _ZN11PrintfAgentI13ResizePrinterEC1EPS0_PN3frg9va_structE isascii _ZN3frg4swapERNS_8optionalIiEES2_ realloc _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ windowCount towupper _ZN5mlibc7fd_fileD2Ev _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZN5mlibc7charset8is_graphEj __cxa_atexit _ZNK3frg17basic_string_viewIcE4sizeEv _Z8DrawRectiiii10RGBAColourP7Surface _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ _ZN13StreamPrinter6appendEPKc _ZN3frg9_redblack15null_aggregator9aggregateINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ strtok at_quick_exit _ZN3frg8optionalIiED2Ev mouseDown _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic fdopen _ZN3frg7mt19937C1Ev _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface isalpha _ZN5mlibc13utf8_charcode12decode_stateC1Ev wcscspn _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE15_construct_slabEi wcstoul _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ strncat _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ wcschr _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN3frg10escape_fmtC1EPKvm _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev fread _ZN3frg3minImEERKT_S3_S3_ _ZN3frg8optionalIiED1Ev _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN5mlibc7fd_fileC1EiPFvPNS_13abstract_fileEE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic lastUptimeSeconds _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ strtoull _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN14LimitedPrinterC2EPcm fopen __bss_start wcsncat _Z8DrawRect4Rect10RGBAColourP7Surface _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm putwchar _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ main wcsspn _ZN11PrintfAgentI14LimitedPrinterEC1EPS0_PN3frg9va_structE ftell _ZN5mlibc7charset8is_lowerEj srand strxfrm _ZN5mlibc8code_seqIKcEcvbEv vfwprintf font_default _Z5floord _ZN13AllocatorLock4lockEv clearerr _ZN3frg15aligned_storageILm32ELm8EEC1Ev _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm _ZN5mlibc7fd_file8io_writeEPKcmPm _ZdaPv _ZnwmPv _ZN3frg15aligned_storageILm1ELm1EEC1Ev fclose _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ getchar _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN5mlibc10infoLoggerE isgraph wcsncpy _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ fgetpos isalnum _ZN3frg8optionalIiEC1Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14size_to_bucketEm tmpnam isprint _ZN4ListIP8Window_sED2Ev _ZN4ListIP8Window_sED1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ _ZN5mlibc16current_charcodeEv _ZNK3frg17basic_string_viewIwE4sizeEv _ZN3frg14format_optionsD2Ev fread_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ strcmp _ZN3frg17basic_string_viewIcE10sub_stringEmm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN5mlibc7charset9is_xdigitEj _ZN3frg8optionalIiE13storage_unionC1Ev _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE _ZN14LimitedPrinter6appendEc memset64_sse2 _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _fini _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic _ZN13AllocatorLockC1Ev _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg15aligned_storageILm32ELm8EEC2Ev _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic fgetc strerror_r _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE7reallocEPvm _ZN5mlibc13abstract_file11_write_backEv strtof strtod_l __cxa_guard_release strcspn _ZN3frg17basic_string_viewIcEC1EPKc _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ _ZN13ResizePrinter6expandEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic flockfile _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8freelistC2Ev iswdigit _ZN4ListIP8Window_sE10get_lengthEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE11_find_frameEm _ZN11PrintfAgentI13BufferPrinterEclEc stderr _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _Z15UpdateFrameRatev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj _ZN5mlibc11panicLoggerE _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ srandom _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC1Ev _ZN16VirtualAllocator5unmapEmm _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ _ZSt7forwardIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZN14LimitedPrinter6appendEPKcm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv putchar_unlocked _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg9_redblack11hook_structC2Ev _ZN13ResizePrinterC2Ev fputc _ZN14LimitedPrinterC1EPcm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv _Znam feof_unlocked _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC1ERS1_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _Z24CreateFramebufferSurface6FBInfoPv _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ getchar_unlocked _ZN11PrintfAgentI14LimitedPrinterEclEc fwide iswupper __ensure_fail _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ _ZN5mlibc13abstract_file5flushEv fflush_unlocked _ZN3frg14format_optionsC2ERKS0_ _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic fputws _ZN3frg14format_optionsC1Ev _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate fwrite_unlocked wmemcmp _ZN11PrintfAgentI13StreamPrinterEclEc lldiv _ZN3frg11unique_lockI13AllocatorLockEC1ERS1_ _Z12getExitQueuev wmemmove _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN5mlibc13abstract_fileC2EPFvPS0_E isdigit _ZN5mlibc13sys_anon_freeEPvm fwrite _edata _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _Z19__mlibc_do_finalizev _end _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _ZN5mlibc9sys_closeEi _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic vfscanf _ZN3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1ERS5_ _ZN3frg14format_options15with_conversionENS_17format_conversionE rewind _ZN3frg9_redblack11hook_structC1Ev freopen _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic fgetc_unlocked _ZN3frg14format_optionsD1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ ungetwc lemon_seek _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg7mt199374seedEj _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc13abstract_fileC1EPFvPS0_E _ZN5mlibc20polymorphic_charcodeD2Ev _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE towlower _ZN5mlibc7charset8is_upperEj llabs _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc9sys_writeEiPKvmPl setbuf _ZN5mlibc20polymorphic_charcode7promoteEcRj iswalnum wcscmp _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev _ZN3frg9_redblack11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ atoi _ZN11PrintfAgentI13ResizePrinterEclEc iscntrl _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ _Z10DrawWindowP8Window_s _ZN3frg11unique_lockI13AllocatorLockED2Ev ferror_unlocked _ZN5mlibc13abstract_fileD0Ev _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ fileno _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE fgets_unlocked getline _Z10surfacecpyP7SurfaceS0_8Vector2i _ZN5mlibc13utf8_charcode12decode_state6cpointEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ wcscat _ZN3frg15aligned_storageILm456ELm8EEC2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ strspn _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc strlen _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC1EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ program_invocation_name _ZN3frg10escape_fmtC2EPKvm toupper lemon_close _ZN5mlibc13utf8_charcode12decode_state8progressEv atoll _ZN5mlibc7charset8is_punctEj _ZN3frg8optionalIiEdeEv _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD1Ev _ZSt4moveIR11ExitHandlerENSt16remove_referenceIT_E4typeEOS3_ wcsxfrm _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1IJRS2_EEEDpOT_ _ZN4ListIP8Window_sE9remove_atEj _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE strchr _ZN5mlibc8sys_exitEi _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev fputs _ZSt4swapIPcEvRT_S2_ _ZN5mlibc17sys_anon_allocateEmPPv _ZN3frg3maxIiEERKT_S3_S3_ font_old _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN5mlibc8sys_readEiPvmPl _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE5frame8containsEPv _ZN3frg8optionalIiE13storage_unionD1Ev fgetwc vfwscanf _ZSt4swapIiEvRT_S1_ vasprintf fbInfo fputc_unlocked strchrnul _ZN3frg11unique_lockI13AllocatorLockED1Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZdaPvm lemon_readdir _ZN5mlibc7charset8is_blankEj memcpy_sse2 _ZN5mlibc7charset8to_lowerEj _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ aligned_alloc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ __cxa_guard_acquire posix_memalign _ZNK3frg17basic_string_viewIcEeqES1_ _ZN5mlibc7fd_fileD0Ev windows _ZN13StreamPrinterC2EP17__mlibc_file_base _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE mbtowc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic vfprintf strpbrk _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN3frg17basic_string_viewIcEC2EPKcm _ZNK3frg6vectorI11ExitHandlerNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv fputwc _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13abstract_file5writeEPKcmPm _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ free _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_14slab_allocatorI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ _ZN5mlibc18generic_is_controlEj  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .tbss .init_array .ctors .dtors .data.rel.ro .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                     � @     �                                     !              @            q�                            '             q�A     q�                                   -             ��A     ��     B�                              5             șB     ș     \                             ?              C                                          E               C                                         Q              C                                         X             ( C     (                                    _             8 C     8                                    l             `C     `     `                              r             �C     �     �                              w      0               �     +                             �                      �     �6                             �                      {D                                   �                      �D     D�                            �                      �1     C[                             �                      �     �y                            �                      �                                   �      0               �     �)                           �                      y0	                                   �                      �0	     `:                                                   �j	     �g         (                	                      ��	     S�                                                   ۗ
     �                              