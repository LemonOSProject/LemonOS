ELF              ��4   TD      4    (  
         � �T(  T(            0   � ��	  
                    �<  ��U������u��  ����U������u��  ����U������u��  �����U������u����������U������u�  �����U������u����������U����E�@�E�E�@�E��E�    �E�@9E���   �E�P�E)�9E�}|�E�    �E�@9E�}a�E�P�E)�9E�}O�E�@�E��E�Ѝ�    �E��U�E�E�@�ЋE�EЍ�    �E���E�딃E��c������U����E�@�E�E�@�E��E�    �E�@9E���   �E�P�E)�9E���   �E�    �E�@9E���   �E�P�E)�9E�}~�E�@�E��E�Ѝ�    �E�Ћ ��=�   vK�E�@�E��E�Ѝ�    �E��U�E�E�@�ЋE�EЍ�    �E�����E��a����E��,������U��S���E�@x�E��E�@|�E�E�@������  �E���   �H�E�P|�E�@xh��j j j QjRP�  �� �E���   �H�E�@|�U�Zx�U���   ڃ�h��j j j QjPR�}  �� �E���   �H�E�P|�E�@xh��j j j jQRP�M  �� �E���   �H�E�P|�E���   ЍP�E�@xh��j j j jQRP�  �� ���9Eu5�E���   �U�R|�J�U�Rx��h��j0j0j0jPQR��  �� �<�E���   �U�R|�J�U�Rx��h��h�   h�   h�   jPQR�  �� �E�@|���E�@x����h��h�   h�   h�   RPh���  �� �E�@x�P�E�@|���U��E�E��U�Rt�Ѻ����j j PQRj�  �� ��]���U��WVS��  ����E���j j j RPj�w  �� ������������P�t  ������������  �����j j j j Pj�-  �� fǅH���@fǅJ���� ǅL���    ���   ���   ���@�����8���P�A  �������j j j j Pj��  �� ��4��������j j j PRj�  �� ��0��������4�����j RjQPj�  �� ��0�����t^�X�������УX��X���y
�X�    �\�����ȸ    )��У\��\���y
�\�    �����t`�X�������)щʉPx�\�������)щʉP|����@x��y����@x    ����@|��y����@|    ������h��h�   h�   j@RPj j ��  �� ��,�����j j j j Pj�h  �� �E�    �U䋅,���9��Z  ��d����E��j j j RPj�2  �� �E�    ����8���P�  ��9E�����t�������E���P��8���P�e  ���@t9�����tN�E���P��8���P�C  ��ƀ�   �E���P��8���P�&  ���Í�d����   �߉Ɖ���   �E��e�����h�   �  ���EԋEԉÍ�d����   �߉Ɖ����d����ЋEԉPx��f����ЋEԉP|��h����ЋEԉ��   ��j����ЋEԉ��   �E�ƀ�   ���uԍ�8���P��  ����E���������������Z  ������K  �������8���P�  �����E܃}� �A  �E܃�P��8���P�  ���EЋX��EЋ@x9���  �X��EЋHx�EЋ��   �9���  �\��EЋ@|9���  �\��EЋH|�EЋ��   �9���  �E܃�P��8���P�  ����P��8���P��  ���E܃�P��8���P�]  ������EЋ@|�P�\�9�|B�EЋ@����u5�X��EЋ@x)\��EЋ@|)��ȉ���������	  �EЋ@����txǅ���   �X��EЋ@x)ЉE̡\��EЋ@|)�f�EʋE������E�Љ�����EЋPp�@l����������������������P�r  �� �   ǅ���   �X��EЋ@x)Ѓ��Eġ\��EЋ@|)Ѓ�f�EE������E�Љ�����EЋPp�@l�������������� ���������P��  �� �	�m������������u�����t
��� �������tQ���������u@��� ǅ����   ����Pp�@l��������������������������P�k  �� �E�    ����8���P�X  ��9E�������   �E؃�P��8���P�@  �����   ����t�E؃�P��8���P�$  ���E؃�P��8���P�  ����P��������E؃�P��8���P��   ��ƀ�    �E��^����������P�z  ��������t[��$���=� u�ǅ����   ��(����� �����������Pp�@l��������������������������P�N  �� ��5\��5X�h��h���>���������E���j j j RPj�  �� ������e�[^_]�U��]�U��E�@]ÐU����E�@��t�E�@9Er	�    � �+�E� �E��E�    �E�;Es�E�� �E��E���E��@�ÐU��E�     �E�@    �]ÐU�����j�,  ���E��E�    �E�    �E�    ���E�P�������E�U��U�P�U��P�E�U�P�E� ��u
�E�U���E�@�U��E�P�E�P�E�U�P�E�@�P�E�P���U����E�@��t�E�@9Er�    � �   �E� �E��E�    �E�;Es�E� �E�E���E�@�E�E� ��t�E� �U�R�P�E�@��t�E�@�U���} u
�E��E��E�@�P��E�P�E�@9E����t�E�P�E�P���u��	  ���E���U����'  L!  �E�    ��U�E�ЋU��E��E�;Er�E��U�����  !  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���  �à   �E���E�E���d  �E�    ��Ѕ�u��d  �E�    ���E����d  �E�    �����E䋃h  9E�s	��h  �E���u��A  ���E��}� u%���	  ���	  ���� ���	  ���	  �    �l�E��     �E��@    �E��U�P��d  �E�E��P�E��@   �E��@    �E��@�ƿ    ��ȹ�P� ����ȹ��Q�E��e�[^_]�U��WVS��L�Y  ��z  �E�    �E�    �E�    �E�    �E�E��E� �,  �}� u5���	  ���	  ���� ���	  ���	  �  ��j�������  ���	  ��u-���u��K��������	  ���	  ��u��
  �    �{  ���	  �E��E�    ���	  ���C  ���	  �P���	  �@)ЉE��E�    �E����    ;E؉�E��
  ���	  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ��	  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u���	  �E��E�    �|  ���u��9������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��й�P� ����й��Q��ع�0�x��й�P� 9Ɖ��s�Ɖ���ع�0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ��й�P� ����й��Q��ع�0�x��й�P� 9Ɖ��s�Ɖ���ع�0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���W  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    ��й�P� ����й��Q��ع�0�x��й�P� 9Ɖ��s�Ɖ���ع�0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    ��й�P� ����й��Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u���	  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������X  �    �e�[^_]�U��WVS��,�%  ��F  �} u#���	  ���	  ���� ���	  ���	  �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx���	  ���	  ���� ���	  ���	  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u���	  ���	  ���� ���	  ���	  �b  �  �E��@�E���й�P� �M��I�ο    )����й��Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ���	  9E�u�E܋@���	  ���	  9E�u
ǃ�	      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋���ȹ�P� �M܋I�ο    )����ȹ��Q�E܋@��P�u��y  ���G���	  ��t=���	  �P���	  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉��	  ��  �e�[^_]�U��S���  �  �U�U�U�U��R���%������E��E��Pj �u��?������E��]���U��S���^  ��  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E���   �E���E�E�@=���tz���	  ���	  ���� ���	  ���	  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u���	  ���	  ���� ���	  ���	  �   �    �_�E�@�E�E�;Er�E�U�P�a   �E�;�W   ���u��������E���u��u�u����������u��������E�]��Ë$Ë$�U�������  �    ]�U�������  �� ��  �    ]�U��S�������  �M�U��j j j QRj���   �� �E�]���U�������  �    ]�U��WVS�r����  �E�]�M�U�u�}�i�[^_]�U��S���G���l  �M�U��j j j QRj�������� �E�]���U��S������6  �U�U�U�U���j j �u��u��uj���j����� ��]���U���������  �E�������E����	��E����	��E��	ЉE�E�@�E��E�    �E9E�}G�E�    �E9E�}2�U�E�E�@�M�U��Ѝ�    �E�E��E��ƃE�뱐��U��S���0���U  �U��j j j j Rj �������� ��E�]��� U��������  �M�U�E �M�U�E�} y�EE�E    �} y�EE�E    �E������E���	��E�	ЉE�E$�@�E��E�    �E�;E}k�U��EE$�@9�}Y�E�    �E�;E}D�U�E�E$�@9�}2�U��EE$�@�M��U�Ѝ�    �E�E��E�봃E�덐��U�������6  �} y�EE�E    �} y�EE�E    �E�������E����	��E��	ЉE�E�@�E��E�    �E�;E}k�U��EE�@9�}Y�E�    �E�;E}D�U�E�E�@9�}2�U��EE�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��� �1���V  �E�E�E�E��E��}��E��f�E��m��]��m��E��E�������v�E�����E���U��S��4�7  ��  �U���������P��H����E��Eԃ��d$��$���l��������E��E�    �E�   �E�    �E�;E��   �E�    �E�;E��   �U�E�E�@�������U�E���E�ȉE��U���ЉE�E��E�P�E�����U���ЉE�ЍP�E��E�@�U�������U���ЉE�ЍP�E��E�@�U�������E��F����E�E�E��$�����]��Ë$�U��WVS��<�����û  �u�M�U�}���EԈMЈỦ��E��E�    �}���   �U�������E��� ���E��E�    �}�]�E�   �����#E܉E������Ѕ�t7�}��u��MЋE� �EE�EċE�E��u WVQjjRP������� �E�띃E��f�����e�[^_]�U��WVS��,�����  �EȋM�U�E�MԈUЈE��E�    �E� ��tC�}��u��]ԋM�U�EЉE� �����u WVSQRP�]������� �E��E볐�e�[^_]�Window /shell.lef /fm.lef /dev/mouse0        zR |�        ����    A�BR�     <   ����    A�BR�     \   ����    A�BS�     |   ����    A�BS�     �   ����    A�BS�     �   |���    A�BS�     �   s����    A�B��    �   ����    A�B��       �����   A�BD����,   @  �����   A�BI�����A�A�A�      p  ����    A�BB�     �  t���    A�BG�     �  `���Q    A�BM�    �  ����    A�BU�     �  �����    A�B��      ����    A�B��    0  ����7    A�Bs�     P  ����r    A�Bn� ,   p  "���&   A�BF����A�A�A�   ,   �  ���4   A�BF���'�A�A�A�   ,   �  ���~   A�BF���q�A�A�A�          j���K    A�BD�C��     $  ����f   A�BD�^��   H  ����          \  ����          p  ����    A�BP�     �  ����    A�BY�      �  ����6    A�BD�n��     �  ����    A�BP�  (   �  ����*    A�BC���`�A�A�A�        ����6    A�BD�n��      D  ����?    A�BD�w��     h  �����    A�B��     �  W���7    A�BD�m��     �  j����    A�B��    �  3����    A�B��    �  ����Q    A�BM�       $���C   A�BD�;��   0  C���       (   D  3����    A�BF�����A�A�A�(   p  �����    A�BF���x�A�A�A�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     �                               �             �   �            �����   �           ���������   �          �������������   �         �����������������   �        ���������������������   �       �������������������������   �      �����������������������������   �     ���������������������������������   �    �������������������������������������   �   ���������������������   �   �   �   �   �   ���������   ���������   �����      �����   �    ���������   �      �   �     ���������   �����      ����   ���������   �          ���������   �       ����   �   �����  @  �                                                                                                                                                                                                                                                                                                       <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;              GCC: (GNU) 8.2.0                        ��          ��          ��           �           �          ��                                ���  ��       
            ���            ��   �        �     '   d�     2   h�     >   �     M   �     Z   ��     m   ��7     }   ��r     �   R�&    �   x�4    �            ���            ���            ���            ���            ��             ���    �      �   3�       ȹ       ��7     /  ЌQ   "  F  X�     O  "�   "  j  ع     v  ^�*     ~  ��     �  ��6     �   �     �  ��     �  ��   "  �  й     �  ��?     �  ��     �  ΁�     �  x�4      ۛ       ��     )   �     6  ؍�   "  U  ��     ]  ��     d  Ă�    {  ��     �  �     �   �     �  ��     �  *�K     �  ��     �  7��     �  ��      �  ��   "  �  @�    �  �6       ʀ       u�f      ���     9  ߛ     O  ��     Y  �C    |  ֝�     �  ��     �  ��      �  ���     �  `�     �  ��     �  ��Q       �       Č   "  0  <��   "  P  "�   "  k  J�     y  ���      ��     �  ��      �  �      �  ��     �  ��     t  ��~     init.asm main.cpp l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 _liballoc.c syscall.c ipc.c graphics.cpp text.cpp _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx l_allocated _Z12GetVideoModev _ZN4ListIP6WindowEixEj mousePos _ZN8ListNodeIP6WindowEC1Ev l_max_inuse syscall liballoc_unlock ReceiveMessage _Znwm _ZN4ListIP6WindowEC2Ev l_inuse SendMessage dragOffset _Z12surfacecpy_tP7SurfaceS0_8Vector2i malloc __x86.get_pc_thunk.ax mouseSurface transparency _ZN4ListIP6WindowE9remove_atEj surface _ZdlPv _Z10DrawWindowP6Window drag liballoc_lock keymap_us active calloc mouseData _Z8DrawCharciihhhP7Surface _ZN4ListIP6WindowEC1Ev mouseSurfaceBuffer liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface testKey font_default _Z5floord _ZdaPv _ZN4ListIP6WindowE10get_lengthEv _ZN4ListIP6WindowE8add_backES1_ _ZN8ListNodeIP6WindowEC2Ev liballoc_free pmain _Znam _edata _end _Z10surfacecpyP7SurfaceS0_8Vector2i _ZdaPvm  .symtab .strtab .shstrtab .text .rodata .eh_frame .got.plt .data .bss .comment                                                     ���   "                 !         ���"  &                  )         ���"  �                 3          � 0                   <          � 0  `	                  B         ���9  �                  G      0       �9                                 �9  �  	            	              D?  �                               D  P                  