ELF              ��4   $`      4    (           � ��@  �@           �@  ����h
          �W  �2  �                 �    UU���&  VW�����_^�  �    �i���f�f�f�f�f��(�=(�t$�    ��tU���h(��Ѓ��Í�&    f�Í�&    ��&    ��(�-(����������t(�    ��tU���Ph(��҃��Í�&    �t& �Í�&    ��&    ��=@� ugU�D���V���S�����������9�s�v ���D����D�9�r��'����    ��t��h��Q~�����@��e�[^]�Í�&    ��&    ��    ��t'U���hH�h��~������	�����&    f������U�� �i�mN�A90  � �� ���%�  ]�U��S���t����9�sz�U��E��j j j RPj�E/  �� �E���    �h��l�)�Ӊȉ�i��  �M��p�)щ�¡t�Уt��E��    �h��l��E�p��w����t�    ��]���U��WVS����j�a  ���ǃ�W�/  ���=|��|��E�   �E�   ���u��u�P�B  ���|��	   �   ��VSP�%  ���`�    ��������������e�[^_]ÍL$����q�U��WVSQ���  �ȋ ��T�������p���P�c
  ��fǅt��� fǅv��� fǅp���@ fǅr���  ǅx���    ��j�v  ���Ã�S�D
  ���|��|��   �   ��WVP�_
  ���|�ǅ���	   ǅ���   ������������P�.
  ���E�    �}�.�E�    �}��E����E�����  �E��߃E��̃���p���P�  ���E������`���tR�����t+��������������� ��� ������`�    ����������������\���P�R,  ����������   ��d�����ui�x���t�x� ������h���=  t)=  w	=
  t�=  t=  t��E�    �>�E�   �5�E�   �,�E�   ��"��d������^������u��  ���<,  �F����x����C  �E�    �}�.�E�    �}��E����E�����  �E��߃E��̡����t�   ��   �����������E�    �|���P��  ��9E�����t[�|��EЍ�������PQR�  ���������|��EЍ�������PQR�  ���������������� �E���E�    �}���   �E�    �}���   �Eč��   �E����E����� ���������E����E����� �������؋E����E����� �������ЋE������E���WVSRjjQP�  �� �E��[����E��A����}���   �}��}� t�  �}��W  �}���  �  �|��|���P�`  ������������RSP��  ���|��|���������j RP�2  ���������� ����|��������j RP�  �����������$�������$����� ���S�  ����  �|��|���P�  �����������RSP�9  ���|��|��������j RP�  �����������(����|��������j RP�d  ���� �����,�������,�����(���S��  ���D  �|��|���P�  ������$�����RSP�  ���|��|���,�����j RP��  ����,�������0����|���4�����j RP��  ����8�����4�������4�����0���S�<  ���   �|��|���P�t  ������<�����RSP��  ���|��|���D�����j RP�F  ����D�����8����|���L�����j RP�  ����P�������<�������<�����8���S�  ����|���T�����j RP��  ����T����|���\�����j RP�  ����`����������� <��   �|���d�����j RP�  ����h�����xq�|���l�����j RP�^  ����l�����xL�|���t�����j RP�9  ����x�����&�|���|�����j RP�  ����|�����~�   ��    ��t]�x��E��   ��Ph�   h�   h�   j j h̲�/  �� �E��   �Eċ@��j j j RPj�:&  �� �~  �|��E���j RP�  ���]��|��E���j RP�h  ���U��������� <������   �|��E���j RP�1  ���]��|��E���j RP�  ���U���������  ���������������������������������t���   �
���    �|�ǅ@���    ǅD���    ����D�����@���P��  ���B  �|��E���j RP�r  ���]��|��E���j RP�W  ���U��������� <������   �|��E���j RP�   ���]��|��E���j RP�  ���U���������  �`�   �����������������������������������������������������)Ѕ�����t���   �
���    �|�ǅH���    ǅL���    ����L�����H���P�   ���E��   �Eċ@��j j j RPj�#  �� ����������U��Ef�   �Ef�@  �Ef�@  �Ef�@  �]ÐU��E�     �E�@    �E�@    �]ÐU��E�     �E�@    �]ÐU��S����j��  �����    �C    �C    �C    ��S�������]�E��     �M�E�U�A�Q�E� ��u
�E�U���E�@�U��E�P�E�P�E�U�P�E�@�P�E�P��]���U��E�@]ÐU����E�@��t�E�@9Es	�E� ��u�E� �M�P�@��Q�J�E� �E��E�    �E�;Es"�E�@9E�s�E�� ��t�E�� �E��E��֋M�E��P�@��Q�E�� U���(�E�@��t�E�@9Er�M�E��U��Q��   �E� �E��E�    �E�;Es"�E�@9E�s�E� ��t�E� �E�E��֋E�P�@�E�U�E� ��t�E�@��t�E� �U�R�P�E�@��t�E� ��t�E�@�U���} u
�E��E��E�@�P��E�P�E�@9E����t�E�P�E�P���u��  ���M�E�U��Q�E�� �U��S����j�  �����    �C    �C    �C    ��S�`������]�E��     �M�E�U�A�Q�E�@��u�E�U�P��E� �U�P�E��E��E�U��E�@�P�E�P��]���f�f�f�f�f��UWVS��
  ��w?  ���D$(�|$$�ƃ�)����ŋD$ ��	��t>��QW�t$,�   ����u	��[^_]Ð���/VR�D$,�P��  ����[^_]Ð��QW�t$,�  ������&    ��    UWVS�P
  ���>  ���t$ �|$$�T$(��   t*�B���t�v ���>�����u��[^_]Í�&    �t& ������R��WV�m  ����tӉ>��t̉~��tĉ~��[^_]Í�&    �t& ���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���|$$�L$,�D$4�\$8�t$(�T$0�|$�L$��y��D$    �L$��y�1����ȁ�   ���	���% �  ���͉���	�k	ǅ�~u;s}p�D2��L$�D$�D$�D��$��&    �D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�  ��)=  ���t$j j j j Vj ��  ��$��[^� f��`  �<  UWVS��,�|$@�t$D�D$�L$L�D$P�\$T�T$X�l$\��y|$H1���y�1�����������	�	E�T$�D$��~\;u}W�D$H��D$�D��D$�
f���9u~9�]������)�;\$OT$H��R��t$�L$ ��P�\$�X�����;t$u���,[^_]Í�&    �  +<  UWVS��,�t$@�l$D�D$�L$L�D$P�|$T��yt$H1���y�1��؉������� �  ��	�	G�T$�D$��~i;o}d�D$H��D$�D��D$��t& ���9o~C�G�_������)����;\$OT$H��R�t$�L$ ���P�\$�~�����;l$u���,[^_]Í�&    ��    UWVS�  ��G;  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$�������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�@  ���9  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�,����� 9t$h�_�����L[^_]Í�&    UWVS�p  ��8  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�\����� 9t$l�_�����L[^_]Í�&    UWVS�  ��76  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�)�����9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$Ë$�f��S�   ������Å4  ���D$��D�P��
  ��[Í�&    �S�������Z4  ���t$��
  ��[Ív S������:4  ���t$�  ��[Ív S������4  ���t$�������[Ív S�c������3  ���t$�H  ��[Ív S�C������3  ���t$�(  ��[�f��UWVS� ����÷3  ���D$<�|$8�t$0�D$�G�D$�D$D���� ��D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�M����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�~����� 9|$�b�����[^_]Í�&    f�UWVS�������W1  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��S�C������0  �� j j j �t$4�D$$Pj�  �D$,��8[�f�S�����ê0  ��j j j j �t$(j!�^  ��([Í�&    f�S�������z0  ��j j j �t$(�t$(j�,  ��([Í�&    UWVS������G0  ��(�l$<U�T����$�   �D$�����+   �T$����1����FjtUPǆ�   ����ǆ�   �����V�  �}�m����    ���� ��f��� vf��� wd���   ������P�/  �����   ���   ���   ��ǆ�       ǆ�       Ɔ�    Ɔ�    ��[^_]Í�&    ��&    �ȃ���P��  ��롍�&    ��    S������:/  ���D$�p�u�����[��  ��/  UWVS���l$0�T$�Eu(�����   S�����   �EP�EPj j ������ �E���   ��~?1����   �v 9�v\�M ��t1��v ���	9�u��A�������WP��E��9�̋��   ��t	��S�Ѓ���S�u�\$�������,[^_]Ð�    ��&    f�UWVS���D$0�l$4�|$8�p��~G� 1ۉD$��&    ��&    9�t<�D$��t1�f���� 9�u��@�P�H9�~9�|&��9�uσ�[^_]Í�&    �    ��&    f�H9�~�P9�~̅�t�T$1���&    ����9�u��T$�D$���@�P�R�D$@�����   ��[^_]Í�&    ��&    S���\$���   ��xn;CsY���t1Ґ���	9�u��A���P�R���   ��;Ss-���t1��t& ����	9�u��A��[Í�&    ��&    ��    ��&    f�ǃ�   ������1�[Í�&    ��&    �VS�2������,  ���t$ j�%����T$ ���     �P��@    ��t�V��P�F�F��[^Ív ��F�F��[^Ë$�f�f�f�f�f�f��U��E�]�Mfof ��������]�U��E�]�M�o� ��������]�U��E�]�M��~4fn�fo �f��fs�f��fs�f��fs�f��f ������]Ð������                U��01�WVS�����ò+  ��(��T
  �����9�P
  C�P
  P����  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p��1���T
  �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � ������  ���   �g�����&    �t& ����+*  ǀ�      ��ǀ�      �    �B    ��ǀT
     �    �B    ��ǀP
      �    �B    ǀ�      ǀ�      ǀ�      ǀ�      ǀ�      ǀ�      Í�&    �UWVS�������w)  ���|$0� ��&    ����  �   ���   �
  �w �
  ��t܋��  �t$�|$0����  �|$0���  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s���  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ����  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$���������B1ҋD$~Q��@�����   ��   �E��  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,�����E$���~�ƈ�Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ��������������  ���K����  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~�ǈ��N,�����ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��4  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS� ����×%  ���D$ ����   �P���)փ� C��  �N�A=����~   �y�Ő�1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o���  ����   ��t�J+J�ʋO)�9�|W�B  ��[^_]Í�&    �v ���  ���   ����� ���� t
f=��t<�u����  ���   뱍�&    ����  롍�&    ����  ���   ��[^_]Í�&    �v �G9��  tU9�ta���t�B�G��t������G1�)Q���wW��  ���4�����&    �t& �o�������&    ����  룍�&    �ǃ�      듍t& WVS�t$�M������#  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS�`������"  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��  �G�P�������   �P9���   �T$��  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ��  ���   %��� =�� tDf����t=���t8�3  1���[��^_]Í�&    �p���  ����[^_]Í�&    �t& ����  ���   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ�����f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f�S������Ê  �� j j j �D$ P�t$8j�;   �D$,��8[�f�S�������Z  ��j �t$0�t$0�t$0�t$(j�   ��([�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��S�c������  ��j j j j j j������ ��&    ��    ���f�f�f�f�f�f��1�Í�&    ��    �����  �����  1�Í�&    �v S������Ê  �� j j j �D$ P�t$8j�;����D$,��8[�f�1��f�f�f�f�f�f��������t6U��S�������&    �v �Ѓ�����u��[]Í�&    ��&    ������     Game Over, Press any key to Reset          zR |�        ����'    A�Bc�      <   �����    A�BD���� (   `   x����    A�BF�����A�A�A�   �   r���)    A�Be�  ,   �   �����
   D Gu Fupu|uxut   �   L���#    A�B_�     �   P���    A�BU�        J����    A�BD����    @  ����    A�BG�     `  �����    A�B��    �  ���   A�B�    �  ����    A�BD���� �   �  �����    A�A�A�A�N c$A(A,D0H G
A�A�A�A�BC$D(A,G0H C
A�A�A�A�BC$A(A,D0H    \   H  �����    A�A�A�A�N n
A�A�A�A�LC$F(D,A0H YA�A�A�A�   �  ����?    Cy 8   �  �����    A�A�A�A�C$�A�A�A�A�8   �  ����.    A�A�NFB B$B(A,B0HC�A� H   8  �����    K�A�A�A�C@�DAHFLHPL@IA�A�A�A� H   �  (����    K�A�A�A�C@�DAHDLJPL@IA�A�A�A� <   �  ����b   A�A�A�A�NPL@�A�A�A�A�X     �����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   l  `����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   �  �����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8     8����    A�A�A�A�C(�A�A�A�A�   P  ����          d  ����           x  ����(    A�SJ HA�     �  ����    A�ND HA�     �  ����    A�ND HA�     �  ����    A�ND HA�       ����    A�ND HA�     ,  ����    A�ND HA�   P  ����W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   d  ���s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�  0   �  @���.    A�N(B,B0B4D8E<B@LA�  0   �  <���'    A�NBB B$B(D,B0HA�  0   $  8���)    A�NBB B$D(D,B0HA�  `   X  4���   A�A�A�A�N<E@a4M8A<A@g0g<G@H0y
A�A�A�A�OE<D@H0      �  ����     A�NG HA� x   �  �����    L�A�A�A�C0Q8G<H@EDEHBLBPH0w8H<A@H0Q<A@E0C8A<C@LA�A�A�A�B0����X   \	  0����    A�A�A�A�C0]
A�A�A�A�HD<F@J0IA�A�A�A�0   �	  �����    A�CkC La
A�P]C� <   �	   ���_    A�A�NF Lh
A�A�DLA�A�      ,
  ?���       D   @
  �����   A�F�A�A�N<Z@J0�
A�A�A�A�M      �
  $����       T   �
  �����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `   �
  H����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   X  �����    A�A�A�WA H��A�A�  �   �  L����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0<      l���   A�A�A�A�C �
C�A�A�A�A 8   `  <����    A�A�A�A��
�A�A�A�P   0   �  ����.    A�N(B,B0B4E8D<B@LA�  0   �  ����-    A�NBD D$D(D,B0HA�  (     ����!    A�A�A�[�A�A�,   0  ����3    A�NBB B$B(B,B0H     `  ����          t  ����       0   �  ����.    A�N(B,B0B4E8D<B@LA�     �  ����           ����    ����                        `�`�@@@�@@@�@@ �`�`�S   S      d                                                                                                                                                                                                                                                                                                <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              p��                           >        p��    src/gfx/sse2.asm NASM 2.14.02 �p�     %  . @   l    '   �       src/gfx/sse2.asm      p�!0==?LL==0/!$!0==?LL==0/!#!0==>=0K�KYKYKYMK>1/""u�                                               t�          ��          ��          ̲          �          ��          ��          ��          ��     	     @�     
                                                                                                                             ��   ��         ��      (   �      ;   ��      =    �      P   P�      f   @�    
 u   D�    
 �   Ё      �   H�    
             ���   ��      �   ��      �   ��      �            ��  ��                  ��           ��#           ��/           ��8           ��C           ��L           ��]  |�       n  ��       �  �       �  ��       �   �     ?           ���  ��    �  $�    	 �   �    	 �  ��    
 �  ��    
 �  ��    
 �  ��    
   ��    
            ��'           ��-           ��7           ��>           ��             ��J  ��      `  ��    
 l  ��.     ~  ���    �  |�    
 �  �.     �  ���   "  �  @�   "    ��    
 !   �'     6  ��    
 C  ��!     K  ���     Y   �     i  @�.     �  ��    
 x  @�(   "  ~  ��    	 �  ��    �  ���     �  ��    
 �  (�    	 �  p�-     �  ��     �  ���       P��      ��    	 "  Z��   "  C  5�     Y  ��    	 f  p�    
 s  ��   "  z  ,��     �  _�     �  ���     S  t�      �  �     �  ��    	 �  @�   "  �  `�    
 �  �)   "    ���     -  ��     4  ��      J  P��     d  x�    
 m  �#   "  �  �W    �  �)   "  7  ��&     �   �_     �  �    	 �  @�.     �  ��   "  �  Э�    �  ���       9�     4  ��    
 B  ��    `  �    	 t  ��b    �  Г�     �  ��      �   �    	 �  p�s     �  ��  "    ̂�        h�    
 2  (�     
 >  ���     d  ��    k  _��
    p   �    	 }  p�?     �  М   "  �  t�    
 �  ��      �  �#   "  �  P�)     �  �'     �  p�     �  ��    
 �  p�   "  �  ��    	 
  ��   "  '  (�     	 .  ��     
 3  `��     M  б3     R  ��   "  t  ���     �   �    	 �  ��      �  �   "  �  p�      �  @��     �  0��     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp graphics.cpp runtime.cpp text.cpp window.cpp font.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset_sse2.loop memset_sse2.ret bigzero allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns memory.c ipc.c syscall.c exit.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface snake _Z13_CreateWindowP10win_info_t _ZN4ListI8Vector2iE9add_frontES0_ _ZN8ListNodeI8Vector2iEC1Ev l_max_inuse _Z14_DestroyWindowPv powerUpTimer syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm bgColourDefault _Z12DrawGradientiiii10RGBAColourS_P7Surface memcpy l_inuse __TMC_END__ SendMessage __DTOR_END__ _Z11PaintWindowP6Window malloc frameWaitTimeDefault _ZN4ListI8Vector2iE8add_backES0_ __x86.get_pc_thunk.ax __dso_handle lastUptimeMs _ZdlPv _Z4Waitv __x86.get_pc_thunk.dx _Z15HandleMouseDownP6Window8Vector2i liballoc_lock frameWaitTime _ZN8ListNodeI8Vector2iEC2Ev powerUp _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm calloc memcpy_sse2_unaligned _Z16memcpy_optimizedPvS_m gameOver _ZN4ListI8Vector2iEC2Ev _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev _Z9AddWidgetP6WidgetP6Window applePos liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx snakeMapCells _Z12CreateWindowP10win_info_t powerUpTimerDefault _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window rand_next _Z10DrawStringPcjjhhhP7Surface _ZN4ListI8Vector2iE9remove_atEj _Z5Resetv lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main font_default _Z5floord _ZdaPv msCounter _fini _ZN4ListI8Vector2iEC1Ev _Z12_PaintWindowPvP7Surface _Z4randv liballoc_free fruitType _Znam snakeCellColours _ZN4ListI8Vector2iE6get_atEj _edata _end _Z13HandleMouseUpP6Window exit _ZN4ListI8Vector2iE10get_lengthEv _Z10surfacecpyP7SurfaceS0_8Vector2i font_old memset_sse2 _ZdaPvm memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                   t�t                     !         ���   12                 '         ���2                    -         ̲�2  "                  5         ��2  �                 ?         ���@                    F         ���@                    M         ���@                   V         ���@  H
                  \         @�(K  �                  a      0       (K  +                 j              SK                     y              sK                    �              �K  B                  �              �K                    �              �K  p                  �              XL                    �              \L                                  lL   
     @         	              lV  �                               \_  �                  