ELF              ��4   �      4    (           � �@[  @[            `   � ��
  �        �W  ��A  �                 �    UU����'  VW�����_^�g  �    �i���f�f�f�f�f����=��t$�    ��tU���h���Ѓ��Í�&    f�Í�&    ��&    ����-�����������t(�    ��tU���Ph���҃��Í�&    �t& �Í�&    ��&    ��=�� ugU�����V��S���������9�s�v ����������9�r��'����    ��t��h���Q~��������e�[^]�Í�&    ��&    ��    ��t'U���h��h���~������	�����&    f������U��S��   ������L���Pj R�m;  ���E��E�    �E�    �E�    �}� ��  �E����EԋE���E��E�`   �E�H   ��hp  �  ���Ã��u��u��u��uԍ�L�����PS�\  �� �]�E�ƀ�   /�E�ƀ�    �E��   ����L�����RP�o5  ���E��   ��P�4  ���P��E����   <fuy�E��   ��P�[4  ���P��E����   <euS�E��   ��P�54  ���P��E����   <lu-�E��   ��P�4  ���P��E����   <.u�   ��    ��t�E��@a�E�ǀ�      �EЃ�u�E�ǀ�      ����P�u���!  ���E��E���у���L���RPQ�9  ���E�E�d�E��Pc�$���9��F����E�L�E�    �6�����]��ÍL$����q�U��VSQ��<�ȋ �E�f�$��f�&��f� �2 f�"�2 �(�    �,�File�0� Man�4�ager�8� ��h ��  ������j h����7  ������h��h���!  ���E���u���"  ���E����u��E&  ��� �� ��u�j�u�P�
"  �����u���!  ����h��h���P!  ���E���u��"  ���E����u���%  �������u�j�u�P�!  �����u��h!  ����h��h����   ���E���u��1"  ���E����u��%  �������u�j�u�P�J!  �����u��!  ���4������E�P�9  ����������   �EЃ�u��y�EЃ�u����P�  ��뾋EЃ�u2�E���f�EދE�f�E��Eމ��E܉ơ���VSP��  ��넋EЃ��x�������P��  ���'9  ���[�������P��  ����D���U����}u�}��  u��h ��!   �����U�����h��  j��������ÐU��Ef�   �Ef�@  �Ef�@  �Ef�@  �]ÐU����E���u�u�u�u�uP�U  �� ����E��Eǀ�       ���U����E�@ �E�@a��t�E�   ��j j j j Pj�8  �� �E���   ��uP����P�.5  ����    �E�   ��j P��4  ��������t����P��  ����ÐU��VS�E�@���r  �E�@��������X��E�@�H��E�@�P�E�@���uh�   h�   h�   SQRP�  �� �E�@��������X��E�@�H��E�P�E�@�������E�@���uh�   h�   h�   SQRP�+  �� �E�@�H��E�@�U�R���uj`j`j`jQPR��  �� �E�@�H��E�P�E�@ЍP��E�@���uj`j`j`jQRP��  �� �E�@�H��E�@�P�E�@�uj`j`j`QjRP�  �� �E�@�H��E�@�P�E�X�E�@؃��uj`j`j`QjRP�]  �� �E���   ��u@� ��E�P�E�X�E�@�������؃����uQj0j0RP�  �� �   �E���   ��u=���E�P�E�X�E�@�������؃����uQj0j0RP�g  �� �I�E���   ��u;���E�P�E�X�E�@�������؃����uQj0j0RP�  �� �E�P�E�@Ѓ��ËE�P�E�@�������E�@X��)ЉE�����uj j j SRP�  �� ��e�[^]ÐU����E� �E�E� ��t�E� �E����u��'  ���E��E��ًE�     �E�@    �E�@    ���f�f��UWVS�
  �ÓU  ���|$$�D$ �l$(	��t��UW�t$,�+  �������)�����RW�t$,��  ����u
��[^_]�f����VW�t$,�V�]+  ����[^_]�f���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�ÐUWVS���D$4�|$,�L$$�\$8�T$0�t$(�|$�ǉL$�ȁ�   ���	���% �  ���͉���	�k	ǅ�~o;s}j�L$�D$�T2��T$�D��$��D$��~<�C�L$9�|�/��&    �t& �C��9�~�S�������ʉ|� ;$u�9t$t��9s���[^_]Í�    VS�~  ��T  ���t$j j j j Vj ��2  ��$��[^� f�UWVS���|$�t$ �l$(�D$,�\$0�L$4�T$8��y|$$1���y�1�����������	�	��B�D$��~j;r}e�D.��$�D$$�\���&    f��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS���|$�t$ �\$(�D$,�T$0��y|$$1���y�1���������� �  ��	�	��B�D$��~m;r}h�D��$�D$$�\���&    �t& ��B�j������ƃ|$$ ~'9�~#�l$�l� �����&    ��9B~�L� 9�u�94$t��9r���[^_]Í�&    �t& UWVS�  ��3R  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$��������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�<  ���P  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�<����� 9t$h�_�����L[^_]Í�&    UWVS�l  ���N  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�l����� 9t$l�_�����L[^_]Í�&    UWVS�  ��#M  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�������9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$�f�f�f��S�   �������qK  ���D$��D�P��  ��[Í�&    �S������FK  ���t$��  ��[Ív S������&K  ���t$��  ��[Ív S������K  ���t$�������[Ív S�_������J  ���t$�  ��[Ív S�?������J  ���t$�  ��[�f��UWVS�����ãJ  ���D$<�|$8�t$0�D$�G�D$�D$D�������D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������� ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�]����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ�*����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��������t$H���t$�t$�D$PjjW�D$P����P������ 9|$�b�����[^_]Í�&    f�UWVS������CH  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��Ð��&    ��&    Ð��&    ��&    �D$�@Ð��    �D$�@Ð��    �D$�@ Ð��    UW1�V1�S�������oG  ���l$0�t$4h�   h�   h�   �u�u�u�u�b����E�D$,�� �l$0���|$0�D$    ��t& �|7
t^�����t$��  ��9�~S���t$8��  P��  P��  P�D$GP�G��P�D7P�����G�� ��9���D$1��f��|$0��l$0�O�t$4j j j jj�t$ Q������ �t$4h�   h�   h�   �ujj �E��P������ �t$4h�   h�   h�   jjj�E��P�Z����� �t$4h�   h�   h�   jj�E��P�E��P�-�����<[^_]Ð�t& U1�WV1�S�h������E  ���|$0�D$    �G���&    f��<0
tN����P�  ��9�~G���t$8j j j �D$ GP�G��P�G�0P������G�� ��9�G��D$1�멍v ��[^_]Í�&    �UWVS�������SE  ���t$ �l$$�F ��~J1���&    ��    �F����    ��R�V(��P�F�U��EF����P�-  ��9~ Ń�[^_]Ð��&    �t& ���  ���D  �D$ǀ     ���(�����T$�P�T$�P�T$�P�T$�PÐ��&    ��&    WVS�|$������ÀD  ��W�M  �T$ ���r=   $��h   j V�L  XZWV�T  ��[^_Ít& ��W�  YZPV��  ���Ő��&    �WVS�t$������D  �|$����<����W��  �FXX�FZWP��  �D$(�F�D$,�F�D$0�F�D$4���F[^_Ít& WVS�t$�)����ðC  �|$�F�N�P��F���|$ ��   Wh�   h�   h�   jRQP������ Wh�   h�   h�   j�F��P�FF��P�F��P�d����� Wh�   h�   h�   �F��Pj�F��P�v�9����� Wh�   h�   h�   �F��Pj�F��P�FF��P������ [^_�Wj`j`j`jRQP������� Wj`j`j`j�F��P�FF��P�F��P������� Wj`j`j`�F��Pj�F��P�v������ Wj`j`j`�o�����t& UWVS�������cB  ���t$0�|$4�F�n�N�P��F���l$���~ ��   ���n\�L$�N�L$����  ����  ����  ��Wh����h�����t$RP�t$ �������j WV������Wj j j �V�������F��P�V����ЋVX��F��)�P�t$(�P����� ��[^_]Ít& ���W��h�   �h�   ��h�   ��QRP�t$ �����V�� W��h�   ��h�   �h�   ���P�R�N�Q�RFP�F��P�N����� Wj`j`j`j�F��P�v�F��P�,����� Wj`j`j`j�F��P�FF��P�F��P������ Wj`j`j`�F��Pj�F��P�v������� Wj`j`j`�F��Pj�F��P�FF��P������ ��[^_]Í�&    ��    ��Wh--��h22���t$RP�t$ �c�����jWV������Wh�   h�   h�   �k�����&    ��&    ���Wh��-�hȠ2�뮃�Wh�77�h�<<��VS�~�����@  ���t$�T$,�V��P�����D$ �F�D$$�F�D$(�F����P�^
  �V�F(�F�V�F ��[^Ít& WVS�t$�����à?  �|$����d����W�^  �F�$�
  �FZYWP�x  �D$(�F�D$,�F�D$0�F�D$4���F[^_Í�&    �t& ��G   ��7?  �D$�@    �@    �@    ��x�����T$�P�T$�P�T$�P�T$�PË$�S�_������>  �� j j j �t$4�D$$Pj�  �D$,��8[�f�S�/����ö>  ��j j j j �t$(j!�z  ��([Í�&    f�S������Æ>  ��j j j �t$(�t$(j�H  ��([Í�&    UWVS�������S>  ��(�l$<U�T����$�   �D$�����+   �T$����1����FjtUPǆ�   ����ǆ�   �����V�-  �}�m����    ���� ��f��� vf��� wd���   ������P�T  �����   ���   ���   ��ǆ�       ǆ�       Ɔ�    Ɔ�    ��[^_]Í�&    ��&    �ȃ���P��  ��롍�&    ��    S������F=  ���D$�p�u�����[��7�����'=  UWVS���l$0�T$�Eu(�����   S�����   �EP�EPj j ������� �E���   ��~?1����   �v 9�v\�M ��t1��v ���	9�u��A�������WP��E��9�̋��   ��t	��S�Ѓ���S�u�\$�������,[^_]Ð�    ��&    f�UWVS���D$0�l$4�|$8�p��~G� 1ۉD$��&    ��&    9�t<�D$��t1�f���� 9�u��@�P�H9�~9�|&��9�uσ�[^_]Í�&    �    ��&    f�H9�~�P9�~̅�t�T$1���&    ����9�u��T$�D$���@�P�R�D$@�����   ��[^_]Í�&    ��&    S���\$���   ��xn;CsY���t1Ґ���	9�u��A���P�R���   ��;Ss-���t1��t& ����	9�u��A��[Í�&    ��&    ��    ��&    f�ǃ�   ������1�[Í�&    ��&    �VS�N������:  ���t$ j�E����T$ ���     �P��@    ��t�V��P�F�F��[^Ív ��F�F��[^Ð�U��S���v  o:  ��h   ����  ���E�}� u�    �%�E�U�P�E�   �E�P�E��@   �E�]���U��S��������:  �E�    ���u��u��  ���E��}� y�    �$���u�u��[������E�}� t�E���    �]���U��S���  �9  �U�R�U���u����  ���    �]���U��S���  {9  �U�R�U�U�U��R�u�u���  ���E��E��]���U��S���B  ;9  �} t,�U�R�U�U�U��R�u�u���  ���E��E�����]���U��S����   �8  �M�U�R���uQR���  ���]���U��S����   �8  �U�R��jj R���v  ���]���U���   �8  �    ]�U���   �8  �    ]�U��S���q   j8  �URjj�UR���������]���U��S��������>8  ���u�	  ���E�E��ujP�u��������E�9�u�    �������]��Ë$�U��������7  ǀ$      ǀ(      ǀ4
     ǀ8
      ���    �B    � ��    �B    �¨��    �B    ǀ,      ǀ0      ǀ4      ǀ8      ǀ<      ǀ@      �]�U����D���=7  �E�    ��U�E�ЋU��E��E�;Er�E��U�������7  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���
����Ñ6  �E���E�E���4
  �E�    ��Ѕ�u��4
  �E�    ���E����4
  �E�    �����E䋃8
  9E�s	��8
  �E���u��  ���E���jj �u���������}� u%��,  ��0  ���� ��,  ��0  �    �l�E��     �E��@    �E��U�P��4
  �E�E��P�E��@   �E��@    �E��@�ƿ    �����P� ��������Q�E��e�[^_]�U��WVS��L�������Y5  �E�    �E�    �E�    �E�    �E�E��E� �X  �}� u5��,  ��0  ���� ��,  ��0  �C  ��j�������  ��$  ��u-���u��9�������$  ��$  ��u�  �    �{  ��$  �E��E�    ��(  ���C  ��(  �P��(  �@)ЉE��E�    �E����    ;E؉�E��
  ��(  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ�(  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u��$  �E��E�    �|  ���u��'������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ����  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ���)  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ���
  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u��$  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������  �    �e�[^_]�U��WVS��,������%.  �} u#��,  ��0  ���� ��,  ��0  �9  �E��� ���E�}�w	�E+E�E�  �E���E��E��@=���tx��4  ��8  ���� ��4  ��8  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��<  ��@  ���� ��<  ��@  �  �  �E��@�E������P� �M��I�ο    )��������Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ��$  9E�u�E܋@��$  ��(  9E�u
ǃ(      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋������P� �M܋I�ο    )��������Q�E܋@��P�u��  ���G��(  ��t=��(  �P��(  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉�(  �  �e�[^_]�U��S�������+  �U�U�U�U��R���%������E��E��Pj �u��-������E��]���U��S���������^+  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E��(  �E���E�E�@=���tz��4  ��8  ���� ��4  ��8  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��<  ��@  ���� ��<  ��@  �  �    �_�E�@�E�E�;Er�E�U�P�  �E�;�  ���u��������E���u��u�u����������u��������E�]���U���� ����)  �E�E���E��P�U��U��E�P��U��u�E��U��� ������)  �E�E��E�E��E�E��"�E��P� �M���Q�E��E��m�E�E�}�w؋E�E���E���E���E��E��m�E�E��}�wދE�E���U��E�ЋM��U��� ��m�E�E�}� uۋE��U���� ���)  �E�    ��E��U��E�� ��u�E���U��S���`������(  �E�    �E�    ��U�EЋM�U�� ��E����u������9E�|ԋU�E��  �E�]���U��������(  �E�    ��U��EЋM��U�� ��E��E�9EwߋU��E��  ���U��S��������>(  ���u�	������EЃ��uP�$������E�]���U������(  ��E�P�U� ��u�    ��E� �U8�u܋E]�U���������'  �E�    �(�E� �U8�u�E�E��E�P�U� ��u�E���E� ��u΋E��U��S���������x'  �E�    ��E��E� ��t"�E�P�U� ����P�u�4�������uЋE�]���U��S��������%'  �E�    �)�E� ����P�u���������t�E���E�E��E� ��u͋E�]���U��VS�J������&  �} t�E��D  ���D  ��u
�    �   ��D  ��D  ���uP�
�������E���u�u�G������EЉ�D  ��D  9EuǃD      ��D  �/��D  � ��t��D  �  ��D  ����    ��D  �E�e�[^]�U������&  ��E�E�E��E� 8�u
�E� ��uދE� �ЋE� ��)�]�U���������%  �E�    ��E��E�E�E��E� 8�u�E� ��t�E�9EwҋE� �ЋE� ��)���U��VS�������c%  ��E�E�E� ����P�\  ���ƋE� ����P�E  ��9�u
�E� ��u��E� �ЋE� ��)Ѝe�[^]�U��VS���h������$  �E�    ��E��E�E�E� ����P��  ���ƋE� ����P��  ��9�u�E� ��t�E�9Ew��E� �ЋE� ��)Ѝe�[^]�U��S���������i$  ���u�4���������P��������E���u����������Pj �u�� ��������u�u�� �������]���U��S�������#  �M�U��j j j QRj���  �� �E�]���U��S��������#  �U��j j j j Rj���  �� ��]���U��S�������#  �]�M�U��j S�uQRj���T  �� �E�]���U��S���d���]#  �]�M�U��j S�uQRj���  �� �E�]���U��S���+���$#  �]�M�U��j SQ�uRj����  �� �E�]���U��S��������"  �]�M�U��j S�uQRj���  �� �E�]���U��S�������"  ���u�u�u����������]���U��S�������"  ���u�u�u���������]���U��S���a���Z"  ���u�u�u���������]���U��S���5���."  ���u�u���������]���U��S������"  ���u���������    �]���U��S���S������!  ��j �u�������E�}� t���u���������    ��   �]���U��S�������!  �M�U��j j j QRj���Q   �� �E�]���U��S���a���Z!  �U�U�U�U��U�U��j �u��u��u��uj���	   �� ��]���U��WVS����!  �E�]�M�U�u�}�i�[^_]�U��S��������   ��j j j j j j�������� ���U��������   �}/~�}9~�}`~�}z~�}@~�}Z�   ��    ]�U�������   �}`~�}f~�}@~�}F�   ��    ]�U���V���O   �}z����]�U���=���6   �}@����]�U���$���   �}/~�}9�   ��    ]�U��������  �}/~�}9~�}`~�}f~�}@~�}F�   ��    ]�U��������  �E�E����U�������  �E��!��]����]�U�������  �} t�}	u�   ��    ]�U���`���Y  �]�U���P���I  �]�U��S��������5  ���u�~�������t���u�I�������u�   ��    �]���U��������  �E��_]�U��������  �E�� ]�U��������  �    ]�U�������  �����  �    ]�U��S�������  �M�U��j j j QRj���T����� �E�]���U���h���a  �    ]�f�f�f�f�������t6U��S������&    �v �Ѓ�����u��[]Í�&    ��&    ��ʾ���     / r /file.bmp /binfile.bmp /folder.bmp          Ї�8�       zR |�        ����)    A�Be�     <   ����>    A�Bz�     \   ����    A�B�� (   |   �����   A�BB����A�A�       �   ����   A�BG���(   �   {���z   D Gu Eutu|ux    �   ����U    A�BQ�      ����(    A�Bd�     8  ����    A�BV�  |   X  ����~    A�A�A�A�N U$A(A,D0H E$K(A,D0H G
A�A�A�A�CC$C(A,G0H CA�A�A�A�     �  ����?    Cy 8   �  �����    A�A�A�A�C$�A�A�A�A�8   ,  ����.    A�A�NFB B$B(A,B0HC�A� 8   h  |����    A�A�A�A�C�A�A�A�A�8   �  ����    A�A�A�A�C�A�A�A�A�<   �  ����b   A�A�A�A�NPL@�A�A�A�A�X      �����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   |  H����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H   �  �����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   $   ����    A�A�A�A�C(�A�A�A�A�   `  ����           t  ����(    A�SJ HA�     �  ����    A�ND HA�     �  ����    A�ND HA�     �  ����    A�ND HA�       ����    A�ND HA�     (  ����    A�ND HA�   L  ����W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   `  ���s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�     �  <���          �  8���          �  4���	          �  0���	            ,���	       �     (���{   A�A�C�C�N0H4E8E<E@CDCHCLCPO0e<D@H0G4D8H<H@HDHHILFPK0c4B8B<B@BDBHDLAPH0D4E8E<E@CDBHBLGPH0D4E8E<E@BDBHBLGPH0D4E8E<E@BDBHGLGPHA�A�A�A� \      �����    A�C�A�C�N0f<A@H0G4D8B<B@BDHHILHPK0YA�A�A�A� H   `  ���s    A�A�A�A�N d$K(G,V0H HA�A�A�A�     �  8���A       d   �  t���g    A�A�A�RA LMEBA FAAA HA
�A�A�ECA FAAA H@   (	  |���\    A�A�A�VL IDAA aD�A�A�   �   l	  ����K   A�A�A�nEEE B$A(A,A0HAEEE B$G(J,G0HAEEE G$B(G,C0HAEEE G$B(G,J0HA
�A�A�AABBB B$A(A,A0HABBB B$G(J,G0HABBB G$B(G,C0HABBB �  d
  ����`   A�A�A�A�N0Z4A8E<E@DDAHALDPH4B8A<A@H4A8B<B@BDSHXLDPH0C
A�A�A�A�FC4H8G<G@DDAHALDPK0A4G8H<G@FDGHDLGPH0A4B8B<B@BDGHCLGPH0A4B8B<B@BDGHJLGPH0A4B8B<B@GDBHGLCPH0A4B8B<B@GDBHGLJPH0C
A�A�A�A�NC4A8E<E@DDAHALDPH4B8A<A@H4A8E<E@EDT0C
4A8E<E@BC4A8E<E@ (   �  ����\    A�A�Nr WA�A�@     ����d    A�A�A�VL TAAA aD�A�A�      \  (���L          p  `���       0   �  P���.    A�N(B,B0B4D8E<B@LA�  0   �  L���'    A�NBB B$B(D,B0HA�  0   �  H���)    A�NBB B$D(D,B0HA�  `      D���   A�A�A�A�N<E@a4M8A<A@g0g<G@H0y
A�A�A�A�OE<D@H0      �  ����     A�NG HA� x   �  �����    L�A�A�A�C0Q8G<H@EDEHBLBPH0w8H<A@H0Q<A@E0C8A<C@LA�A�A�A�B0����X   $  @����    A�A�A�A�C0]
A�A�A�A�HD<F@J0IA�A�A�A�0   �  �����    A�CkC La
A�P]C� <   �  0���_    A�A�NF Lh
A�A�DLA�A�       �  Q���]    A�BD�U��       ����c    A�BD�[��     <  ����4    A�BD�l��      `  ����@    A�BD�x��      �  ����J    A�BD�B��     �  ���1    A�BD�i��      �  (���.    A�BD�f��     �  2���    A�BP�       &���    A�BP�      0  ���,    A�BD�d��      T  "���Q    A�BD�I��    x  O���          �  ?����    A�B��    �  ����7    A�Bs�     �  ����r    A�Bn� ,   �  5���8   A�BF���+�A�A�A�   ,     =���4   A�BF���'�A�A�A�   ,   L  A���~   A�BF���q�A�A�A�       |  ����K    A�BD�C��     �  ����f   A�BD�^��   �  ����8    A�Bt�     �  ����    A�B��      ����1    A�Bm�      $  ����a    A�BD�Y��    H  ����H    A�BD�     h  ���>    A�BD�v��     �  (���8    A�Bt�     �  @���P    A�BL�     �  p���S    A�BD�K��     �  ����V    A�BD�N�� $     �����    A�BB����A�A�   <  o���I    A�BE�    \  ����_    A�B[� $   |  ����q    A�BB��i�A�A�$   �   ����    A�BE��|�A�A�    �  ���k    A�BD�c��     �  ����6    A�BD�n��        ����2    A�BD�j��      8  ����9    A�BD�q��      \  ����9    A�BD�q��      �  ���9    A�BD�q��      �  %���9    A�BD�q��      �  :���,    A�BD�d��      �  B���,    A�BD�d��        J���,    A�BD�d��      4  R���)    A�BD�a��      X  W���+    A�BD�c��      |  ^���J    A�BD�B��     �  ����6    A�BD�n��      �  ����F    A�BD�~��  (   �  ����*    A�BC���`�A�A�A�      ����-    A�BD�   0  ����?    A�B{�     P  ����3    A�Bo�     p  ����    A�BU�     �  ����    A�BU�     �  ����'    A�Bc�     �  ����?    A�B{�     �  ���    A�BU�       
���    A�BZ�     0  ���'    A�Bc�     P  ���    A�BL�     p  ����    A�BL�      �  ����G    A�BD���     �  ���    A�BQ�     �  ���    A�BQ�     �  ����    A�BP�       ����    A�BY�      4  ����6    A�BD�n��     X  ����    A�BP�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������    ����            ��ИИ        ���И         �� �        0�ИИ        ��ИИ        ��ИИ                                                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              �                           >        ��    src/gfx/sse2.asm NASM 2.14.02 ��     %  . @   :    '   �       src/gfx/sse2.asm      �                                         t�          ��          ��          ��          ��           �          �          �          �     	     ��     
     ��          ��                                                                                                                                  ��   �         �      (   ��      ;   ��      =    �      P   P�      f   ��     u   ��     �   Ё      �   ��                 ���   �      �   <�      �   @�      �            ��  ��                  ��  ��(     F  ��     d           ��q           ��}           ���           ���           ���           ���           ���           ���           ���  ��     �  ��     �  ��     �  ��     �  ��     �  ��       ��       D�7     *  {�r     :  �8    L  %�4    `           ��i           ��r  ��     y           ���           ���           ���           ���           ���           ��             ���  ��     
 �  ��     �  ��a     �  ��.     �  ���       ��     E  ��.     d  Ї�  "  �   �`    �  ��     �  С'     �  l�*     �  ���     �  ��     �  �6     �  ��     �  �(   "  �  �9       +�       ���    :  ��A     3  ���     N  p�\     c  ��     k  ��     w  &�F     �  �     �  ��6     �  5�     �  ��     �  �     �  `��     �  %�4    �   �t     �  ��     �  ��     �  K�G       �{    !  �'     )  �     0  МK    Y  <�   ! 	 e  &�,     k  �     n  `�   "  u  (�   ! 	 �  ���     �  ��     �  0��     �  ��U   "  �  ��?     �  t�      �  ��     �  ��>   "    �	     /  І)   "  C  ��P     K  p�\     `  ״K     �  ��,     g  �     x  ��~     �  ���     �  B�>     �  �    �  ��1     �  #�9     �  ��W    �  І)   "    И        �     �  ��&     $  �     1  x�   ! 	   ν,     G  ��A     [  N�     c  ��_     k  ��_     �  ��6     �  0�s     �  ��   "  �  ��H     �  �q     �  "�f    �  ���     �  ���       �       0�    5  �]     <  P�b    _  ���     {  @�      �  �3     �  �   ! 	 �  @�s     �  �@     �  �k     �  n�c     �  ��      �  ���     #  ��8     	  �z    	  ��.     	  ��     %	  p�?     /	  P�   ! 	 U   �     ;	  ��   "  B	  P�L     _	  Ѧ4     f	  ��     n	  ÿ?     v	  ;�     ~	  w�I     �	  ��\     �	  ��   !  �	  ��      �	   �g     �	  [�V     �	   �)     �	  ��     
  #�     
  ��\     '
  �,     -
  @�   "  3
  8��   "  O
  И     f
  g�'     n
  E�J     u
  ��J     |
  ��      �
  ��      �
  �d     �
  ��     �
  \�9     �
  ��-     �
   �	     �
  ��     �
  `��     	  �S       h�1     �  R�)       ��       ��2     +  �d     ?  ��8     F  B�Q     L  ��     U  d�   ! 	 `  ��	     {  ��   "  �  ��9     �  �      %  {�+     �  ��>   "  �  ��     
  Y�~    �  P�L      crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_fileIconBuffer graphics.cpp runtime.cpp text.cpp widgets.cpp window.cpp font.cpp src/gfx/sse2.asm fileio.c l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 memory.c string.c p.1056 filesystem.c ipc.c syscall.c exit.c ctype.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated strcpy _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN15ScrollContainer5PaintEP7Surface _Z13_CreateWindowP10win_info_t _ZN10FileButton5PaintEP7Surface _ZN6Button5PaintEP7Surface l_max_inuse _Z14_DestroyWindowPv syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm lemon_read isblank _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN7TextBoxC2E4Rect _ZN6ButtonC1EPc4Rect l_inuse __TMC_END__ SendMessage __DTOR_END__ lemon_open islower tolower feof _Z11PaintWindowP6Window malloc windowInfo __x86.get_pc_thunk.ax __dso_handle ispunct _ZN7TextBox5PaintEP7Surface isspace fflush _ZN6Button17DrawButtonBordersEP7Surfaceb _ZTV6Button lseek fd _ZdlPv _ZTV7TextBox strncasecmp __x86.get_pc_thunk.dx _Z15HandleMouseDownP6Window8Vector2i _ZN4ListIP6WidgetE5clearEv isxdigit liballoc_lock _ZN10FileButtonC2EPc4Rect _ZN6Button11OnMouseDownEv _ZN10win_info_tC2Ev strrchr _ZN6ButtonC2EPc4Rect calloc folderIconBuffer _Z16memcpy_optimizedPvS_m _ZN5Label5PaintEP7Surface strcat _Z12RefreshFilesv fseek lemon_write _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev _ZN6Widget11OnMouseDownEv win exIconBuffer _ZTV15ScrollContainer _ZN7TextBoxC1E4Rect isupper strncmp _Z9AddWidgetP6WidgetP6Window liballoc_alloc _ZN6Bitmap5PaintEP7Surface _ZdlPvm strncpy strcasecmp realloc _Z8DrawRectiiii10RGBAColourP7Surface strtok __x86.get_pc_thunk.bx _Z12CreateWindowP10win_info_t fdopen _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window isalpha _ZTV6Widget _Z10DrawStringPcjjhhhP7Surface fread strdup fopen __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface main ftell font_default _Z5floord _ZTV6Bitmap _ZdaPv _ZN15ScrollContainerC2E4Rect fclose isgraph isalnum isprint strcmp _ZN6BitmapC1E4Rect _ZTV10FileButton _fini _ZN7TextBox8LoadTextEPc strcspn _Z12_PaintWindowPvP7Surface _ZN6Widget5PaintEP7Surface liballoc_free _ZN6BitmapC2E4Rect fputc _Znam _ZN10FileButton9OnMouseUpEv _ZN6Widget9OnMouseUpEv isdigit fwrite access _edata _end _ZN5LabelC2EPc4Rect _Z13HandleMouseUpP6Window lemon_seek exit _ZN6Button9OnMouseUpEv iscntrl _Z10surfacecpyP7SurfaceS0_8Vector2i strspn strlen toupper lemon_close _ZN5LabelC1EPc4Rect strchr fputs font_old _ZTV5Label _ZN7TextBox11OnMouseDownEv _ZdaPvm lemon_readdir memcpy_sse2 _ZN10FileButtonC1EPc4Rect _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN15ScrollContainerC1E4Rect  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .data.rel.ro .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                   t�t                     !         ���   �A                 '         ���B                    -         ���B  <                  5         ���B  x                 ?          � `                   K         �`                    R         �`                    Y         �`  x                  f         ���`                   o         ���`  (
                  u         ���j  �                   z      0       �j  +                 �              �j                     �              k                    �              %k  B                  �              gk                    �              �k  >                  �              �k                    �              �k                                  �k  `     H         	              4z                                 7�  �                  