ELF          >     @     @       ��=         @ 8  @                   @       @     d�     d�                   �      �K      �K            �                    �      �K      �K                           �C  �+ �             H��    UH���������  ��+ H��   �i���f.�     � �K H= �K t�    H��t	� �K ��f��ff.�     @ � �K H�� �K H��H��H��?H�H��t�    H��t� �K ���ff.�     @ �=y�  uwUH�w� H��ATA�(�K S�0�K H��(�K H��H��H9�s%f.�     H��H�=� A��H�2� H9�r��0����    H��t
��J �����[A\�� ]��ff.�     @ �    H��tU�@�K ��J H������]����D  ����UH��H��   H�E�A�    A�    �    �    H�ƿ   �nS �E��� �E�    �0�K ��  9E�������   �E� �E�    �`� 9E�}kH��`���H���^  �E�Hc�H��`���A�    A�    �    H�ƿ   ��R H�E�H�E�E��ƿ0�K �  H� H9E�����t�E���E���E�����t�E��ƿ0�K �|  ��� �E��=������UH��H��   H�E�A�    A�    �    �    H�ƿ   �fR �E܉�� �E�    �{� 9E���  �E� H��`���H���q  �E�Hc�H��`���A�    A�    �    H�ƿ   �	R H�E�H�E��E�    �0�K �  9E�����t)�E�ƿ0�K �  H� H9E�����t�E���E����E�������   ��   �v H�E�H�E�H��`���H��h���H�PH�HH��p���H��x���H�PH�H H�U�H�M�H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�U؉��   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�E�H�ƿ0�K ��  ��� �E��c������UH��AVAUATSH��   H�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸��K A�    A�    H�ƿ   �]P �Y  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H���  H��P���H�E��@����H��X���H�    ����H!�H	�H��X���H��X�����H�       H	�H��X���H��P���H��X���H��H��H�й��K ��H��H���/E �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H���L  H��`���H��h���H�    ����H!�H��H��h���H�E��@������H�� H��h�����H	�H��h���H��`���H��h���H��H��H�й��K ��H��H���uD �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H���  H��p���H�E��@������H��x���H�    ����H!�H	�H��x���H��x�����H�       H	�H��x���H��p���H��x���H��H��H�й��K ��H��H���C �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H���  H�E�H�U�H�    ����H!�H��H�E�H�E��@������H�� H�U���H	�H�E�H�E�H�U�H��H��H�й��K ��H��H����B A�    A�*�2   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H����  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A���K D���H��H���F H�E����   ����H�E����   ����H�E�H��H��h��K A��   A��   ��   H����K H���E�   �E�   H�E�H���   H�E�H��H���   H�E�H�E�H�U�H����K A�    A�    H���   ��K H�e�[A\A]A^]�UH��H���   ���K ��< H�Y� H�R� H��H��H�L� H��K� �H�E� f�HH���@ H��H�E�H�E�H�H�HH�+� H�,� H�PH�HH�%� H�&� H�@ H�#� �� �� ��H�H���.p H��� H�E؋PH�E؋@�u�h�   A�    A��   �щ¾    �    ��? H��A�    A�    �    �    �    �   ��J � -H �-H �� H�E�H�Eк   �    H���O� H�H�E�H�Eк    �    H���3� H�E�H�H���uo H�E�H�u�H�U�H�E�H�Ѻ   H���$$ H�Eȋ@��H��H��H�H��H��H�E�H�H�E��J�    �D�    ��  �o H�?� �-� �#� H�M�A� �K I�ȉщ¾    �    �? �-H A�    A�    �    �    H�ƿ   ��I �    �-H ��: �E��E��   ���K ���; ���K �3  ������t(�#-H A�    A�    �    �    H�ƿ    �oI H�K� ���K �    �?-H H���ı  �E��}� t(�E�H��P-H A�    A�    �    H�¿    � I H�� �   �    H���Z9  H��� �A   H���&=  �E��M�H��� �    ��H����S  ��� ��t,�u� �k� A���K D��� �щ¾    �    �> �E�    ��� 9E�}%�E��ƿ0�K �.  H�E�H�E�H�������E����M�  �E��   ���K ����9 �+� �� ��Љ� �� ��� ��)Љ� ��� ����   ��� ��� ��� H�>� )щʉ��   ��� ��� H�!� )щʉ��   H�� ���   ��yH��� ǀ�       H��� ���   ��yH��� ǀ�       �L� �������#  �:� �����  �(� �0�K ��  ���E��}� ��  �E��ƿ0�K ��  H�E��
� H�E����   9���  ��� H�E����   H�E��@���9���  ��� H�E����   9��  ��� H�E����   H�E��@���9��Z  �E��ƿ0�K �u  H�ƿ0�K �  H�E�H��� �p� H�E����   �P�Y� 9�|LH�E��@����u>�=� H�E����   )/� H�E����   )��ȉ� �� ��� ��   H�E�   H�E��@����t0��� H�E����   )ЉE��� H�E����   )ЉE��4��� H�E����   )Ѓ��E��� H�E����   )Ѓ��E��E�H�� H�E�H	�H�E�H�E�H�@|H�E�H�E�H�@tH���u��u��u���x�����p���H���A H��0�	�m������� ����t�
� ��t���  ��� ����  ��� ��������  ���  ���  H�B� H����  ��� H�,� ���   9���  ��� H�� ���   H�� �@���9��h  ��� H��� ���   9��M  �n� H��� ���   H��� �@���9��"  �F� H��� ���   �P�,� 9�|H��� �@������   H�p� H����   H�E�   H�X� �@����t6��� H�A� ���   )ЉE��� H�'� ���   )ЉE��:��� H�� ���   )Ѓ��E��� H��� ���   )Ѓ��E�E�H�� H�E�H	�H�E�H��� H�@|H�E�H��� H�@tH���u��u��u���x�����p���H����> H��0H��@���H���> H�������  H��P���H=�  ��   H=� u�H�L� H����   H��X���H����   H��X���H��H��t0H��X�����H��t!H�E�   H��X���������K H�H�E��H�E�   H��X�������K H�H�E�H��� H�@|H�E�H��� H�@tH���u��u��u���x�����p���H���> H��0�(H��X���H��u�����H��X���H��u������������������5�� �� h��K j A�    A��   �   �   ���6 H���E�    �}��E�    �}��E���E���A� �?� ������H�\� H�E�H�@H��H���5 �5o� �e� A���K D�a� �   �   ����6 ����UH��H���}��u��}�u'�}���  u�0�K �   ���K �0�K �t@ �(D ���UH����  �   ����]�UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]�UH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H��H�}��u�U�H�E���H���   ��UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H����b H�E��ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �: H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H�� H�}�H�E�H� H�E�H�E�@��tH�E�    H���'�������@ U��@H H��S��-H H��D  H��H�����  H�3H��u�H��[]�ff.�     f�USH���-H H��  �y� H���A  ����6  fD  �� �7  ��	�.  H��1��$�    ��:t"�H��H��H���   �  �Hc���u��< �>:��   H9���   H��1�H���(�     ��=t%���   H��H��H=�   ��   �Hc���u�Ƅ<�    �9=��   H9��|   H��1�H���!���	t'��   H��H��H=�   �|   �U Hc����u�Ƅ4    �E ��t<	u0H9�t+H��$   H��$�   H��H���>  �UH�E�������H�ĸ  []�fD  H���� ��   �������   �>�����   �ff.�     f�AUATI��USH��� H��tiL��H��H���;u  A�Ņ�uDI�,$��-H ��@H fD  H��H����  H�3H��u�I�<$����H��D��[]A\A]�D  H���h ��fD  H��A�   [D��]A\A]�ff.�     �H��tSH��2>  H���* 1�[�fD  �!   �f.�     H�71�H���t# H��H��H��H)�H�
H���u��D  �ff.�     @ Hc��H��H��H)���H�H��H��H)�H��H��H��H����H�H��H��H)�H����H���     �9����     ATUH��SH��L�f H�|$H�|$�V�M1�H��I���     H�;H��t'H�t$�U��uH��I9�v�E��I��H�;H��u�H��H��[]A\�D  ATI��UH��SH�FH��H��tH����I�D$H�@xH��tH����H�sPH�EH��t	H����H�EH�CP    H��H��[]A\���     H�wPH��t\HcGHH��H��@ H��H9�w;H��zcinuu�D�BA�� 
 t	A��   u�H���   1�� H��xcinutH��H9�v�&   �D  H���   1��fD  SH�7H��H��t
H�G8H���PH�    H�C    H�C0    [ÐH���   HcNH��H��H��?H�� �  H���   H��H��H��?H���H�FH��H��?H�� �  H�����H�H�F H���   H��H�H�� �  HcVH��H�� H���H�F(H���   H��H�H�� �  H��H�� H���H�F0��     ������f9|�����ff.�     �H�6H�?�8t1��H���E� ����H���ff.�     f�H�H�USH��  ��|�   f.�     L��H��H��  Z I��H��H��  ��|�H��1���� A�   � f�H��L)�M�H)�M�H��t4H�,� 0H �HO�M�I��I��H��y�H��L�M)�H�M�H��u�H�[L�]�H��  - �&f�H��H��H��  Z H��H��H��  - �I���k���H��I���`����L�H�USL��H��I9���   H9���   I�ӻ  Z H��1���� A�   �$fD  H��M�L)�H�M�H��t4H�,� 0H �HN�O�I��I��H���H��M)�L�H)�M�H��u�H��xQH��L�H���H�[]�1�H9�}�H��H��  ��L��H��I���l����H�һ  � H��  L�I��HN�H���M���f��   L�H)�H��H���H��H�[]�D  L�L��   D��D����M��AI���M��AI�	��҃�)эB�����I��I��L�L��@ �   )�I��I��L�L��@ H���  H��A��H����A���   H����   AWE��AVL�wAUI��ATI��USH��H���GD�L$I�,�I9�r�&�    I��L9�vI�H��H� H�x�s� ��u�L9���   I�>H�H�@@H��tB�8.H ��H��t6E��t(H� H��t)I�>�L$H��L��[L��]A\A]A^A_��f�H�@H��u'�   H��[]A\A]A^A_� �   �f.�     I�>H��L��L��[]A\A]A^A_���    �!   �f.�     �   �f�     H�H����   H�x(��HDx ��t`�B��    H�T��#D  H��H��xGH�� H��H��H�F�H9�t.H�H��y�H��H��x�I��I)�L��H��H��H��H�F�H9�u�1�ÐI��I)�L��H���ݐ�$   �f.�     SL�^A�ҋFM�م�t&H�9��8��8I��L�@$L��I��?H��H��I��M)�H�^�FI�؅�t&H�9��8��8H��H�p$H��H��?H��H��I��I)�M��uwH��ME�I�� I�� I���I���tTM��tO�G8��~HH�w@�P�1�H��� H��H�FH�� H���I9�uH�H�� H���L9�t,E��u'H�GH�� H9�uʸ   [� H��MD���    1�H��t�H�9[�ff.�     �L�WfE��teH�GI��H�8H�HI�H��I��I��I9�v0@ H�H9�HO�I9�LL�H�PH9�HO�I9�LL�H��I9�w�H�>L�NH�NL�F�@ E1�E1�1�1�H�>L�NH�NL�F�fD  HcHcWSHcLcNLcFH��L��L��HcNH��H��?H��M��H�� �  I��?M��[H��I��?Hc�K�� �  H��H��H��?H�H�H�K�� �  H��Hc�H��1 �  H��H�H�H�G�@ ATUSH�oH�_H��H�H9�s I��@ H��tL��H���@���H��H9�w�[]A\�f�AWI��AVAUATUSH��(H������H�$H�D$H9��6  H�t$H�T$H9��#  ��A�   I�k��H��E��Hǉ���H��H�	�1�����A)�DH�)���A���A)�DH�f����   I�C��L�m1�L�XM�$S1�D  H�D��H��H��H�H�0L�pH��D��I��9�|UA��Hc�A)�H��I�H��I��H�M�fD  H�D��L�xH��H��D��I��H�L��M)�I��I��H�H��I9�u΍SL��M9�tI���r���f.�     �   H�������H��([]A\A]A^A_�H��(�   []A\A]A^A_�ff.�     SH��H�wH�[�� H�G    �����[H�H��H��H�H�GH��H��H�G�@ AWAVI��AUATI��USH���GHH�wP��~T1��    H�,�L�,�    H�E L���   H�EH�@H��tH����H��L��H��A�WI�t$PJ�.    A9\$H�H��tL��A�VI�D$P    A�D$H    H��[]A\A]A^A_�H�GH�F    H�H��tH�pH�w� H�7H�w��     H�H�VH��tH�PH��tH���    H�H��u�H�G� AWI��AVAUATUSH��H�H��t6I��H��I��fD  L�cM��tH�sL��H��A��H��H��L���UM��u�I�    I�G    H��[]A\A]A^A_� H��H��H��?H��8�  f1��f.�     H����  f1��D  H��f1��f�     I��I�й   H��yH�߹����H��yH����I��H��yH����I�и���M��tI��L��1�H��H�I��H��H�ڃ��HD��@ I��I�й   H��yH�߹����H��yH����I��H��yH����I�и���M��tH��1�I��I��H��H�ڃ��HD��f.�     Hc�Hc�H��H��H��?H�� �  H��H��H��A�   H��y	H��A�����H��y	H��A��H�ٸ���H��tH��H��1�H��H�H��H��H��A���HD��H���G  H���>  LcHcNAWAVAUATLcfUHcnSLcLcOHcWL��M��M��L��I��L��M��L��L��I��?I��H��?I��O��* �  H�D$�I��?M��I��I��?L��J��; �  Mc�H��?O��3 �  H��I��H�D$�I��HcGHc�Mc�I��?H��L�J��" �  H��H�H�\$�H��Hc�H��M�� �  H�\$�H��?H��I��H��?M�� �  H��9 �  [H��( �  I��H��Mc�H��Mc�Hc�M�H�L�]L�NH�A\A]H�NA^A_H�F��    �ff.�     @ H����  L�GH�7L�OH�WIc�Hc�H��Lc�Ic�I��I��I��I��?I��?J�� �  N�� �  H���   I��Hc�Mc�L)���   I��H����   H��H����  I��I��J�1�H��H��H�GM����   I��1�K�I��I��H����   H��H�GM���a  I��1�K�I��H�H���0  H��1�J�I��H�G1��@ ��    H��H��H����   I��I��J�1�H��H�GM���r���I��L��1�L)�I��I��H��y?L��H��H�GM��y=I��L��1�L)�I���2  f.�     I��L��1�L)�H��I��L�OM����   I��1�K�I��H���/���H��H�H����   H��1�J�I��H��yH��H�G1��I��M��I��J�1�I��H��H�GM�������I��L��1�L)�I��I���:����    H��L��1�H)�I����    I��L��1�L)�I���i���@ H��L��1�H)�I��H���n���H�G1�ÐI��I��M��I��J�1�I������fD  I��L��1�L)�I��H������H�H������H��L��1�H)�I�������     �   �f.�     H���  H���  AWI��H��AVI��AUATUSH��H��(L�H�/L��H��L�L$�]���L�sM�cL��H�$L��L���C���H��M�{L��H�D$L���,���L��M�kL��H��L������L�sL�L$L��H�D$L��L�������H�[L��L��H�D$H�������L��L��L��H�D$ �����L��H��L��I�������Hl$L�$$H�T$Ld$I�I�kHT$ M�#I�SM�sH��([]A\A]A^A_��    �ff.�     @ H��t{H��tvAVI��H��AUI��ATUSH�/H��H�6H���C���L�kI�sL��I��L���-���H��I�sL��I��M�����L��I�sL��H������L�#H�H�k[]A\A]A^� �ff.�     @ H�H�WA�   A�ɉЅ�y	A��A�����A�   ��y
��A�������E���T  ���<  AUATUSA9��U  ����D��ھ����A��1����A��H��I9�@�Ń�A)�E���@  D��A����A9��  D����¹   )�f�     A�ȉ�E����A����E��D��A��A��D��A�A���  AI�D��   A����	��A�Յ�D����  DI�A��D����  �D��H��H��A���HD�H���H��H��A���HD�E����H�WD�D����  AH���   E���~   A�L$��   []��D��A\A]����@ A��D��Mc�L��f���tA��Mc�L�_���    D���������@ ����D������@ ��)�A������������     ��)�[]��A\A]� H��1�H��H)�H����H��?)��fD  I��H�L�I��?L1�L)�I��I��?L1�L)�H9���   H�4vH��H�H��H��?H1�H)�H��H��?H1�H)�H9�~kH�IH��H�H�H1�I��L��H��?I)�I1�I)�M9�~#K�@H��L�H�H)�H��H9������@ K�IH��L��� H�<H��H��v���H�RH��H�� �oO(H�GX�G    �GP    �oG�oW8�o_HOpG`��   ��   H���   �ff.�     �USH��H��H�w H�/H��tH���UH�s(H�C     H��tH���UH�s0H�C(    H��tH���UH�s@H�C0    H��tH���UH�sXH�C@    H��tH���UH�CH    �oK(�C    �oS8�CP    �oC�o[HH�CX    H�C    �C    C`Kp��   ��   Hǃ�       H��[]�USH��H��H�/����H��H�EH��H��[]��ff.�     f�H��t��f�     �ff.�     @ H�GH�O �G`    Ǉ�       H��HG(H��H�GpH�G0Hр H�OhH�OH�HH�GxtH�G@H�HWHH���   H���   �GPH�@H��HGXH���   �f�     H��tS�O�Wb�G`fG�f�W���   WPf��~&H�Wx�p�H�BH�4p�
fD  H��f
H��H9�u��,���@ ��    H��tsAUI��ATUH��SH���GH�_ ��t2��L�d��     H�3H��tH���UH�    H��L9�u�I�] H��t	H��H���UI�E     H��[]A\A]�D  ��    H������H�H��H�B�    HD�H���ff.�     @ H�����e���H�H��H�B�    HD�H���ff.�     f�H��tSUH��SH��H��t5H��H�?H��u�(H��H�;H��tH���� ��u�H�CH��[]�D  H��1�[]��    1��D  H�w@H�WH�OP�GT    �ff.�     f�������f.�     H���wT�   ��4 ff.�     @ H��t;ATU��SH�G0H��L�g8H��t�Ѕ�uI�D$H��L��[]A\��fD  []A\� �ff.�     @ H��(  H��tL�P��tDSH���   H��H��tH�GH���   H���PH��(  �PHǃ�       ����P[�fD  HǇ�       �ff.�     �ATUSH�GH��H���   H�EL�eH���   H��t��H���`���H��(  H��tH�E H� ��tL��A�T$Hǃ(      []A\�H�>H��t����H��(  H�    �� AVAUATUSH��H���   H�� H��(  H��t
�@��   H���  H�*L�ZA��H����   L�4$L�T$L�l$L�L$I�.K�4I�D- K�H�$H�t$H�D$H�T$A����   A���  A�   �   A���8  H��?H��?H���H���H���H���I��I��H)�H)�I��I��H��H�����K  ���Z  H����tj�   D���   D���   D���   f���   ���   ���   ���   H�� []A\A]A^�f.�     H����������� E1�1������fD  H�HH��H�� H�t$H��H��耒  H�$H�t$A�   H�D$H�T$�   ����D  H�t$H�|$H���F�  H�$H�t$A�   H�D$H�T$�   ����� M)�I��?��   H��?H���H���H�$H�D$M)�I��?MH���H��?H���H�$H�D$A�   �   ����H�@H�HH��������    H�RH������@ H�� H�� H����f.�     H�� H�� H���H���H�$H�D$�t���f�UH��SH��H���o���H���   H��[]ÐH���   USH��H�WH���   H���   H�hH��t"H�AH9�u�T H�PH9�tH��H��H��u�H��[]�D  H�QH�G(H��H��t��H���^���H�EH��H��H��[]��@ �H���   ��ff.�      AVAUI��ATUH��SH���   H��L�bH��tH���   ���	@ �+���H���   H��u�H��tH���   L��H��p@ �s���Hǃ�       H�C`H��tH����H��H���O���I�D$hH��tH����L���   M��t!I�D$0L�kM�t$8H��tL����A��   tCH���   H�EHǃ�       H��tH����H�EHǃ�       H��H��[]A\A]A^��@ L��L��A�V�@ H��tNH���   �@0    H��t@�o �oNHH�NHNtH�@0   H��tR�oP H�JH
t�H0�@ H�    H��H�@    H�@    H�@   H�>   u�H�~   u�몐H�@     H�@(    �ff.�     @ H��tH���   �@x1��D  �#   �f�H����   ATUSH���   H��twH���   �Px�J��Hx1���~	[]A\�@ H�M H��u�MD  H�IH��t?H;yu�L�eH��H��H�} �V���L��A�T$H��H��L������[1�]A\�f�     [�#   ]A\�fD  �#   �f.�     H����   AUATUSH��H�/H����   L���   M����   H���   H��u�[ H�IH��tOH;yu�M�l$H��H��H���   ����L��A�UH9��   t:L��H��L���\���1�H��[]A\A]��    H���$   []A\A]��     H���   Hǅ�       H��t�H�@H���   �@ �$   �f��#   �f�     �"   �f�     �Gt���u�������@ �#   �f��   �f.�     H�WH�GI��I)�H��y
H9�HM�I��H��u&H�gfffffffK�@H��H��H��?H��H��H��H)�H�W H�OH�w8H��H��?H�H��H��L)�H)�H��H��?H�O(H�H��H�G0�H��Hw@H���   H�VL�NL�B I��fD�AM�A I��fD�A�G��   ���   H��xIH����   H��H��H��H�1�H��H�A M����   H��I��1�H��L�H��H�qH�A(����f�H��  �H��tH��H��H��H)�1�H��H��H�A M��xv����H��t^�f.�     �H�A    H�A(   ��L�I0H�H�A8    H�A@H�QH� L��H�A ���H�   ����H��?H!�H���H�A(H�q�����H��  �H��t�H��I��1�H��L)�H��H�qH��H�A(�����f�AUATUSH��H���   L�e�Gt%D�.H��H��H�~L�FA����  D���$� /H f��EAD$AD$ I�D$0    H�E    H�E(   H��[]A\A]��     D���   ���   H���   A)�Mc�H��H��?H1�H)�L��H��?I1�I)��AI����t&H�9��8��8H��L�P$L��I��?H��H��L)�I�ӋAM��t&H�9��8��8I��H�H$H��H��?H��H��H)�I��H���P  M����  ����H��tH��L��1�H��H��H�H��H��H�M M���X  M����  ����M���	  H�}(A���   E��tfH�} L�E(�!�H�} L�E(H����  L�E L���     ���   Hc�Mc�H��L��H��L��H��?H��?L�� �  M��  �  I��I��I�� I�� L��H��I��I��fD�]fD�UH��[]A\A]�����fD  ���   ���   )�Hc�I���b���D  ���   I���h����H�sxL���   H+shL+Kp�5����     M��x[����M��tL��L��H��H��H�1�I��H�E(H�E L��L���9���I��������H�M(H��L��L������I������fD  H��  �M��t�L��L��H��H��H)�1�I��H���f.�     H��  �H���;���L��H��H��H��H)�1�H��H��H������H��  �M���/���L��L��H��H��H)�1�I��H��H������M���G���H�}(I���;��� L��L��1�H��H��H�I��H������� H9�}H�M(H��I������@ H�} I�������1�E1������f.�     H��tK�GtE��x19w8~,H���   Hc�H�@H���   H��t2H���   ��f�     �   �f.�     �#   �f.�     H���g���1�H���H��t[H��tfH�~ x_H�~ xX��   ��wASH��H��H���   H�GPH�@    H���   H�@H���   H��t*��H��[�f��#   �f.�     �   �f.�     H�CH����H��u@�t,�   ��u�H�L$H��������u��t$H��������@ �#   �f�     H�������1��y����H��(H��toH��HDָ@   H��@HL�H��@HLЅ�t7E��DD�H�t$H���$    H�T$�L$D�D$�����H��(�f�     E��uA�H   �H   �fD  H���D���ff.�      H��(��t(��Dց���  ���  G�������  G����@ ��u1�@   �@   H�t$H���$    H�T$H�D$    �0���H��(É���    H���g  M���n  H���   I�     I�@    H�@H���   H���,  ATA��L��UL��SH���Љƅ���   A����   L���   HcE IcQ H��H�H�� �  HcUIcA(H��H��Hc�H�M H�H�� �  H��Hc�I��H�}A����   A�Af��w6H��H����   H��G�z�GL�PL��H��L��H)�H��H�H��H�M A�Af��w2H��H���   H��G�z�GH�xH��H��H��H)�H��L�I��H�� I�� H���I���H�M L�E[��]A\� 1�[]��A\��    1���� �#   ����     �   ��f�     H��G�z�GA�   I)�L��H��I)�I��I�I��I���x���f�H��G�z�G�   H)�H��H��H)�H��H�H��H������ H��tkH��tvL���   I� H�@@H��tsAUI���C.H ATI��U��SH��L��H����H��tH� H��L���L��H��[]A\A]��D  H���   []A\A]ø#   �f.�     �   �f.�     �   �f.�     H��t[��tH��cinut_H�GPH��t^HcWHH��H9�s*H�;ruH���   1���    H�9rt�H��H9�w�   �f�     �#   �f.�     ���� �&   �f�H��tFH�H��t>�PH��~4H�pPH;>t+�J��   H���D  H��H9|��t��H9�u��D  1�ø�����ff.�     @ H��t+H���   H��tSH�PH��H���R;C r1�[��     1��ff.�     f�ATI��USH��H��t@H���   H��H��t1H�  t*�t$fD  H�CH�t$H���P ;E s�1҅�t
�T$�1�1�M��tA�$H��H��[]A\��    UH��SH���D$    H��tJH��H���   H��t;H�{  t4H�G1��P;C r�D$    H�T$1�H���?����D  �D$��t�1�H��t�T$�U H��[]�ff.�     ��t	H����   ��tz�N�E1�H��H��H��<@ H=fdcl��   H=deesutH�BH���   H��tD� ��AH��FtH��H9�t+H�H=kradu�H�BH���   H��t%�8�FpH��H9�u�1��f��Ft������    �Fp��f.�     �   �f.�     �   �f.�     H��tK�GtEH��t@H���   H�BPH���t/UH��SH��H��H��t&H�@H��t8H��H��H��[]���    1��D  H���   H�H�@@H��uH�BP����H��1�[]�@ �K.H ��H��tH���   H�BP��    H���   H�@P������ff.�     @ H����   H��tj��tf� ��H;G }c�GtUL���   I�@PH���tDU��SH��H��H��t\H� H��tH����H��[]���    I�@P����H���   []�@ �   �f��   �f.�     �#   �f.�     H���   H�H�@@H��t��L$�K.H H�$��H�$�L$H��tH���   H�FP�e����H���   H�@P�����t���ff.�     �H��tkH���   H�B8H���tZSH��H��tH� H��t$H��[�� H���   H�H�@@H��uH�B8����1�[Ð�V.H ��H��tH���   H�B8��    1��D  H���   H�@8�������    H��t[�GtUH���   H�H�@@H��tBU���k.H SH��H��H����H��tH�@H����H��[]���    H��1�[]��    1��ff.�     f�H��t[�GtUL���   I�H�@@H��tbAVM��AUI��ATI��UH���k.H SH��L����H��t,M��L��L��H��H��H� []A\A]A^��#   �f.�     [�   ]A\A]A^�f��   �f.�     �#   H��tv�Gt}L���   I�H�@@H��teAUI��ATI��U���k.H SH��L��H����H��t!M��H�L$L���H���PH��[]A\A]� H���   []A\A]��     ��    �   �f�H��t[H�H��tSH���   H�H�@@H��t@S�v.H H��H��H����H��tH��H�����uH�$H��[� H��1�[��     1��ff.�     f�H��tTSH��H��H�H��t;H���   H�H�R@H��t(�v.H ��H��tH��H�����uH�D$H��[�D  H��������H����f�H��t{ATUSH�_PH��tNH��tII��H��H���{���H��t#IcD$HH��H9�sH;+u�0H9+t+H��H9�w�[�   ]A\��     [�&   ]A\�fD  I��$�   1�[]A\Ð�#   �f.�     H��tTUHc�SH�,�H��H��H9�w�4@ H��H9�v'H�;�   u������H��u�H�H��[]�fD  H��1�[]�1��@ H��tH���   H��t	�xcinut1�� ATI��UH��SH��H�wP�H�g���H��t"H�PH���   D��H��[L�B(��]A\A��@ [1�]A\�f�     H��t<UH��SH��H��H�wP�H����H��tH�H���H���Q0��H��[]ø���������ff.�     H��t3SH��H�wP�H�����H��tH�PH���   H��[H�R8��1�[�@ 1��D  H��tKUH��SH��H��H�wP�H����H��tH�PH���   H��H�J@H����[]��f�H��1�[]��    1��ff.�     f�H��tKUH��SH��H��H�wP�H�#���H��tH�PH���   H��H�JHH����[]��f�H��1�[]��    1��ff.�     f�H��t+H�H��tH���    tH���   1���    �#   �f��$   �f.�     H��tEH��  H��tH�H��tH�HH�    H��t!H�A;p u�@ H�A9p tH�IH��u�1�� H��tH�
��    �ff.�     @ H��t-H��  H��t!H�B;p u�@ H�B;p tH�RH��u�1���f.�     ���   =stib��   AUI��ATA��UH��SH��=ltuo��   H����   H��  H��u�   �    H�[H��tzL�CA;@ u�D  1�D��H��L��A�Px��th<uYD���   M��tMI��  H��tH�KH��u�6fD  H�IH��t'L�AE;H u�H���L��(  H��  M��u��   H��[]A\A]�H��1�[]A\A]�1��ff.�     f�H��H��t(H�OH��tH���   H�z��H�������f.�     �   �f.�     AUATUSH��H��tQH��tL�GH�_I��L�,�L9�r�7�    H��I9�v'H�+L��H�E H�x袨 ��u�H��H��[]A\A]�f�H��1�[H��]A\A]�H������H��tH� H�@(H���fD  1�H���f�     H����   AUATI��UH��S��H��H�H�@@H��ta��H����tF��tBH�EH�X�@L�,�L9�s,D  H�;H9�tH�H�@@H��t
L����H��uH��I9�w�1�H��[]A\A]�@ �   1���    1��D  H����  H��t0�WH�GH��H��H9�sH;wu��    H90tH��H9�w�"   �@ AW��AVAUATUSH���OH�z�H9�v H�HH��H�H�H9�w�L�6L�fH��H�B�    L�nI�M��tI;�$0  ��   �uW�u3I�F8H��tH����H��L��A�UH��1�[]A\A]A^A_�f.�     H�SH��t�H�{ H�پ ;@ ������@ I��$  H��u뚐H�mH��t�H;]u�H�CM�<$�xHltuot~I��$  H���`���L��A�WI��$  H��u�qf.�     H�@H��t^H�P�z ltuou�H�I��$(  H� � ����    IǄ$0      �����    �!   �H�{hH���u���H�@p�P(�i���1��D  E1�A�   �����f�E1�E1������D  A�   A�   ����ff.�     @ H��t��X  1�Ð�!   �f.�     H��t+D�OD�G�GH��tD�H��tD�H��t���     1�E1�E1���fD  H���=  ��X  �P�1���X  ���  AWAVAUATI��USH��(H�D�H�D$.H H�T$H�D$    H�$H�D$D��E����   H�$1�L�(��    H��D��A9�vOI�\�L�3M��tI�~L��衤 ��u�A�t�H�C H��t�H�x����H�C H��u�E�|$H��D��A9�w�H�$H�$H�T$ H9��s���E��t���L��I�t�����A�D$��u�H�D$L��H���PH��(1�[]A\A]A^A_��     �H�$H�$H�L$ H9�u��ø!   �@ H����������tH��u�f.�     ��H���8  �D  H��t;H����.H ����H��t 1Ҿ�.H H���I���H��t� H���D  1�H��Ð1��ff.�     f�H��t{L���   �   M��t���   pmoct�D  9��   v��H�vH��I�A��AoB�A�B�A�BA� A�BA�H�D$ �AoJ H1�)L$��f�     �   �f.�     H���  H���f  AWAVAUATUSH��   f�? �n L�~(�J  H�G� f�D$f���  H�T$E1�H�4$H�|$H�D$(    L�D$L��H�|$��H��I�PI��I��L�4I��AoI�)L$@L�L$HH��H��L��L)�H��H�t$@L)�H�D$HI�$M�L$foT$@I��L��M�HI��)T$0H��M�A�
�����b  ����   H�$L�T$ H�|$@H�t$���uuM9���  L�T$ M��L��M��A�WL�pI�_����   ����  H�p��H�|$pH��H�t$H��L)�H�T$pH�PH��H��L)�H�D$xH�$�P���c  H�Ĉ   []A\A]A^A_�f.�     A�9M)�L)�������  I�H�L��H��H��?H��?I�H�I��H��L�\$@H�D$HI��I������f�H�p��H��H��L)�H�T$0H�PH��H��L)�H�D$8M9�wq�n  @���'  HT$0HD$8L�|$0H��H�t$pL��H��?H�H��H�T$pH��H��?H�H�T$H��H�D$xH�$�P������foD$`)D$0M9��T  I��I���H���3H��H���L)�H�T$`I�~H��H��L)�H�D$h@���W���H�$H�T$H�t$`H�|$0�P�������I��L��L9��0���M��H�$H�t$H�|$@�P��   �H�P I9��3  A�W�����"  H�p��L�p0H��H�pH��L)�H�T$PH��H�p H��L)�H�T$XH��H�p(H��L)�H�T$`H��H��L)�H�T$hM9��  H�p0H�|$PH��H�t$`H��L)�H�T$pH�P8H��H�T$pH��H�L$L)�H�D$xH�$�P�������I��L�������     M��M��H�$H�T$H�t$@L���P�������H�D$D�T$��D$(A����9�~_H�\$H�D$(H�SH��H�D$(�Bf�\$f�������     �   �*���fD  L�\$@I��H�\$H�n���D  �   �1������ �   �M��L�t$0�K���H�$M��H�L$H�T$@H�t$`H�|$P�P�<���f�H��t[�wD�1���fD	�tN��~EE��~@H�1������D  �G9�~(9�~$H����A9����    9ֺ   E��fD  �   �f.�     H���g  AWAVAUATI��USH��(H���    �(  H���   H���  H�߉�L���   A���t���f��C0C@CPC`��   AEI�E     ƃ�    I��$�   Hǃ�       H�Bǃ�       Hǃ�       L��0  ��ǃ�         ��   Hǃ�       E�Hǃ       Hǃ      Hǃ       ǃ�       H�Cp    H�Cx    Hǃ      Hǃ      @��t�����
������  @ E�M��t$���  uH�H� H����   H��   �!  H�BI��$�   ��D��H�����   ����  ���   ltuo��  A��A��A��A��   E����  Hǃ�       H�SPH���   ��    ujA�D$tbI��$�   H�SpH�y H��H��H����  H����  H�V H��H�SpH�SxH�q(H��H��H���z  H���z  H�Q H��H�SxE����   M��$�   A�t$0��tzH�S���   H���   H�RH��(  H��t;O t+H��  H��u�4  @ H�RH���#  H�z;O u�H�GI�L$ L��H���PXH���   L��D$�u����D$��ug@��ua���   ��pmoctS��stibtK������u1���   @�����tH��(H��[]A\A]A^A_�^���fD  1�H�߉D$�z����D$H��([]A\A]A^A_��    H��(�#   []A\A]A^A_�@ Hǃ�       H�ShH���   �F���D  I�L$�� �����A��A��   u&I��$�   H�~ H�>��  H��������    @�� u	����  A��I��$�   A����tK@��uEH�B��D�L$D��D�T$��@H�����   D�T$D�L$��u���   stib�|���I��$�   I�D�L$H��A��M��$�   D�T$H��L��H�@(A�K0L�\$A�C0    �L$D���P�L$L�\$D�T$D�L$A�K0����fD  L��������������A��A��A��A��   @�������H�K0H�s8L�{XL�s`H�{@H�L$H�KHM��M��H�t$H��I���I���H�Q?H���H���E���  H�L$H�SHH�s@H�t$J�T9?L�[XH���L�C`L)�H�S0J�T6?H���L)�H�S8H�KPH�Q H�KhH���H�SPH�Q H���H�Sh�@���fD  �#   �f.�     H���y����    H)�H��H���m��� H��������    H)�H��H���z��� ��ltuo�����@���:  ����������   M�D$(M�L$ H���   �������1��    ��L
��LBH��9������fD  L�C`L�D$H+L$H�SHI�|8?H���L�[XH���H)�H�s@H)�H�S8H�{0�����H��������X�����L��D�T$��H�T$���D$��c  �/hH H���ޚ I�L$H�T$H��D�T$t�z8t�|$tq�������I��$�   �����fA��$�   �����I��$   �t���I��$(   �e��������f�     L��L��D$豼��A�t$0�D$����H�H� ��u����� H���g  AWAVAUATUL��SH��M���]  H�G A��A��1�A�A��I������9���D9������   ����   E����   H���   H�@H���   H��t*A����   I��D��D����L���Ѕ���   <��   �   A��    uuA��   �   E��A��DD�Mc��"@ H���   I��H�ȃ�H�E H��A9�tPD���L���������u&I��$�   A��u�H���   I��H���� �   H��[]A\A]A^A_�@ A��tRH��1�[]A\A]A^A_ÐD���������@�������f�     �#   �f.�     �   �f�     H��D��D��H��[I��$�   ]A\A]A^A_����ff.�     �H����   H����   ;w ��   AUA��ATI��U��SH��H��H���   H�@H���   H��t<��t,M����   D��H���Ѕ�tN<tH��[]A\A]��    ������t�H��M����D��H�ߺ   []A\A]����fD  �   �f�@��u�H��H���   ��L��[�   ]A\A]�*���f.�     �#   �f.�     �   �f.�     H��t;U��SH��H��H���   H��tH�G�P;C �Ƹ    C�H����H��[]������#   �f.�     H��tSH��tN�   �9uSH9�tFUH��SH��H��H�Wf��uXH�f��u7�C �U �����	ЉE H��1�[]�D  �   �f�1��D  ��    H�}H�sH��� �fD  H�~H�sH���� H�}H�SH�s��� � H����   H����   UH��SH��H���F t:H�vH��t�WH�sH�C    H��tH���UH�sH�C    H��tH���U�    1�H�C    H�C    H�C    �C     H��[]�@ �   �f.�     �   �f.�     H��tH�?�C��� �!   �f.�     H��tH��t�Ѷ����ff.�     @ H��t)D�GH�GE��~1� ��H0��HPH��D9�|�ÐH����   f�? ��   1�E1��     H�WA��Hc�L�BH�GH��H��L��H�M��H��H�H9�s%L�H�rH��H���o@B�L�PH�pH9�r�H�WH�
L�H9�s ��2H��H��@�p��JH9�r�A���A�IA��9��g����w �f�H����   H����   H����   ATI��UH��SL��(  H��  H�rM��ttI�xhL��A�Pp��tN<uJH��  H��tH�KH��u�3f.�     H�IH��t L�AA�x ltuou�H��I�xhL��A�Pp��u�[]A\ø!   ø   ø   ø   ��f�     H��t;H��h�BH�$�P��D$    ��v<u�D$   H������H��h�fD  �   �f.�     H��tH��t�A�����ff.�     @ H��tH��t鱵����ff.�     @ H���  AWH��H��AVH��?H��?AUH�H�ATH��H��USH��xH�L$8H	�H�D$Ht0f� H��H�|$P~2茵���D$\��u,f�; �   u
�     1�H��x[]A\A]A^A_��D$\    H�D$Pf�8 L�p~�H�D$(    E1�E��f�     H�D$PH�|$(E1�D��D�|$XE1�M��M��H�@H�D$    H�D$     D�xH�D$    �D$����H�D$    D��E���lD  Hc�Hc�H�|$`H��H��L�L�H�
H�RH+H+PH�L$`H�T$h�*���A��M��tH�D$`H�|$hM��uP��H�D$I��M�ՍED9�MD$X��9��  ;\$��  ;l$u�H�D$ H�|$L�T$H�D$`H�|$hM��t��L$��yH�L$L�|$�\$H�L$ L�l$HcT$Lc�Lc�L��M��H��H��H��?H�L$0Ic�L��H�L$@L��H��?M�� �  H�L$0I��H�� �  Mc�H��Hc�I�I�����|  H�L$@HD$I��L�H�D$0I��   I��H��H��?H�� �  H��Hc�H��H��?H�� �  �T$\H��H����<  H)�H��H�D$M9�L�L$8Lc|$Ic�MO�Ic�Ic�I��H��H��H��H��?H��?H�� �  L��2 �  H��I��A9��   L��L��L�D$@�X���L�D$@H�|$HH�t$8Hc�H��I��L�<0H��H��?H�� �  H��A9���   I��H��H�|$0L������D�L$XL�@ Hc�H��L�L:HB�SA9މ�AN�9�u�H�D$`H�|$h�����H�D$PH�D$(E��M��H�t$(E�y� 9����������fD  H�D$HL�|$8D�L$X��    H)�H�\$0H�L$����fD  H�T$H�|$0L���^���D�L$XHD$H�O����    H�T$L��L�D$@�6���L�D$@������   �fD  H��������     H��tf� ~鏱���    1��D  AVI�։ʹ   AUH��ATI����.H USH��0��À� �ۅ��4  ��txH�l$L�m�
   H�t$L����� �E H�D$�8,��   L9���   H��L�pI9�u�L���
   H�t$�� �ǉD$,H�D$� ���   L9���   L�t$�A�~A�A�F����   ����   A�NA�v��xy��xu9�q9�mE�F9�eA���  w\E�NE�VA���  @��A���  A��D�u9���  w1A�T$@E�D$DA�D$HE�T$LA�L$PE�L$TA�t$XA�|$\��    �   H��0��[]A\A]A^�@ ��.H �   H����À� �ۅ�uL����   ��.H �   L���   ��� ��u�A�D$8   �   H��0��[]A\A]A^�f.�     ��.H �   H����À� �ۅ�tD��.H �   H����À� �ۅ�uX����   A����    H�A�D$`�.���f�     ��uLA�A�D$<����fD  A�>t"�   ������     �   �����fD  A�D$8   �����f�1��
   L���� H��A�D$<���� �
   1�L���f� �_���ff.�     �I���   ��.H I����� ����tR��.H �   L����� ����t'��.H �   L����� ����u\A�H<�
�@ A�H8�
�f�     A�H@�
A�HD�JA�HH�JA�HL�JA�HP�JA�HT�JA�HX�JA�H\�J��     �   �f.�     AWI��AVI��AUM��ATM��UH��S1�H��H�T$�ef.�     I�F(H��t1�1�1�L����H��u_I�F    A��    H��M�D� H��H�T$H��L��L��H�����0H A��H��H��	t3H�E     M��u�A��    �fD  A��U   H��H��H��	u�H��[]A\A]A^A_� 1�H��t�Gt��0  �ff.�     H�7H�WH�G    H�G@    H�G(    H�G0    ��     H��tH�G0H��t���ff.�     @ UH��SH��H��H�G(H��t1�1���H��uH�kH��1�[]� H9ws�H���U   []�ff.�      H��xSUH��SH��H�_H�G(H�H��t"1�1�H����H��uH�]H��1�[]��    H;_v�H���U   []�fD  �U   �f�H�G�ff.�     AUATUSH��L�gI9�v=L�G(I��H��H��H��M��t8A��I��I�41�H�uM9�rH��[]A\A]��     H���U   []A\A]�I)�H�7H��L9�LF�H�L���`� � H��H��H�w�q����U1�SH��H�GL�OL9�s"L�W(H��I��H��M��t!H��H��A��H��HkH��H��[]��    I)�L9�LF�HL��H��L��L����� ���     SH��H��tH�( tH�6H��t
H�G8H���PH�    [�D  L�G(H�WM����   �U   H9���   AUATUH��SH��H��H��~lL�g8L��A�T$H����   H�sH�H��H��H���S(H�3I��H9�vXH��tL��A�T$1�Lk�U   H�s@H�H�    H�sHH��[]A\A]�@ H�    �   u�H�w1�1�A��H�3I��H�s@H�1�H�sHLkH��[]A\A]�D  H�O�U   H9�s*H)�H9�r"H�H�H�G@H�H�H�GH1�H�w��    ��    H�    �@   �`���ff.�     @ UH��SH��H��������uH�S@H�U H�C@    H�CH    H��[]�ff.�     �SH�( H��tH�7H��t
H�G8H���PH�    H�C@    H�CH    [�f.�     H�W@1�H;WHsH�BH�G@���     H�W@1�H�JH9OHv�H�������B�	�H�W@�f�     H�W@1�H�JH9OHv�BH�������B�	�H�W@��     H�W@1�H�JH9OHv��JH������	��J�	�H�W@�f�H�W@1�H�JH9OHv
�H��ȉ�H�W@ÐH�W@1�H�JH9OHv�H��H�W@�D  UH��SH��H��H�G(�    �D$ H�wH��tL�   H�T$��H��t�E U   H��1�[]�f.�     H�s�D$H��H�sH��[]��     H9wv�H��0�ڐUH��SH���    H�wH�FH;GsKH�G(H��H��tW�   H�T$��H��u-H�sH�T$������B	�H��H�sH��[]��    �E U   H��1�[]��     1�H��Ht��@ AVI��AUM��ATI��USH��H��0H�F(H����  1�1�L��H����H����  L�c�   L��H��H�T$�D$    �����ŉD$���4  �|$ �k  �D$���^  �T$���Q  D�L$E���B  �L$�����t$D�D$A�����Hc�	��D$I�u 	��D$��	��D$Hc���	��T$	��T$��	��T$H���D	�E��D	�D�L$A��D	�Hc҅���  H9���  H��H)�H9���  H��������L�I��M)�M9���  L�L)�L9��{  L�H�KH�H9��h  I�L�H9��Y  H�C(I�u H���  1�1�L��H����D�D$H���  L�cA���   L��H�T$ H��D�D$/�D$    �4����ŉD$����   1��   �   1��     �T ��E�:TE�H��H��u�	���   H�CH�hH�C(H����   1�1�H��H����H����   H�k1�H�t$H�߉D$�����l$��u1H��H��xjI�H�C(H����   1�1�L��H����H��u$L�cM�&H��0��[]A\A]A^�@ L;c�����H��0�U   [��]A\A]A^�f�H��H)�H9��X���H��0�   [��]A\A]A^�D  H;V�8����H;k�?����U   �;���L;c�t����ff.�     �UH��SH���    H�wH�FH;GsKH�G(H��H��tW�   H�T$��H��u-H�sH�T$�B�����	�H��H�sH��[]��    �E U   H��1�[]��     1�H��Ht��@ UH��SH���    H�wH�FH;GsSH�G(H��H��tW�   H�T$��H��u5H�sH�T$��J�R����	�	�H��H�sH��[]��     �E U   H��1�[]�1�H��Ht��@ UH��SH���    H�wH�FH;GsCH�G(H��H��tG�   H�T$��H��u%H�sH�T$�ȉ�H��H�sH��[]��    �E U   H��1�[]�1�H��Ht���@ AVAUATI��U��SH��H��H�t$�b����T$��u	9�t�   H����[]A\A]A^�f�H�t$H���3����T$��u�H�CH�hH�C(H����   1�1�H��H����H����   H�kH�t$H���D$    �����T$��u�f��t�D��E1��,f�1�1�H��H����H��uNH�k�D$    A��E9��P���H�t$H�������T$���<�����t@H�CH�hH�C(H��u�H;kv�H���U   [��]A\A]A^�D  H;k�M�����@ H�t$H���;���H�ŋD$���y���H�t$H�������T$���`���Hc�I�,$�����    H��H�    H��tL�¾  �d���@ �Q   �f.�     H��H�    H��tL�¾ �4���@ �Q   �f.�     UH��SH���    H�wH�FH;Gs;H�G(H��H��tG�   H�T$��H��uH�sH�T$�H��H�sH��[]� �E U   H��1�[]��     1�H��Ht���@ H���G  H���N  AUE1�ATI��UH��SH�^H���s�H�W@�F�<��   ���$�H/H f.�     �C�L�L;EH��  �U   E��t:H�}( t#H�u H��tH�U8�D$H���R�D$H�E     H�E@    H�EH    H��[]A\A]��    �B�JH������	��J�	ȹ   f�     ��tH����H��K��s�L�@���/  @���  @����   H�H���s��F�<����H�U@1��1���f.�     ��JH������	��J�	ȹ   뀋1�H���s��� �1�H��ȉ��_����    �BH�������B�	ȹ   ���8����     �H�������B�	ȹ   ���������   H��������    �s�H���������k���H�U@A�   ����D  �����f�     ������f�     f�������     @��t L�������f��   �f.�     �(   ��K�L��s&�uT��t��2@�1�t��T�f�T��fD  H�2H�1��H�|2�H�|1�H�yH���H)��H)���H�։��H��|����2���1�T��T��i��� H��H��H���q���H�$H����     H��H��H���Q���H�D$H����    H��H��H���1���H�$H�T$�   H��H��yH�ھ����H��yH����H������H��tH��H��H��H�1�H��H��H�ڃ��HD�H����     H��H	�u1��D  H��L�T$H�<$H��H�t$L���s���H���k���H�D$H��ÐH��t醝��fD  �ff.�     @ H���/  H���&  USH���oH�)$HD$��   L�\$I��H��H��L�������H��L�҉�����H�$H��xv�[��H��H��   @H�T$H�� H��x~�[��H��H��   @H�� ����   �M��   ��H�H�0H�H��?H��?HΉ�H�H��H��H�3H�SH��[]�D  H��&$����H��H��   @H�T$H�� H��H��y�H��&$����H��H��   @H�� H�څ��z�������H��H��H�3H�SH��[]�fD  ��    H����   SH���o)$H�$H��tiH�|$ uH�H��H1�[H)�� L�T$H��L��踕��H���讔��H�$H��xM�[��H��H��   @H�� ��U�ى�H����[����    H�T$H�D$H��[H��?H1�H)��fD  H��&$����H��H��   @H�� H�څ�~��K��   H��H����[H�H��H���@ 1��D  H��H�<$H��H�t$�����H���fD  H����H�������   H��tATUSH���o)$H�$HD$tUL�T$H��H��H��L��覔��H��A��蛓��H�<$H��xB�[��H��H��   @H�� E��xJD��H��H�D$H�;H�E H��[]A\�fD  ��    H��&$����H��H��   @H�� H��E��y�D�������fD  H��tH�7H��H�G    ������     �ff.�     @ H��H)�H= L�}f�H  hH= L�|�ÐH-  hH=  � �ÐUH��SH��H��H��~/�WH��H��tDH��1�H����� H��1��E H��H��[]�D  1�H����Ѓ��E H��H��[]�fD  �@   ��f�     UH����   SH��H��H�T$�u����T$��uH�H�E H����[]�ff.�     f�AVAUATI��UH��SH��H��H���D$    �y� L��I���n� H�T$H��I�t�����T$��un�/   H��H����s I��H��tNI��H��H��I)�I�mI�V�-o B�D3 L��H���o H��H���o H��H��[]A\A]A^�f�     � �� H��1�H��[]A\A]A^�fD  UH�ֺ�.H H��SL��H��H�?����H��tH�E 1�H�    H��[]� H���@   []�ff.�     �UH�ֺ�.H H��SL��H��H�?�����H��tH�E 1�H�    H��[]� H���@   []�ff.�     �AWI��H��AVI��AUM��ATI��U�
   SH���� H=���wI�?H�pH�T$H�������l$��tH����[]A\A]A^A_�@ H��L��H���� H�H���c   �/rsrf�CI�I�E     �AWI��H��AVI��AUM��ATI��U�
   SH���w� H=���wI�?H�pH�T$H�������l$��tH����[]A\A]A^A_�@ H��L��H���-� fo�� H�H���c   f�CI�I�E     �ff.�     H��t[H��tVUH���`  SH��H��H�T$����H�D$��u&H�   	   H�H�J�B    ǂX     H�U H��[]� �   �f.�     AVAUATUSH��H�    H���  H����   L�7I��H��H�T$�P   L��� ���D�l$H��E��uBL�p8��tIH�CH�SH�E    H�E@    H�U H�EH�E(    H�E0    L�u8I�,$H��D��[]A\A]A^Ð�u<I�V���   H�{  ��   H��L���ҋD$H�k ��t�H��u(A����    H�sH���$� H�S�D$H�U ��t�I�VH��L��1���D�l$�w���@ H��A�   [D��]A\A]A^�f�H��A�!   [D��]A\A]A^�f.�     �D$   �fD  ATUH��SH��PH�t$(H�T$H�t$�D$   �y����Å�u@H�|$H��tIH�� �����H�l$��H��tH�E0L�e8H��tH����H��L��A�T$H��P��[]A\��     H��P�Q   ��[]A\�AVH�ֺ /H M��AUI��ATUH��SH��L�'L�������H��tSL��H��H��H���2�����t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      AVH�ֺ/H M��AUI��ATUH��SH��L�'L���8���H��tSL��H��H��H��������t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      AVH�ֺ/H M��AUI��ATUH��SH��L�'L������H��tSL��H��H��H���������t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      H����   ATUSH�� L���   M����   H��I�|$H�T$H���������unI�D$L�d$H���   �   H��tL��H����L�d$1�H�{  t�+���M��t1I�T$0I�\$8H��t�D$L���ҋD$��u�D$L��H���S�D$H�� []A\��    H�� �"   []A\�f.�     �#   �f.�     H��t+H��HH�t$H��H�D$     �$   �����H��H�D  �   �f.�     ATI��USH��H��H�GH��(  H���   �B�tIH���   H��tH���UHǃ�       H�T$L��H�������H���   �D$H��[]A\��     ���B���     H���'  H���   H���  AWAVAUATUH��SH��H��(L�hH�@H�T$H�pXL������I�ċD$��tH��tH�E     H��([]A\A]A^A_� I�\$H�T$�H   L���   �D$    I�GM�wH�$I�GL��I�$�&����T$I������   I��$(  I�H� ��ttH�$H���   H����   L���ЉD$��uvH���   I�T$L���   H���U���L�e H��([]A\A]A^A_�@ �   �f.�     �#   �f.�     H�T$��   L��L�D$�y����T$��t!�T$L�������L��L��A�U�D$�����f�L�D$L�0I� �D$    �4����     �D$�D����    AWI��AVAUE��ATI��USH��8H�oH�_H�D$,�T$H�uHH��H��H�L$L�L$������T$,I�ƅ��0  L���   �|$ H���   I�$I���   tI�N   H�T$,��   H������I�ǋD$,����   M���   I�Gh    E��~<H�L$A�U�H��H��H��fD  H��I�h uH�8rcniuH�HI�OhH9�u�H�E`A�Gt����H����   �T$L�D$D��L��I�<$��I���   �D$,I�$����   H��L������H�EhH��tL����M��t	L��H���SM��t	L��H���SH�D$pH�     �D$,H��8[]A\A]A^A_�f�H��tsH��H��E1�轍��H�EhH��u��f�I���   I�$L��蝃����t<&t�D$,�f���@ H�D$pL�0�D$,��t�H��L���m���H�EhH���N����S��� H�EhH���Z���1����Q���f�H���  H���  H���   H����   AWAVAUATI��USH��H��L�pH�    H���   H�T$I�vPH�������t$I�Ņ�t$M��t	L��H���U�D$H��[]A\A]A^A_� H�T$�   H���v����L$I�ǅ�tM��t�L��H���U� I�] H�T$�H   H���B����T$��u�I�EPI�FpH��tL���ЉD$��u�M�,$H���   L��M�o�ٌ���D$���c���� �"   �f��#   �f.�     �   �f.�     H���O  H���N  H�~ 	  �   �+  AWAVAUATUH��SH��(�GH�4$�D$���f  ��L�fH�_L�l� �D  H��I9�t?L�;L��M�7I�~�cc ��u�H�$�   I�VH9Q��   L��H��菻���E�D$�|$L�m �0   �D$    wxL�4$H�T$L��I�v�����H�ËD$��uXI�H�kL��L�kL�3�uq�tH��0  �tH�SH�$H�@0H����  H���ЉD$���?  �U�J�MH�\�H��([]A\A]A^A_�f�     ��    �!   �f��   �L�e H�T$�   L���T���I�ǋD$����   H�M��A�ƋBHH�S�C =ltuou@H�BpH�T$H�@H��t.H�shL���ЉD$����   H�T$H�BpH�@ H�CpH�BPH�CxI�_H��  L��觊��H��  H��u�   fD  H�@H����   H�P�z ltuou�|$H��(  ��t	E����   H�3�|$H��H����������    M��ua�D$H�3�t"H�CH��t�xHltuouH�{hH��tH�@p�P(H��L��A�U�D$�����D$�{���L�/�D$    ����1��d���L��L��A�T$�|$�h���fD  SH��H��~�W1�H�������[�D  1�H����у��[�ff.�     @ SI��H��H��H��?H��H��?��H���uH��y�   A�H��L��[� H��tKH��tF�����
   H�H��H9�|�H��H��H��uNL�$H��L��1�A�RL�$H��I�������@ 1�M��t�L�$L��L��A�RL�$E1�L��A�H��[�H��L�L$L��L��L�$A�RL�$L�L$H��LE�H��ۃ�@�D���ff.�     AVAUI��ATM��UH��SH��H��L�L$�D$    �����I�ƋD$��uI9�|A�$H��L��[]A\A]A^�f�L)�1�H��H��I��I�<.�\� �D$�ːSH��E1�1Ҿ   H���GH�?L�L$� �k���H��H�C@�D$��uVH�sL�C �C�SH��Hs(H��H��H�spH�s0I�H�H�L�ChL�CH�SHH�J�4FH���   H�sxH���   H��[�AWAVAUATA��USH��H��(�G�WbD�L�/�D$    ��D9�w,�G�O`�W�A�1�D9���   H��([]A\A]A^A_�f��n������  �N  D��L�G A��   L�L$L��H��L��H�D$�g����t$H�C ����   L�C(H�T$L��L��L�L$�   �9����L$H�C(����   �{ �  H�s�C`�k�S�H��A�D9���   �    A��A���A���  ��   L�C0L��D��L�L$�   �����H��H�C0�D$��uWD�cH�KH�SL�C H��HS(H��H�SpH�OI��{ H�SxL�ChtH�S@H�HsHH���   H���   �������H���L����D$H��([]A\A]A^A_�f�     H��(�
   []A\A]A^A_�@ �D$H�{0�i��� L�C@C�?�L- L��L�L$�   ������T$H�C@��u�H�T$I��J�<0H��H�4�9� Ls@L�sH�����    AWAVAUATI��USH��H��L�nL�~D��D����������tH����[]A\A]A^A_�L��E���D$H�{ L��I�t$ H��H��H�D$�d� H�{(I�t$(L���S� H�{0D��I�t$0H��?� �{ �L$tZA�|$ ��   H��H�S f�kH��Hk(fD�kH�H�kpH�ShH�S0J�jH�SxH�S@H�HCHH���   H���   �@����H��f�kHk(H��HC fD�kH�ChH�C0H�kpJ�hH�Cx�����    L�|$H�{@I�t$@L���� H�{HI�t$HL���|� H��H�S f�kH��Hk(fD�kH{ �L$H�kpH�ShH�S0J�jH�Sx�E�������ff.�     @ USH�����   �WGPL��D$    �1�9�wH��[]�@ �^L�GXH��L�L$����0   L�׉������H��H�EX�D$��uŋMP�]H�IH��H�H���   H��[]ÐSH��E1�H����   1Ҿ   H�P   �   H��H��C    L�L$H�C�@ H�C�@ �X���H�C �D$H��[�f.�     H���  AUATUSH��L�'IcT$H��~3M�D$PI;8t4�J��   ��H����    H��I9|��t��H9�u�H��[]A\A]�1ۍJ�fD  H��Hc�L�L$�   I��$�   M�l�������T$I�D$P��u�A�|$H�SD�G�9�~8Hc�H���H���H��H�9�tI�D$PH�t�D9�u߃�L�.H��9�u�E�D$HI9�$�   t:H�E H���   H�EH�@H��tH����H��H���SH��[]A\A]Ð��    IǄ$�       �f.�     AWAVAUATUSH��(�D$    H����   H����   L�*M����   M���   H��H��I��H�t$H�7H�T$L���g���I�ƋD$��uf�oE H�CI�^AH��tH�t$L���ЉD$��utIcUHM�EPL�L$L���   �JHc��T���H��I�EP�D$��uEIcUH�rA�uHL�4�M��tM�4$H��([]A\A]A^A_�fD  H��(�   []A\A]A^A_�@ I�H���   I�FH�@H��tL����L��H��E1��S�D$M��u��ff.�     f�H����   H����   �    H�A    H�A    H�A    �A     ����   9���   �
   ���  ��   AVA��E1��   AUATA��1�UH��SH��L��H��L�L$�9����T$H�C��u&L�L$E1�L��1Ҿ   H������H�C�D$��t7�K H��H�������D$H��[]A\A]A^��    ��    �   �f�Ic�L�L$E1�1Ҿ   H������H�C�D$��u�fD�sfD�#�K �ff.�     H��tH�?����� �!   �f.�     AWAVI��AUI��H��ATI��USH��H���ns���D$    I��H� H��tL�h1�H����[]A\A]A^A_�@ H�T$�   L��������l$��u�I�L� L�h�C;s���C�D  D�c�����E1�L��L�L$�   L�{ �D$    C�$�ȉK����1�����H�C �D$��uaE��tcA�D$�M��M�l��    I�$H��tH�8H���r��I�$H�I��M9�u�M��t
L��L��A�V�D$��u�C�P���D  ������M��u���f�����ff.�     ������f�     AWI��AVM��AUATUSH��H��8H�H�L$H�D$H�F(D�L$H����   1�1�L��H����H����   L�{H�t$,H���D$,    �<����T$,��ux�D�`A���  ��   1�E��G�   fD  H�t$,H�������T$,f�D$��u:H�t$,H��������T$,��u%M9�tl��A9�tTH�t$,H�������T$,I�Ņ�t�H��8��[]A\A]A^A_� H;V�I����U   ���    �   ��f�     �   �f�     �T$H�L$xH��Iǃ�Hc�H�H��H���
  w�H�C(H���l  1�1�L��H����H��u�H�D$xL�{1�L�L$,H�|$E1��   �D$,    H��n����T$,I�Ņ��3���H�D$xH�0H���  L��E1��    1�1�L��H����H����   L�sH�t$,H���D$,    �����L$,I�ǅ���   H�CL�pH�C(H����   1�1�L��H����H��umL�s�D$,    M���  H�D$xA����� I��H��L�}�H�0L9�~wH�t$,H���+����t$,f�E ��u'H�CL�pH�C(H���:���L;s�E����D$,U   M��tH�D$L��H���P�T$,� ���L;s�e�����L;{������#����|$ u{H�D$xH�|$1�E1�L�L$,�   H��	����T$,��u�H�L$x1�H�9 ~#H��H�|$H��I|H�L$xH�<�H��H9�H�T$p�D$,    H��T����D$,   �G����0@ �   L���� �n����     AWAVAUATI��UH��SH��H��   H�L�D$H�L$`L�D$hH�$�{���A��tH�Ĉ   D��[]A\A]A^A_��    L�t$xA�   H��H��AVA�TSOPL�l$xAUH�L$xH�T$p�����AYAZ���  AVE1�A�tnfsH��AUH�L$xH��H�T$p�����A��XZE���y���L��H�L$xH�t$pH�H��I��I��?I1�L9��`  H�E N�,�H�D$H�C(H����  D�T$1�1�L��H����D�T$H���?  L�kH�t$\H��D�T$�D$\    �����D�t$\D�T$I��E���  H���M  H=��� �1  H�L$L��H��H��D�T$�.  D�T$��A�ƉD$\�:  H�C(I��H����  1�1�L��H����D�T$H����  L�kH�|$H�T$\L��D�T$�D$\    �l���D�t$\D�T$I��E���v  H�sL��H��H��D�T$����D�T$��A�ƉD$\�F  A��.H I��~A�<$OTTO�/H LD�L�L$1�L��L��H��D�T$�  D�T$A��H�t$pH��tf�H�$D�T$H���PD�T$E���L  H�D$H�T$xH� H�����fD  I��L�|$xL�t$p�D$\   I���h  M����  H�E E1�E1�H�l$H�D$�xf�     1�1�H��H����H��uqH�kH�t$\H���D$\    �����D�T$\E����  H=��� ��   ���� I�L$H)�H9���   N�d I�EI9���   I��H�C(K�,�H��u�H;kv�L�t$pA�U   M��tH�$D�T$L��H���PD�T$E�������H�D$H� H�    ����f.�     L;k�W���A�U   H�������E���[����    L�t$pA�	   � I�D$H�l$H�D$0H���o  H�t$0H�|$H�T$\�+���D�T$\I��E����  E1�� �  1ɾ   fD�@�   1�L�d$@I��L�t$(I��L�l$8I��H�l$HH���D$$   �e  �1�1�L��L�D$H����L�D$H���e  L�CH��H�t$\�D$\    �H����|$\���@  H=���H�D$�/  H�t$\H���>����t$\�����  ���D$\
   ��   H�T$H�J�H���    HF�;D$$�n  H�|$0I�uH9���   L��G�4/H��C�T/L��H��C�T/L��H��C�T/���1  H�UH9��I  A�/�L�mI��A�D/A�D/ A�D/ A�D/ A�D/ �D$$H�D$@H9��  H�,H9��  H�sL�H��������D$\��u3I�D$L;d$8�  I��H�D$(N��H�C(H�������L;C������D$\   H�D$L��H���PD�T$\L�t$p�T����    A�   M���C��������@ A�   �}���L;k�d��� H�t$pA�U   �`���H�t$p�V���fD  L�t$pA�
   �����I�H������H�t$pA�	   �%���H�t$pA�   �����L$\���E����8���@ H�t$pH�����������H��H�|$0L��L��H�PH�l$H�D$\
   H9������I�uA��A�DH9�r�H��A�L�L$H��H��A�/H A�DH��H��A�DH��1�H��A�7L���
  L�t$pA������M�������H�D$D�T$L��H���PD�t$\D�T$�����H��H��L��L��H�l$H�D$\
   H�PH;T$0�F���A�?�A�D?�Q���f�AWH��AVH��AUATUSH��  H��H�D$X    A��H��?H�D$`    A����  H����  E��E1��tE1�H�~  A��H�T$H�T$XH��H��D�D$(H�L$H�|$�����D$T����  H�H�D$ �E ��p  L�](M���c  I���A  ��l  D�E0L�M8H��L��D��H�D$hPH�L$H�t$hL�\$ �s������D$dA[[L�\$�  M��H�|$ H�T$T�   �h����|$T���%  L�D$`I���   L�@H�� tH���q��L�D$`H�|$ xH1�L���W����D$T���{  H�|$`H��$0  ������D$T���]  L�D$`H��$0  I���   I�@�t+A���   f��y
��fA���   � uA���   fA���   ��  A�P8���  I�@@�z�H��H�H H��$fD  H�x xIH�x xBH��H9���  H�� �f��y��f�H�pH��yH��H�pH�pH��yH��H�pf��y�1�1�H�@    f�Pf�0H�@    H�@    � H�D$     ��E1�H�\$X��Qtg��tb��Ut]H��t4H�C0H�k8H��tL�\$H����L�\$E��uL�\$H��H���UL�\$H�t$`H��tH�|$ L��������D$T�	  @ �|$( ��  �T$T��u��D$T   널H�D$�D$T   H�X�@L�$�L9���  E1��   �    D�E0L�M8H��D��L��H�D$hPH�L$H�t$h������D$dAYAZ���������E��t1H���.H �	   H�H�r��� ��u=�   tjf.�     M���������H��I9��'  L�;I�� t��E �b���E1�E1��_����    �   H�ĸ  []A\A]A^A_�f�     L�D$XI�@(H��tZ1�1�1�L��L�D$0��H��uJH�t$XL�D$0I�@    H�L$H�T$H�|$�D$T    �  �D$T����  ���;��� L�����D$TU   H�\$XM��H���  H�C(H��tL�\$(1�1�1�H����L�\$(H���X  1���   H��L�\$(H�C    H��$0  H��H�D$0����L�\$(����   ��$0  
�$z  
�$�  ��  ��$1  �P��� ��  ��$o   �  ��2   �q  ��$�   �c  ��$�  L�D$H��L�\$(H�L$H�|$�Hc�H��H��H������L�\$(�Ѓ��  ����  ��U��  �D$TH�\$X���H���H���"���H�C0H�k8H��tH����E������H��H���U�����fD  �D$T�����D$T    H�\$XH������������E u�D$TU   H�\$X�f���E1�E1�����H��$0  H�D$0H�D$H�UH��E1�L�D$0L�L$pL�\$@H��$�   L�0H��H��A�   H�D$h    �h���1�1�D�l$(L�t$8��L�l$0D��I��M��I�����   F�D�pE����   J����   Ǆ$�      H����  H�T$hH��$�   L��H��$�   �I�����t<Q��  ��utH�t$hK�T� L��L�D$H�L$����H�t$hH��t<H�N0H�V8H��t!�D$LH��H�T$0H�t$�ыD$LH�T$0H�t$�D$H���R�D$���  �۹   E�I��I��	��   L��H�����0H ��1ۃ�����@��uһ   �����L�D$H�L$1�H��H�|$L�\$(�_���L�\$(������f�H�|$`���������I���   H�|$ H�    H�@    H�@    H�@   H�@     H�@(    �@x   �@p���   H�D$L� ����H��u�M���v���f.�     I�G�q����E �4��������L�\$@H��$�   D�l$(A��L�t$8H�]HM���    H�u H��tL��A�VH�E     H��H9�u�M��H�\$XE���3����D$T    H�\$X������   ����L����~�������H�\$XE1�����H�\$XH�������H�C0H�k8H��tH����E�������H��H���U�D$T����ff.�     f�H��t3H��HA�   H�t$H���$   H�D$     ����H��H��    �   �f�H���7  AWAVI��AUI��ATM��UH���P   SH��XL�?H�T$L�D$L��H�$����H�ËD$����   L�D$H�+L�sH�C    H�C@    H�C(    H�C0P@ �D$   H�\$0M��tL��L���D$
   �o���H�D$8H�$E1�L��H�t$L��������uI�$H�b����H��X[]A\A]A^A_�@ H�S0H��t�$H���ҋ$�$H��L��A�W�$H��X[]A\A]A^A_�D  �$H��L��A�W�$H��X[]A\A]A^A_�f�     �   �f.�     AWI��AVAUI��ATUSH��H��HH�H��L��H�L$H�D$��HO�H�FH�t$<H�$�����T$<��uUH=1pytt]�D$<   I�G(H����  1�1�H�4$L����H����  H�$�T$<I�GH��H��[]A\A]A^A_�D  �T$<��u��f�H�t$<L��購���T$<A�ą�u�I�GH�hI�G(H���c  1�1�H��L����H���>  A��I�o�D$<    �D$ ����  H��H������L�l$(1�H���D$' I��H��?H�D$�- I��1PYT�#  �|$ t	L9��K  ��;l$ �.  H�t$<L��������T$<I�ą��"���I�GL�pI�G(H����   1�1�L��L����H����   M�wH�t$<L���D$<    �����T$<I�ƅ������H�t$<L���s����T$<�������I�� DIC�B���I��I��H��H����  �D$'�0��� H�$I;G�X���f.�     �U   �P���fD  I;o�������@ M;w�N����U   �&���@ I��I��H��H���t  �D$' ����f�     ��   �����fD  L�l$(I��I�G�D$<    �   L9������H�ƺ   L)�L9������M�G(L4$M����   L�\$1�1�L��L��A��L�\$H���)���M�wH�|$H�T$<L���D$<    L�\$�v����T$<H�����k���L�\$I�wH��L��L��轵��L�\$���D$<u^�|$' �/H L��H��A�'hH �    L�L$L��LD�H��HN������D$<��������D  L9��V����z���f.�     H��t�H�D$H��H���P�T$<�������I��L�l$(�D$'����I��L�l$(�D$' ����ff.�     f�H��t;H��HH��L��A�   H�t$H��H�T$H���$   H�D$     �����H��HÐ�   �f.�     A�   ����D  AW�   AVAUATUSH���D$   H��thH��tc�Gt]��0  9�vR��H��H  H��1�H��H��CL�sf��tM��tC���f�E �Cf�E�Cf�E�CL�u�Uf�E1�H��[]A\A]A^A_�f�     L���   1���E1�L���   L�L$�   L�������T$H�C��udM�E(L�{M��tI1�1�L��L��A��H��upH�CM�}�KH��L��L���D$    苳���D$��u@L�s�S�6���M;}v��D$U   H��tH��L��A�T$1�H�C    1�f�C����H�C���D$U   H�C��ff.�     @ AW�   AVAUATUSH���D$   H��tfH��ta�Gt[f��8  �   uL�   �� �  v?�� �  ;�P  s1H��X  H��H�vH�,�1��E L�uf��tM��t��L�31��SH��[]A\A]A^A_�L���   1���E1�L���   L�L$�   L���3����T$H�E��uJM�E(L�}M��to1�1�L��L��A��H��umM�}�M L��L��H�U�D$    �����D$��t)H�EH��tH��L��A�T$1�H�E    1�f�E �F���L�u�U �9���M;}v��D$U   ��D$U   H�E�ff.�     f�SH��E1�H����   1Ҿ   H�P   �   H��H��C    L�L$H�C`@ H�CP@ �8���H�C �D$H��[�f.�     H��t�g�     �ff.�     @ AUATI��UH��SH��H��H��~@H���WI��H��tJE1�H��tL��H��H���ϡ I��E�,$H��L��[]A\A]��    A�    A�   t����     A�@   ���     ATI��1�UH��SH��H��tH���r� H�PL��H��H��[]A\�N���ff.�      H��v:���t3H�T��@ ���t!H��H���G�H9�u�� 1��> ���D  H��1�� �> ��ÐH��t#H�H��tH;pu� H9ptH�@H��u��1���@ H��tH��t�A^����ff.�     @ H��tH��tH�H�    H�FH��tH�0H�7�@ H�w��f�H��tH��t�!^����ff.�     @ H��t1H��t,H�H��t$H�VH�PH��t!H�H�H�    H�FH�0H�7�f�     H�G��f.�     H����   AUATUH��SH��H����   I��A��H�˅�t
�   H��ttI��  I��  H��u�}D  H�vH��toH;nu��L����} ltuotsH�EL�hhE��t>E�a�I��I��I��D  H��L9�tH�SH�3H��A�Յ�t�H��[]A\A]� H��1�[]A\A]� H���   []A\A]��     H�EI��(  L�hhE��u���f.�     �!   �f.�     H��tKH��tFATI��UH��SH�?H��u�"f�H��H��tH�_L���Յ�t�[]A\�fD  [1�]A\�f�     �   �f.�     H��tH��t�q\����f.�     D  H��tH���   H�H�@@H��t�`1H ���1��ff.�     f���f.�     @ H�/H���    �   �f.�     �   �f.�     H��p  H�    H�A    H��tSH�����   H�H�1�[�f�1��ff.�     f�H�H���   H�@hH��t}H�L�BM��tqSH��H�� HcW`H�D$    H��H�$HcWdH�D$    H�xH�T$1�A�Ѕ�u'�$�{l Hǃ0      �C`�D$�Cdu�Cl�ChH�� [�f�     �ff.�     @ H��X  �   H�J
H9�`  rw������B	�f�G<�B�����B	�H��H�G@�B�����B	�H��H�GH�B�����B	�H��H�GP�B�����B	H��X  	�H��H�GX1��ff.�     @ HcG`H�w@H�HcOdH)�H���   H��H��H��zx(tXH�Gp1�H�Gx    H���   HǇ�       H��8  Hc�0  H��H  Hc�4  HGXH��@  H)�H��P  �fD  H��  H��t���)   A����.   H�Gp��H�Gx    H���   HǇ�       A��t�������Hc��s���1��l���@ H��pglh�s  vqH��srts�T  �.  H��oxps�1  ��   H��r  H��sxbs�  ��   H��x  H��oybs��  H��t  �    H��sybsHD��D  H��7psg��  �e  H��dlch��  �
  H��9psg��  ��  H���  H��csah��  H���  �    H��alchHD�� H��v  �    H��oxbsHD��H���  H��oyps�C  ��  H��|  H��syps�)  H�Ǆ  �    H��ortsHD��f.�     H��nrcv��   ��  H��  H��sdnu��   �S  H��   H��csav��   H��  �    H��focvHD���    H���  H��nrch��   ��   H���  H��srcht}H���  �    H��csdhHD��fD  H��2psg�S  vY1�H��4psg��  ��  H��5psg��  H��6psg�  f���  vH���  H���@ H��  ��     H��0psg��  �  H���  �    H��thpcHD��D  H�Ǫ  �    H��fochHD���     H��z  �    H��sxpsHD���     H��   �    H��odnuHD���     H��  H��csdv�S���v2H��  H��pglv�=���H���  �    H��tghxHD��fD  H��  �    H��srcvHD����    1�f���  �����H���  H���@ 1�f���  	�����H���  H�� �@ 1�f���  
�����H���  H��$�@ f���  �����H���  H���fD  f���  �q���H���  H���fD  f���  �Q���H���  H���fD  1�f���  �/���H���  �H���  ��     1�f���  ����H���  H���@ H��~  ��     H���  ��     H���  ��     1�f���  �����H���  H���@ Hc�Hc�H��H��H��?H��    H���f����  ��     H���  H���@ H���  H���@ H���  H��@ H���H���   �@x��(t��#tHV(�
�fD  ��+   u�H��HV(H��HFH�
�f�     H���H���   �xx(tH��H��HFHHHV(�
�fD  ��+   tڀ�,   tр�-   u��� ��H��HVH
Ð��H��HVHJ�H��H��xHк    HH�� H)к    H��HO���     �Љ�%�   ��@t��   =�   �)  =�   �  H��H��H  �Ѓ�0����   ~k�� ��   ��0ucH�vH��H�HHI�H��
����   ��Hc�H��H��H�BHH�H��H��H��H��P  H��H  H��X  �f.�     1Ʌ�t�H��P  H����u��@�     ��udf����H����0H��H  ���S���H��H�NHI�H��
���g���H�V��w����    H��H��?H�H��	���@������    H��H  �����@ ���Hc�H��H  �����@ H��"  H��$  Hc�Hc�H��H��H�H��H��?H��    H��H���     H��  H��   Hc�Hc�H��H��H�H��H��?H��    H��H���     H���ff.�     �H���ff.�     �H��&  ��"  f�� @�N  ��(  L��$  f�� @��   H��H��H��I��H�H��H���  f�� @��   f��$   @�$  HǇ�  ��@ f��   @��   f��    @��   HǇ�  ��@ H���  HǇ�   �@ HǇ   `�@ H= @  tkH�  H=�  wHǇ�   @  HǇ�      �fD  L���  f�� @�[���f��   @HǇ�   �@ �j���HǇ�   �@ �t���@ f��&   @tef��(   @u�HǇ�  ��@ HǇ    �@ �}����    H��H���  ������     HǇ�  0�@ ����HǇ�  0�@ �����HǇ�  P�@ HǇ   ��@ HǇ�      �ff.�      H���  Hc��  H��  H���  H9�}-H���  ����  �� >H ���  ��xHc�H�H9�};�G�   �   �D  L�@L9�~��t��   )򉗜  Hc�H�H9�|�1��@ AWAVAUATUSH��H��L�.��  fD9��   �/  H�vH���  H�NH�WH9��  f9CT�	  H��H  H��8  H�|$H���  H����  H��X  I��H)�H�H1�H)�H;�P  ��  }H��H��M��HH�I��A��L���   H��HCXH��H��L�L�PI�f��n   I��uF��&  D���g�����(  D��H�I�M��P���H�I�H���   M�P�Ao L�RL�
I�PI�0H��L)�L)����  H���   H��I����  L�H��HC`H�QH�1H+PH+0���  ��D   H��tL��L��H��L1�LH����  H����H����  @���  ��n  f9�l  uL��L)�H��H��?H1�H)�H;D$MO�H�L$L��H�����  ���  H�L$��tM����   H9�HL�H)�A��H��H��H���   ���  ��  f��  ���  tfD��  fD��  H��[]A\A]A^A_�fD  ���   t��C�   f��  ���  t��fD  L��X  L��H��?H��L1�H)�H;�P  LM�����f�     L��M��x(Hк    HH��$����    H��H9�HO��#����H)к    H��HO������ff.�     �AVAUATUH��SH����  L�m M����  I��H�s8A�   �   �E H�����  H��H����<q��   L�F <rID���`  H�H��I9�tWI��M9�r=H����   H�C0H�~�H�{8H�T��f9STw����   H��t�I���C�   M9�s�H�s@[]A\A]A^�@ ��H�A�H��H�Ή�HI�H�*�b  H���   H��H��xx(tXH�sH��H�����  H�s8�`����    H���>����    ���   t�C�   1�H�C8    H�s@[]A\A]A^Ð��+   t���,   u6���   tf��(   ����L�Cp��H��A� ������e���D  ��-   H��������H�s8����ff.�     f������Ƈ�    H���   1�HǇ  �����ff.�     @ �Gx(   1��fD  �ff.�     @ H���  A��I9���   f���   L���  t<��M��LƋL�^ȉ�I��M9���   H��h  H9�sb�    1���    �L��L�^��A���FD	�M�H��I��M9�wD�FE��D�FA��E	�E��H��h  H�M�H9�r�L9�sH��I9�u�)Ɖ2� 1�1��2ÐL9�w�D����fD  �v�A���W��� USH��H�/��x   ��   H�GH�WƇ�    �oG�oO(�oW8H���   ��   G`Op��   f����   �Obf����   H����P  ��   HcOpH���   H��H��H��?H��8 �  H���� ���H�H�CxH���   H��H��H��?H��8 �  H���� ���H�H���   H���   ƃ�   H��H��H��?H�� �  H���� ���H�H���   @����   1�H��[]��    Ƈ�   @��u�����f9�sIH�Spf���   H��H���   �oI��Hǃ�      H���   ǃ  ����H�C`H�CX1���    H�Khf���   H��H��Hǃ�      H���   �I��H���   ��    H�����   H������? ��H���{b���   H�Ch��Hc���H��HcSh�KbH�CpH���   H��H�H�� �  �S`H���� ���H�H���   �����    SH��H�?H���   �Gu,H��p  H�S���   ��t�����H���   [�f�     �+^��H��1�����1�[�ff.�     f�H��H��   �^���1�H����    �����   AW�   I��AVE1�AUI��ATI��U1�S��f�� @H��L�D$�>�    H��H��HN�H9���   H��H��HI�H9���   H����F��A��E97vWD��I�T� H��t�I�wH�4�H��tgH9�t�f��t�I�<�H9�|TL�L$I��H9�FH9�~)H)�H)�H��A���gF��E97w�H��[]A\A]A^A_� H��H)�H)�H��H���r���@ H��1�[]A\A]A^A_ø   ÐAWAVAUI��ATI��UH��S��H��H��&  H��u!H��(  H��uMH��[]A\A]A^A_�D  I�D$D��H���  H��I��N�48�E��I�T$H��(  I�N�4:H��t�I�D$H��H���  L��L�t�E��I�T$L�H�DH��[]A\A]A^A_�fD  AWAVAUATI��UH��S��H��H��&  H��t.H�D��H���   �@x��(��   ��#��   I�D$(L�H��(  H��tSH�E H���   �xx(u��+   ��   I�D$I��H���  H��I��N�l0��D��I�T$L�J�D2I\$(�H��[]A\A]A^A_��    ��+   �r���I�D$M��H���  H��I��N�48H�L$�gD��I�T$H�L$I�N�4:�8������,   �`�����-   u��R���D  AWAVAUATUH��SH��(��  ��  ���  �  �_VD�_TH�WHD�PD�wRL�OXf�\$H�_hL�W`L�gxD���   H�\$H�_pH�\$fD9��%  H��T$H��fD�yf�QH�T$fD�q
H�Q H�T$L�QH�Q(L�a0fD�i8fD�YL�IfA� H��I�L�H�t$I�RI�2H+PH+0���  H���  H��&  H��I���6C��H�t$L��H�H��(  H���  �C��H�E H��(1�[]A\A]A^A_�f����   D���   H���   D���   f�D$H���   D���   L���   H�D$H���   L���   L���   H�D$��D���   fD9���������   t�G�   1�fA� H��(�   []A\A]A^A_�f�     AWAVAUATUSH��H��(H��0  H9W ��   f��l   ��  �GT��   f9���   L�cXH����  I�Hk`f;��   �a  H��H��   H��A�   H�PH�0I+T$I+4$���  H�D$��  H��H��H��   H�PH�0H+UH+u ���  H��0  H�D$�   �    ���   H�C8��   Hǃ0     H�C@H��([]A\A]A^A_�f�     f��n   ����f��p   ����f9�s�L�ghH����  I�Ho`f;��   �  H�D$    E1�H�D$    H�C8H���s���H�S0H��H�C8L�<����   D9�wV���   ��   �C�   H��([]A\A]A^A_� �C�   �%���@ H�D$    A�   H�D$    �fD  D��I�$M�T$H��L���  E����   H��H��   H�L$H�VH�6L)�H)�H��A��H�L$I��H��   H��H�QH�1H+UH+u ���  1�I��M��tH�|$ L����   L)�A��H���   H�����  H�C8H��0  H�W�H��0  H��������D��� H���   L���  H�L$H���  H�H�2H�RI9�t_)�D)�Mc�Hc�Hc�Hc�I��H��H��H��H��?H��?H��0 �  H��: �  H��H��H��Hc�Hc�A��H�L$I���	����    L)�������     H�T$H�t$L��H�D$�	?��L�T$H������@ H���  H���  H��H��   M�$H�0H�PM�D$H���  H9�t[D)�D)�Hc�Hc�Hc�Hc�E1�H��H��H��H��H��?H��?H��> �  H��H��
 �  H��H��Hc�Hc���H�D$���� L)�L)�H��E1���H�D$����USH��H��H�oH�w0Ǉ       H���m���H�C0    H���  H��H�C(    �N���H���  H��Hǃ�      Hǃ�      �)���H�C    H��H��Hǃ�      ǃ�      H�    H��[]�����@ USH��H�/H��tvH�w0H��H�������H�C0    H�s(H������H�C(    H�sH������H�C    H�sH������H�C    H�s H������H�C     H�    H�C    H��[]�D  USH��H��H�H��  H���   H��t����Hǃ      H���  H���"���H���  H��Hǃ�      Hǃ�      �����1�H���  Hǃ�      f���  �����H��   H�������H��  H��Hǃ       ����Hǃ�       Hǃ      Hǃ      Hǃ      Hǃ  ����H��[]�fD  SH������ƃ�    [�ff.�      AUATUSH��H��H�vL���   H��tl���tVE1�f.�     D��L��A��H�,@H��H�t.����H�CL��H�H�@    H�p�����H�sH�D.    D9#w�L�������H�C    H�sH��tA�C��t*1�D  A��L���J�4�����H�sJ��    9kw�L������H�C    H��[]A\A]�f�AVAUATUSH���  H����  L���   H�CI��H�sL��(�<���H�C    H�sL���(���H�C    H�s(L������H�C(    H�sL��� ���H�s8H�C    H��tJ��t6D�m�1�I��I��D  H�t.L�������H�s8H�D.    H��L9�u�L������H�C8    H�sHH��tLL���D���H�CHL��H�p0����H�CHL��H�@0    H�p(�l���H�sHL��H�F(    �X���H�CH    H�sXH��tLL�������H�CXL��H�p0�/���H�CXL��H�@0    H�p(����H�sXL��H�F(    ����H�CX    H�s`H��t8H��L������H�C`L��H�p(�����H�s`L��H�F(    �����H�C`    H�spL������H�Cp    H���   L������H��L��Hǃ�       []A\A]A^�y���f�     []A\A]A^��    L�1�M9�r�D  ATI��L��UH��L��SI��H��   H��M�$L�L$�A���I�$�D$��uH�+H��[]A\�f�     UH��SH��H��H�7H�WH���6  ���   �o��   f���o��   �o��   ���  ���   �o��   �o��   ���  ��  ���  ��  ���  H��   H���  H��  H���  H���   ��  H���  H�BX��  �o��  ��  ��  �oX�  ��  �o` ��  H�@0H���  ��  �o�   �o�0  ���  ��  �o�@  �o�P  �  ���  H���  �o�`  �o�p  �  �o��  �o��  �(  �o��  H���  H���  �o��  �(  �8  H���  ���  �  f��8  H���  �H  �X  �h  H��@  �H  �o��  �o��  �o�   GH�X  �h  �x  GXGhGx��   ��   ��   ��   ��   ��   ��   ��   H�C(H�{�   H�K0H�t$H�D$���  L�@ �#���H�T$H�S(���
   H��[]� ���  H�{�   H���  D���  H�t$H�D$������T$���  ��u��o�  �o�(  ǃ      �o�  �o�8  ƃ`   ��   ��   ��   ��   ��   ��   ��   ��   [HSXKhCxH��[]�ff.�     �AUH��A��ATUH��SH��L�'H��  L��H���x������f  ƃ`   D���  I��$(  I��$0  H�C     ǃ�      H��  H��   Hǃ(      Hǃ0      H���  1҉�  H�       @H�   @   @f��(  ���  H��  �   �o�8  H��   �o�H  f��p  �o�  �o�X  �o�  ǃl    �o�h  �o�  Hǃ0     �o�(  ���   ���  �P  �o�(  �`  ��  ���  �p  ��  ���  ��  ��  ��  ��  �   �0  �@  H��[]A\A]��    H���  H��H���  Hǃ�      ǃx     A��$H  ����D  AVAUA��ATUSH�H��H���   H���   H�GL��  M��~���   H���   H���t H���   H�SH��  �o�P  �o�`  �o�p  �o��  �  �o��  �(  �o��  �8  �H  �X  �h  E���e  H�RXH�JH�RH���  H���  ���   H��H�L�H�9H�W H���H�H�L�H�9H�W H���H�H�L�H�yH�W H���H�QH�T�H�BH�� H���H�BM��[�}x(��  ���   H���   H���ot�)sp�o|�)��   �oD��8  �oL�1��H  []A\A]A^� H��  H�CL�ppD���  fo��   H���  L��0  �  fo��   H��(  �  fo��   �(  fo�   H���  �   �8  L���  HǇ�      Ǉx     _HWXOhGx��   ��   ��   ��   ��   ��   ��   ��   Ǉl    f��p  H�Ǉ"   @  Ǉ&   @  Ǉ   @  Ǉ@     HǇ0     H�G     Ǉ�      ��H  H��  ��t���   �������h  ��A
��A��}x(�E���H��  1���+   �/���[]A\A]A^��    ���   H���   Hǀ�     Hǀ�     H���q H���   �|����    ATH��A��UH��SH�_0H��������t[]A\�fD  D��H��譁����u�H�S@H��X  H�SH[H��`  ]A\�ff.�      H�0������    AWAVAUATI��UH��SH��H��(L�o8�    �D$    ����H�$��������   D���\  D��H9���   A�NL�L$E1�1Ҿ   L��补��H�$�D$����   D�31�1�E��tD  L��蘂��H�$A�ǉ؃�L�,BE����   A��L��D$�o������fA�m E��thH�4$D�l$��L�<FA��@ I��D9�t?L����4������fA�/A9�w�H�$H��([]A\A]A^A_� H�$    ��fD  D���X���A9��O�����D  A��L��A�ǉD$�����fA�m E��t�H�$D�l$��L�<BA��@ I��D9�t�L���輁���fA�/A9�w��f���A��L��聁��A����A��A	�D��H9�������R���f�AW��AVAUATUSH��(H�G8�D$    H�D$H9��&  ��I��L�L$E1�1Ҿ   H��������L$I�Ņ���   1ۅ�tbD  L�������A��A��?����   �@uU9���   E1�f.�     L��A���Ā���Kf�fA�D] ��E9�r9�wމ�E9�v9�r�H��(L��[]A\A]A^A_Ð9�vdE1�f�     L��A��蔀���KfA�D] ��E9�r�9�w��fD  9�v,E1���C1�A��fA�T] ��E9�r9�w�������    H�|$L��E1�������p��� E1��e����     H���  H��u��$  f��uH���  H���  H���fD  ��"  H���  f��uH���  H���f�SH�����  �������A������Hc�Ic��َ��H���  [�ATI��UH��SH���n���L��H����,��H���  H�[]A\� ATI��UH��SH���>���H���  H��H��J���,��H�[]A\�UH��SH��H������H���  H�Hc�H��[]H��H�H�� �  H��H���    SH����������  [H�H��H�H�� �  H���f.�     AWAVAUATUH��SH��(D�<H��X  L��`  L�gE��E����  A�D$A�T$`�D�A;D$�   A���  ��  M�D$xI��I�<@C�D?H�H�I9���  ������A	�E��~fA� f����  I�PH�YH9�sP�qH�Y��A���qD	�fA�pf9�|(�p  f�H���C������C�	�f�f9��O  ��H��H9�r�E����  D�z�A���,  D��A�L$A�D$b�D�A;D$�n  H�EL�SHǀ      Hǀ       M9���  ��[��	�D���E ��   L��L)�L9���  H��  �   M��H�t$L�T$���  H���  L�$H�|$H�x�V���H��  �L$���  ���o  H�EL�$f��H���  L�T$L��  H��   t%L��L��L�L$L�$�j L�L$L�$�     M�D$pM�Mc�O�M9��v  I�qI9���   A�I�@A����_  L��L��L)�L)�L�I��' H�~I9���   �W�H���P����/  H��H9�u�I�T$hI��M��N�I9���   I�t$pL9���  1��4@ L�AM9�wm�	�uGH)�L��H�:���H��H���F�I9��  ��uɨu�L�AM9�w2D��IA��D	�H��H�L���f�     H�AM�D$xI9�s�   H��([]A\A]A^A_�fD  �L�������A	��&���f�1�D��L��H�$����H�$�������봐1�E1��{���fD  1�A�wL���������|����H��L��f�L�NM9��q����7H��H�I9��_�������   ����L�DfD  H���P�L9�u��&����   �0���I�T$hI�t$pI�I9�vo1��8�    L�AM9������	� uHH)�L��H�z��H��H���F�I9�v3��uȨ u�L�AM9������D��IA��D	�H��H�L���fE�|$b1�fE�t$`H��X  ����L�������I���q���f�H��(  H�8�1����H���  AUATUSH��H��H��X  L���   H���   L��p  H��t	H��P  ��M��tH��A�T$H���   H���  �w��L���   Hǃ�      H���  I�|$8����H���  L��Hǃ�      �Sw��H��@  L�������H��   H��Hǃ@      Hǃ8      �w��H��0  H���w��H��Hǃ      Hǃ(      �2���Hǃ�      H��[]A\A]�@ ��    AWAVAUATUSH��xL���  H�^8�D$d    M��t+H��@   H��tH��I��H�L$h�ravc��@  �D$\��t_�D$\    E1�E1�E1�H�$    L��H������L��H��� ���H�4$H�������L��H��������D$\H��x[]A\A]A^A_�fD  H�t$hL���Cv���D$\��u�I�D$@L��H�D$I�$H�D$�x��H=   t(L���D$\    E1�E1��w��E1�H�$    �\���f�A�M H��L�L$\E1�1Ҿ   �u����|$\I�ƅ�t"L��E1��?w��E1�H�$    �����    A�M �   L�L$\1�E1�H���-����t$\H�$��tL��E1���v��E1������fD  A�M H��L�L$\E1�1Ҿ   �����L$\L��I�ǅ��8  �w��L��T$�w���T$H�t$h��A��fA���A���D$4��H�H9���  H�D$H+D$H�H�D$f����  E1�fE���E  H�D$     �D$    L�T$HH�\$8H�l$@@ L���v��L��f�D$�{v����f����  ��%�  A;Eh�P  A�U L��H��H����I�MpH�4��d ��@��  H�$��M��L��L���S����l$Hl$H��H�l$H���5  I�$I�T$@H�|$H)�H�T$(I�T$HH��H)�H�H9�H�t$hHG�I�T$@�� ��  �T$dH�\$H�T$`��uH�D$@��8  L��H�L$�!���H��H���  H���  H�|$ ��D$`H�L$�  ��tXL�T$@D�@�1�Hc�M��8  �@ H���SL9�s(H�DU I��@  H��I��I��?J�� �  H��fNH�BL9�u�H�t$ H�|$8����H�D$     H�|$8H������I�D$HI�$H�\$(H��H)�H�H9�HG�I�D$@H�T$�D$�D$H�T$9D$4�&���L�T$HH�\$8L��L�T$�?t��L�T$I����%������� H�|$ ��a���H�D$ �����k���fD  A�E ���$���1�f�\$(��H�,$�    L���@t���ك����H�H�D� A�E 9�w��\$(�������1�f�     L���t��������H�I��A9m w������D$\   L���~s��E1��`���H�T$`L��H�L$�t����T$`H�t$hH�D$ H��H�L$�����A�U 1���Z��� L���s��������H�I��A9m w��5���H�T$@L��8  L9������M�������H�D$@Hc�1�H��@  1�D  H�TE H��I��I��?J��
 �  H��fG�FH��I9�w�����L�T$HH�\$8�D$\   �^���I�T$HI�$D�D$H�|$M�L$@H��H)�I)�H�H9�L��L�L$HG�I�T$@H�T$d�f���I�T$@L�L$I��I�$D�D$H)�H�T$I�T$HH��H)�L�L9�HG�I�T$@fE������������L��L�T$�r��L�T$������     AUH��ATI��USH��H��H�n8� tvcH�L$��@  �D$��t)Hǃ8      1�Hǃ@      H��[]A\A]�fD  H�L$L�L$E1�1Ҿ   H��H��H��8  蒔��H��@  �D$��u�H��8  L��H�4 ��o���D$��u�H��@  H��8  L�lE L9�sL��H���q��f�E�I9�w�L���q����y   �D$�Y���L��H���w����I���f�AW�ravaAVAUATUSH��(H���   L���  �D$    H�L$L�k8H��A�D$0��@  �D$��tH��([]A\A]A^A_��     H�t$H���o���D$��u�H���cq��H��H���Xq��H��H�D$H��   tH���Op��H��([]A\A]A^A_�I�D$� H9�u�H��L�L$E1�I�־   1�L���7����T$I��I�D$8��u�M��t�H�$    f.�     H��Hc,$�Dp����fA�H��    H;D$��   L�L$E1�1Ҿ   L���Ӓ��I�G�D$��ul1�fA�? tFfD  H��I��H����o��I�OI��H�ߘ��H�J�1��o��I�O���H�J�D1A�9��H�$I��H�$H9D$�P���������E�I�t$8���tBLc�H�$I����H)�H��H�� D  J�t>L������I�t$8J�D>    I��L9�u�L������I�D$8    ����fD  AWAVAUI��ATI��USH��8H���   L���  H��H�k8�2k���D$,��t*E1�L��H��茺���D$,H��8[]A\A]A^A_�f�     H�t$,H���p���T$,��u�f��t�D$,   � H�t$,H����t��H�D$�D$,��u�H�t$,H����o��D�|$,��A�U E���r�����t���L�L$,E1�1Ҿ   H������D�\$,I��E���F���E�U E��tA1�f���H�t$,H�߉T$I��H�$�Et��H�$D�L$,H�E���	����T$��A9U w�H�t$H��L��j���D$,�������H�t$,H���o��D�D$,fA�EE�������H��H�t$,��n���|$,��A�U�������I�VA�M;
t�D$,   ����E1�1��Ⱦ   L�L$,H���#����|$, I�E�]����D$    �D$A9E��   D�t$I�EE1�1�A�ML�L$,�   H��N��L�$�я��L�$�|$, I�����I�EfA�} N�4���   �$    H�t$,H���'n���t$,f�D$�������H�t$,H���	n���L$,f�D$�������H�t$,H����m���T$,�������H�T$H���$I��H���$H��I�F�A�EI�V�H�T$H��I�V�9��k����D$�����A�M E1�1�L�L$,�   H�������|$, I�E�$����$    �$A9E �����$H��I�4�Lk�MuL��h���D$,�������H�t$,H���$m���|$, ��A������H�t$,H���m���|$, ���D$�����H�t$,H����l���|$, ��A�V�����;T$�����A;U�����E1�1��Ⱦ   L�L$,H�������|$, I�F�Q���1��:H�t$,H�߉T$�l���L$I�v�����|$, H��� ���A;E�������A�F9�w���A�E1�1�L�L$,�   H��襍���|$, I�F�����1�A�A�F9�vPE1��>H�t$,H��D�D$�L$�T$��k���|$, ������T$I�vD�D$�L$f�VA��B�D;D$r��A�$�[���H�t$,H�߉L$�T$�*k���|$, �X����|$I�vf��L$f�~H������)�A9Fw����R���fD  AWAVE1�AUATI��USH��L��X  H��`  H�_�   D  ��L�H9��1  A�M����  fE����  E�E��D	�M�E�ɉHA�M��A��A�MD	��ɉHf���  A�M�hE1�E1҉�A�H��	�H��H��H�σ� H�HE��L�PL�H H�x(�1  E�~H��D�������ƅ���   M�EL9�rK�vH��H��   H�@    A�U A�M��	�f�PA�}A��A������A�}	�fA����ɉ8����׃�f���������@��   ��L�H9�������    �   H����[]A\A]A^A_�f.�     ��@��   A�M�hE1҉�A�H��	�A�xH����H��A��A�xD	�E1�H��H�������D  ��fE����   E�E��D	�M�E�ɉHA�M��A��A�MD	��ɉH�e���D�Q�IE������HA�MM�E�H�A���@ ���   A�E�HM�hE�P��A�H��	�D��E�H��H��A	�D��E�PH����M��A	�A�xI��M����I��A��A�xD	�H��H�������D  �HA�MM�E�H����@ M��E1ɿ   E1ҹ   �����     D���   I�|$0�t$��c��M��$X  �t$L�H)�I��$   �A���ff.�     �I���   �l1H ��� ����t�   ��    A�Hx�
Ð���   tH��p  ��   H���   ��f��h  �t6���  )�f����  ���  ����)�)�9�H�fA� �f�     ���  )�f����  ���  ��@ AV1�1�1�AUA��1�ATUSH��H��L�g0H�/f�T$
L��f�L$f�t$f�D$��b��1�L�D$D��I��H��p  H�L$H�����   H�SXD��H��L�D$H�L$
����L��L����a����u3�T$�L$
�{l �S`�T$��0  �L$�Sd��4  u�Cl�ShH��[]A\A]A^�f�     AWAVAUATI��US��H��H�G%  ���toH����   �   A��$�  t?��t9L��D�<L�t$L�l$���M��L��1�L���H���G����D$H�E�D9�u�1�H��[]A\A]A^A_��     H��t{�   A��$�  tԅ�t�L��D�<L�t$L�l$fD  I��$p  ��M��L��1�L���H�����   �D$H�E�A9�u��fD  �G��(����3���f�     �G��{����@ H���  H��t4H��t�8�>H��tH�pH�2H��tH�PH�M��tH�@I� 1��@ H��t�    H��tH�    M��t�I�     1��f.�     Hc�H��H�H���  H��t:H��   H9�|H���  1�H���  H���  ��x  ��G�   �   � �G�   �   � ���  H���  H��H��H9���   ���  �f�     H��(H9�vw:Hu�x t�Hc��  ;��  }e�JH���  H��I�����  ��x  H��  �
H�N�0H�JH�B   H�B�V���w)H�P� ���Aƀ�   ��    �G�   ��G�   ��G�   ���    H�B H��xH�    H���HH��fD  H)�    H���H��H��HO��f�     H��xH�2�    H���H�� HH��D  H)�H������H���H��H)�H��HO��@ H��xH��    H���HH��f�     H�к    H)�H���H��H��HO��fD  H�B?H��xH�    H���HH��fD  H)�    H���H��H��HO��f�     H�BH��xH�    H���HH��fD  H)�    H���H��H��HO��f�     L��P  H��X  H��H  L)�H��H�H��H��xH�1H!�L�IH�� H)�H��H!�H��L)�I��H��IO��ff.�      L��P  H��X  L)�H�H��H  H��xH�H�H��H��L�IH�� H)�H�H��H��H��L)�I��H��IO��ff.�     H�H��uH�8 tAH��  H���  x1Hc��  ��~H��H��  H�R�H;BƇ�   H�> x� �G�   ��     H��@  H��H��@  H;�H  v��G�   �ff.�     f�f��&   t3H�H���   �xx(tf��H��H��   HE��t��H��   �f��(   t4H�H���   �xx(t9��H��H��   HHE��t��H��   ��@ ��+   u��D  ��+   t���,   t���-   u�� AWAVAUI��ATUSH��H����  f;��   �h  f9GT�^  ��H��L��8  H���  H��f��l   tf��n   �}  H���   HCXH��H�H�VH�6H+PH+0��I��H��P  H��~-H��X  H�L9�~H��H)�I9�~H��H��M��HH�I��f����  H��H����  ���   L��H�����  I�����  tM����   I��M9�MO���  H��   H��H�UH�u H��HC`H+PH+0���  L��A��H��H)�H���   ���  ��  f��  fD��  ���  tfD��  H��[]A\A]A^A_�f.�     ���   t��C�   �fD  ��M����   M��Iֺ    LH���=���M9�ML��1���f�     H���   HGhL���  H���  H�L�L�HH�2H�RI9��}   D)�D)�Mc�Hc�Hc�Hc�I��H��H��H��H��?H��?H�� �  H��: �  H��H��H��Hc�Hc���I���!���f.�     I)׺    M��M��LO���~����o����L)�L)�H����Hc��  H�H��H�L�� �  I��Mc������f�AWHc�A��AVH��I��M��AUA�Չ�H��AT)�E��UH�D1�SH��8�t$H�|$H�D$D�\$Ic�Ic�I�I�H��H��I�I�<I�M�$I��I��I)�M)�L9���   H��H)�L�L$(L)�D�T$$D�D$ H�$�A	��H�$L��t$D�D$ D�T$$M��I��H��H��L��L�L$(I��D��E��A��9t$|^H�t$H�H�$I�6I�1H�t$H��L��D  L�H��H�H��H9�t%H�H9�~�L9�|`L�H��H��H�A�H9�u�@ H��H�������H��8[]A\A]A^A_� uH9�u�L9�uB1��t$9t$�f�����f.�     )�H�H�$I��I��?J�� �  H��H�H��]���L��M��I��H��H��H��L��I��H��D��E��A�������AWAVAUATUSH���   L���   ��y   L���  Ǆ$�       M�}8��   M����   1�A9vx��   M���   ��nI�4�I94�t~A�̉L$@E1��   H�T$L��$�   L��1�H�|$ L����|��D��$�   H�D$E��tjH�$    H�D$    H�t$L��謥��H�t$L��蟥��H�4$L��蓥����$�   H���   []A\A]A^A_�f.�     �   ��f�     L��$�   E1�L��1Ҿ   L���c|��D��$�   H�$    H�D$E���l���E1�L��$�   L��1Ҿ   L���(|��D��$�   H�$E���:���I���   L��H�4��pU����$�   ������I���   L��H�4�H+4��:W����$�   �������A�L��L��$�   1�E1��   I�]@I�m �{����$�   H�D$(����  A��   E1�1�L��$�   L���u{����$�   H�D$0���I  A�L��$�   E1�1Ҿ   L���D{����$�   H�D$H    H�D$8���!  L���_X��L��T$D�QX���T$DI���   D��A��fA���A����$�   ��L�H9��G	  H)�I�f���]	  �|$@ t1H�D$H�t$H�H�D$@�P�1�H��H���oH��H9�u�fE���:  �\$@H�,$L�|$pH�D$X    �C��D$D    ��$�   H��$�   H��H��H��$�   �C���$�   �C���$�   �C���$�   L���hW��L��f�D$P�[W����f���[  ��%�  A;Fh�w  A�H�|$(H��H����I�NpH�4���D ��@�c  L�D$8H�L$0��L��H�T$(�-���D�|$PI��K�'H�D$PM���.  I�E I�U@I���   H)�H�T$xI�UHH��H)�L�L9�HG�I�U@�� ��  ��$�   H�\$H��$�   D�|$@��L��L��$�   AD��������$�   I���   L��I��H�D$`��AD������H����M��H��H�D$h����(  H��L��$�   �  H����@  1��|$@ H��t+H�L$H��$�   H�|$� �oH��H��H9�u�1Ƀ�$�    Ic�tyL�L$L�T$`L�\$hD�D$@���<sH��D9�sK�D= I�<rH��I�4sL�H��H��I��I��?J��' �  H��H:H��H��?H��> �  H��Hr��9�$�   w�H�D$f�8 ��   H�\$E1�E1�L��$�   L��$�   E��H��H��$�   H�HI���QD9�|AIcր|  H��$�   ��  A�VHc��f�     H���|� ��  A��9�}�A��A��fD;|�L��$�   L��$�   1�1҃|$@ ��   H�|$L�D$D��$�   D��$�   H�\$ L�T$D�\$@�I�JH�H1Ly��H��A9�tUH�LI+L H�4I��I+4 D9�r��  A9���  9�$�   �@  9�$�   u����  u�I�JH�Ly�H�|$X�tH�t$XH�|$p蝟��H�D$X    H�\$pH�t$`H��肟��H�t$hH���u���I�EHI�U H�\$xH��H)�H�H9�HG�I�E@�D$DL�d$P�D$D9�$�   �)���L�|$pH�|$H�uFH�t$(L������H�t$0L������H�t$8L������L����R���?���H�D$H    H�D$8    H�t$HL���ٞ���H�D$H    H�D$8    H�D$0    ��E��E�UE��Mc�D9��r  fD��$�   ��D��H��I��L��A��� L�L$L�D$���7�����H��A9���   �<+ t�u��z9�~Љ���A��������E1�L��f�\$`H�\$0I��D��I��L���R��������H�H��A�9�w�L���\$`M�����H���E1�L��H�\$8I��D��I�� L���@R��������H�H��A9.w�L���\$`M������H��L��D��A��D��$�   E�T$D9��g  �zA9�|EL�L$L�D$D��D��H��$�   D��$�   D��$�   �$���H��$�   D��$�   D��$�   E����  A�u�A9���  L�L$L�D$D��D��D��H��$�   D��$�   D��$�   �����D��$�   D��$�   H��$�   E���o������  �����I�JH�H1����H��$�   L��L�D$`�������$�   L�D$`H�D$XI���   H���^���A�E1��������f�D$`H�\$(L��I��D��I�ǐL����P��������H�H��A9.w�L���\$`M���������  �W����Y���Mc�H�T$L��H��H�HL$H�2H+1H�zH+yH��H	�tjE9�~:L��$�   A��G�>L��M�H��I��HL$L�$�   H1HyH��I9�u�A9�}&�K�D)�L�H��H�$�   HrHzH��H9�u�E���������   �����������|$@ �����Ic�1�L�L$`L�T$hL��$�   D��$�   H�|$ H�t$�$I��I��LfI$IL$H�JI9��v���H��I�QH��H��H��?H�� �  I�RH��H��I��I��?J��! �  A��H��A9�w�t;D9�$�   tMD9�$�   tND9�$�   u����  u�H��H��H^HK�s������  u�H��H��HNH�W������  u������   u��Ǆ$�      ����Ǆ$�      L�|$p����I�EHI�U I�]@H��H)�H)�L9�vJ�"I�E@H��$�   L��D�D$D�,���I�U M�e@H�D$HI�EHI)�D�D$DH��H)�H9�vH�I�E@�;���ff.�     AWAVAUI��ATA��U��S��H��h  H�GL�7Ǆ$�       H�D$A���  9�sfA���  A�](A�E u_I�EH�@XH�HH�@H�D$I���   H�L$H�@hH��tWH�xH� H��$�   �����$�   ���c  H��h  []A\A]A^A_ÐH�D$   I���   H�D$   H�@hH��u�I�U8��L��E1�����A�M8���y  �D$  ����  fA�}< ��  L���p������)���fA�}< �-  L��A��`  ��$�   ���  L��A��P  M�efAoMpI�L$bI�T$hH��H��fAo��   T�Ao�8  \ �Ao�H  d0I�T$p�
 I�T$p�D
 I�T$p�D
 I�T$p�D
 I�} ��H�G  �u�G�tPA�u(I�T$`����I�} ���  ��uI�t$hH�L+A�Mh��uI�L$hH�T0+T A��4  ���^  I�E I�t$hH�Ń���  H�K@�uqI�EH�H�@XL�HL�@H9�vYMc�Mc�H��@ HcH��I��I��I��?J�� �  H��Hc�H�P�HcP�I��I��I��?J�� �  H��Hc�H�P�H9�w����  ��  H���  ���  fA���   1�L���B�����$�   ����    H�|$����   �Hc�$�   L��$  H��$�   f��L��)�$  A�U8)�$   )�$0  )�$@  )�$P  ��F��A�M8M�}01�A�   �������I��p  H����  H�L��A��H  ��$�   ��u#L��A��X  ��$�   ����  L��A��P  E��tI���   H��$�   H�@hH�xH� �P��$�   ����D  I�E@    ��L��I�EP    I�EH    I�EX    �������$�   ���/  A���%  L���M���������I�F  ��x  A�F��m  A�E ��   Hct$IcEpH��H�H�� �  H��H�I�EpIc��   H��H�H�� �  H��H�I���   Ic�8  H��H�H�� �  HcT$H��H�I��8  Ic�@  H��H��H��?H�� �  H��H�I��@  Ic�H  H��H��H��?H�� �  H��H�I��H  Ic�P  H��H��H��?H�� �  H��H�I��P  Ǆ$�       �     �|$  �P����U���I���   H�~h ����Ǆ$�      �3���fD  ��L���~�����$�   ���
���A��� ���A�M8�D$ �;����    H�     I�} �   ��H��$�   I�EpH��$�   Ǆ$�   H��$�   I�ExǄ$�     H��$�   I���   H��$�   I���   H��$�   I��8  H��$�   I��@  H��$�   I��H  H��$   I��P  H��$  H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   �������$�   �������H��$�   H��$  H��$�   H��$�   I�ExH��$�   I��P  I�M I���   H��$�   H��$�   ���  I�}pI��@  H��$   I���   I��8  I��H  ��u)�A�Uh������)�A��4  ����������I���   �����A��I��h  fA�M<M��h  H�D$(H��t"����  ���
f�����  H�R��H��u�L��L��L�D$0�\���L�D$0H���P  Ǆ$�      �~���fD  �o,A)mp�otA)��   ���   �o| A�8  �o|0A�H  H�������Ǆ$�       �����A�T$`A�D$bE1�I��$�   fA���   I��$�   fA���   I���   I�T$pI���   I���   I�T$xI���   I��   H�PfE��  H���m3 I�E I�t$hI�} H�Ń��}���H�������ol A�8  �ot0A�H  �=���H��$�   H���F���苄$�   ����  I�U f;��  �[  �ո   A;U8�U  I��  �   I��H��$�   ���  H�xH��$�   H���  �$���I��  ��$�   ��$�   ���  ����   H���  H��H���B����$�   ����   I��  I�E�\$Z�|$xH���  H��  H��   I�U�BH�r@)�fA���   �B)�fA���   �D$\H��HB(H��H�I���   H�r H�HJHI���   ��H�HB01�I���   I���   I��   fA��  �I���   H�H��� �A���   ��9�w���   L��fA���   褼����$�   �-���H��H������fD  H�pH�@H��u�L��L��H�T$0�[���H�T$0H�������L�bH�D$L���H�@f�L$Zf�D$xA��h  ��$�   ���Y���I��   L��H�D$`A��P  I�F  �uA�F��y  H�D$1�E1��   L��$�   ���   HǄ$�       HǄ$�       �ωL$ HǄ$�       �GH�|$(H��f��$�   f��$�   �ve����$�   I�ą���  H�|$(E1�1Ҿ   H��$�   L��$�   �?e����$�    H�D$0�_  H�|$(E1�1Ҿ   H��$�   L��$�   �e����$�    �,  �L$ H�t$L�T$0f��A��H���   �A	  L��1�Hc~H��H��0H�y�Hc~�H�y�A�f�PH��fA9���T$ H��I�}pD�D$0H��H��L�H�9I�}xH�y�zA�2M���   f�pH��H��H��L�L�	M���   L�IA�2M��8  f�<p�z��H��H��H��L�L�	M��@  L�IA�2f�<pH��I��H  H��H��L�H�9I��P  H�yL��A�2f�p��$�   H��$�   ��L��$�   L��$�   H��$�   �)�����$�   ����   H�D$H���   �D$ f����  ��D�D$0L����H��Hk�0H��Bt�1�r�q�rH��0H��H9�u�I��H��I�I�LH�:H�RI�t I�UxI�}pH�H�II���   I���   H�H�vI��8  I��@  I�t0H�H�vI��P  A���  I��H  @��u)�A�Uh@��u	)�A��4  H�\$(H��$�   H��蘋��H��$�   H��HǄ$�       �|���H��$�   H��HǄ$�       �`�����$�   HǄ$�       ������I�E ���   Hc|$IcUpHct$H��H��H��?H��
 �  H��Hc�I�UpIc��   H��H��H��?H��
 �  H��Hc�I���   Ic�8  H��H��H��?H��
 �  H��Hc�I��8  Ic�@  H��H��H��?H��
 �  H��Hc�I��@  Ic�H  H��H��H��H��?H�� �  H��Hc�I��H  Ic�P  H��H��H��H��?H�� �  H��Hc�I��P  ����  H�D$I�M0D���   H�ǋXPH�L$pA�M8�L$|�����E���C  A�D$��L$ZL�[D�|${H�DI��L�t$hL��H�@�L$\�ML�t$H���L$LM��H�D$P�kA�D$E�T$\D9��K  A9��B  I�t$ ��L��H��H��H�H�L� L�hL+"L+jL��L	��s  Ǆ$�       I��0L;|$P�  H�CxH��H  L��P  H���   H��@  D�KhH�D$ I�FXH�T$8D��4  �T$LL�\$@B�48E�^H�L$(1�L�kpH�|$0H��L���   H��8  D�L$D�D$D�\$�������$�   ���W  I�NXD�\$L��A��u`H�t$ H�|$0L�kpH�T$8D�L$L���   H�sxH�t$(D�D$H��8  H���   H�t$@H��@  H��H  H��P  D�KhD��4  A�nA9������L�cD��A��H��IT$ H��$�   A�T$D)�f��$�   A���   ��   �QLci��;�����D	������Lc�E��t	����  H�S ���W���H�CH�pXHcFL��L��H��?M�� �  HcFI��L��Mc�L��H��?M�� �  I��Mc��A�	������ ���H�H���   �xx#uI�� I���I�� I���������ol A�8  �ot0A�H  ����H�qH��$�   D�D$D�\$H�L$�d.��H�L$D�D$D�\$�A�����L��L��H�L$H��$�   �,��H�L$Ǆ$�       �k���H�|$(�   L�D$0H��$�   �K����$�    ����L�D$0L�`H��L��������r���H�|$�A���I�Eǀ�   pmoc�C���D�|${L�t$h�3���D�|${L�t$hǄ$�      ����H�D$pD�|${I��L�t$hH�C0�D$|�C8H�D$`H��   �C ������A�����9l$\�����H�[�Cf���t�Sb�TB;S�<  Ǆ$�       H�KH�S fAo}pH��H��<fAo��   |�Ao�8  | �Ao�H  |0H�C(� H�CH�S(�D H�CH�S(�D H�CH�S(�D I�]0I��   H����5����$�   ���9����������H�qH�yH�L$�H��H�L$H�D$H�q H�y(�H��HcT$H�L$H�L��L��L��L��H��?H��?M�� �  M�� �  I��I��Mc�Mc������H�D$pI�E0�D$|A�E8H�D$`I��   �u����p1�H���\����$�   ��� �������E1��?���1������f������I��  �����ff.�     AW��AVH�@AUATUSH��8H�FL�Љ�A�@M�P��H�T$����  I��I��1�E1��    I�@E��fA�} B��I�EH�,��Y  E1�   �H�E H�uH9��  H�}H9��  H��H��A��H��?A��t	H����   H����   I�H�RJ��H9�|H9�~p1�fD  A�EI��H��D9�w�Lt$A��K�rH��H��H��H��?H�� �  H��H�H�E;x�.���H��8�� �  [��]A\A]A^A_�fD  H9�tcL�L$(H�L$ L�T$L�D$~wH��H)�H)�����L�D$L�T$H�H�L$ L�L$(H��H��H��?H�� �  H��Hc��:���f.�     H��H��H��?H�� �  H������@ �   ����H��H)�H)�H���H��81�[]A\A]A^A_��    AW��E��AVH��I��I��AUATA��US��H��8H�L�N�M9�~H��L��I��L��M��I��I�vI�N�L�<L�,J� L��M��L�$L)�I)�M9�tvM9�tqH�D$    E1�A9�rML��L�T$I��E1�H���D  Hȃ�H�.A9�r&I���H��H�(I9�}�I9�jL���H�.A9�s�H��8[]A\A]A^A_�@ A9�r��H��L�8M9�|"@ IɃ�L�>D9�wƉ�H��L�8M9�}�O�L9�MO�M����f�E��t;�/Mc�D)�H�I��I��I��?J�� �  A�   H��H�H��<���f�     H�t$H�<$L�D$(H�L$ L)�H)�L�L$H�T$�h���I�~I�vI��L�D$(H�L$ L�L$H�T$�y���@ AWAVAUATUSH��HH�H���   �xx(��   f��   �  ���  �  H��  A�   H��H�D$ H��   H��H�D$(H��(  H��H�D$0��  I��E1�E1҉T$8f�     I��8  I���,AA��@  )ōB�9�F�A9�w0I��0  E��D��F�,t�   f���D�,��   ��9�v�A��A��fE9�  ~IA��  뒀�+   ������,   t	��-   u ��  ���  ��  Ƈ,  f��uH��H[]A\A]A^A_�H��  A�   H�D$ H��   H�D$(H��(  H�D$0�����D  �CA��A��9�vb�   fD  �L$8D9�vdD9�v_D��E��H�|$ �D$L�\$E��D�L$D�T$�t���D�T$D�L$L�\$�D$A��A9�w)I��0  D��D�,
t�A�T$�A�w9�v�E��A��A9�v�A9�t|A�w��9�w3�D$89�v+A9�s&A��D����D�L$H�|$ D�T$�����D�L$D�T$��tX�S�D9�rP�D$89�vHA9�sCD��A��D��D�L$H�|$ ����E��D�L$�T���H�t$(��H�|$ H��H�H+u@ E���.���A9�s@A��L��A�<H��I�H�I��J�|fD  H
H��H9�u�9�r���H��H9�s�E�������Ƈ-  f���$�������f�ATI��USH��H��H�?�GtIH��p  H�T$���   �Ņ���   �����H�;H���   L������H��@uH����[]A\�f�1���@ 1�H�������Ņ�u�H�CXA�T$�Hf9AGT$A�<$t��u�H   ���   �Ҿ   ����H���   H����[]A\�D  H�t$H��軕��H����[��]A\�ff.�      AWAVI��AUATUSH��H�oH�|$�M H�]9�F�t$��t|I��D�f�E1��$fD  �"  K��    H��0I�GM9�tLI��H�sK�D� H��H9�H9CHMCH��H�CH9�~�H�sH)�H��0H)�����H��K��I�GM9�u��M H�D$�\$L�`89��  ����)�I��H�I�T�fD  H�     H��H9�u�M��teE1�E�$A��vIM�T$D��A�   1�M�<�I�?I�RI�B I�JH9�~�e H��H�@H�P�H9�HA��A�pA9�u�A��I��D;m r�H��[]A\A]A^A_��    H)�H)�����K�������@ D��H��I�I�H�qA��I��I+rH)�H)�����I�T$�HDI�D;m �1����M��t���t������AWAVAUI��ATUSH���   H���   L���  H�t$H���   H�D$Ǆ$�       M����  �D$@ E�'E1�D��A�MH�DH����L$8H�D$ H�[H��H�D$(��H��H�D$��A��H��H��    H�D$0M���u  H�|$ �*  I���  H�|$H��$�   H�p ��>��H����$�   ���  I���  H��H�P H�p�� H�T$(H�|$H��H�D$ D�AH�D H�H�AH�QH�E��t,A��H��H��I��N�Df�     H�>H��H�L9�u�H�t$Ht$0H�E��tpA�t$�H�|�H��=H��htdw�{  H��zspo�~  H��tnlsuH� �1H fD  H��H��0H9�t$H�p H�H��thgwu�H��H� �1H H��0H9�u�H�D$H���$�   H���   []A\A]A^A_�fD  H��$�   H��ravg��@  ��$�   ��t%H��$�   H��2FFCL��A��@  ��$�   ��u�H��$�   H��ravfL��A��@  ��$�   ���y���H���)��H��$�   � 7H H��I���5����$�   ���J���H�|$H��$�   ��   ��$�   D��$�   ��<��I���  ��$�   ������B��   D��$�   9��D$@�a����    H� %DH ����@ H� �1H ����@ H�|$C��H�L$HH��$�   H�t Ht$(Ht$ I���  Ht$0H�|$H�p �I<��H��H�D$P��$�   ���r���H�T$ L� H�L$(I���  D�T$8L�L�
H�xE��H�L$HD�'�G����D�WH�WL�_H�|$I�4;t3�|$8L��    L�؃�H��H��L��    H�0H��L�H9�u���$�   H�D$HD$0I�L�E���!  E�D$�K�D�L� L�I��H��0L9�u�H��H�L$XL�D$H�'��L�D$HH�L$X����$�   �����H�D$PH�L$XH��$�   D�d$HM��L�pJ�D@"H�\$`I��L��I��@ L�� 7H H���3����$�   ���1���H��$�   H�C H��$�   H��H�SH��$�   H�SH��$�   H�S��$�   �S(H��H�C H�H���BH�C H�H���BH�H�S �PH��@ ��$�   fA�$H�CH9CH;C~H�CH�CI��H��0M9��:���D�d$HH�L$XH�\$`H�|$E1�1Ҿ   M���  L��$�   �XL��I�F(��$�   ���E���f��$�    �6  1�9D$8�  I��p  L��$�   �   L��L�t$8L��H��$�   ���   ����  L��H��$�   �   L�����   ��tpA�   H�L$8H��$�   �   L�����   ��tK��$�   H�|$PH��HGH�WD�p�@   H� E��tA�L$�H�t�H�JH��H��0H�H�H9�u�I���   M���  �RAVML��H�L$8L�u8H��A��@  ��$�   �������H���H%��H��$�   H��H�D$8�)����$�   �T$@��������   H���$���T$@��$�   f��������������H��$�   �0   L���8����$�    I�G`�p����   H���`$����$�   ���T���I�W`H��$�   H��H�T$@�)��H�T$@��$�    f��%���H��$�   H����(����$�    f�D$@����H���W$��I�`�t$@Ht$8H�D$HH�WL���(�����$�   �������M�W`E1�1Ҿ   L��$�   L��A�
L�T$8��I��L�T$8��$�    I�B(�����H�t$HH���.#����$�   ���r���I�G`H���0��Hc���$����$�   ���N���I�O`H�\$8�L�q(H��H��L�H�D$@�OH���2'��H��I��&��H��fA�F�&��A�vfA�F
��;s�*  ����Hk�HC;0�  I��L9t$@w�H�\$8�  f.�     I���  �x0 �f  H�|$PH�@(H�H���|$@L�l$`I��H�H�\$xE1�H���D�d$HH�D�H�D$XH��    H�D$hA�D$�I��H��   H�D$pf�H�t$XH����#����$�   ���t���H���%��H����A�F�%��M�.H�D$p�T$HI�\ ��t�     H��I���&��I�E�L9�u�|$@ udA�F��  H�D$`I�L��A���t$HI��H���  �I���H��Ld$h��$����$�   D9��K���D�d$HL�l$`H�\$x�����    H����$����A�F�H��H�L$H�!��H�L$H����$�   ���������H���!��L��I���f���L��H���� ����$�   ���\���f��$�    H�D$PH�@H��I���  H�@(H���T��������fD  A�   �K���H��$�   H�D$8����Ǆ$�      H�\$8H����#����$�    �����I�G`�H�P(H��H��H�2L���&v��H��t� f�BH��H9�w�A���     �d����AWAVI��AUATI��U��S��H��xH���   L���  Ƈy   �D$0    H�$M���^  M�}A�79�Fޅ�tFI�H   H=   ��  I�F�S�H���@ H�8H��H��   H��   ��  H9�u�A��$x   uI���    ��  I�} �D$ �0  I�}H���Z  ���i  I�H9�i  D�S�L�G�   I��� L�HI��M�<�L99��  L�ȉ�L��L9�u��D$    E1�M�D$A��  ��  A��D��L�M�E(I��9���  D�F�A�   A)�N��   E1�fD  N�< N9<EE�I��M9�u�E����  H�9 ��  �BH��H���@ H��H�x� ��  ��9�r�A�u ��L��H���� @����  �|$ M�uI�MtA�] I��$�  ��9F(H�D$���0  �u�1���H��H��I��H�PH9�u��9�v&����)�I��H�I�T� H�     H��H9�u�H�D$L�h8M���>  ���N  �]��l$M��L��H��H��L�fD  E�A��vLM�WH�} �   E1�I�RI�B M�JH9�~#��   �     I��H�@H�P�H9���   �΍ND9�u�I��H��I9�u�H�D$�l$H�@H�H1��>�:  �q)�Hc�Hc�H��H��H��?H��2 �  H��Hc�H�I��H��H��09�vzI��H�yH��y���+q�fD  �   H��x[]A\A]A^A_�@ A��I��M�I�BI�1I+2H)�H)�����I�WJ*H�E �>���H�D$H�@H�H���G��� I��$@  AƄ$y  H��t;�D$����   ��u)H�<$�k��I��$�   L��IǄ$@      苭���D$0I��$`  H�<$�fk���D$0IǄ$`      H��x[]A\A]A^A_��    I�<�������    9���  �F�A�   )�L�T�H��D  H�8 EE�H��I9�u������f.�     �D$   �!��� 1������D$0�������M��$�  ����A�   �D$   �R���D  I��$�   L�������D$0����H�<$��L�L$0E1�1Ҿ   �A��I�E�D$0���B���A�7�D$����H�<$��L�L$0E1�1Ҿ   �^A��H��I�E�D$0������A�7�D$   �Y���I��$�   H�L$8�ravgH�x8H�D$H��H�|$L��A��$@  �D$4�������H�|$���H�|$H�T$@��6H H�D$�.'���D$4�������H�|$@   �   �{���I�M�T$Hf;�i����L$JH�|$8H��H��H��H��H9��I����L$ZD�D$X��f��H�H���H��I��H9�����A�uhH�t$`A�H1�I���   H�|$L�L$4E�ExE1�H�t$ �   �,@��I���   �D$4�������A�ExH�t$ Ht$H�t$ �p�D$Z��   H�|$H���J���D$4�������1҉l$,�݉�H�|$���I���   ��HD$ ��H��A;]xv�H�|$��l$,���A�Eh����   �D$4�D$0���@���A�7���������E���*�������1������H��1�1������H��1�1�A�   �D$   �������������H�|$H�����D$4�������1҉l$,�݉�H�|$�F��I���   �ك�H�%�� HD$ H��A;]xv��/����L$HH�|$E1�1�L�L$4�   ���>��I�Ep�D$4���j���H�|$H�t$Ht$P�	���D$4���J����t$HA�uhH�|$H������D$4���'���1�L�t$M��A�܉l$��A;mhs<1�f�|$H t-H�|$�}���T$H�������H�D�I�}p��J��9�wӃ��H�|$D��l$M��L�t$�����d����    AWI��AVAUI��ATUS��H��L���  L���   �D$    M����  I�nI�F�M 9�F�H����  ����  D�C�1�1�M�H�@ H��I�4�H94�t	H�4п   H�rL9�u�J�ȉ�I�UA����  ���   ��H��HUH�R�N��9�v5�Q�)�L��   1�f.�     I�4H94t	H�4�   H��I9�u�@���d  L�L$E1�1Ҿ   L����<��I�ǋD$��uNI���  �0 ��   I�VL�����
����u 1�L��L���
����D$��uI�EH�̀����HD�I�EL��L���`e���D$H��[]A\A]A^A_�D  K�@H��HU9��P���D�A�E��A)�N�D�D  H�rH90tH�0�   H��H��0I9�u�����D  L��� ���I���  �<���@ 1������D$��uAM���  �*���D  1�L�L$E1��   L����;���T$I�F��u�M ����D  E1������     1�1��4������������ff.�     f�AV�   AUATU��SH��H��H���  H����   �K9�rA��tNL�jI�UH��tA��L���   H��H��L�t�H��p  H�T$A�v���   ��tAH��[]A\A]A^�@ 1�1�H�������S��H�c���H	�H�kH��[]A\A]A^ÐH�s0L���c��H�D$I�H��A�u H�C0������t��fD  1�������u�H���  �/���f�     AUI��ATI��US��H��H���  H����   H�} ��   9] ��FM A��y   t`��t H�}�q�1���H��H��I��H�PH9�u�9�v(����)�I��H�I�T�D  H�     H��H9�u�1�H��[]A\A]� ��t��Q�L��I�T��H�     H��H9�u��fD  1��������u�I���  H�} �H��� 1�1��   L����������,����ff.�     f�AUI��ATI��US��H��H���  H����   H�} ��   9] ��FM A��y   t`��t H�}�q�1���H��H��I��H�PH9�u�9�v(����)�I��H�I�T�D  H�     H��H9�u�1�H��[]A\A]� ��t��Q�L��I�T��H�     H��H9�u��fD  1��������u�I���  H�} �H��� 1�1��   L����������,����ff.�     f�U�   ��SH��H��������uH�SH�р΀����HD�H�SH��[]�f�     AWAVI��AUATA��USH��8H���   H���  H��@  L�k8@��t6�EPH�L$(H�ھRAVV��A�D$ E��t6H��8D��[]A\A]A^A_�D  �E@H�L$(H�ھRAVH��A�D$ E��u�H�����H�t$ H��H�$���D�T$ A��E��u��   H���&��A�D$ ��u�A�   fA���{���H�t$ H�����D�T$ I��E���]���H��H�t$ ���D�T$ H��E���?���H�T$ �8   L��E��tw�$��D�T$ I��H�EXE������H�$L��L��J�48�ߤ��A�D$ �������H��uQA���  E��t���EQA���  �����@ ���EAA���  �����@$��D�T$ I��H�EHE��t�����M���   H�4$�D$I�G8H�L��H�D$����ƉD$$��tA���f���H�t$$L������t$$�؅�u�H�t$$L������t$$��A�U ��u�f����D�T$t�   �H�|$�   ��E1�L�L$$1�D�T$��5���t$$I�E0��u�A�M H�|$�   1�L�L$$E1��5���t$$I�E(���W����ٸ   ��D�T$����E1��������$E;E ��   E1�1�H�t$$L��D�T$D�D$D�L$�T$�L$�N���t$$��������T$D�L$���L$D�D$��A��D�T$	�A9�r�����A;E ����I�}(D��#$��Hk�IE;�����I�E0A�����^����    �D$$������A�������@ 1���y   ��   AUATUSH��H��L���  M����   ��I�Մ�t;A�|$P ��   A�|$Q ��   I�t$XH�F0H��uFH�V�   9*vc1��K@ A�|$@ u1�����A�D$DL���  A�|$A tUI�t$HH�F0H��t��V �J�9�H�V(HF���,�H���  ���{���AE 1�H��[]A\A]�f.�     ��    A�D$D�ܐA�D$T��f�     �   ����A�D$TL���  �&���D  �   �����fD  1������f�     ���  �#  AWAVI��AUATUSH��L���  M�D$`A�(I�X(H��H�H9�sOL���  �f�     M�D$`H�3L���pb���K
�SL��I��I�p����M��tfCfA�H��H9�w�fA��h  �tIH�  ����  I���  ��   A���  A���  fA���   fA��  )�fA���   fA���   A��  A��   �0�@ ��fA���   f���1�f��)�fA���   H��I���   []A\A]A^A_�Q^�����    A���  A���  ��fA���   ���fA���   fA���   �v���D  AWAVI��AUM��ATA��USH��H���   H���   ��1H �T$H�x����H���  1�L��I���$���Ņ���   M��D��T$H��L��A�W�Ņ�upH��  �dbk�H9���H=eurt��!ʹtsl�H9�����tH-   H�������  H���   �T$H�K   H�D$��xM��D��H��H��A�W�Ņ�tH���   ��[]A\A]A^A_�@ L�c(M��tOA�@<H A�>H �
�I��M9�t7L��L���u� H��t�H�D$PL��@  H�D$ �  ��   �f�     H�|$P1��   f��    H��H�|$ L��@  �H��  1�H�Fh�D$: �D$; �D$9 f�|$H�$�l$<D�d$H��(  I��J� H��mgpf�x  H��perp��   H�� tvc�F  f�D$�D$f;�   r��l$<�T$PH�L$ �h7H �H<H �|$9D�D$;D�L$:��     H��0H��H9���   �@��uH�8 u���E��uH�x u���E��uH�x  u�����u��q@ �D$:��  A�   I��L�|$ 1�M��� I��I��0L9<$�8���H��(  I��h7H L�H9Pu�H���f  A�I9�`7H u��A���u��l$<H�K    L�|$H�L$ �xmdhH��M�g8L��A�҉D$L��uH�t$PH���8  H�C���   H���   H�xh ��  H�t$H��譙���Ņ�t<������H�L$ H�T$�mgpfH����@  ���e  Hǃ       Hǃ      H�L$ H�T$�perpH����@  ����  Hǃ0      1�Hǃ(      H���   H�xh ��  H�C�t$����t����  HǃH  `�@ HǃX  ��@ Hǃ`  P�@ Hǃh   A HǃP  ��@ ���� M�������1�H���   H�0H��A�҅���   H��(  N�l H���   L��H��L�l$(H�D$��������   I���+  H�\$0L��L�l$1�@ L��H���,���H��w�H�d$(H�\$0H�D$(H��tCA�   �   H�\$(A)�D��A���H�|$�:
����    ������A�9�u�H�\$(D��H�|$��	��L��@  ����fD  ��  E1��D$9�N���fD  �ć  A�   �D$;�3��� L���  L��L���>	���D$L���  L���  A�GE�w��AΉ�A�G	�A��A������DG�f=� ��   D��E��f���T  I�V�H����  ��   H�L$P1�E1�L�L$L�   L��D�T$H�$���,���T$LD�T$H���  ����   H�<$O�D7L�L9��  E�J�1�1��!f.�     L�H��I�H9�rH���  A�t@�4�rI9�u�H�D$P���  L���  H���  �D$L����������[��� �   �N���fD  �D$L   H�|$L�����Hǃ�      �fD  H��h  H�T$�fylgH����@  ��<���  �������H���   H�xh ��  Hǃp      H�L$ H�T$�acolH����@  ��   �������f���   H�D$P�a  H=�� �  H��H���  �   H�S H�rH9�t	H9��  H�t$PH�|$H���  ���H��h   ��t<��C�����������6���fD  1�� ���H��������Ņ�����H����������H�t$PH�|$H��   H��  ����Ņ������<�������}���L�L$LE1�1�1Ҿ   L����)��H���  �D$L���j���1�����H�t$PH�|$H��0  H��(  �F���Ņ��[���<��t����N���Hǃh      Hǃp      �}���1��D$: �D$; �D$9 �T���H=�� ��   H��H���  �   �����s8������H���   �����H���   �����E1�E1�E1�fD  H�T$LD��H����g���L$L��tA�������M��A�   I��L;��  r�A�������M����   H�CH���H�C����H�D$P�� ���  �����H�D$P�� ���  �7���D��   H��(  H��H�|$I��I��I����L9�sk1������   �    H�UH)�H��~
H9�HL�L�H�� I9�w�@��t4I9�wAH�C L�l$PH��H���  �y���H�|$���H��p  �����H�L$H�IH�$H)��H���  1�H��tH�B�H�C �6���H�T$ �   D��H���������w����|$P.�l���H�|$ ��1H �Z� ��������P���ff.�     @ ATI���@AH UH��S�<���H��H��tH��[]A\�@ M��t�I�|$H��t徙1H ����H��t�H� H�@(H��t�[H��L��]H�@ A\��ff.�      U��H���   S�l1H H����À� �ۅ�t�   H����[]�fD  H�ׄ�u1���#t��(t�   H����[]��    �ExH����[]�@ �
   1��I� ��f�UH��SH��H��H�<$H��H�t$�#���H�4$H�T$H��H�FHI�H��H��f�E H�BHI�H��f�H��[]�ff.�      f9��   v_f9��   vVD����I��L��   H��H��   M�M�@L+H�@L��L��H)�H	�t5���  tIL)�H��L��H	�uC1�� ���   �   t&�G�   �f�� @  H��H��H�I����1�H����H��L����L����fD  AW1�I��AVAUATUSH���   L�I���   �zx(�  M���  1�A��  A��+  fA��,  �   A��T  H��L�H�H��HC�H9�vH��   ���  HC�fA��T  IǇ0      IǇ@      f���  ���2   �2   Ƀ�2L�Hc�I���  �  H�I��8  I�P H��H��H��H9�s
I��8  H��I��H  A���  IǇ�      fA9��  ��  IǇ   �@ IǇ  ��@ IǇ  ��@ IǇ   ��@ L���[��A��@  <w���$��1H @ IǇ�  �A D  I���  I���  E1�A�   I���  �Lc���A���  A�� >H A���  ���  H�H�H9��T  A�� ?H I� ����H)�I�8�~  I�(����)  Hc�I�W8�� ?H ��H�I�G@H9��.  M�G0AƇ�  A�G    I�,Ѐ���$  D��B�$� 2H H�E H��~	H9���(  A���   �3%  H�E      I�G@A���  I�G ���|   I��I��@B �8$  I���  I���  H9��^  A��`   �����1��    L�JI9��J  D�LD�ȸ   D)�A���  �����H�U I��H  f�I�G Ic��  I��  �q���f�     I�H���  H���5  �IG8I�G@H9��j   A�G�   ��   H���   []A\A]A^A_� A���   �_$  ��t1I�01�H��    A���  H��Hc����� ?H ����f9�w�I�G8    �2����     J��,  I��8  � ���@ H���������L��H��H��������    IǇ  �@ IǇ   �@ IǇ  0�@ IǇ   @�@ �����    ��)  �������1�A�@ �������d  ������������    I�G@������    IǇ�   A ������     IǇ�  �A �����IǇ�  �A �����IǇ�   A ����IǇ�  @A ����IǇ�  �@ ����IǇ�  �A ����L���H���A�G@ ���h���=�   �@���A���  I���  H��H��H9�r� ���D  H��(H9������z t��rA8��  u�Ic��  A;��  ��   A��x  I���  H��I��  �H�N�2H�HH�@   H�P�F�����   H�RL���+���<�����A�G����f.�     H��L���U\��A�G�����} ��"  A���   �t���A�G�   ��   �E���A���  1����4���A�G�   ��   �"����    A�G�   ��   �	���H�} �����H��L��谛��A�G����H�EH9E ����H�E I�G@A���  �����H�U A�OTL�Ef9���  fD9���  H�}A���   H�uf9���  f9���  H�M fA9��   ��  I�G`��E��H�L$hI��H������H�T$ H��H�L�H�L�JH��H�|$XL�`L�D$`H��H�\$(H�I���   L�L$HH)�H�:H�H�\$H��H�8H�rH�@L��@   H�t$0H)�L��L)�L�T$PL)�H�|$H�t$8H�D$脧��H�t$H�|$�@   H���m���H�t$H�|$�@   H��V���L�L$HH�|$�@   H�D$@L��L)��7���H��H�L$hL�T$PH��?H��L�\$XL�D$`H����H1�I��H)�I��H��H�4PH�D$@H�H�H1�H)�H9��'  I���   I�W`M��   H�I�J�4HT$ I�HHHH�xHH�H��I�I�CHCHFHBH�PHH�H��I�AI��   �	A�G�f���fD  A��"  A��&  L���T��A�G�A���I��(  I��&  H�EH�U I�G@A���  ����I��$  I��"  H�EH�U I�G@A���  �k���HcU Ic��  H��H��H��?H��
 �  H��Hc�I��X  ����H�U I��P  ����I�G H�E I�G@A���  ����H�E H�UH�EH�U I�G@A���  �����I�G@    1��e���H�E H�EI�G@A���  �����������f% @f�� @��w fA��"  fA��$  fA��  fA��   �������fA��&  fA��(  ����H�E H�u��f	������I��(  I��&  H��H�������t���H�E H�u��f	�tI��$  I��"  H��H������A��"  A��  �7����U �uI��&  L���������� ��������U �uI��"  L�������������A��"  L��A��  � R��A�G�'���H�E A��8  H9���  I��@  H��H�E I�G@A���  �n���H�U A��8  H9��m  H�MI��@  H��I�G@A���  �9���L���e���A�G����H�m fA;oT�-  1ɀ�.t9��L��H��IG`H�PH�0A���  I���  L��H��H��A���  H)�H����I�wHL��A���  fA��  A�GfA��  �3���A���  ����  �Q�A���  Hc�H��I��  H�rH��H�rAƇ�   H����  H�RA���  H�RI���  I�G �X���A��x  ����  A���  M���  H�U H��H��I��I9�r�  f�     I��(L9���  A�AH9�u�H����  ��  I���  �   A�9fA�IH��A�QI�AA���  I�A     H9�vA���  L����Q���������A���  <-��  <�t<,u�A�G�   ��   �K���A���  H�M ��H��H9������A���  I���  9���  ��H��H�4�H9�r��  @ H��(H9���  �PH9�u�x �����A���  A;��  �����A��x  Hcу�H��I��  �2I���  H�B   H��H�BH�r�0A���  �V����!  H�PL������A�GAƇ�   ����H�U fA9WT��  fA��&  Ƀ��fA��(   t�����IGp A�G�����AǇ@     IǇ�  �A ����I��0  I9G ��  A�wTfA9�  ��  I���   H��;��  f�     A���   �n���I��0  H��I��0  H���r  M�G0H��I�W8I�,�fA;��   s�A��  ��L��H��I��   H��IG`H�QH�1H+PH+0A���  ��H��L��H��H��A���  I�W8�v���H�] fA;��   �f  A��  fA;WT�S  ��D��I���   D��H��I��H�t$fA��n   ��  I���   L�IG`H�QL��H�1H+PH+0A���  H�UL��I���   H��D��H)�A���  A��  fA��  fA��  A���  �����fA��  A�G����L����\��A�G�	���fA��l   A�   tfA��n   tE1�fA��p   A��I��0  I;O ��  L�M A��&  D���8I��A��(  D��Lc��%I��Lc�H��:��  �     A���   �~���I��0  H��I��0  H����  M�G0H��I�W8I��fA;��   s�I�H���   �yx(��  A��+   ��  E��u=A��,   t
A��-   u�A���   tfA��(   uI���   ����g���1���A�   L��L���s���I�W8�H���fA��p   H�] �   tA���   f9������L�D$~H��$�   L��H��$�   H��$�   �`Y�����.���1�f��tI���   H�Ӹ   fA+�   fDQ�fA��p   ��  E���   D��fA9�w:�����fD  H��$�   A�   D��L��H��$�   觐��A��fE9������I���   H9�$�   u�fD9L$~u���H�U I��8  �����AǇ@      IǇ�  �A ����AǇ@     IǇ�  �A ����H�U H�������I��0  ����H�U ����  ����  �Ao�  �Ao�  �Ao�(  �Ao�8  AgHAoXAwhAx�Ao_H�AoWXfA��l  �AoOh�AoGxfA��n  A��   A��   A��   A��   A��   A��   A��   A��   fA��p  ����H�U ���x  ���8  �Ao�  �Ao�  �Ao�(  �Ao�8  A��   A��   A��   A��   �H�U ���f  ����  �Ao�  �Ao�  �Ao�(  �Ao�8  A��   A��   A��   A��   fA��n  �����H�U ���I  ���w  �Ao�  �Ao�  �Ao�(  �Ao�8  AgHAoXAwhAxfA��l  ����A���  H�u�SH��H9������A���  I���  9��  ��H��H�<�H9�r�  fD  H��(H9���  �JH9�u�z �5���A���  A;��  �k���H�}  ����A��x  Hc���H��I��  �0I���  H��H�pHcu H�PH�p�2A���  �F����  H�RL��褉��AƇ�   H�E I�0  I��0  I;�8  �S���A�G�   ��   ����� A�   �<Y����A)��%���L���I��<����A���  <Xu�A����I���  ��A+ D�DL��A9��s���A��f����  �   �f�     I���  H��LH�L��H��f9�s���IG@A���  I�G@�W���L�e D��fE;gT�{  H�uI;��  �j  I��H  L��H�D$A��  H��A��H��fA��l   H���L  IG`H�PH�0L��A���  H��A���  t.H��L��H)�H�H1�H)�H9D$I���  HL�H��A���  H��H)�A��I�wHL��H��A���  A�GfE��  fE��  ����I��0  I9G ��  L�D$~H��$�   L��H��$�   H��$�   �S�����|���I��0   I�W81��   A���   �����I��0  H��I��0  H����  I�G0H��I�W8H��fA;��   s�H��$�   ��A�   L��H��$�   ����I�W8�I���  ��A+ D�DL��A9��l���H��A��I���  f��tG�G���H�|� �D  I���  H��H�BI���  ��T���H��H�E H9�u�I�G@H�AƇ�   I�G@�����H�EH9E ����H�E I�G@A���  ����H�EH9E ����H�E I�G@A���  �����H�U fA��  �`���H�U fA��  �O���H�U fA��  �>���H�EH9E ����H�E I�G@A���  ����H�EH9E ����H�E I�G@A���  �t���A�G�   ��   �9���AƇD   �����AƇD  �����I�H���   �xx#�b  I���  H�E I�G@A���  ����L��A��  H�E A�G�����A�H�u L��H�I����  A���  H�E A�G�]���H�E H��?H���H�E I�G@A���  ����H�e �I�G@A���  ����H�UH�M H�EH�MH�Uf�H�E I�G@A���  �w���AǇ@     IǇ�   A �����AǇ@     IǇ�  @A �����H�uH�V�H���C	  H�} �N��   ��H��tHc�H9��$	  ��A"�d  	�A��d  H���x���I�H���   �zx(�d���H��A��+  �S��� AǇ@     IǇ�  �@ �5���H�} �*����z���H�U �A-  L����?��A�GAǇ@     IǇ�   A �����H�] I�G@A���  �\���H�U H�������H��H�U I�G@A���  �7���H�uH�} �@   蹓��H�E A�G����H�UH����  A�G�   ��   �����H�EH)E I�G@A���  �����H�EHE I�G@A���  �����H�U H���u���fA��b  �0���H�U fA��`  ����H�UH;U ����H�U I�G@A���  �x���H�}  �C���H�}  �   �����H�} ���������H�E H���������I�H���   �����H�E    I�G@A���  ����H�}  �����A�   �     L���B��<�&���A���  <X�G
  <Y�3
  <u�A������t������1�H�u L��A���  �����H�E A�G����1�H�u L��A���  ��H��@����H�E A�G�����H�EH9E ����A��x  ���  A���  M���  H��H��I��I9�s$H�U A�AH9�u�5 A�AH9�t)I��(L9�w�L9�uA;��  ��  ��A���  H�U H���   ��  I���  A�QA�AA���  H��A�9I�AH�E H9�v
��A���  L����@���������A���  <-��	  <�����<,u������H�E A���   H9��E���H����F�r  I��   L��H�PH�0A���  H��A�GH�U ����H�u I;��  �	  L��A��  H�E A�G����I�H���   �zx(�:  H�uH�} E��  ���fA9���  fA9���  f9��L�����I�0  �f9�s������I�H���   �xx(�Q  I��0  I9G �M
  H��5�`   A���   �����I��0  H��I��0  H����  M�G0H��I�W8I��fA9�  v���I�0  �0I�W8�H�UH;U ���������L�e fE;��   �  H�mfA;oT�  ��A��L��H��H��IO`I��   H�QH�1H+PH+0A���  I���   L��H��H��?H�H��A��H��H��H��A���  H����L��I�wHA���  A�G�����H�U I;��  �{  Ic��  HcEH��I���  H��H��?H��0 �  H��H�H��I�G@A���  �'���H�U � @  L���j:��A�GAǇ@     IǇ�  �A �{���L���   A��  H�m I�W8I��H��u*�  �    A���   �>���H��H��H9��x  H���w  I�G0H�J�I�O8H�t��I;��  s�H�<�A���  H��H������t��  L�@ ��uID�A��`  H�H��I9�u���D��H�G�H��H��L��HI�A*�b  H��A��   I�W8�`����A�H�I����  H�E H����  Hк    HH��d���H�U fA9��   ��  H�MfA9��   ��  ��I���   ��H��H��H�I��I���   H��H�H�H�NH�zH+H��H��H)�H	���
  ����  H)�H��H	��  M��   I��   I�L$H�}I�$H+E H��H��H)�H	��u
  ����  H)�H��H	���  L���o:��A�G����H�E fA9GT�����H�UfA9��   ���������H��H����I�O  I���   IG`L��H�0H�H�PH+1H+QA���  H��A�G�j���H�] fA;��   ��   I���   D��L��I��L�H�PH�0A���  H�M��L��I���   H)�A���  fA��p   �����I���   I���   �Bo"B �e���H�u I;��  s2H�UL��A��  A�G����H�M H9�|H����	  f�     A���   �b���A�G�   ��   ����I�O8I�G0AƇ�  A�G    H��H��������wA+w 9��`������;  �p�H�z1��H��H��H��H��H�PH9�u��Z���I�7H�U H���   ���Hx�    HE���tA��   t����tA��   t����tH���   t���� tA��(   t����(�l���A��)   �^���H���� ��@HE���tA��*   t�̀H��H��   ��HE�H��H��   ��HE�������A��.   ����H   ����� H�U H�����������  A��h  �����I�H���   �zx(��  H�uH�} E��  ���fA9��G���fA9��=���f9��������I�0  � �f9�s��@���H�U �ʁ��   ��  ����   ��tA���  9�|AƇe  H�U ��tA��   tAƇe  H�U ��tA��   tAƇe  H�U ��tA���  9�}AƇe   H�U ��tA��   tAƇe   H�U �� �����A��   �����AƇe   ���������M  �����  ����"  ���������ˍGA+G f�� ��9�������   H�I��  �H�T��H��f9�s������@ L����A�   L��L����{��I�W8����H���K�����   �x���A���������A������A���   tcA�G�   ��   IǇ0     I�W@�8���IǇ0     A�GI�W@�����A��+   �����A��,   �����A��-   �����IǇ0     I�W@�����A���   �}���H�E     I�G@A���  �����A�G�   ��   H�E     ����A���   ��  fE��  fE��  ����A�G�   ��   �l���I���  I�AA�G����H)к    H��HO������L9��n���A;��  �
  ��A���  �R���A�G�   ��   ����A�G�����A���   ��  A�GI�G8    1�����L�D$~H��$�   L��H��$�   H��$�   �KB��������A��p  f����  E���   fE�������E1��/ H��$�   E1�D��L��H��$�   �y��A��fE9������I���   H9�$�   u�fD9L$~u���A��+   ����A��,   � ���A��-   ����������f�A���   ����A�G�   ��   IǇ0     I�W@�����H�} �@   ����H�E A�G�v����Ao�H  �Ao�X  �Ao�h  �Ao�x  AGHAOXAWhA_x�����Ao�H  �Ao�X  �Ao�h  �Ao�x  A��   A��   A��   A��   �&����Ao�H  �Ao�X  �Ao�h  �Ao�x  A��   A��   A��   A��   �����Ao�H  �Ao�X  �Ao�h  �Ao�x  AgHAoXAwhAx����H��L���4��A�G�V���L��A��  H�E �����A��+   �����A��,   �����A��-   ���������@ H)�I��H�E I�G@A���  �p����2�F�������H�RL���s��A�G�����A�G�   ��   ����H9���������H9��e�������A�G�   ��   �����fA��  fA��  ��   A�G�   �����I��   L��H�PH�0A���  H��A�G����A�G�   ��   ����A��&  ���-��I�OXA��(  ��H�H�H��-��H�H�AI�G`�oH��u���H�u L���:w������H��H�ЋzH9��	���H���.���I�OXL�L$L��I���   I���   �oB
D��H�MA��   I���   L�L$I���   �BoA��  L�	H�������H��H��D�AL9������H������� @  I��$  I��"  �"�������1ۿ @  I��   I��  ��������A�G�   ��   I�G8    I�G@    �?���AƇe  �����H��H������H)�H��I�< I�t H��� I�G0I�W8H�\��A�G����I���   H��A�   fE+�   fDZ�F�����I����GA+G ��9������I���  f�� H�P��H�L� �I���  H��H�BI���  ��T���H��H�E H9�u�AƇ�   I�G@�6���fA��l   M���  ��   fA��n   ��   M���  I���  IGhI��   L�H�0H�HH�RI9���  ����Mc�Hc�D)�)�H�Hc�I��H��L��H��H��H��?H��?H��0 �  H��
 �  H��H��Hc�Hc�A��H��A�G����f������I���   f�������I���   D�TB�A�������L�I�G@I�G �#���A�G�   ��   AƇ�   �X���I���   IGXL��H�0H�H�PH+1H+QA��H��A�G����I�G@�   �E���A�G�   �����H�|$(H�t$8�@   L�L$HH�L$@L)����H�t$L��@   H+|$0H�D$ ���L�d$ H�t$H��I�L���w��H�t$H��L��H�D$�b��L�L$HL�D$I��   M��   LHCM�H�L$@I�A����H)�L)�L��H��A��Ic��  H�H��H�H�� �  A�GH��Hc��*���H������H��H������H������H��H������fD  USH��H����   H�oH�T$�P  H��������L$H�Å���   H�h1�L�L$E1��    �    H��ǀ�      ������T$H���  ��uKǃ       H��H�C(    ǃ�      H�C0    Hǃ�      H�    H�C    H��[]� H����?���D$��t
�     1�H��H��[]�@ AWLcٹ/   I��AVAUE��ATUH��SH��H��XL�bD�D$I��$�   M��$�   H�D$1��H�A��uEE��txL�[ 1�L�#H�kL�SL�s0Hǃh      Hǃp      H��X[]A\A]A^A_�fD  E��u�I��(  D�\$L�T$L�(L���?���L�kLc\$L�T$��    D�؃���D$��  ���0  ��  ���  ��u��Ѕ�u�L��  M���8
  D��H�t$�����~x(��	  AƇ*   ��D�l$(�D$H��L��L��D�\$8L�T$ ��C�����&���H�t$A��(  L�T$ D�\$8�~x(��	  8D$��   �D$A��(  H���   tPM��$@  H���  1�1��    I�PHc��   H��H��H��?H�� �  H��H�׍VH��H;��  r��t$H��D�\$L�T$�F��L�T$D�\$���l���A��d  �tA��D�ރ�@�t$���   1ҹ   H�       @IǇ0     I��  H   @I��   1�fA��(  H�      IǇ8  @   AǇ@     AƇD  IǇH  D   IǇP      IǇX      AǇ`  	  fA��d  I��h  fA��p  �D$A���  I���  L��  H��  ���� ���s�����   L�>H��   D�\$8H�T$ I���   H��H�D$����H��  H�|$Hǅ       ����H���  H�|$Hǅ      ����H�|$Hǅ�      H���  ���L�T$ D�\$8Hǅ�      H��  H��tD�\$8L�T$ ��;��D�\$8L�T$ H���  D�\$8H��L�T$ H�D$(�\<��I���   Hǅ  �����%���1�H�|$E1�H��  L�L$H�(   A���  H�����   A���  ǅ�       ��  I��8  ǅ      H���  A���  Hǅ      f���   1�f���  Hǅ�       Hǅ�       Hǅ�       Hǅ�       �����L$HL�T$ H��   D�\$8����  ��  H�|$E1�1�L�L$H�(   �i���L�T$ D�\$8H��  �D$H����  H�|$E1�1�L�L$HH���  �   �,���L�T$ D�\$8H���  �D$H���O  H�|$E1�1�L�L$H���  �   �����L�T$ D�\$8H���  �D$H���  H�|$f��E1�1�A���  L�L$LHǅ      H���  �p��  ��f�t$8�   ��  H����  D�\$<L�T$0H�D$ �i���L�T$0D�\$<H���  �D$L��uEH�L$ H�|$E1�1�L�L$L�   D�\$<L�T$0�(���L�T$0D�\$<H���  �D$L����  H�|$(D�\$ L�T$��9���D$LL�T$D�\$ ���D$H�  �D$8D�\$(E1ۺpyA ƅ|  H��  f���  H�       @H��P  H��H   @H��X  H�      H���  �   fD���  f���  I���   L�T$ E1�H�@H�L$fD��`  H��8  Hǅh     Hǅp  @   ǅx     H��Hǅ�  D   HD�H��Hǅ�      Hǅ�      ǅ�  	  I��H  L�} L����=��������H�L$�D$L�T$ D�\$(Ɓ`   ���  I��  I��   ǁ�      H��H�A     HǁH  @   HǁP      HǁX      Hǁ�   @  ǁ�      Hǁ�      Hǁ�      fǁ�    Hǁ�      Hǁ�     H��  H��  Hǁ      Hǁ       Hǁ(      Hǁ0      �  ǅ      ���  �o�  �o�  �o�(  ���   ���  ��  ���  ��  ���  �   ��  �0  �@   ��  ������f�H���   �t$H�E tKL��@  H���  1�1� I�PLc��   I��I��I��?J�� �  H��H�׍QH��H;��  r����  ��tJ�x�H���  H���  1�H��H��@ H�    H�D    H�    H�D    H��H9�u����  ��t-H���  �H�H�BH���
fD  H��H�    H��H9�u�1�E1�A�   D�\$ H�       @L�T$H��P  H   @H��X  H�      f��`  H��Hǅh     Hǅp  @   ǅx     ƅ|  Hǅ�  D   Hǅ�      Hǅ�      ǅ�  	  fD���  H���  fD���  �>��L�T$D�\$ �e����H��D�\$ L�T$�.6���D$HL�T$D�\$ ���������� ����   A��   D���D$(����A��*  �   D�l$�D$�=����     A��.  �t$A8�)  t4A��)  8T$(tJ�t$(A��.  8D$�G����N���f���   �1���8T$(u��!��� AƇ*   D��D�l$(�}���8D$�	�������D�\$8H��L�T$ H���  H���  Hǁ�      ǁx     H�L$A��H  H�L$L�T$ ����  D�\$8���������H�L$ H�|$E1�1�L�L$L�   �X����|$L L�T$0H���  D�\$<�1���H�L$ H�|$E1�1�L�L$L�   �����|$L L�T$0H���  D�\$<�����H�|$E1�1�1�L�L$L�   D�\$0L�T$ ������|$L L�T$ H��   D�\$0������D$8�D$H    fǅ�    f���  �����ff.�     @ AW�����A��AVI��AUA��ATUH��SH��  H���   H9��  ���  H�}H�G  ��  �G���  H��H��p  L���   L���   L��$�   AT���   AXAY�Å���  ��$�   ǅ�       ǅ�   stibH��H�E0��$�   H��H�E8H��$�   H��H��H�E@H��$�   H��H��H�EH��$�   H��H�EPH��$�   H��H��H�EXH��$�   H��H��H�E`��$�   H��H�EhA����  ���   ���   H�E�@��   A�   D��H��L��L�������1ҹ   D��L���u��H��$�   1�1�I��$h  H���   �a��Hc�$�   H�}P Hc�$�  H�UpH�Exu+H��t&I�NXHcIH��H��H��?H��
 �  H��Hc�H�UPH�}h u%H��t I�VXHcRH��H�H�� �  H��H�H�EhH��  ��[]A\A]A^A_��    L�MI�A������J  H��t��    D�����D$��  �   A�� @  u�E1�D��H��L��L��$�   L�������Å�u�1�1�D��L��ǅ�   ltuoǅ�       ǅ�       ��s���Å��  ���   pmocH��$�   ��  �o@�oH(H��$�   H�@8��   H���   ��   ���   ����H���[  A��uEH��$�  ��e   �@  ��h  ��t%��  ����  ���  ���   fD  L��$�   L��$�   H�D$   H��$�   I���   ��$�   uH�qXH�VH�T$A���   pmoc��  I���   H�t$@H�L$(H�D$ L�D$許��L�D$H�D$ H�L$(Hc�$�   H�|$@L�L$XI�ppH��$   H+�$�   �xx(I�x@M�HHI�pP�m  H��$�   %   I�  uWH�AXD�A���  ��tDM���  A�fA9��  ��H�P�   ��A�H�pfA9���  H��H9�u�D  H�D$PH)�L��H+|$HI�@0I�x8A���   tfA��   �O  H�t$L�D$�@m��L�D$fA��h  �H����  A���  A���  )�Hc�H��H)�I��I��?I�I��I���   H�PhH��tNH�H�@H��tBL�D$H�zD��   H�L$pH�L$`H�D$`    L�L$h��L�D$���$  L�L$hH�L$pI�Hx��$�   u?Lc|$Mc�Hc�M��L��L��H��?M�� �  L��H��?I��I�� �  Mc�H��Hc�I�PPM�H`I�HhH��H��?H�I�P@H��H)�I�PXH��$�   I��$h  1�1�H���   ����D$���
���I�FXf�x��������      ������    A���    �$   ����������     fo�$�   fo�$�   )T$@)\$P�v����    ���   �����@ ���P����H��$�  H���������+   ������p���D  �PPH�@X���   H���   �L����    A���  A���  )�Hc�����fD  ���x������    �\���@ H��$�  H�t$L�D$L)���j��H��$�  1�L�D$L��H��$�  H9������H�t$H)�L�L$ �j��L�D$L�L$ ������fD  H��H���   1���������H�������1�1�1�1�I���   f�T$>f�L$@f�t$`f��$�   �Q���I��p  L��D��1�L�D$`H�L$>L�L$1����   L�L$M��1�H�L$@D��L���V��H�D$>H�E0    H�E8    H�E@�D$`H�EH    H�EPH�D$@H�EX    H�E`��$�   ǅ�   stibH�Ehƅ�   Hǅ�       ǅ�       ����1�fD  I���  A�uH9������H��H�DI��  ������ ��I�@P������    ���   ���   �w����    ���   0����ff.�     �H��H�wH����   H����   ;V rL���   I�xh ��   ��t[H�vA��A�����    AE�A��A��  �ŀuWE��tA�ȃ�A��	H��AE���t$H�pH�pXH��H������f�     ��  u(H�p`H�pXH��H���e���D  ��E��u��fD  H�v��    �@ �$   �f.�     �#   �f.�     �   �f.�     ��G�H��H	��FH��H	�H9��H9Ѻ   G���    H��  ��     �o��   �o�  N�o�  V H��(  H�F01��ff.�     @ ��0  f�1�� �   �f.�     �o�8  1��o�H  N�o�X  V �o�h  ^0�o�x  f@�o��  nP�o��  v`�o��  ~p�o��  ��   �o��  ��   �o��  ��   �o��  ��   �o��  ��   �o�  ��   �@ H��P  H��t\D�I�1҉F1�D�E��tA�    H�|�H��H�|H���   L�L�DD���   J�|��H�|H��A9�w�1�� �   �f�H��S1�H��1�1�H���Ph��`  [�D  ���  ��     AWAVI��AUI��ATA��USH��H��H�o�W8H�H9�vW� ��0��	wLH���SHH��I���S@H�H�PI�M��x.H)�L9�~&�SI�GH1�M�} ����H��[]A\A]A^A_�f�1�E��u��C   H��[]A\A]A^A_� H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ USH��H�GH��p  H��t.H���   H���`BH H�x����H��tH���UH��(  H�B@H��1�[]� AWI��AVAUA��ATUSH��H���	  H�oH�L$L��  �o��  �o��  �o��  I�FH�$H���   L�`h��
  ��
  ��
  M���m  I�$I�|$����"  ���    �-  �   H��H��$�  A�V0H��8  H�T$H��A�V8H�D$IcWI�7H��$ 	  H�$H��$�  �P<�u/H�CH��$�  ƀ0   H�D$� H�$IcWI�7�PfD  ����   M����   I�$H�z t|H�{@�;b��H�{PH�D$    H��H�D$� b��H�{XH��H�D$ �b��1�I�|$D��H��H�L$H�D$(I�$�PH�T$H��H�S@H�T$ H��H�SPH�T$(H��H�SXH���	  []A\A]A^A_�fD  H�$A�WH��I�7�P�:���f.�     H���  ��H��I�H���  ��A�G���    ������ SH��H��0H�L$H�T$ �D$ �������u+H�SH���   H�RhH��tH�zH��D$H�t$ �R�D$H��0[�ff.�     @ AV1�1�AUATI��UH��SH���  L��  H�    H��L��P  L���  I�Fh��A j j H�|$ �H�� A�Ņ���   ��`  Ƅ$�   1�Ƅ$�    ��$�
  H��h  H��$�
  H��p  H��$�
  H��x  H��$�
  H��h  H��$�  ��`  I�$    ��$�  ���  ��~+ ��H������H�D$P��tI;$~I�$��9��  �I�FH���PH���  D��[]A\A]A^� AUATA��USL��H���  ���  H��  H��I����L��P  H��1�1�H�@L���  h��A j j H�|$ �H�� ����   A��`  Ƅ$�   Ƅ$�    ��$�
  I��h  H��$�
  I��p  H��$�
  I��x  H��$�
  I��h  H��$�  A��`  ��$�  E��tIA��D  ��H�    H��A9�t,��H��������u�H�|$P��H����^��H��H�C�A9�u�1�H���  []A\A]�f�     ��t�B�I�D�@ H�    H��H9�u�1���ff.�     �AWAVAUA��ATA��UH��SH��H��P  L���   �D$    H����  E���y  ���t#D9��j  H���   []A\A]A^A_�fD  E��L�L$E1�1�L��8   L������H��   �D$���_  L�L$E1�L��1Ҿ�   L���n���H���  �D$���2  L�L$E1�L��1Ҿ    L���A���H��8  �D$���  1�C�$L�L$E1��   L������H��H��  �D$����   J��H��  H���   H��  H��8  H���  H���  H��0  A��vTA�T$�H��   H���(  fD  H�8H��H�W8H���   H�H���   H��  H���   H�W H��  H9�u�D�# �k������E��tA9�t���z���D�kD��   D�#E��t��tH�{( tU�D$H��[]A\A]A^A_�f.�     H�T$�   L������H�ËD$��u�ǃ�      H��P  �����D  D��   L�L$E1���1�L������H��H�C(�D$��u�A���y���A�L$�H�S0L�D�8���H�s(��H���H�4�H�r�I9�u��I���f�AW�   AVAUATUH��SH��H��  L��P  H��H�t$ H�L$�Sx�t$��   ��x t6��1M��t4A���t-�   9���   �CH�Ĩ  []A\A]A^A_� �   ��1�H���������u�H�CL��P  L�3H�D$�D$��~GL�d$ 1�I�$1�H��I��H�I�D$�H�CI��  L�,��SPI��  I�E H��H��9l$�H�D$L�3H�C1��]���D  H�CL�3H�D$�f.�     AWI���   AVAUATUSH��H��(  H�|$H�L$8L��H��$�   A�Wx�T$8��   ���2  �R  ���I  I��D$    �D$    H��P  H�D$ I�GH�D$(H��$�   H�D$fD  H�L$�   H�t$@L��H�I�H�AH�L$<I�GA�Wx�D$����   �T$<�B��T$����   H�\$�t$8H���F�������   H��P  �D$<LcT$H�l$@E1�M�r��~:fD  H�E 1�L��H��I�H�E�I�GJ�D�N�$�I��A�WPI�$D9l$<̃D$�D$H�D$9D$8�+���H�D$ I�H�D$(I�G1�A�GH��(  []A\A]A^A_�f��D$9D$<�_����   ��ff.�     AWI���   AVAUATUSH��H��  H���   L��H�L$8�D$4    H�t$@H�D$A�Wx�T$8��   ����  ��  ����  I�1�H��H�D$ I�GH�D$(�������D$4���[  �D$8H��P  ���7  H�D$@�D$    H�Ũ   H�D$f.�     H�|$H�L$<�   H��$�   H�I�H�GL��I�GA�Wx�L$<�A����  H�} ��   �H�|$L�L$4E1�Hc�1Ҿ   �{����L$4H�E����   HcL$<H��H��H�M�U ��~gL��$�   E1���    H�EI�u I�ML��I��N�$�    I��H�VJ� I�H�Q�I�WA�WH1�L��H�H�]A�WPL�H�D9t$<��D$H���D$H�D$9D$8������L$4H�D$ I�H�D$(I�GA�OH�Ĉ  []A\A]A^A_�D  �   ��f�     UH��SH��H��H�vH�[���H�CH    H�s8H���CP    �@���H�C8    H��H���C@    H��[]� ���AWAVAUATUSH��H��P  H���o  L���   D�3I��H�s(�kL�������H�C(    A���T  A�V�H�C0H�T�8�    H�     H��H9�u�H���  L������H��   L��Hǃ�      ����H��8  L��Hǃ       �m���1�Hǃ8      HǄà      HǄ�      HǄ�0      H��A9�w�H��  L���$���Hǃ      Hǃ      ��t]D�}�L�sJ�l�I�6L��I�������I�F�    I9�u�K�H���   H����   H�u L��H������H�E�    �E� H9�u�I��P  L������IǅP      H��[]A\A]A^A_�@ H���  L���q���H��   L��Hǃ�      �W���H��8  L��Hǃ       �=���Hǃ8      E�������Hǃ�      Hǃ      Hǃ0      ����� AWI��AVAUATUH��SH��8L��  H�^H���V8M�7L9��  A��PЀ�	vK<[tGI�FH9��2  �iBH �   L����� ���  ǅ      H��8[]A\A]A^A_�D  I�O H�$<[��  L��A�   A�WH�D$ =   �D$DN�L��A�W8I9s�H��8  I���   H�D$H��tDH�<$����H��@  H�<$Hǅ8      ����I��   Hǅ@      H��t	I���   ��D��(  Mc�H�<$1�L�L$,E1�L�Ѿ   E���   L�T$�����H��8  �D$,����   A�GH��8[]A\A]A^A_�f.�     I�FH9�vG�zBH �   L����� ��u/ǅ      �����A�G   H��8[]A\A]A^A_�f�     I�FH9���  ��BH �   L����� ���w  ǅ      �l����     L�T$H�<$L�L$,1�E1��   L�������H��@  �D$,��� ���I�E H�$D��I���   ��D$,��� ���E1�E��~7H�$D��M���   �    �ރ��   ��1H L��A��  A9�u�H�$L��A�W8M�/L9���  D�t$H�l$L���$    D�d$�]�    <]��  ��0��	waE����   L��A�WHL��I��A�W8M�/I9���   I�EH9���  L��A�W8I�/H9��b  �E <du�L�mI9�s
�}e�  E��ubL��A�W@A�G������I���f.�     A�G�   H��8[]A\A]A^A_�f�     I�F�D$A�   I��D$   �����H�EI��H9�v�} /u	�$9L$A�G   �����     A��I��L��M�/A�W@I�H9��w���A�W���k����$9L$~;L)�L��D��H�|$H�ōHA��  A�G���;���I���   Mc��J��� �$�����f.�     �}f������E<>wLH�6  !� PH�������f.�     H�l$M��ǅ      M�7�����fD  I��H�l$M�u�ڃ�߃�[���}�����A�} /�B����$9T$�5��������D  AWA��AVA��AUI��ATUSH��H��H  H�o�D$/ H��  H�@H�D$;U rH���   H�xh ��  A��   �v  A������M���t  I�M H��8  I�M(H��@  ��0  D��H��H��ǃ�       ��H��ǃ�   ltuo����1  D��L��P  ��L���  h��A ��PRH�D$(L��H��$�   �H�� A�ą���  ��`  D��H�L$/H�T$0��   H��$�   ��$  H��h  �t$D��H��$   H��p  ��$  H��$(  H��x  H��$0  H��h  H��$  ��`  ��$   ����A�ą��<  ��0  H�D$H��$�   �o�$8  L��$`  �o�$H  �L$H��$X  )D$@)L$PH�L$�P���   �T$�������   ���  H��$�   �M��H��$�   H��H�CP�M��H��H�CpH��(  �@ D�����D$�5  H���  H+��  H��H�ChH�Cxǃ�   ltuoM��tfA�}w
���      H�|$@   L���   uH�|$X   �  H�t$@L���ē��HcCPHcT$@H��H�H�� �  HcShH��H�H�CPHcD$XH��H�H�� �  H��H�H�ChH�t$H��L	�tL��L���J���H�D$LshHCPA��t�|$/ tj�|$ Hc�@  Hc�8  ��  H��$   ��  HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$`L��虐��H�T$`H�D$pH)�H�S@H�C0H�D$xH��H�CH�D$H+L$hH�K8����   H�shH�{0�Fb���   �A��1�1�M�������Hǃ8     Hǃ@     ����@ H��$�   L��(  �|K��H��$�   H��H�C@�gK��H�L$foT$@H��fo\$PH�CPI�M0M�u8A�EAUA] H�D$0H��   HcD$8H��  H���   H�@hH��t%H�xH� H�t$0�PHǃ       Hǃ      H��H  D��[]A\A]A^A_�D  H�D$H��$�   �P��fD  A�   ��H��$�   �Pf���C����z�H�@H��H��H�f�     HcH��H��I��I��?J�� �  H��Hc�H�P�HcP�H��I��I��?J�� �  H��Hc�H�P�H9�u�������    H��$�   �J��H��$�   H��H�Ch�J��H��H�Cx����f�     H�D$HHD$P�.��������ff.�     H���G  USH��H��H��h  H���   H��tH���#���Hǃh      ǃ`      H�������H���   H��HǃP      �����H��   H��Hǃ�       �����H��  H��Hǃ       ����H��  H��Hǃ      ����H��  H��Hǃ      ����H���  H��Hǃ      �j���H���  H��Hǃ�      �P���H���  H��Hǃ�      �6���H��h  H��Hǃ�      ����H��p  H��Hǃh      ����H��x  H��Hǃp      �U��H��x  H�������H��H  H��Hǃx      ����H��P  H��HǃH      ����H��X  H��HǃP      ����H��8  H��HǃX      �q���H��@  H��Hǃ8      �W���H��  H��Hǃ@      �=���H��  Hǃ      H��tH������H�C(    H�C0    H��[]��    �ff.�     @ ���  ��~cAUD�h�ATUH��S1�H��L���  �f.�     H�CL9�t'H��I�4�H��� ��u�H����[]A\A]��    H��1�[]A\A]�1��AWI��AVAUATUSH�
H��8H�H�|$H��H�^�F    �V8M�7L9���   I�6  !� PE1�1��xD  <c��   I�F
H9�tv=A�F	<>�(  I��s*f.�     ��BH �	   L����� ��tx�     I�W@L����A�G��ucE1�L��A�W8M�7L9�vMA�<eu�I�FH9�tv�A�F<>��  I��s��    ��BH �   L����� ��u��     A�GH��8[]A\A]A^A_�D  <FuiI�FH9�t#�e���A�F<>�h  I���N���fD  ��BH �   L����� ���,���A���  �t
��A���  I��M�7�����Ѓ�0��	w(L��A�W@A�G���a���L��A�   ������    <RudI�FH9������A�~D�����E�������H�D$I�/1�H�T$(H�t$ L��H���   H�xh ���������������   �����fD  <-uI�FH9��_���A�~|t��S���I�W@</�K���I�FH9��>���M�fL��M�'��A�G�������I�H��L)�J�������H9�����A�F��A�x1H A��FH H�t$�D$�v   ��I��0M�M�������A� 8D$u�L��L�D$�ǆ H9D$L�D$u�H�T$L��L���� L�D$��u�A���  �Ѓ���A�F(�������t��BH �   L����� ���k���H�D$H��P  1�H��t�
��HE�A�v��t^A�~��   A�N�$��DH ��߃�[���b�������D  ��߃�[������������D  ��߃�[������������D  L��H�|$A�VA�GA�G�������<��(���A�G    E1�����H�T$(1�H�T$(H�: tރ�	E1�L����L��v	A���   �A���   �H�D$H�   H�D$(1�H�T$(�H�L$H���   H�T$(H��t�H��  ��H�D$1�H�T$(H0  H�D$(�H�D$1�H�T$(H�D$(�n���L�|$(1�H�T$(�]���H�L$H���  H�T$(H��t�H��0  ��9���H�L$H��8  H�T$(H���X���H���  �����f�     AU1�ATI��UH��SH��H��f�H�    H�t$����A�ŋD$��uA���  f��vfD�+H��[]A\A]�H�t$H������H�D$��u�I�$��f�AW�   AVAUI��ATUSH��L��H��x�D$    H�L$H�t$A�Ux�T$��   ����   ��   ����   1�H�������D$����   �T$L��P  L���   ����   L�|$1��YD  I�t�H��tL���n����sH�T$L���>���H��I�D��D$��uC��I�7H��H��H��I���a� � 9l$~<I��8/uH��I�I�_H)Å�u�f��   A�EH��x[]A\A]A^A_��     �D$��f.�     AWAVI��AUATI��USH��hH�F L�.H�^H�D$H��  H��H�D$�VH���B  H�ډ�H�L)�H��H9�O����  A�v����  I���  A��(  H�D$(I��0  H�D$ I���  H�D$8���  �D$3 E1��D$4    �    L��A�V8M�>L9��  I�GH9�v<A�G<>�g  H�6  !� PH��sA�<d�e  <euA�n��  @ L��A�V@M�I9��e  A�V����  A�?/u�I�GL�D$H9��A  1�H�T$XH�t$PL��I��$�   H�xh �����������  A��(  ���6���L�D$I�WD��H�|$ I)�A�HL�D$A���  �D$L����  I��X  Ic�L�D$H��E��B� A�.u?I��X  ��1H �   H�<��L$4�t$3�� �����   AD�D��L$4@�t$3Ic�$<  H�L$P����  �UD9���  H9��K  H�|$H�T$LH���y���I�ǋD$L���/  H�T$PH�t$XL��� H�D$��  L��H�t$P�P H�L$PD��H�|$(Ic�$<  H)�L�H�L$PA���  H�|$L���D$L�+����D$L�r  f�A�d�=���D  E����  I��X  �|$3 E��(  H��  I��`  H�\$8�D$\1��D$X���H�ߋA��@  �D$L���]  I���  I���  �   H�ߋ
H�A��@  �D$L���/  H�\$ �   ��1H 1�H��A���  �D$L���  L�|$(�   H�T$X1�L��A���  �D$L����   I��   I��  D��H�ߋ
H�A���  �D$L����   I��   D��L���HI��  H�PA���  ����   A��(  H��h[]A\A]A^A_��    H�T$XD��H�|$(A���  �D$L��uQA���s��� ��߃�[�������A�<d�����A�e�����A�f�����E��������[���f��   A�FH��h[]A\A]A^A_��     L�|$D�mH�T$I���  D��I���D$L��u�I�H�T$D��I��0  ��D$L��u�I�H�T$�   I���  ��D$L�������뀾�1H �   H����� �������I��`  L�|$81��L��A��@  �D$L���>���I���  I���  �   L���
H�A��@  �D$L������Hc\$4I��`  �   L����I��X  H��A��@  �D$L�������I���  �   L����I���  H��A��@  �D$L�������I��   I��  ��L�|$ �
H�L��A���  �D$L���{���I��   ��H�\$(�HI��  H��H�PA���  �D$L���I���I��   1�L���HI��  H�PA���  �D$L������I��   1�H�ߋHI��  H�PA���  ���p��������f�     AWI��AVAUATUH��SH��HH��  L�v H��H�D$�V8I�L��I;Gs	�8[�y  A�WH�D$����  I�WI�H9�r H)�H�H��H9�~I���   �T$��  L��A�W@A����  I��X  L��H�D$A�W8A��P  ��u$H�D$L��t$I��X  H� ��D$,���  I�7H�FI9G��  E1��   �    H9���  H�T$,L������I�ŋD$,����  H�T$0H�t$8L���Dz H�D$��  L��H�t$0�P H�L$0��H�|$Hc�<  H)�L�H�L$0A���  L��L���D$,������D$,���q  I�7A��H�FI9G��   �   ��BH ��� ����   L��A�W@L��A�WH1�H�T$8H�t$0H��H���   L��H�xh �����������   L��A�W@A�O����   L��A�W8I�7H�FI9Gv#��BH �   ��� ��uL��A�W@L��A�W8I���  H��tE���L��L��L������A��P  ������Hc�<  H�t$0���~�����H�T$8��H�|$A���  �D$,�����A��P  ��u�D$A��P  H��H[]A\A]A^A_� A�W@L��A�W8I�I;Gs�8]t�A�G   H��H[]A\A]A^A_ø   A�GH��H[]A\A]A^A_�L��H�T$,�(   ����H��I���  �D$,��u�L��蔲���D$,���C����fD  UH���   �   SH��H��H��8H���Uh��~|H�T$H��trH��H��?H��H1�H)�H��   uiH�D$(H�$H���  H��H�T$ H���  H���  H�L$H��H���  H�L$H���  H���  H��8[]��     �E   H��8[]�f�H���  ��6��H�<$H��f���   ��6��H�|$H��H�$�6��H�|$H��H�D$�6��H�|$ H��H�D$�6��H�|$(H��H�D$ �6��H�T$H��?H��  ��H��   ����ff.�     f�L�GL�WI�H9�}PD�A��v<I�HH9���   A����H�<�   �   � H�PI�L�H9�}"H��H9�u�K�D��H���I�H����     I�T �M�L�UH��H��SH)�H)�H��I�I�,��5��H��H)�H��H��H�[]�M�Ѹ   ��f�     � PH ��A��fD  AWAVAUATUSH��L��  M����   A�D$@I��A��I��1ۅ�u�M@ H�EI���A9\$@v8��H�<�I�D$8H�,�D9m u�H�EL9��H�UH�u L9�}$I�7��A9\$@w�H��1�[]A\A]A^A_�fD  L��H)�H+uH)��4��HEI��D  H���   []A\A]A^A_�@ AUATUS�    H��M��II؃�-w��I���$�EH 9�`  ��  D  H������H��H��[]A\A]� H����  H����  ��0  �   f���@ H���g  H���]  ��,  �   f��@ H���?  H���5  ��*  �   f��x���f�     H����  H����  ��(  �   ��J��� H�L$L��  @ L���>u H�L$H�hH������H9�����H��L��H���t ����f�H�L$L��  �f�H�L$L��  �f�H�L$L��   �f�H�L$L���   �f�H����  H����  H��   �   H�����f�     H����  H����  H��  �   H��h���f�     ���O���H����  H����  �н   ��G  f��,���D  H����  H����  ���  �   ����� H����  H����  ��<  �   ������ H���_  H���V  ���  �   ����� H���O  H���E  ���  �   f�����f�     H���  H���  ���  �   f��X���f�     H��x  H���'�����H�L$��=��H���#����H�L$��I��$p  ���jH��t"H9�rI��$h  H�U�H�4�H����q �D(� H�������H��H��[]A\A]�fD  H���  H���u  ��`  �   ����� ��   �����H�L$9�(  �����H��@  ��L�,�L���r H�L$I��H�hH���_���H9��V���H��L��H���Tq B�  �>����    H����  H����  ��   �   ����� 9��  �������H���  ���jH�������H9������H�U�H���  ����� H�L$9��  �����H���  ��L�$��u���D  H���W  H���M  ���  �   ����� H���/  H���%  ��8  �   ��Z��� H�L$L��  �����    H����  H����  ���  �   ����� ������H��t-H��v'����  ����  ����  H���  f�H��   ����� H���W  H���N  ���  �   ����� H��t�H��v�H��   �   H�����f�     ���o���H��t�H��v����1  ���  ���+  H���  �e���D  H����  H����  ��C  �   ����� H����  H����  ��B  �   ������ ��A  9������H����  H���v  �н   ��G`  f������    H���7  H���.  ���  �   ����� H���7  H���-  ���  �   ��b��� H���z���H���p���H���  �a������C  9��)���H����  H����  �н   ��G�  f������    H����  H���~  ���  �   ������ ���  9������H���h  H���^  �н   ��G�  f������    ���  9������H���(  H���  �н   ��G�  f��^����    H����   H����   ��A  �   ��2��� H����   H����   ���  �   ��
��� ��@  9������H����   H����   �н   ��GD  f�������    H��tSH��tN��@  �   ����� ��B  9������H��t<H��v6�н   ��Gt  f��v����    H���   [H��]A\A]�D  �   �M���fD  �   �=���H���  �R���H���  �F���H���  �:���H���  �.���H���  �"���H���  ����fD  H��H�Љ�H���  ��H��H�4�����1�H���ff.�     H��  H�    H�A    H��tlL�@H�@P����H��H��H	�L��H��H�s�H�L�@I9�w>H��L)�H��H��H��?H�H��H��L��8D�HH��L	�H9�tH9�w�H�p�I9�v�1��fD  HcPHc@H�H�A1��ff.�      H�O����   L�G����   L�W8L�O(����   H�GhHGxHGXHGHL�L�L�H�H�H�GpHGxHGXHGPHG8HG0HGHGH�FH�GpHGxHGhHG`HG8HG0HG(HG H�FH�GpHGxHGhHG`HGXHGPHGHHG@H�F�f�     I�H�H�GHGH�F�@ H��@ K�L�H�H�H�G0HG8HGHGH�FH�G0HG8HG(HG H�F�f.�     USH��(H��P  H��t~H��H��  �UA��H������D9]D��FU��t1�D  H��H��H��9�w�A9�v+A����A)�H��I�J�T�fD  H�  �  H��H9�u�H��(1�[]��    H��(�   []�@ AVAUATUSH�� H��P  H����   I��H��  �UA��H��E���	���D9eDFuE��t)H�Ũ   1�f�H�4�H��H������I�D� H��A9�w�E9�v-A��D��E)�I�D� I�K�T�fD  H�     H��H9�u�H�� 1�[]A\A]A^ÐH�� �   []A\A]A^�ff.�      AVAUATUH��SH��   L���   H��P  H�t$0�����D$��tH�Ġ   []A\A]A^�fD  �D$0H�T$L��H�4@H��H�� �ۊ��I�ċD$��uT$4�L$0A�D$    I�D$    A�T$I�T$ A�$I�T$����   ��L�D$0H�IH��M�TPfD  I�HM�H�����H��L�
H�JI�x�B(����H��H�r H�H�zH��H�JM��t!�   ��1H L������� ��u9H�B thgwH��0I��L9�u��K�   ��93tfL�e H�Ġ   []A\A]A^�f��   �%DH L������� ��uH�B htdw�D  �   ��1H L������� ��u�H�B zspo�D  H��  ��H�t$H�è   E1������D$0��t.J�t�O�tm H��I��I��Mt$H������I�FD9l$0wҋD$�>���@ H����   AW�����AVAUATUSD�w�A9�AF�A�����   �A��D$� 1�A�   H�D$�A�^�E1�A�   L��  �    A��1��   E��u�Z�    H�ǉ�� �  A9�vH�<�   L��HN�H��IH�E��A��L��H)�E��HD�H��H �  H��H��H�GH9�u�I9t� t
I�t� �D$�H�EH9l$�t	H���q�����D$�������[]A\A]A^A_ø   �f�AWAVAUATUSH��   L��P  M���v  A��A�vI��H�|$D9�DF���%  I���   1��     L�ML�]D�} A9���   I�|� E��E����   I;9��   ��   �   E1�� �    I�H9�toH��H9���   Lc�A�@D9�u�K�D��H�D�H��H��9�w�H�\$H�T$H��P  �
�����uH�SE����   �΀H�SH�Ę   []A\A]A^A_�I�I���     A��I�D��I+H��H��?H�H���-���f�K��I��I�4�K+4�H)�H)��"��A�v�[���1�H�T$L���}����������H�D$H�PH�D$��H�P1��g����   �]���ff.�     @ AVAUI��ATU�   SH�� ��F�I���t(I��1�I���    I�<���!��H��I��H��9�w�L���L�������H�� []A\A]A^�ff.�     f�U��SH��H��P  ������uH�SH�р΀����HD�H�S[]�ff.�     @ 1�1��f.�     SH���   �`BH H��p  H�x��N��H��tH��tH�H��t	H��[�� 1�[�@ ATI��USH��H�?����H�;L��H���`9��H��tH�CPH�S(E1�1�H�s H�8�U[1�]A\�ff.�     f�SH��H��H�?�`���H��1�H��t(H�H�T$H��8  H���   ���uH�SPH�L$H�
H��[��     H�GPH�8 t.SH��H�?�
���H��t
H�SPH�:�PH�CPH�     [�fD  ��    AWAVAUATE1�USH��H����  wk���  ��~aH�t$I��D�x�1�L���  �D  H�CI9�tWH��I�l� A��H��t�A�8E u�H���b H9D$u�H�T$L��H����� ��u�H��D��[]A\A]A^A_�f�     E1���ff.�     AWI��AVAUATUSH��H��hL�f8H��  �D$(   H��tL���l���Hǃ      H�T$(�X   L��蟃���L$(H�Ņ�t$H����   �D$(H��h[]A\A]A^A_��     I�wL���q���D$(��u�H���  �o��  �o��  L��  H�E(H���  EH�E0I�EHMH����   I�OHI�W@H�|$0I�w8��D$(��t?<uI�GH��vI�W@�z�   L����q��H��L���}����=����     H���   H�|$0H�l$@H�D$PI�EHH�D$H B �PH�|$0�D$(I�EH�P�D$(<t���u�H�E�oU�o]H����  H�ChH�E��  H��H�CpH�EH��  H��H�CxH�E H��  H��H���   H�E(H �  H��f���   H�E0H �  H��f���   �EP������H�K@L��H��  ��p���N���f�     �JH9������I�G8I�OH�D$,    H�D$H�BeH9���  �Bd�����Bc	���H�DuH�pH9���  �p���0��	�f���i  �@H�H9��Z  L�pL9��Z  �P�����	��EP��L�H9��7  f���!  H�|$��E1�1�L�L$,�   �B����|$, H��H�EHH���	  �EP�KHD�,�    H���   M�H�D$��~6H�CPH�0f�~��   H����H���H�0H��f�~��   H9�u�M9�sVA�6H��H�T$I���>��H�T$H�߉A�v���=��H�T$�BA�F�H������A�F��B�    	Ș�B�M9�w�H�|$ tH�t$H���fD���D$,�|$, H�}Hu3�uP�   �@�A �eg �T$,��u`�D$(    �r����D$,   H�}HH��H�|$������D$,H�EH    �EP    �D$(�9���H��H�T$��C��H�T$���D$,����H�}H��    ATI��1�UH��SH��H�� �(k����tH�� []A\� H�T$H�t$H���������u�f�|$�t1�H����j����u�H��H����l����u�H�{@H��L���� �   H�߅�ED$�'n���D$H�� []A\�f.�     AW1��Y   1�AVI��1�AUATUSH��H  H��  M���   IǆX  ����H�\$pM���   Aǆ`      Aǆ<     H���H�L��H�      H��I���  Iǆ�  \  H�EIǆ�   �' �E1Һ   ��BH L��L��$   HǄ$      HǄ$      HǄ$      HǄ$       fD��$(  Ƅ$*   �o����D$`���1  <�  ��$)   �D$`��  �D$XH��$�  H��$�   H��t	H���   ��H��$X  H��t	H���  ��H��$�  H��t	H��0  ��H��$�  H��t	H���  ��H��$   H��t	H��X  ��H��$(  H���%��H��$(  H���_���H��$�   H��$  HǄ$(      H���;�����$)   HǄ$      ��   H����$�   �D$XH��H  []A\A]A^A_Ð�
   ��BH L���>����D$`�������1�L���hh���D$`�������L�l$hH�t$\L��L���7����D$`�������f�|$\���   1�L���$h���D$`���}���I�t$H�t$h�y@ H��$  H���h���HǄ$      �6����    H��$  L���@����D$`HǄ$      �D$X���/���H��$  1��   D  Ƅ$(  H�t$hI�|$( ��  H�D$`L��H����{��D�L$`H��$  E�������H�T$hH��L���h���D$`�������H�L$hH��$  H��$  �D$X    H�
H�T$xH�T$pH��$�   H��L��������D$X���v�����$(   L��$   �D$\    L��$�   �U  H��$  H��$  I��H�1�@ I��L9��  A�<$eu�I�T$	H9�v�A�|$eu�A�|$xu�A�|$eu�A�|$cu�I��
H��H�L$pL��$�   L9�r<�  @ H����$�   D��$�   E����  H����$�   H�D$pI9��r  �8eu�H�PI9�v��xeu��xxu��xeu��xcu�H��$  H�$  H��H��$�   ��$�   L��$�   L�l$p�
   L��L��L)�H��H�L$�d� H�L$H����  H�ʾ   L��H�D$�A� L�D$I9�������M9���  A�U �J����q  �� �h  ��u���[  H��$  H��L)�H�$  ��$)   H�D$`�o  Ƅ$*  H��$  H��$   HǄ$      HǄ$      I�EI9��  A�E �PЀ�	v��߃�A<��  A�E�PЀ�	v��߃�A<��  A�E�PЀ�	v��߃�A<��  A�E�PЀ�	v��߃�A<��  H�EH��L�l$pE1�H��$   H��$  H�L$h�P0H�D$hH��$  H��$   � H��$   H��$  �q�  �U H��$   ��  H��$  �  H��$  �@ H��$  �@ H��$  �@ H��$  H��$   H�T$xH�
H�T$pH��$�   �D$\�D$X���.���H��L�������D$X������I��P  A��@  �H���$  ���  ��t;Pt
ǀ�      ���t�P��uL��覼��I��P  H����  �P��t5���    ��  ��H�RH���D  H�����    ��  H9�u�A��`  ����  H��$�   ��$�  �D$8A���  tb��$�  HǄ$�      A��`  H��$�  I��H  H��$�  I��h  H��$�  I��p  H��$(  HǄ$(      I��x  I���   H�xh �J  H��$   A��   HǄ$      I��P  H��$(  I���  H��$0  I���  H��$�  HǄ$�      I��X  H��$�  HǄ$�      H��I���  �e�����$X  ����  I��8  ��L�t$HE1�H�D$(�D$8H�L$I��@  I�փ��D$<    H�L$H��$`  H�D$@H�L$ �D  I�D$L9d$(�(  I��H�D$1�fB�4`H�D$J���1H H�D$ N�,�A�D$�D$M��t��L$8��~�E1�L�d$0M��L�|$@� I�D$M9��B  I��K�,�L��H���f� ��u�M��H�D$L�d$0H��   ��1H fF�<`H�D$J�,��L$<�� ��D9��=������D$D��D$<�+���H��$  H��$  H�1I9������fD  �   �����fD  L��L�l$h�#a��H�l$H�D$H�D$`HǄ$       H��H�D$�*fD  H�t$`L��H�H��$   �`���D$\�������H��L��L�������D$\�������f�|$h�H��$   t�H�l$H���+  �D$X   �Y���fD  L�d$0�F���fD  I�D$L��I$H��$  H��$  Ƅ$)  ��_���D$`�������H��$  �N���fD  L���ȸ��I��P   �`���f.�     Aǆ`      �U���L�t$HAǆ,      �D$<A��0  ��$0  A��(  ����f�H��$   ������D$X   ����@ L�L$XE1�1Ҿ   I���   �u����|$XI��h  �������Aǆ`      �=���f�H�t$L���^���D$\������H��$   H�T$\L����r��H��$  �D$\�������HǄ$       L�|$�5 f�|$h�uOH�T$`H�L���_���D$\�������H�D$`H�$   L��L��L������H��$  H��$   �D$\��t��D$\    ������D$<    ����I���l����   �_���H��$  H�T$`L����O H��$   H��$  ����H�pH�T$\L����q��H��$  �D$\������H�D$`H��$   ����f�AVAUATU�պ   SH��H��H�   H���   ��BH �b;����BH H��  I��H���   H�x�;��H��  H���s  I��H���   �`BH H�x��:��H��H��p  �\���A�Ņ���  ����  ����  ��  Hc��  H�C    H�C H�CH��H��
  ��(   H�St
H
  H�CH��P   tH�K   H��  H�C0    H�K(H���G  H��  H���G  �@ ��t4�1@8��x  < ��  <-��  @�� t
@��-�   H����u�H�C0�BH H��    H�C    H��  tH�C   H��t:�DH �   H����� ����  H�ƿCH �   ��� ����  �H���  H���  �C8    H�C@    H��H��H�ChH���  H�{pH����  H���  H��H����  ���   H�sxH��H���   f����  �@A���������A����A������D��f���   )�D)�f���   H��9�f���   H��AN�f���   ��������  ���   f���   ��*  ���   M����   M�f@1�H��1�H�cinu  H�$H�D$I�|$�>���A�Ņ�t<�uZ��   �   f�|$����  �  ����  ��u*�   �D$EBDAI�|$f�L$H��t1�H��1��އ����A��H��D��[]A\A]A^�f�     H��  H��tH�C(H��  H��   H���  H�C0H�C    H�������������    H�K����fD  �BH��H���g����    �BH���S��� H��A�   [D��]A\A]A^�f.�     A��  ��  fD���   A��  �8���f��������   �D$CBDAI�|$f�T$����� H��A�   [D��]A\A]A^�f�H�<$�	��H��f���   �����    @�������H�S0�����fD  1�H��H�C0�BH ��H�C�����    �   �D$1talI�|$f�D$�]���@ 1��D$BODAI�<$f�t$�A���H�H��P  H  H�G1��f�     H�G    ��    1����   w
H�G���p�ff.�     �1��    ���   w"H�O���    �Q��uH����   u�� ��D  L�H��I��P  I���   H��    H��`  t�P$E1�H�A�@6B ��f.�     ��   �f.�     H�H��P  H��`  �`ff.�     �H�H��P  H��`  �`ff.�     �H��p  H�    H�A    H��tSH�����   H�H�1�[�f�1��ff.�     f�1��G���fD  H��P  � H��t��L  ��  t�1��ff.�     @ H��P  1�H��t2��L  ��  �   t!9q$r1�H��tH��   ���q�
�D  �ff.�     @ H���  �`fD  H���  �`fD  H���  �` fD  H���  �`(fD  H���  �`0fD  H���  �`8fD  H���  � �    H���  �`8fD  1����   w
����? TH �ff.�     H�WH��t�����   <t1��D  ��+G;G��   D�D�WD��D�BI���A	�E��D9�r�D�J�BH�JE��D�JA��E	�E��D9�s-�Nf�     �H���Q���A���Q�D	���9�r,A��I9�w��l���@ ���2�f�     �G�D��E��D)�D�O�W�G��    H���  �`@fD  H���  H��t�`H��ff.�     @ H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ SH�H��H�w H���   蹣��H�C     �C    [��     AUI��ATUSH��H��H�wH��t2�W��t+1�fD  A��L���J�4��f���H�sJ��    9kw�L���M���H�sH�C    H��t6���t0E1� D��L��A��H��H�t.����H�sH�D.    D9#w�L�������H�C    H��[]A\A]�ff.�     USH��H�GH��P  H��X  H��t.H���   H���`BH H�x�0��H��tH���UH��(  H�B@H��1�[]�ff.�     �H���   1�H���H���H  @�~��t�H���P  f�LFH��9�w���I  @�~	��t!1�f.�     H����  f�LF(H��9�w���J  @�~
��t!1�f.�     H���  f�LF<H��9�w���K  @�~��t!1�f.�     H��  f�LFXH��9�w�H���  H�FpH���  �FxH���  �F|H���  f���   H���  f���   ���  @���   ��t1�@ H���   f��F�   H��9�w����  @���   ��t1�@ H���h  f��F�   H��9�w����  ���   Hc��  H���   ���  �F�ff.�     H�H��tHUSH��H��H�8 H�h8tH�w8H���S��H�s0H��輠��f��CC C0H��[]�f��ff.�     @ H�GH=@gH tlH=�gH tdUH����1H SH��H��H�H���   H�x�X.��1Ҿv.H H����.��H��tH� H��tH��H��H��[]��fD  H��1�[]��    ��   �f�USH��H��P  �Gt
H��p   uH��8  H��[]�D  H���   H����1H H�x��-��1ҾV.H H���Y.��H��t�H� H��t�H��H��[]���AWAVAUATUH��SH��H��tH�    E1�E1�1�E1��   A�   D  ��t	H��H9�s;�E��A)���D������tM��	�|   I�����~CI����t�H��H9�r�f�E1�L��H�؅�LE�H��[]L��A\A]A^A_��    �   뉐��uM��uE1��w����    O��H�I��N�@�]���D  E1��
��   ���  ����  E1�M���y���L�N�,O�4+H����  M�I����  I���  �8  M��M)�M��~RI���   IN�H��L)�H��~:L�� dH I)�M��I���  ~"L��I��?I��H�gfffffffH��H��L)�I��I��L�U �����fD  A�   f���tH��H9�������E��A)���D�����	������uM��uI����t���f�I������I���O��H�I��N�@롐�D$   E1�E1�A�   @ ��tH��H9��G����E��A)���D������	1I���  O��H�N�P��t����     A�   ��     �D$��t'E�������I��M��������h����D$    �i���M�������E���I���A��������L��J�4��cH H�H��H=�  ~tJ�4��cH L��I���H���L�u I������I���I����l���M����   M)�I��
tmM����   I��N�� dH L��H��I�� �  A����LL��+���L��I�������L�u I������L�Ǿ
   �����I��L��L)�H��H�E �����L��I��?� ʚ;H�gfffffffH��H��L)�I��L��H�H��H=�  �����L���n���I������L��I��M�H�J�<� dH I���+���J�4� dH 뷐AUATUH��SH��H��L��P  H���   A�}(��   �   ��BH �*��H��H����   A�E$����   E1��8 ��  A;�H  sI��P  H�4�H��tH���� ��t`A��E9e$vSI��   D���<Bf���w��U(H����fD  H���1H ��(��1ҾK.H H���s)��H��tH�@H��uD  E1�H��D��[]A\A]��    H��H��H��[]A\A]��fD  AT1�USH���O �D$    ����   I��A��H������   H�G�V�1�H�4P� H���f9�B�H�HH9�u��˾   E1�H��L�L$1�L���=q��H��H�E�D$��u)D��H�EH�� �Pf�NH��H���u�] 1�D�e$H��[]A\�@ L�L$E1��   1Ҿ   L��1���p��H�E�D$��t���ff.�     ��? �   t9wt�9Wu�1���t�H����H�wH��H����� ����H���D  AWAVAUATUSH��XL�w�D$L    I�F� H�D$��t&A���  9�t�   H��X[]A\A]A^A_�fD  A9��  v݉��T$(�W I��H��I��  L�G(�t$,�(H�L$ H��L�L$LH�|$�   H�D$�MH��H����o��I�E(�D$L��u���A�] L�\$��   ��M��1�M��H�D$�D$(��L�L@I��M���Lf�     I�S�E���A9��  �/���I�H(�t$(L�4�    J�1��ui�    H�EH9l$tH��H��u�I�@(�    H�EH9l$u�M�ŋD$,�|$(A�E���  �D$(A�E A�E�D$LH��X[]A\A]A^A_�@ I���  L�d$ �   1�L�T$L�<� I�?�   H�H�H�wH9�AH�H9�8H��I��A��I��?E��tH��u �   H��tM�$L9�L9�}H1�fD  J�41H��I��HcH��H��H��?H�� �  H���L9��w���L�T$�����D  L9�t�L�D$8L�\$0~!L��H)�H)�����L�D$8L�\$0Hc�I�H(�H��L)�H)�H���ڋ\$(A�UL�L$L�   H�|$M�EH��H��H����m��H��I�E�D$L���}���H�t$ H����8 ����AWI��AVI��AUATUSH��H��HL�?H�0 H�$D�oM�g8�D$8    H�    ��  E��u�D$8H��H[]A\A]A^A_��     1�A�ML�L$8E1��   L��L�T$H�k(�,m���T$8H�D$ �Ѕ�u�L�T$I�t- H�t$(M����  H�T$8L���Z���T$8L�T$I�ǅ҉��{���H�D$ �KL�K8L�8����  H�D$ 1�1�A�   L�`�zfD  H9k(HFk(M���  H�T L�I�$H9�tAI�|$�L�L�T$H�L$H)�L�L$�y7 I�$H�L$H��L�T$L�L$�  H��I�$�CI��I��L9�r:H�C0J�,�H��H9��w���M����  H�1I��I��L�I�D$��CL9�s�H�D$ �T$8I�M��tM�:H�<$��H���x���H�L$(H��k���f�H�T$�D$<    E���O����GA�mE1�1Ҿ   L�L$<H��L��D$�k��D�D$<L�T$H��H�C0E��t>fD  L��L�T$�K����D$<L�T$H�C0    ���D$8�����D�k�����D  �sL��Hs�D��L�T$���D$<��   �D$L��L�T$H��H���gF��L�T$���D$<ueI�G@�|$H�S0H�4(@����   @����   @����   H9�s�H��H��ɉ�H�z�H9�w�L��L�T$�G���|$<L�T$��tUH�s0����@ H��I�1I�$�,����     L�K8H�D$ E1��sL��������H�D$ I��[���f�     D�k�D$8    ����I��6���H9��o����H��H�����H���	���H�J�H9�w��H���1�H9��=����4H�4�H��H9�u��'���H9�������xH��H������	��x�	���H�z�H9�w���������t`��t���   #��u���H��f�H�W1�H9�r5�Gȉ��D  H�O1����   ~JH9�r��   )��W��)Ѓ�lH���    H�W1�H9�r��G�����G	�H���f�     H9�rˁ��   �G���DlH���    ����  t@���  wH��`  H��t,H�@(����@ ��  1�;�H  sH��P  H���@ 1��D  H��P  ��H��   �4p�f.�     AUATUSH��H��P  H��tP��L  ����  tTH��I��I��H��tH��x  H��tBI�E M��tH���  H��tEI�$H��t
H��X  �E 1�H��[]A\A]�D  �   �鐉�H������H��x  �D  ��P  H�������H���  뤐AT1�USH��L��P  �D$    M��t2I��$p  H��H��t2�oE �oMK�oU S H�U0H�S0H��[]A\��    H���   H�T$�8   �U��H�ŋD$��u�A��$h  L���O���A��$l  L��H�E �;���A��$t  L��H�E�'���A��$x  L��H�E����A��$|  L��H�E�����H�E I��$�  H�E(A��$�  �E0I��$�  f�E2I��$�  f�E4�D$I��$p  ����f.�     AU1�ATUSH��L��P  �D$    M��tI��$�  H��H��t�f�U H��[]A\A]�fD  H���   H�T$�   �T��H�ËD$��u�1�A��$H  L��f��2���H��t}�pQH H���� H��tkL�h��1H L���� H��tUI9�tPH� $     �,@ �f���w0���f�fA�M �T
�f�I��L9�tA�U �JЀ�	vˀ� v1�f��I��$�  �D$�����    H��r���SH��P  �`BH H��X  H���   H�x�<��H��tH��tH�H��t
H��[��@ 1�[�ff.�     �AWAVAUATUH��SH��H�wXH�?�s��H�} ����H����   I��H�E H�U(E1�H�u 1�L��P  H�EPL�8M���  I�?A�UA��0  ��tv�X�H���RD  L��H��L��H�L$�E���H�L$H�}(L��H�$H���-���L�$H��I�|H��E1�1�L��A�UH���tI��8  L�M H�HhI9�u�H�U(��H��1�[]A\A]A^A_�ff.�     @ AUATUSH��H�GPH�(H��tjH�?L���   H��P  ����I��H��t-H�} �P��0  ��t��H�\� H�;H��A�T$H9�u�H��H��L��[]A\A]隌��f.�     H��[]A\A]�D  AWAVAUATUH��SH��H��(H�?�Gt'H��p  H�T$���   ����   �����H�} H�EXH�����H�} �����I��H����   H�E H�U(E1�1�H�u L��P  H�EPL�8M���  I�?A�UA��0  ��tw�X�H���SfD  L��H��L��H�L$����H�L$H�}(L��H�$H���m���L�$H��I�|H��E1�1�L��A�UH���tI��8  L�M H�HhI9�u�H�U(��H��(1�[]A\A]A^A_��    H�t$H���;���H��([]A\A]A^A_�ff.�     �AWAVAUATUH��SH��  H�?�D$    ����H����   I��H�E H�T$�  H���   L��P  �O��D�t$I��H�D$E��tH��  D��[]A\A]A^A_��     I��h  H�t$ ����H�E L��H�t$ H���   A�$A�ƉD$��u�A��0  ��tr�X�I��H���D  H��H���tVI��8  H�t$ �����H�E I�H�t$ H���   A�$�D$��t�A���O���@ D�t$�����H�EX�8���D  H�EPH�L$H���f�UH��SH��H���H�t$�;��1҅�u%�;��t1��     �tH��H��H	�9��E H��H��[]�ff.�     @ AW�   AVAUATUSH��(�D$    H����   ���wH��9���   H�G0I��L�?H����   ��L�$�M����   �}���H��H�H�t��D  H��H9�tjH�H��t�I�WH�s H��H9��J  H��H)�M��tSL9�vNL)�H��H�H�C8H����   J�D �I��D$H��([]A\A]A^A_�f�     E1�I�WH�s H��H9�w�I�    �D$H�    H��([]A\A]A^A_� �wH�GH�L$H��wL����H���8���D$��u�L�kH�;H�T$L���K���I�ċD$���d���M��H�L$�n����@ 9k�b���H�;H�T$L��H�L$������H�L$H��t�������     H�C L��I�t��_8���D$�������L��H��L���u;�������H��H)�H9����������ff.�     �USH��H��(H�W8H��tfH�j8H��8H�L$H�T$������D$��uGH�D$H��H�T$H�p�)L��H�ŋD$��uH�T$H��uD�D  H�{p t H��(H��[]�fD  1�H��(H��[]�@ H�{8H�t$�J9��H��(H��[]�H�t$H���) H�T$�ff.�     �AWf��AVA��AUATA��UH��SH��H��L�n8H�7H�G8    L�|$GGG(H����7��L��H��H�CE��tk�A���|$��u.A���C   E��ul�D$H��[]A\A]A^A_�@ �D$   H�s0L���4���H�C0    �D$H��[]A\A]A^A_�f�     �;���t$��u�D���C   E��t�L��H���;���L$��u��P���w��CA�t$���SH��HSD�cH��H�H)�H�S �6���D$���`���H�;L��H�s�����T$���E���H���4���H�p�H�s(E��t'H�S8H���#9���D$������H��[]A\A]A^A_�H��� 6���D$��f.�     UH��SH��H��H���   H�@hH��t$H�xH� H���H�$H�HcT$H�U H��[]ÐH��P  H��8  �M���H��[]�fD  H��H���   H�@hH��t$H�H�x�T$H��H� H�$�PH����    H��P  H��p   u�H��8  ��6����f�     AWAVAUA��ATI��U��SH��H��x  L�wM��P  A��L  ��  t<I��(  H��t0E��t1E;�0  ��  A�   H��x  D��[]A\A]A^A_� E9o$v܉����   E�I���  H�D$H�@PHǃ8     H�D$Hǃ@     M��tLI�D$ I�t$XH��8  I�D$(H��@  �����H9�t%I�$H��p  H���    t@����  fD  �� @  �F���E��0  E����  I���  �D$( �Ao��  �Ao��  H�D$I���  )D$PH�D$ )L$`��A��L��L��ǃ�       ��A����A��ǃ�   ltuo������ЈL$0A�ȉD$<��A��h�BB h�BB ��1  H�D$��0  H��H��$�  �_AX��   tƄ$
  H�L$pH�T$HD��L��Ƅ$   �L���A�����Y���H�D$D��L��H��$�  �PA�����8���H�L$1�H��$�  H��$�   �Q0H�D$H�T$pH��$�   H�t$H�PA��<���  H�T$pH�t$HL��D�L$�*���D�L$E�������I���   H�xh ��  Hǃ       Hǃ      D�L$H��$�  ��$   I���   D�L$H�@hH����   H�L�BM����   H��$�  H�xD�L$D��H�D$x    H�L$pH�T$pH��$�  H��$�   H��$�  H��$�   1�A��H�T$pD�L$��H��$�  H��$�   H��$�  H��$�   H��$�  �I  A��A��   ��  H��$�  H��(  H�t$fod$PH�S@H��$
  fol$`H�SPH�p0H�t$ `h H�p8�@���� I��8  D������A��0  ��9�r�B���I���8  I���  �D$( �oP@�oXPH�ppL�@hH�@x)T$P)\$`H�t$H�D$ L9�����H��8  L��H��L�D$0H�L$(�����L�D$0H�L$(H��8  H��@  L��H�������D$(H��@  �����fD  H��L���   ��L��H��$�  L���   RD�����   AZA[A�����8�����$�  ǃ�       ǃ�   stibH��H�C0��$�  H��H�C8H��$�  H��H��H�C@H��$�  H��H��H�CH��$�  H��H�CPH��$�  H��H��H�CXH��$�  H��H��H�C`��$�  H����H�Ch�+  ���   ���   I��p  1�D��L��D�L$L�D$pH��$�   ���   �D$pD�L$H�CpA���   ��  fA��   ��  D�L$L�D$pD��L��I��p  H��$�   �   ���   �D$pD�L$H�Cx�H���F�,hE���X����/���D  H�D$ƃ0   H��$�   H�T$pH�t$H�P�D$(A���D$0 ����D  fA���   �I  I��p  1�1�D�L$f�L$HD��L�D$pL��f�t$pH�L$H1����   �D$pD�L$H�T$HH�CPH�S@H�CpH��(  �@ A���   �2  fA��   �#  1�1�D�L$L�D$pf�D$HI��p  H�L$HL��f�T$p�   D��A�   ���   H�D$HD�L$H�C`�D$pH�ChH�Cx�   ǃ�   ltuoǃ�       M��tfA�|$�%   ��H�|$P   ���   L���   uH�|$h   �f  H�t$PL��D�L$�$��HcCPHcT$PD�L$H��H�H�� �  HcT$hH��H�H�CPHcChH��H�H�� �  H��H�H�ChL�t$L�l$ L��L	�t L��L��L��D�L$�!��LsPD�L$Lkh�D$<u�|$( tj�|$0 Hc�@  Hc�8  ��   H��$   ��   HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$pL��D�L$�� ��H�D$pD�L$H��$�   H�C@H)�H�S0H��$�   H��H+L$xE��H�SHH�K8��   H�KPH��H��?H�H��H)�H�CX�V���fD  fA��h  ���   A���  A���  )�H�H�Ch����@ ���   f�������z�H���   H��H��H� HcH��H��I��I��?J�� �  H��Hc�H�P�HcP�H��I��I��?J�� �  H��Hc�H�P�H9�u������    H��$
  H�CPH�Cp����� ������H�shH�{0D�L$����D�L$�c��� H�D$XHD$`��������� A���  A���  )�H�H�Ch���� I��h  H���l���D��H��I��p  H�D�H��   H�D$pH��  �A���D  fA��h  �tEA���  A���  )�H�H�Cx������     ���   ���   ������    A������A���  A���  )�H�H�Cx�{��� H��tKH��t&��uH�GH9u(���� 1������f�     ��������     �#   �f.�     �%   �f.�     AWAVAUATI��US��H��(H�GL���   ���   H�w% �  ��  �H	�����   H��t�   ���  t^A��$�   ti��tML��D�<L�t$L�l$@ I��$p  ��M��L��   L���H�����   �D$H�E�A9�u�D  1�H��([]A\A]A^A_��    ���L��A��A�͉D$A����u"�� E��I�GxIDGp��H��H�E�;\$t�I��$�   D���L��������t�H��([]A\A]A^A_� H��t�   ���  �k���fA��$�   �q������Q���L��D�<L�t$L�l$I��$p  ��M��L��1�L���H�����   �D$H�E�A9�u�1�����f�     UH��H��x  SH��H���x���H���  H���Yw��H��8  H��Hǃ�      �?w��H��H  H��Hǃ8      �%w��H��`  H��HǃH      �w��Hǃ`      H��[]�f�     H����  AVAUATUH��SH��p  L���   H��t�PH��P  H���4  H���   L�c����H��x  ����H�{8����H��8  ������0  ��tGE1��     J���8  H��tL�������I��D9�0  w�H��8  L���?v��Hǃ8      H�Cǃ�       Hǃ       H��(  ǃ      L�h8L����u��H��   L��Hǃ(      ǃ0      ��u��H���  L��Hǃ       ǃ      Hǃ      ����H��h  L������H��@   tH�{H��@  ��'��ǃH      H��p  L��ƃ8   ǃ<      �Xu��H��8  L��Hǃp      �>u��H��@  L��Hǃ8      �$u��H��P  L��Hǃ@      �
u��H��X  L��HǃP      ��t��H���  HǃX      H��t#H���  ��H���  L����t��Hǃ�      H���  L���t��H��P  L��Hǃ�      �t��HǅP      H���  H��tH���PHHǅ�      []A\A]A^�@ ��    �>H��tpH��H��H��I������H��M��u.����H���  H��H��  �H��H�� ���HN�H���f�H��H��?H��H1�H)�J;ŠcH J�� dH � H��1�H���+��� H��H��  �����HO�� AT��   USH�o H�U H9W(��   L�g8H��H�u 1�H��/���H�������H�uH�{1�I��$�   ����H�������H�uH�{1�I��$�   �����H������H�uH�{1�I��$�   �����H������I��$�   1�[]A\�ff.�     �H��<t><�tH�7H���g����    �F�N�V����	�	Ѓ���H����    H��H��H�71�1�H������H��H���f�     AWH��AVAUATI��USH��(H�wH�T$H�W H�GH�W(H�wH9���   I��I���ff�=�   ��   D9��  H�rI�t$(L�2���v  ����  ���[  I�VI�N=�   HG�I��L9t$��   I�T$(M�l$ A�H��E�L$0L)�H����A����@��A���r���D9���  L�2���-  AD$4�   � ZH =   u��   f�9Ct3�S H�� ��u�I��M�l$(L9t$�v���1�H��([]A\A]A^A_� I�D$8D�CJ�, ����   ���  ����   �$ՠQH f.�     I�|$I�u �   �����S��tM����  ����  H�E fD  I���;�����M�l$ �U����I�|$I�u 1��p����S��u�f�E �ɐL���S��t��7����I�l$8���k  I�u I�|$�����s���I�VH9T$�I  A�FI�ր������I���V����    9s�SFs@�4���R���I�D$E1�H�D$�F�I�D�H�D$� fD  <tTL�} �CH�L9l$����I��I�u�H�|$�����I��C<t<u�D�} ���    fD�} �f�     D�} �I������H�L$I�FH9��3���A�FI�v������tx��<tqI�FH�y�* �P�I�Ɖ�@��@���`�����H�����P���H9�u�1������D  �E �P����     �E �@���H��(�   []A\A]A^A_�I������ff.�     �AVAUATU1�SH��`H���    H�_H��(  Ɔ!   t
H���    uH��`��[]A\A]A^�D  I��L��H  I��1�H��P  L��HǆH      H���H)����  ���H�L��X  Hǆ�     Hǆ�     D��4  ǆ�  ����Hǆ�  \  Hǆ�   �' H��  ��P  A�}0 ��   I�U �a   �a   �    L�2f��H�T$I��D$H1�E1��   D$8D�L$PL�L$�|$DL��D$D$(L�T$H��D���T$H�D$0����   �l$@H�D$8I��$�   H��Iu�,���Ņ�uI��$�   H��� ���Ņ���   H�t$0I��$`  AǄ$p      I��$h  H�D$H�8�Nm��H��`��[]A\A]A^��    A���  I�U � P  �HH������D  H��L���m���D$H�D$0    ���H���1�1��x����    H�SHH�s@H�|$�F���H�߉��� �����H���I��$�  H�t$0A��$H  �H��x�,���IǄ$�  �h�:����f�H��I��$�  �	���SH�_8H��t6H���  H��t*��!   ��   uH�G H��H�0�L������  1�[�f��   [�f�     SH�_8H��t&H�G H��H�0����1�ǃ@    [��     �   [�f�     AT��   USH�o H�UH9W(rFH�_H�u L�g8H�������H�uH��A��$�   ����H�uH��A��$�   ����I��$�   1�[]A\�ff.�      H�W ��   H�J(H9O(s�@ USH��H�H��H�2H�o(�O���H�P�H���   H��w'H�S(H+S f��4  1�H����f��6  f�K@f�SBH��[]�ff.�     @ AT��   USH�o H�UH9W(s	[]A\�@ H�_H�u L�g8H�������H��x/I��$�   H�uH������H��xI��$�   1�[]A\��    [�   ]A\�ff.�      H�G8H���K  AWAVAUATUSH��8L���  M���  M��X  ���  I��I��   E��P  H��L���D��������tL��D���H����������  I�G(M�gL��H�p������H��A9G0��  I��(  E��@  �D$,    I�O H�xI�G(D��H�X���   H)�H��A9���  A��p  D�\� A��t  D�9���  D)�A��p  �+�D$���D  ��f�A��I��H  L��T$J�4�H�h�R����T$A��A��A��@  �9  �   )ЉD$fD  I�G ��D�JL��H��D�D$H�4�D�L$�����E�D�D$D�L$A��D$D��D�A;�@  r�I��h  I�W D����J��H�PI��h  � �I��h  H�PI��h  D�����I��h  H�PI��h  D�����I��h  H�PI��h  �(I��h  H�PI��h  D� I�O 9\$t&D�������fD  �   H��8[]A\A]A^A_�@ �D$H��I�G(�D$,AƆ!  H��8[]A\A]A^A_�f�     A�������     M��`  I��h  A�L�L$,�   D�\$M��H�D$L�T$��>��H��I��`  �D$,��u�A��p  D�\$L�T$E�t  H��H�I�O I��h  D�I9������M�������M�G(H��L)�I9������H���    H�:I9�wH9|$vH�H�:H��L9�r�����D  �   �f�AW��   AVAUATUSH��hL� I�W0H9W(�p  L�g8I��E1�H�       �H��������A�D$`�   f�H=�� ��  H=?B ��  H=�� ��  H=�����  H= ʚ;��� �'  ��HL�D����A����	H��H�H��H=�  sMc�N�D40�����J�4H��tJ�D40H9�HL�H9�HO�I��I��0��   K�<7�?��  K�t7����H��H=�  �>���J�D40    H����    ��Hc�H�4� dH J�L40�����fD  H�$H��I�D$@H�D$I�D$PH�D$I�D$HH�D$I�D$XH�D$ I�D$pH�D$(I�D$xH�� dH I�D$h1�H��h[]A\A]A^A_�@ H�C	H��	��   H��H)�H��	��   H��������1�I�      �I�       ��6�     I��I)�I9���   H�H�H��H�D  H��H��0�*���H�H��t�H��H+T0H�4� dH H��H��H��y�N�I9���   H)�H�H��H�� I�D$@   1�I�D$P    I�D$H    I�D$X   I�D$p    I�D$x    I�D$h   H��h[]A\A]A^A_�H�D$0I�u1�J�0����������    H��H�H��H��/����    L��H�H��H������    �
   �   �'�����
   A�   �   ���� �d   A�   �   �h��� ��  A�   �   �P���ff.�     ATI��� eH UH��S����H��H��tH��[]A\�@ M��t�I�|$H��t徙1H ����H��t�H�[H��H��]A\H�R@���    AUI��ATA��UH��S��H��H��P  �(t>H��`   t]H��   �4X1��R���H��tD��H��L����c��H����[]A\A]�f�H���   ��1H H�x�����1ҾK.H H���|���H��uH���   ��[]A\A]�D  H� H��t�H��D��L���H��[]A\A]���AWf��AVI��AUATI��UH���   SA�� ������H��   ��H��$�   �T$HɁ�  L�D$H���  H��`��H�D$     E�E1�H�D$H��$�   A��  A��`H�L�*D$XD$hD�L$dL�L$(H�|$hL��H�T$01�D$8D$H�	9���L$(H�D$P���  D�|$`H�D$XI�~L��1�Iǆ@      H���H)���H  �����H�I�F(  ��H���  ��  I�I�FI�FI���   ��U%�  I�F0  2 ��0A�F<   I�F@   I�FX   Iǆ  "  Aǆ�   ��  Aǆ0  ��  A��@  ����   L�l$ �t$H�L$(H��L���z���A�ǅ��Q  �E����   H�}8 ��  E��uA���   ��  ��   H�t$P�(@ H��L���`��D�|$(H�D$P    E�������1�H�D$0H�8�`��H�Ĉ   D��[]A\A]A^A_�f�H�u L�����A�ǅ�u�L�l$ H�u(L��L�����A�ǅ��{���H�U(H�T$(H�t$ H�|$0H�����A�ǋE���1���L��L���j���,���D  H��$�   1�1�L�������A�ǅ�������t_H��$�   H���   �@t�����   A���  ����   H�l$L��$�   fD  ���U(I���   �Bt��x�A���  ����   I���  H�������H�t$I��   L��H�����A�ǅ������1�I��x  ��L�����   H���n���A�ǅ��`���I���  1�1�H������A���E����     H�} L���T�������    I���  A���  �W���H��$�   H���   �E`A���  ��t�L�l$ ��A�U(�E`��x�����H�T$(�_���@ AWAVA��AUI��ATUSH��H��8  H���   ��1H �$H�hL�D$H�������H���E  I���   �   ��BH I��������`BH H��H�D$������BH H��H�D$����H����   I���  �   �xQH I���   ����1�H��H�D$ �{��A�ǉ�$�   ����   L�D$�$D��L��H��A�T$A�ǉ�$�   ����   I��  OTTO��   E����   1�H�ھdaehL��A��@  ��$�   ����  H��L��A�T$@A�ǉ�$�   ��uI�$1�H�ھ2FFCL��A��@  A�ǉ�$�   ���
  Aƅx  A�   �D$s�P@ A�   H��8  D��[]A\A]A^A_�D  A�   ��1�H���v��A�ǉ�$�   ��u��D$s E1��$I���   H��$�   ��  H��H�D$�!��D��$�   I��E��u�I�{L��I��P  H�C8H���f��H)�H�D$01����  I�    Iǃ�      ��L�\$(�H�H��)�$�   )�$�   )�$�   )�$�   �l��L�\$(H�L$0H�߾�QH H�D$8I�+L��I�[I�KE�c0I�C�j��L�\$(����$�   �v  E���  A�{(��  A�{*��  H��$�   H��L�\$(H��H�D$H�Z��L�\$(��A�C,��$�   ���  A�s*H��Ht$8L�\$(���L�\$(����$�   ��  f��I��x  H��L�\$(A�x  EE E0�x��L�\$(H��I���  A�C,L�\$@I���  H������H��$�   L�\$@����$�   H�L$(��  I���   �   �   H��H��H��$�   �����L�\$@����$�   �U  A�CL��$�   �<$ A��H  �q  A�ΉL$@�L$tE��~9���  A�C E���e  A��AUI��h  H��AS�L�|$HH��% �����$�   D�� 0  M��L�\$P��������$�   AZA[L�\$@�2  I��(  H��L��
��L�\$@����$�   �  A��I��8  1�H�މ�$�   ����L�\$@����$�   ��  A��L  ��  u	E���  I���  H�K8Ǆ$�      H�D$X    H�L$@H���0  Ǆ$�       H�t$XH�|$@L�\$P�jY����$�    L�\$P��  Ǆ$�       H�t$8H��L�\$@I��  ��	��L�\$@����$�   �/  L��$�   ��$�   1�H��L���3���L�\$@����$�   ��  ��$  =   ��  A��0  L�L$H1҉�H�|$0E1���  ��/����$�    L�\$@��  ��$  1��I���8  H��H�  9�w�A��D�d$0I��L��E�D�t$@1�A�� ���A�� @  E���>H���8  AUE���SL�D$HL��L��H��������$�   AXAY����  ��$  9�w�I��L��D�d$0D�t$@E��t	����   H�t$8H��L�\$0I��  A��L  �j��L�\$0����$�   ��   H��$�   H��������$�    L�\$0��   A��8  AǃP      ���i  <�Q  H��$�   H��L�\$0�����$�    L�\$0u?�����"  �@��A��H  A��H  I��@  H��L�\$0��
��L�\$0��$�   ��$�   ��$�   L��L�\$0������$�    L�\$0�H  H�|$(L�\$0����D��$�   D��$�   E�������A��L�\$0�D$@�   fD  L�D$�$D��L��H��A�T$A�ǉ�$�   ���v����$ �(����<$ ��  D  H��$�   H�D$(H�|$(L�\$0�d�����$�   ��$�   ���^  A��E��L�\$0�D$@�
  H�D$H�L$A��L  ��  I��X  H�D$ I��`  I��h  HcD$@I�EA�C$I�E u	H�������A�EtVI���  A��H��tFE��tAL�\$I���  D��L���P8A�ǉ�$�   �������H��L�\$tL���S8L�\$D  A���   u�<$ ��  uA���   I���  I���  I���  H���U  H��H��?H1�H)�H��   �[  I���  H��I���  I���  A��0  ���:  ��L�l$I��0  M��M���8  �    A���   taI���  A�   H��vI�T$hH��v
H9�HF�I��I�t$@L��H��辺��I�|$pL��H���޻��I���  I�|$hL���:���I�D$hM�t$XM����   L��H��?I1�I)�I��   ��   I�D$xH��I��I�|$pI�D$xL9��\  M�'A�|$` �=����Ao��  �Ao��  AL$@�Ao��  A\$pAT$PI���  I�D$h�j����    I�D$PM�t$PH��?I1�I)��e����    I�|$hL���K���I�|$@L��I�D$h�9���I�|$PL��I�D$@�'���I�|$HL��I�D$P����I�|$XL��I�D$H����I�|$pL��I�D$X����I�|$xL��I�D$p�ߴ�������f.�     <�����1�H�ھ FFCL��A��@  A�ǉ�$�   ��������D$sE1��)���D  H��$�   Ǆ$�      H�D$(�p��� M��L�l$�<$ A��L  ��  A�C I�E ����  ��  A��0  ��I�E I���  �����I���  H��I�EhI��   H��D��I�upH��  H��I�ExI��  H����  I���  fA���   H��fA���   ���@I���   ��fA���   ������)�A��x  D)�����9�I���  L�H��fA���   I���  fA���   H��fA���   ���  I�E(L��$�   H���U  A��t  L��L�\$�˿��I�u(L�\$H��tCH��t>���t7�8��  �� ��  ��-��  �� �  ��-��  ���8  H�|$L����BH L�\$��Q��L�\$I�E0�|$s����  A���   t��H�I	EA��|  1�L��I���   L�\$������L�\$H��t1�DH �   H����� ��tRH�ƿCH �   ��� ��t:I�E0H��t4�DH �   H����� ��tH�ƿCH �   ��� ��u��A��L  Hc�I�]����  �R  A�]HI�M   ���q  I�EPH��z  ��   f�z ��   H��1��%f.�     H��y  ��   H��f�y t}��9�wށ���  t
�<$ �  1�1�H��$�   L�$H�cinu  �@gH L��$�   H��$�   ��-��L�$��A��t<������I���    Ǆ$�       �L  @ A��  ����   I��   �   L��$�   f��$�   H���S  Ǆ$�   BODA1�f��$�   1�H��$�   1���gH �9-��A�������H�|$(L�$������$�   L�$����$�   ��  f�     A��������     D��$�   ���� H��$�   H��L�\$(H��H�D$H������$�   L�\$(������A�{(�����A�S*<��������~���H�D$8H��L�\$(H�4�����L�\$(����$�   �����I�{81�1�H��L�\$(�_���L�\$(����$�   �����A�CL��v
I9C`��  I��x  1�1�H��H��L�\$(����L�\$(����$�   �i���1ɺ   H��L�\$@H��$�   H��H�D$(�����L�\$@����$�   �>���I���   �   H��H��H��$�   1�����L�\$@����$�   �	���H�|$(I��`  I��X  I��P  轶��L�\$@����$�   �����A�CLA;��  �t���Ǆ$�      �����     ����  �  A�]H����������� I���  I���  H��?H1�H)����� I���  H��L�\$�\���L�\$H��I���  I���  �A���L�\$H��I���  I���  �&���L�\$H��I���  I���  ����L�\$H��I���  I���  ����L�\$H��I���  I���  �խ��L�\$H��I���  I���  躭��L�\$�����A�C I�E �����I�M   ���  �����H����  Ǆ$�   CBDA�   f��$�   ����A��L  �%���L��L�\$����L�\$H�������L��$�   H�|$H��L�\$L���&L��L�\$I�E(������PH��������PH��H��������t$@L��L�\$����L�\$H��I��I�E(��   L��H���1����׃��m���A�x+�b����   �$M�HD)�L��L��A���fD  ��tH�����A<�v��t4E1���E��t*�W�Lʃ�t�AH���A�H9�u�����~A�x+t�I�}( �����A���  L��L�\$貸��L�\$H���*���H�|$L��H���K��L�\$I�E(����H�������Ǆ$�   EBDA�   f��$�   ����A;]H�����I�EPH��I���   ����H�|$H��L��L�\$�J��I�](I��H���� L��I���� L�\$A9�Hc���   ��~B�P�A�N�Hc�Hc��A8<uw��Ic�L�H��H�1�H���D�D�H��D:D�uQH9�u�D��)��ȃ�t@Hc���r�@��?w+H�(     �H��s��H��H�Hcȅ�~��� ��?v�D M�e0����H��H��r����������D$t    �����$��������$�   H��$�   H�D$(����H�|$(L�\$0Ǆ$�      ����D��$�   L�\$0E��D��$�   ���������Aǃ0      I��(   ��   Ǆ$�      ����H�t$@I���  �٤����$�   L�\$P����$�   �n�������H�L$8H��L�\$PH�4�����L�\$P����$�   ��  �   H��L�\$P�����L�\$P����$�   ��  H��L��$�   �9���L��H��H�D$h������$�    L�\$P��  f����
  Ǆ$�      �>���A��L  1�1�L�\$0H��$�   I��@  A�C$����L�\$0����$�   �����E���;  E�c$E���.  A��L  I��  H�L$PH�K8�D$XI��  H�L$0Ǆ$�       H����  I��  ����  ����  A���   ��  D��H�|$0E1�1�L��$�   H��   L�\$@���L�\$@��$�    I��   ��  H� XH ���  @����  ��t�� �@����  �|$X��  t)�<$ t#H�T$0H�|$PD��L�\$@�ޫ��L�\$@��$�   ��$�    �  Ǆ$�       A��L  ��  t"�t$tL��L�\$0蛾��L�\$0I��8  �*���1�I��    I��   E�c$Ǆ$�       �=  fAǄ    fAǄ    H��H=   u�H����  I��  �E  I��  H��� � TH H���H)�I��  H��� H)�   ��I��  ���H�H�S8H�|$PD��L�\$0Aǃ      �˪��L�\$0����$�   ��   �   �5A;�0  w<I��(  �Qf��t,fA��C
  A��  H��H=  tzA��C
  H�ʅ�u�fAǄC
    fAǄC
    �̋=� ����XH �T(��5�������XH f�T(��"���Ǆ$�      ��$�   ��$�   ����M��L�l$0��$�   ��$�   ���?�������H��� I��  � RH H���H)�I��  H��� ��   H)�I��  ���H�����H�t$8H��L�\$0H�I��   ����L�\$0����$�   �W���L��$�   H��L��� ���L�\$0��A���   ��$�    �'���L��H���������$�    L�\$0�	���A���   �����  �������Aǃ      �D$8   �D$@    L�l$0M��;l$@��   L��H��������$�    �ЉT$H��   L��H���q�����$�    ��ur��A;�  �T$HvA��  �t$8H��H��<�:A9�v+���   w#��M��   H�L�f��  E�0fD��  ����H��9�rD$@�|$8�L���M��L�l$0�	���M��L�l$0A��     vAǃ     A���   ������L��H��L�\$0������$�    L�\$0���D$@������D$8    L�l$0M�݋L$89L$@�����L��H���d�����$�    ���a���L��H���������$�    �H���H�1�I�T- f��  �I��   H�qf;O��   H��A9�w��   �U��H��L�\$0A��  �;���L�\$0����$�   �����H�s@1��   �2H�HA9�v#�I��   H�L�f��  �<Of��  ��H��9�s�H��L�\$0�W���L�\$0����f��  �D$8�����A���   ��  D��H�|$0E1�1�L��$�   H��   L�\$@�(��L�\$@��$�    I��   ��  H���y  @���V  ���;������ �@���(��������VH f�T(�����H�L$8H��L�\$@H�4I��  ����L�\$@����$�   �;  L��$�   H��L������L�\$@��A��  ��$�    �  H�|$0E1�1�D��M���   �O��L�\$@��$�    I��   ��   f�   A��  ����  ���y  D�t$H�   L�l$@A��L��E9���  L��H��������$�    A��uw��  L��H��tV�������$�    ��uV�ƺ��  A��H)�H9�~D������H��   1�D��A�<A����f�<VE9�v�9�v��z���������$�    ��t�L�l$@D�t$HI��L�|$0I��   L�\$@L���%?��L�\$@L��I��(  L�\$0Iǃ       �?��L�\$0Aǃ      ��$�   Iǃ(      Iǃ      Iǃ       ��$�   ��������l���H�� H�xH���H���H��XH H�L�H)�H��H)�����H������Ǆ$�      �1���A��Ww�D��H�|$0E1�1�L��$�   H��   L�\$@�b��L�\$@��$�    I��   �����H� VH H�ǉ������I��L�l$@D�t$H�m���A��$���H��L�\$@��k���L�\$@����$�   �����D�t$@1�M��I��L���L��L�|- L�   ����fA�H��A9�w�H�\$HL��M��D�t$@H������L�\$H������|� �����VH �T(������H�b� H�x��VH H���H���H���VH H�L�H)�H��H)�����H�����I��D�t$@L��D�d$0����L��H��L�\$P������$�    L�\$PH�D$x��  L��H������L�\$P��A���  ��$�    �r  H�|$@E1�1���M���   ������$�    L�\$PH�D$X����L�l$P1�I��D�t$`E��M���*H�L$X��L��L��H���������$�    H��  ��A;�$�  r̋D$hH�t$xL��L��$�   H��E��L�l$PD�t$`H�H��$�   ����L��$�   ����$�   �����L��H��L�\$P����L�\$P��$�    fA���  �W���L��H���z���L�\$P��A���  ��$�    �/���H�|$@E1�1���M���   ���L�\$P��$�    I���  ������D$x    D�d$PL�l$`D�t$hM�ދD$xA;��  �R  �D$xH�|$@E1�M��I���  A���  �   L�,�1��@����$�    I�E ��   E1��   L��Ik�H��Im ������$�    f��$�   ��   L��H��������$�    f��$�   ��   L��H��I���]�����$�    ��   H��$�   H��H��H��H�EH�U H��$�   H��H�UA���  D9��Z����D$x�����H�D$X    �����M��L��E��L�l$PD�t$`����Ǆ$�      ����A��H  �����M��D�d$PL�l$`D�t$h�~���M��H�|$@E1�1�A���  M���   D�d$PL�l$`D�t$hL�\$P����L�\$P��$�    I���  �.����D$`    D�d$PM�܋D$`A;�$�  ��   I��$�  �l$`H��H��$�   H�D$hH�D$XH4��������$�   ����   �   H���$�����$�   ����   L��H��H��Hl$h������ЉU ��$�    ��   H�|$@E1�1���M���   �����$�    H�Eu|1�D�t$hM��M��I�܉�;] sML��L���s���H�M��������$�    u����M��D�d$P����M��L��M��D�d$PD�t$h����L��D$`M��M��D�t$h�����M��D�d$P�����f.�     �Hc��   ��x=;�8  }5H��SH��1�H��H��H�@  H���RPH���   H���   1�[�@ 1��D  H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ H��  H��t1Ҁ8/��H���     �o�8  �o�H  N�o�X  V H��h  H�F01��ff.�     @ ��P  f�1�� H��t
H��   H�H��t
H��(  H�H��t��0  �1��f�H��t�1��D  H��t�21��fD  USH��H�GH��`  H��t.H���   H���`BH H�x�r���H��tH���UH��(  H�B@H��1�[]� AWAVAUATUH��SH��
  L��t$I���   M��p  �D$<    H�$I��   H�D$I���   L�phM����  I�I�~H��$  ��D$<���m  A��(  H��$  @���  �V�1���H�L�     H���P�H��H	�H9�u싔$  E1�H�D$    ����  I�I�~H��$  �P�T$<����  H��H��I�X  �H�@Hǅ�
      Hǅ�
      H���
  H��H�����
  �    H��I�@  �S�o�  �o�  �o�(  ����
  I���
  ��
  ���
  Hc�H;L$�  ��x'�D$ H�D$��  L��H�L$(H�t$�P H�L$(�D$ D���   I�t H�t$ E���  �T$H��E1�)�H�D$H�@�P�D$<M����   ����   I�H�x ��   H�}@�����H�}PHǄ$      H��H��$  蠔��H�}XH��H��$   苔��I�~1ҋt$H��H��$  H��$(  I��P�D$<H��$  H��H�E@H��$   H��H�EPH��$(  H��H�EX���D$<	   E1�H�<$L���3��H�ED��1  �D$<H��
  []A\A]A^A_��     E1��� H�D$H�L$(�   H��H��$  �P0L��L�|$H�D$@H��H��A�W8H�D$@H�\$H�L$(H��$0	  I�GH��$  H)�H�t$ H���P�D$<<������H�EH��H�t$ H��$  A�   ƀ0   H�D$H�@�P�D$<�X����1�����f�     )�H�<$Hc�H�T$<H��H�D$�u����L$<I�Ņ�����H�T$Ic�(  H��H�$  �� �����D  �D$A��,  L��L�D$A�(  I��   ��I�H  H�����L�D$���D$<��  �4L��L�D$�����D$<���k  L�D$Ic�(  I�P@@���]  �F�1���H�Df.�     H���J�H��H	�H9�u�A��,  ����   �z�1�@��H��L�8@ H���P�H��H	�L9�u�H�E1�H�48f.�     H���P�I��I	�H9�u�L��H�L$ L�D$�J���Ic�8  H9���   L�D$M9`��   H�L$ I9���   I)�L�D$(H�L$ tyH�<$L��H�T$<L�d$E1������I�ŋD$<���A���H�L$ I��H  L��L�D$(H�H�L$L�������D$<���S�������L������Ic�8  H9�w�D$<	   E1�E1������H��1������AWA�   AVAUATUSH��(  L�gA;T$ �h  H��I��A�։����n  ������I�M H��E1�E1�I��$   H��8  I�M(��0  ����H�t$�D$����1  ��L�~L����H��@  H��ǃ�       ��ǃ�   ltuohp�B PRL��H��$�   A�H�� A�ǅ���  ��D��H�|$`%   �D$��$�   �?���A�ǅ��  ��0  H�$H�|$`�o�$  L��$@  �o�$(  �D$��1  )D$ )L$0�D$H��$8  H�D$H�A�P���   �������   �D$���G  H��$�   肏��H��$�   H��H�CP�m���H��H�CpH��(  �@ I��$�  I+�$x  ǃ�   ltuoH��fA�}H�ChH�Cxw
���      H�|$    L���   uH�|$8   �a  H�t$ L�������HcCPHcT$ H��H�H�� �  HcShH��H�H�CPHcD$8H��H�H�� �  H��H�H�ChL�l$L��L	�tL��L��L���G���LkPLsh�D$u�|$ ��   �|$ Hc�@  Hc�8  ��  H��$�   �Pf��~_D�B�H�@I��I��I�HcH��H��I��I��?J��
 �  H��Hc�H�P�HcP�H��I��I��?J��
 �  H��Hc�H�P�L9�u�HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$@L���5���H�T$@H�D$PH)�H�S@H�C0H�D$XH��H+t$H��H�CHH�s8��   H��(  D��[]A\A]A^A_�D  ��1�1�����@ H��$�   H��(  �4���H��$�   H��H�C@����foT$ fo\$0H��H�CPH�D$U] H�E0L�u8�E�{���D  H�$H�|$`H�@�P�a��� H��$�    ������X���@ H�shH�{0�+����4���fD  H�D$(HD$0���������ff.�     H����  AUATUSH��H��H��X  L���   H��tw��8  ��~ZE1�f.�     L��H��H�H�EH��t-H�0L���+��H�uL��H�    �+��H�E    H��X  I��D9�8  �L���k+��HǃX      H��8  L���Q+��H��@  L��Hǃ8      �7+��H��H  L��Hǃ@      �+��H��P  L��HǃH      �+��H��X  L��HǃP      ��*��H��@  L��HǃX      ��*��H��  L��Hǃ@      ǃ8      �*��H��   L��Hǃ      �*��H��(  L��Hǃ       �w*��H�C(    H��h  L��Hǃ(      H�C0    �M*��H��p  L��Hǃh      �3*��Hǃp      H��[]A\A]�D  ��    AU1�ATUSH��8Hc��   ����   ;�8  ��   H��L��@  H��H���   �   H���Ph�¸   ��~~H�L$H��H��?I��I1�I)�H��tdI��   ujH�D$(H��H�4$H��H��H��L�H��  H�t$H��   H�L$ H��  H�t$H��H��0  1�H��  H��(  H��8[]A\A]�@ L���  �Ê��H�<$L��f���   谊��H�|$L��H�$蟊��H�|$L��H�D$荊��H�|$ L��H�D$�{���H�|$(L��H�D$ �i���H�L$H��?H��  ��H��   ����ff.�     f�AUATI��USH��H���   H��L���   �D$    �VHH�ø   H��x2H���(\���(I�UH��H��H��D$H��H9�HB�I��$@   tH��[]A\A]�D  H��L�L$E1�1ҾP  H���.���H��I��$@  �D$��u�A��$8  ��~��s�H�QH�<�H�4�H��H��1T  @ �   H��P  H9�u��ff.�     ���iH 馕��fD  SH���   �`BH H��`  H�x胵��H��tH��tH�H��t	H��[�� 1�[�@ SH��H�?�4���H�;����H��tH�{PH�S(E1�1�H�s H�?�P1�[�ff.�     �SH��H��H�?�p���I��1�M��t9H�H�JH���   H��H�4�H��H�@  H�T$A���uH�SPH�L$H�
H��[��    H�GPH�8 t.SH��H�?�
���H��t
H�SPH�:�PH�CPH�     [�fD  ��    AWAVAUI��ATUSH��H��8  H��    H�   �T$8�h  I��`   ��  1�H�������A����tH��8  D��[]A\A]A^A_�@ L�t$P1��   I��   L��I���   I���   HǄ$      �H�L��H��H�t$1�H�B1��H��H��$�   � ����   H��H�D$�.�������  H�u@��hH �   �H���� ���&  �����D$L   H��$�    tH��$�   I���   ����L����$�   D�D$LE�������D$8������f���  I��0  A�EH    I�E    I�E I�EH��H��  A��h   I�Ut
H  I�EI��P  I�E0�BH I�U(H����  I��H  H��t<����t4�
8���  < ��  <-��  �� t	��-�3  H����u� I��`   I�E    tI�E   I��X  H��tB�DH �   H����� ����  H�ƿCH �   ��� ����  f�     I��p  I��x  A�E8    I�E@    H��H��I�EhI���  I�upH��  H��I�ExI���  H����  A���   H��I���   f���c  �@�������������������D��fA���   )�D)�fA���   9�A��j  N�A���   fA���   �/����[���L�l$ H��A�	  L��$   ����H�$    L��I��L�}H���f���L��H��I)�I9�LG�L�����������  O�L<�H��$   C�< I9��;  D��$   �D�@A��s��  H��I9��  A��Su޿�gH �	   H����� ��u�H��$   H)�I�D
H�$L�<$H�t$H��L��H)��
������  I���   H��H��� �������  L��$�   H��$�   L��L��$�   L�L�D$XL�D$PL�D$H�\$`Ǆ$  ������$�   L����$�   L��H�\$P��$�   L����$�   L�d$`L�|$PL�D$M�l$�M9��L  �D$h���h  I��	�Df�A�s�e  L����$�   L����$�   H�T$PL9��  �D$hI��L�����!  I��A�?Su�M9�w���gH �	   L����� ��u��hH �   L��L�l$ ��� ���  �D$L    L��$�   H��$�   �D$h    L�H�C�H�\$`H�$f.�     L�d$PL����$�   H�l$PH9���  H�$H��I9�r�eD  I��I9�sGA�<$%u�hH �   L����� ��u�E��8  E��~�I����$  I9�r�f.�     H9���  �    E��8  E���   �D$hD�T$8�D$LE��������������H�|$H�T$L�P   ����D�L$LI��p  E�������H��$   I���   H��$�   H���I  H�BH)�H9�vH��$   H��H�|$H�T$L����D�D$LH��I��h  E���B���I���   H��$�   L��$   H���,������t  I�L9���  A�   H��$   L�,$H��E���AfD  �N�1�E���*  ��H��M �   D)�A��@���K  H��H��L9��;  H9��  �
�΃�0��	v��N����K  �N�����  �N�1���     �hH �   H����� ������H��$   H)�I�DH�$�)���f.�     L<$I����  J��<  �	   H��$   I��   �� �   H�$	   L��$)  �5����    I�M�6���fD  �hH �   L����� ������L�l$ �   f.�     �D$L�����    �FH��H���?����    �FH���+��� H���   ��BH H�x�C���H����  I��`   I��   �s���D  I���   �`BH H�x����I��`  �M����    I���   H�������H�4$H�������������D  L�l$ �D$L�����f���  ��  fA���   ��  ����@ I��  H�������I�E(�����    A�   �����D  H�E�I9��,��� L����$�   L�d$PL9��h����D$h���t  �} /�����H�EH9������H�EL��H)B��T$����������u�R�A��jH ��gH H�|$H�z�C   L�d$0A��H�\$ L��I��L�l$(I���@ H��0L�+M����   A�E A8�u�L���d� H9D$u׃|$t-�EA8EuƸ   ��    �TH��A:T�u�L9�u�I��L�l$(H�\$ A�W����  A�O����  �@  ����  I��p  ���6  ��	E1�1�H��$   ��L��L��H��$   �K  ��$�   �D$h���[���L�d$P�q����L�d$0H�\$ L�l$(�\���@ A��8  ���)���f�     �D$L   ���� M H�}�����@ H���X���H�SI��H)���  H��   �   H��$   H��HG���������  H������H��$   L)�H��H�����f�1��V���f�     �o �oJH�oR P �oZ0X0�ob@`@I��H  E��(  E���.���E��,  E������A������A���
���M��p  E��8  I�I+�H  E����  I��@  Hc�H  ���������8  u��������������H��@  H9������E�A�H���  K��M��I��I��`D  ��t��H��H)�1�H��H9��n���L9��n  Hcq���Y����u���M������D���H��P  H������H9��-�����y��$���@ �������I�u0������    A�   ����D  @�� v'@��>��   L�,$��   �����L�l$ �   �����H�6     H��s�H������L�,$I��h  I��p  �D$L    H��$   ����IǅH      �=���1��
   H��葽 H���c���H��$   �D$L    �\���I��  �������Hc�$  ����  A;�8  �y  Hi�P  I�@  �����   1��������$�   ����I��   H9������H)�C�1�H��Hc�H��I9�0  �����I���   Ic�E1�1�I��   L��$   �   H�<$H�D$0�������$    H�D$I��X  ��  H�D$    1��D$    I�܋D$A9�8  ��  Li\$P  I��@  Lۋ�8  ���=  �C�L$�D$<�E�D$ 9�vL�E���9���  �T$H�<$M����L��$   �   �D$(�N�����$    I���K  D�T$(D�T$H��@  L��I�H  ������$   ���  �t$ ��H  L���[�����$   ����  D��H  I�G@1�A�y�@��H����M��E����  L�81�D  H���H�H��H	�I9�u��I�L��9�s�L���o���I�4$I;t$��  �U�I�D$I�L��H�H��H;�j  H9�u��I��I�GI+�H  H9��K  H)�L$ H�<$E1�H�T$(L��$   1Ҿ   ������$    H��H�D$H�X�  H��$   H�t$(H�<$H��������$    H���  I�4$L��I�H  �4�����$   ����  H�\$H�T$(L��H�CH�0�L�����$   ����  H�K1�I�T�I+�H�H�T�H���P9�v�|$< �+  H�D$�(H�D$H�D$����L��L��A�W�D$h����I��P  �S���I��8  �G���L�,$�����I��1��e����D$h�   ��   ����Ǆ$      L��I��X   ��   A��8   ��   I��X  E1�L��H��H�D.H��tH�0H�<$���I��X  H�D.H�     H�t.H�<$I���a��I��X  H�D.    E9�8  �H�<$�?��IǅX      H�<$H���(����$   �D$L����1���1��	H�D$H�HH�D$0I�t���  I+4�H�<�H���P 9�w�����I��X  �L���L������I��X   L��Ǆ$   �   �����u���f�     H���H  H��X  �WH�G ��v+�p90s-�J�H��H��H��D  �H��;sH9�u�1��fD  �   �f.�     H�G     �G    ËWE1�A9�sF��L�O D)���B�H��H��A;4t-v#�/D  ��D)���B� H��H��A94tr��A9�r�1�Éȃ�Éȉ�f�D�@����     �D�_D�HD��1�9�sFA��L�W A)�A��A� I��H��E;tHv!�U D��)���H��H��E9
t1r?A��D9�r�E1�D9�s?��t=��H��HW D�
D��D��@ ��u"A���D��A�ȍBD���t���D  1�D�ÍB��D  H�    �   ��t$��H��t9�H  vH��H�X  HcFH�1��ff.�     AVAUATI��USH��H�    H�A    ��t.����H  ����   9�����9�vh�1�H��[]A\A]A^Ð��uD1�1�H��X  H��h  �,0���	�H��t�f�     9kw9ksNH�H��u��@ ��H  ��1�9�w���H��H����u��f�     1�9��x���H��1��fD  L���   H�sL���u������O����s�sL���M������7����SD�[	�   �D�CI�}@��E��A����A�����D����)�tPA��H��
D�rE����   L�R��9�tis*1�E��@��J�|�f.�     �
L�R�9�tAHB�A9�s ���H��
D�rE��u���L�RD	�����OE��tW�L�W�9�u%A�
E��t����A�J	����S
�Hc�I�$L��D$������D$�;�����L�R��D	��H�����L�W	��ff.�     f�AU1�ATUSH��H�zh �D$    tH��[]A\A]�f.�     L�G�   I9�w��A����A��E��A�C�L- I�L9�r�H��H��D��E1�H�} L�L$1Ҿ   �@���H�ǋD$��u�E��H�}hJ��H�UXE���w���A�E�1��@ H���LS���LS��	��ɉ�H�JH9�u݋D$�?���@ AWAVL�wAUATUSH��(H��D$    L9��  I��D�oI���o���   L��M��$�   F�*E;�$�   �   A��1���A��A����������@�����A��A�������@�������@�����A��L�I9���  E���l  ��A�M�H��H�L�I��L���   @ A�M�F��A�N��	��ɉHA��HE����   A�HE�pI�XE�@��A��D	�D	��H@����   �D�sL�C�[��A��D	�	ىH@����   A�H��(I�X��A��A�HD	��ɉH�L9���   �L�sE��tD�C��L�sD	��ɉ@���0���A�M�F�HA��HE���?���A�HI�X��A��A�HD	��ɉH@���E����L�C��A���KD	��ɉH@���J���A�H��(I�X�H�L9��[���D�D$A��$�   H��([]A\A]A^A_�fD  �   H��([]A\A]A^A_�@ A��L�L$�(   H��A���D��D�T$�f���I��I��$�   �D$��u�D�T$A��$�   E��$�   ����f�     USH��H��H��X  H��8  H�(H������H��P  H��Hǃ8      Hǃ@      ǃ4      ���ƃ`   HǃH      HǃP      HǃX      H��[]�H��H��(  H��f��H�:�P  Hǀ`      H��X  �0  �@  �v��1�H����     AUATI���    UH��SH��H��L�*H�T$�D$    L�������H�ƋD$���  H�KI9��  D�D�N�S���S��	�H��f�V
�S�V	D�EH+��   L�A��H�~A����   �F   A�   ��tA��D�VA�щ�A��H�I9���   E����   ���{D�KA��H�E����   �K��D	�����A���KD	���	ω~�
�����J	��z�R����	���	ʉVH���   H�    H�2H���   �V��   H��[]A\A]�fD  L����	��H���   []A\A]��     �F   A�   ����fD  L���	���D$�f.�     ��D	ω~�
�R��	ʉV�`��� AT1�USH��H�zp �D$    tH��[]A\�fD  H��H��H�T$I��H)�H�;�u����H��H�Cp�D$��uƉ�L��H���;� H�Cp�( �D$H��[]A\�ff.�     AUI��ATI��UH��S��H��H�1�D$    H��tH������I�$    ����   �S��|  ��   �E �� <_wj�   � �| H���W���_wO9�w�sH�T$L���K���H���D$��u6H��H��H���}� H��� �D$I�$H��[]A\A]��     �D$1�I�$H��[]A\A]� ��t���h���ff.�     f���vH ��u��fD  AVAUI��ATM��USH��H���   H��t���  �H��t���  �H��tQ�}���  ��Hc��Di���}���  I����Hc��,i��M��tM�u M��tI�$[1�]A\A]A^��    �   A�   ��ff.�     �> ��   D�_bH�G`S1�E��A�K�f��~L�GxH��A�TP�9�~\L�OhLc�Hc�H��I��M�I�I�I9tH�WxD�@fD�G`f�B[� �fD  I�YI9Xu�A��A�K�fD�Wbf�     9�~�� [��    �ff.�     @ UH��SH��H���������  ���  9�tH�} H��u6H�}H��uH��1�[]�@ ���  ���  �g��H�EH��1�[]�f���f��H�}H�E H��t���ff.�     ��   @��tfUH��SH��H��H�Wb�OH�ЍT;Ww-foE H��H��HShH�Sp�1�f�CbH��[]�@ 1Ҿ   �������u�H�Cb뼐�ff.�     @ AWI��AVI��H�4
AUL��M��ATUSH��   H�T$����A�ą�tH�Ĉ   D��[]A\A]A^A_�f�     L��L���ŷ��A�ą�u�I�F@M�W(J�,(I�:H�XM��t	�8 ��   �D$<    H9���   D�(E����   A����   H�XH9���   �@A�����D$A��E�A�WM�GD9���	  D��I��I�GE���0  A�z�1�1�1��7�L�KL9�rw����KL����	���Hc���I��H�BH9���  H����uH�CH9�r<�3H��@��u�H�CH9�r'D�H��D�� A�w�D$@    �t$H9�sS A�   L����������D  A����  A���d  E1�H�CH9�r���\$E�H������D  ���y��փ�?��@@�t$D��t^H�XH9�r��P��tMH�XH9��x����@H�H9�s(�g����    H�CH9��S����H�H9��D�����u��    �D$A�WD�9���  D�hL�T$(A���D�\$ A��@�	���M�G D��L�L$@�    �3����T$@I�G ���)	  D�\$ L�T$(E�o�|$I��H�|$ I���|$ J�(�I	  H�CH9������E�C�I��I��I��   D  L�HL9�������8L���������>  ���U  L�HL9��X����0L�ȉz�r��@�C  H�pH9��6����8�@��	����B���|  H�^H9�����������F	����BH�� A�GL9��  H�CH9�������3H�   ��@��t*H�CH9�������{��A���{D	�����Hc�H�:H�B   �� t)H�xH9������D��@A��D	Ș��H�H�BH���σ�@����  @�������1������f.�     H�XH9��3���D�XA���S���E���D$    �b���@ 1�����f�     H�pH9������� �B������\$@L��L�T$�����L�T$���t  A�G+D$�n���H�|$ ��A�jL��M�O D�d$H�DA��H��H�D$M�H�T$L��L��A�IE�AA����������  M�O �KM��H�C I��K�)A��)�H�2L�H��   uH�z   ��  ��~n��D�ZLcBHc�H���zH��H��HcH��H��H��H��?H��* �  H��D�Hc�H�P�HcP�I��H��H��?H��* �  H���Hc�H�P�H9�u�I�� L9l$�P  E�������     H�^H9��������N����	��N	ȉB�{���fD  I�G�D$    E1�I�GA��thH�SA�   H9��J��������  H�SH9��2����[H�H9�s$�!��� H�SH9������H�H9��������u��D$<    H�D$H    H�؋\$E��H�D$@    foT$@A�G0 )T$pL�`L9������D� D��A������A���N  D���$�`tH ��   H�T$P1��vf�H�D$pH�B�����������   ����  ����  H�D$xH�B��ȅ���   ����   I�D$H9��+���foJ�A�4$�   I��)L$pH��H����������  ����  ���m���M�L$L9������I�$HD$pM��H�B����������W���M�L$L9������A�$��A��A�D$M��D	�H��H�B��ȅ��D���fD  foB�����)D$p9��T���I�O(A���  B�$ŠtH �   �+  ����9��;���H�T$p��H�T$@I�WH��H�D$Hfod$@)d$p�D9�����I�W��H��H�D$@H�D$xH�D$Hfo\$@)\$p�y����   ��  �G���A�w0H�T$@H��������D$<��uL�������H��I�w0�t���I�(�{i��D�d$<����H��I�w0H�L$�P���H�L$A�G0�Q�Ab�D;A��  �Q�A`�D;A�s  I�(A�w0H�T$@�9����D$<�t���M�L$L9��"���A�$��A��A�D$M��D	�H��H�B�����fD  M�L$L9������E�$L��E9������M�WM��I��H�B��N���D  M�L$L9������E�$L��A9������M�WM��I��H�B��A���D  M�L$L9��z���I�$HD$xM��H�B�����@ L�HL9��S����8��A���xL��D	��������     L�HL9��#����0��A���pL��D	��������     A�BL�L$<�   D�\$ ���D�T$���D$����D�d$<I��I�GE��������D$D�T$A�G�D$ I��I��I�G����@ �������HcrHcz�Q�H��H��H�f�H0HxH��H9�u����� A������D�d$����I�G �x����   ����A�0 ��   H�Qb�qH�ЍT;Qwqfol$@H��HApH��HQh*fot$Prfo|$`z �  f��@�D$<    f�Ab�!����   �   H���������s�������A������1Ҿ   H��H�L$�������u$H�L$H�Ab�h����D$<   �����H�������D$<�����L��L�T$耭��L�T$����A��� ���ff.�      AWAVAUATUS��H��XL�o�����M���e  A9�H  �X  H��I��A����	�^  A�� @  �9  H��I�X  ǅ�   ltuoǅ�       A��0  D�CI���   H��X  D�cH�T$L�D$H�4$�c��L�D$H�T$L��ǅH      H�4$H��0  �����A�ą���  H��X  A���o@��   �oH(��   H�@8H���   ��������   M��tfA�w  ���   A���  A���  H�EP    H�Eh    HcC9�tH����X��A���  �@  H�EhL�EPI��L�EpL�UxH�EX    H�E`    E����   ���   H���   Icw(Ic f��~]�J�H��H��H� HcH��H��I��I��?J��
 �  H��Hc�H�P�HcP�H��I��I��?J��
 �  H��Hc�H�P�H9�u�Mc�Mc�I��I��H��H��?H�� �  H��H�H�EPH��H��?H�� �  H��H�H�EhH���   H�t$0����H�L$0H�D$@H�T$8H)�H�M@H�E0H�D$HH�UHH)�H�E8��    A�   H��XD��[]A\A]A^A_�A��   M��(  ����������NH�D�I����     I��(I9��e���A9$u�A�GA9D$u�A�D$I���   A�t$��H�<$���������������I��X  ���I�x  �T$H�D$账����������T$H�<$��A�t$臨���������A�|$��E1�H�$H��HD$A�t$A��D�L�Y@H�D$A�����|$A����A������A�������A���@��@��   ��@�πH�AHA�Љ|$A�|$I�<H9�rVL��H������D��I9�sNL�d$(I��L�l$ ��L�H��H9���   �E��tD�j��D	���H9��L�l$ L�d$(�D$$�D$�D$��@�D$A�D$1��D$�ty9�r�s ��9�vj�7D������L��L�aE��tL�a�I��	���A9�r�vV�z�@ H�EPL�UhI��������LkD$��H��H��L9��  fD  H�<$臨���d���L�l$ L�d$(�Q���A�T$A�$�D$�z  ��I��	���H�D$A�$A�T$�D$�@  ����E�d$	�A	�H�<$����H�|$ �����H�D$A���  A���  Hc@H��9�t��H���T��H�t$A���  HcvA�H�EpH���T��A��0  H�D$L�L�$$L���;����������H�t$L��L�$$����A�ą��i���H�4$H�F@H�NHH�PH9������D�D�҃�����  ���V  ���,  L�HL9�������@A������A��H��M��H�D$D��@����@����  @����  1�1�@���[  D��@����@����  @���~  @���P  A��A������E����  A������L�D$�։�H��I��H��I��Mi��   L9���������   ��L�D$H����H��H�u0H��H��ƅ�   ��H�U8L��H��H�����   D�H�U@L��E��H�����   H�UHH�T$ǅ�   stibH��H�uXH�� H�E`    H���H�UPI�W@D���   H�Uh���   A��  @ �0  Hc�H��D�D$H��L�L$H��D�T$�I���D�T$L�L$��A��D�D$�������   ����  ���   ����  ��H���   ���   ��A��D  u������Hc�H�H�$H�SHA���7  E����  A����  I��A��E1�A��   �   �   Hc��'D�0I�D E1�A��I��A��   A��1�E��@�Ń����0  ���  ��tE	�A��t�A��u�D�0A��   H��E1�뼉։�H��H��H��H��H;|$��������I�qH9������A�I�����������I�yH9������A�A�AA�q��	�A�AI������	����I���I�qH9������A�A�AI���+���L�HL9������L�XH�@H�D$�����L�HL9��_���D�X�P�p��A��A	��P��A	��P�@��	�	�H�D$����L�HL9������PD�X��A	��P�@M����	�H��H�D$�\���I�qH9������A�	I����Hc�H�|$����I�qH9������A�9A�I����	�A�yI��	���H�|$�X���I�qH9������A�	A�yI����	�H��H�|$�,���A��A��A	�E������I��H�D$����I��E�A���E�������L9�w������A���   tD�0H�<$衢�������L)�I��A��A��   ��Hc�9�G�1�E1������I�1�A��I��A��   ����t8����9�uE�)I��A�ŀtD	�E�A��t�A��uшA��   H��1���A���   �l�����e���I��E1���E1�E1�A��   �   Hc�A�   �&D�8I�D E1���I��A��   A��1�E��@�Ń���tc��uOE��u��t�A��u�D�8A��   H��E1���E	�A�   ��L9�v�E�I��E��A��E��E1�A��E��u�E��u�E��A�   ��A���   �����D�8����f�     H����  AUATUSH��H��H���   H���   H��  L�hH�G(    H�G0    H�������H��  H��Hǃ      �����H��  H��Hǃ      �����H��   H��Hǃ      ����H��(  H��Hǃ       ǃ�      Hǃ�      ǃ�      �r���H��X  H��Hǃ       Hǃ(      �M���H��8  H��HǃX      ǃH      HǃP      ����H��h  Hǃ8      ǃ0      H��tD  L�&H�������L��M��u�Hǃh      H�s@L��Hǃp      ǃ`      ����H�C@    H��[]A\A]�fD  �ff.�     @ AWAVAUATA��UH��SH��1�H��X������tH��X[]A\A]A^A_��    H���   �@uH H��质����uҋ�@  �D$<    ���  �   ���   0RFPu����   w���  9v���   
  u�D��  H��L���x����D$@���n���H�t$@H�������ЋD$@���R����ʁ�23  �  H�}�t�I��M)�L9���  k���_H9���  �D$<    H�E���	���E���   I9��������  H��D��@  ������D$@�������H�t$@H�������ЋD$@��������   A9������Ak�H�������D$@�������H�t$@H��襟��D���D$@���w���H�t$@H���أ��H�ƋD$@���[���A�ĉ�h  H�����d  �?����D$@���5���L��H�������D$@������H�U@J�4"L�JL9���  ��J����	��J	ȉ�l  �B�J����	��J	ȉ�p  �B�J����	��J	ȉ�t  �B	�J
����	��J	�1ɉ�x  �zL��A��A��t������Ƀ�@��u��A��A��t@�� A������Dك�L�H9��+  E��tI�JH�B@��tH�B�R��	��ɉ��  @��u��HH������	��H�	ʉ��  E��t#�@�� ��   �H��H��	��҉��  @��@t@H�HH9���   �H���H�HH9���   � H�H9��~   ����u��D$@    H�PH9�rf��H��	��ɉ��  �P�x����	��x	����  E��t8H�PH9�r'�@������  � �   �(���H���E����D$@   H���}����D$@�D$<�������H�M8���  H��H��h  H��p  D���  H���  H�Ɖ��  Hǃh      H�$H�D$貗���D$@�������L��H��苙���D$@�������H�E@N� L�hH���  M9���  ����P��	��҉��  �P���P��	��҉��  �P���P��	��҉��  �P���P��	�H��H���  �P���P	��	�H��H���  �P
���P��	�H��H���  �P���P��	�H��H���  �P�шT$&�����  �L$'u!L�hM9��  �P�@��	И���  �|$& ��  I�EI9���   A�U A�ME�E����	�D	���  A��N�4(M9���   H��  H�l$L��I��H�L$(L�T$�f����  H��L)���  H�xI9���  �D�`��A	�A��fA����  E��I9���  �HJ� �����H	�f���  f��u�H�L$(�r�H�$�#����D$@��t������D$@   H�������H���.���Hǃ�      H��x  �D$@�D$<���^�����H  L�{H�KH��H��H�C ��t0H��X  D�BE��u5H��1��fD  H���z���u��9�u    ��  H�C    ���  ��uH�KH�C��   ��`  H��H��H�� ��HE�H��H����HE�H�C��tH�K@H��  H�C(H����  H��  �����H���  �C8    L���  �o��  H�C@    H�C0���  ���o��  Chf���   ���@Kx��f���   ��fD���   ��A����)։�D��D)�A9�L�f���   ����   ����   ���  f���   ���   ���   �gfff1���vH H�\$@f���   �����H�T$@����f���   i���  1���f���   H�cinu  H�D$H������`  ���|���H�K@�r�����H  H��X  ���2  �r�1�H��H��HƋH9�L�H��H9�u�f���   �C���H���   1҉�L�L$<E1��    H�x8蝹��H��H�C@�D$<��������u�H��(  H��H��H֋G�H�� H��(f�B���f�J���H�B�H�J�H�B�H9�uԉk8���  ����H��  H�C(����H�P$H9��t����P���P��	���A���  �P���P��	���A���  �P�@��	ИA���  �(���I��  �r������   �+���1������L�T$H�l$L��M�nM9��r���E�L�T$C�M��D�\$L�D��0  I9��J���H�<$1�E1�L��L�L$@�   �U���1҃|$@ L�T$H��8  D�\$t"����A�LV����A�LV	��ɉ�H��A9�w�M�M�M�eM9������A�E D�t$&��@  A�EA����D  A�E����A�E	������  A�E����A�E	������  A�EA�U��	�L��H+E@HD$A��H��P  D���D��H  ���|$' t���|$&�������L$�������@��@�|$����� ���L$&���A��L�I9�����H�<$��E1�1�L�L$@�   �����|$@ H��X  �����H��1�D�\$&�n�0H�����p���	����|$�rH����|$ �8�G  H�p�@��	����BE���  ��~L�f�v����	�	��B��H��A9��\���A�4$I�D$E��tA�|$��I�D$	����|$' �2�Z������  �d���I������I�EI9�r~E�u L���  H�\$I��L��E��tiI�}H9�rTA�UE�m I�L9�rB��t��tH �;tH��H�HH��u�A��뽹 �B L��L���х�t�H�\$�D$@����H�\$�   ��I���D$@    H�\$�����L�f�����F	��������H�p@������f.�     @ H��  ��     �o��   �o�  N�o�  V H��(  H�F01��ff.�     @ ��0  f�1�� �   �f.�     �o�8  1��o�H  N�o�X  V �o�h  ^0�o�x  f@�o��  nP�o��  v`�o��  ~p�o��  ��   �o��  ��   �o��  ��   �o��  ��   �o��  ��   �o�  ��   �@ �ff.�     @ ATI��USH��H�/H�X�h��H��(  D���Y����u1H��(  H���   �oBC�oJ(K(�oR8S8H�RHH�SH[]A\ÐATI��USH��H�/H�X�Zh��H��(  L���Y����u1H��(  H���   �oBC�oJ(K(�oR8S8H�RHH�SH[]A\ÐH��0  ��N��@ H�GH���    H��(  t+SH��H��H��H�t$����H�T$H��0  H��[�@ H���   H��0  1��ff.�     @ USH��H��H�H�t$H��(  胭��H�|$��H�{X�sg��H����[]�f.�     H����  USH��H��H���   H��(  H��t�P��H���   H���W���H��   H��Hǃ�       �=���H��  H��Hǃ       �#���H��  H��Hǃ      �	���H��  H��Hǃ      �����H���  H��Hǃ      �����H���  H��Hǃ�      ����H���  H��Hǃ�      ����H��P  H��Hǃ�      ����H��X  H��HǃP      �m���H��8  H��HǃX      �S���H��@  H��Hǃ8      �9���H��  H��Hǃ@      ����H��  H��Hǃ      ����H���  H��Hǃ      �����H�C(    Hǃ�      ǃx      H�C0    H��[]��    ��    SH��H���.H �g��H��tH� H�C81�[�fD  �   [Ð���  ����   AW��AVL�<�   I��AUI��ATUS1�H��L���  �.�D  H��L9�t?I�4@:.u�L��� ��u�I���  �
   1�H�<��} H��[]A\A]A^A_�@ H��1�[]A\A]A^A_�1��@ AWAVAUATUH��H��SH��H��HH�F H�$H�FI��H�D$�V8H�L9��V  H�PH��8[�F  H���S8L�L;\$�2  A�<]�^  �D$ E1�H��E1�H�D$(    D��E1�E1��D$    I��<<�c  ��0��	w`�|$ �$  L��L�T$A�RHL�T$H����   L��I��A�R@L�T$A�J����   I�H�T$H)�L�xL9���   J�D0I�M����  A����  M����  L�d$E1�M+"����  ���@  ����   I��M9�r�L��L�T$A�R8L�T$M�L;\$�6  A�<]����I��M��1  L���    �C   H��H[]A\A]A^A_�H��    �T$H�<$H��I��L�L$4�   L�T$��L�\$ ��Hc������T$4L�T$H��  ����  L9�   L�\$ ��  C�I�UI��B�(I��M9�s1@ L9�   �o  C�H��  I�MI��B�(I��M9�rӻ   ������C�I�EI��C�(I��M9������L��  I��~�A�@A�P��Љ��D$����Hc�H��   I9���   H�<$�   L�L$4�   L�T$L�\$ �&����T$4L�T$H��  ����  L9�   L�\$ ~5C�I�UI���   B�(I��M9��-���I��H��  H9�   ˋT$���e����Pʉ�I9�rW�|$H�p(H��   ��H��H��1�     H�����H�H��   H9��&����H��ʉ�I9�rM��I)�I9�}��D$4   L�Ӻ   �S�|$ �����H�<$L������H��H[]A\A]A^A_� C�|7� I�F��1���I��� ����     L��L�T$L�\$ A�R@L�T$A�r��u�L�\$ I�M��I��L�I��I��?I�I���b���H�T$(H�<$M��L��L�L$4�   L�T$L�\$ 薫���T$4L�T$I�ǅ�uFL�\$ L��H�L$8L��A�   H��M�A�RXL�t$8L�d$(�D$L�T$�R���D  L���b���L�������I��L�������D$4   A�B   ������    UH��1ɾ   SH��H��H��8H���Uh��~wH�T$H��tmH��H�<$H��?H��H1�H)�H��   uhH�D$(H�L$H���  H��H�T$ H���  H���  H�L$H��H���  H���  H���  H��8[]� �E   H��8[]�f.�     H����4��H�|$H��H�$��4��H�|$H��H�D$�4��H�|$ H��H�D$�4��H�|$(H��H�D$ �4��H�T$H�<$H��?H��  ��H��   �.����� |H ��@��fD  H��H�Љ�H���  ��H��H�4�����1�H���ff.�     1�@�� wH�6     ��H����D  AWI��AVAUATUSH��8L��  L�n H��H�^�V8I�H9���  � ��0��	��  L��A�WHA�A��  ����  ����  I�H��H�H)�H��H9�~A��  H9���  I���   ��  I�I���  A��  L��H������r  I�M��   A��  L��L������Q  I�I���  L��   H�|$����0  �D$ E1��D$     D�l$D�l$�Ef.�     <>t|L��A�W@I�H9���  A�W����  E�A��/�^  A��(�T  L��A�W8M�7L9�v6A�<eu�I�FH9�v�A�~nu�A�~du�A�~�M�����t�f�     �D$�|$ A��  �o  I��H  ��1H �   H�H����� ���R  I��P  L�t$1��L��A��0  ���,  I���  I���  �   L���
H�A��0  ���  Hc\$ I��P  �   L����I��H  H��A��0  ����   I���  �   L����I���  H��A��0  ����   I��  I��  ��L��
H�A��p  ���~   I��  ��H��HI��  H�PA���  ��uYI��  1�L��HI��  H�PA��p  ��u4I��  1�H��HI��  H�PA���  ��t� ��<t�   A�GH��8[]A\A]A^A_� L��A�W@A�w��u�L��A�W8M�'L9�v�L��1��% <>t4L��A�W@A�O��u�L��A�W8I�H9�s�� </u׃���f.�     A��  M�'�����A��(�G  I�VH9��_���I�VH)ЉD$$�HD�T$�t$L��A��p  ���;���I��H  J��    D�T$H�D$(�D$$J��� A�~.u?I��H  �   ��1H J�<��L$ �� ����DL$�D$�L$ �   D��D$D�T$L��A�W8D�T$A��(uL��A�W@I�L��H�T$A�WHM�I9������H�T$�t$H��I)�M��A�IA���  ���p���I���  J��    E��I��H�B� �D$���D$E9�  ��������f.�     I�VH9�����I�VH)Љ����D$$����ff.�      AWAVI��AUATUH��SH��8L��  H�^H���V8M�>L9���  A��PЀ�	vK<[tGI�GH9��r  �iBH �   L����� ���V  ǅ      H��8[]A\A]A^A_�D  I�N H�$<[��  L��A�VH�D$ A��=   �>  L��A�V8I9s�H��8  I���   H�D$H��tDH�<$�a���H��@  H�<$Hǅ8      �F���I��  Hǅ@      H��t	I���   ��D��(  Mc�H�<$1�L�L$,E1�L�Ѿ   E���   L�T$����H��8  �D$,���  L�T$H�<$L�L$,1�E1��   L������H��@  �D$,����  I�E H�$D��I���   ��D$,����  E1�E��~9H�$D��M���   f�     �ރ��   ��1H L��A��  A9�u�H�$L��A�V8M�.I9��^  D�|$�$    H�l$L��D�d$�]�    <]�H  ��0��	waE���_  L��A�VHL��I��A�V8M�.I9��]  I�EH9��  L��A�V8I�.H9���  �E <du�L�mI9�s
�}e��  E����   L��A�V@A�F�������I���fD  I�GH9�vG�zBH �   L����� ��u/ǅ      ����A�F   H��8[]A\A]A^A_�f�     I�GH9�v'��BH �   L����� ��uǅ      �4���A�F�   H��8[]A\A]A^A_�f�     A�FH��8[]A\A]A^A_�D  I�G�D$A�   L��I�A�V8I9�$���������H�EI��H9�v�} /u	�$9L$A�F   �����     A��I��L��M�.A�V@I�H9������A�V���{���L)�L��D��H�|$H�ōHA��  A�F���T���I���   Mc��$J��� �.��� �}f�O����}�]������>���H�l$M��ǅ      M�>����� I��H�l$M�}��A�} /������$9T$������0���ff.�     f�AW��AVAUI��ATA��UH��SH��H�GH���   L�p8H�1�H���  H�<к
   �3m H��0  I��H���<7��f��D��D��C0��C@CPC`��   ��   Hǃ�       ��   ��   Hǃ�       I�uXHǃ�       H��0  ǃ�       Hǃ�       Hǃ       Hǃ      Hǃ       ǃ�       H�Cp    H�Cx    A���   ����   H��0  �oJ0�o��   �o��   M0�oR@U@�oZP]P�ob`e`H�JpH�MpH�JxH�Mx���   ��   �o��   ���   ��   H���   ��   �o��   H���   ��   H���   H���   ���   ���   ���   ���   ���   ���   H���   H���   H��   H��  H��   H��  H��[]A\A]A^A_�ff.�     �SH�H��H�wXH��(  H���   ����H��tH�{X�<��H�CX    [�f.�     AWAVAUATUSH��H���  H�   H���   Hǆ(      ��BH �T$�   �L$@L�D$�T����BH H�D$H��  H���   H�x�6T��H��  H����  H��$�   I��1��H   H��H�T$|�   L���   �H�L���e���D�d$|H��  E����  H��$�  H��t	H���   ��H��$x  H��t	H���  ��H��$  H��t	H��   ��H��$�  H��t	H���  �Ѐ�$H   ��  H����$�   D�t$|E����   �D$����   A��A����  ��   Hc��  H�S�CH    H�C    H�C H��H  ��(   H�Ct	H��H  H��  ��H�C0�BH H�CH�S(H���F  H��  H���F  � ���8  �
8�t1< �a  <-�Y  �� t	��-�
  H�����  �
8�u��FH��H���f�A�   H���  D��[]A\A]A^A_�D  L���   I�EL��1�Hǃ      1�H��Ǆ$�       �1�L��L��$0  HǄ$@      HǄ$8      Ƅ$H   �!t����$�   ����  ��$H   ��$�   ��  �D$|�����@ H��$8  H��$�   �K���HǄ$8      �0���f.�     H��  H��tH�C(H���   �C8    ��.H H�C@    Ǆ$�   	   H�x��P��H��$�   H��  H��$�   H��   H��$�   �D$@��t��$�   H�D$��$�   H��$�   H���   1�H��(  H��H�x�+�������  H��(  H���   �@8��H��(  H��    �o@h���   Ch�oHxf���   ���   Kxf���   ���   f���   ���   f���   ���   f���   ���   H�C    f���   ��*  ���   tH�C   �@tH�K�@ tH�K H�|$ �����M�m@1�H��1�H�cinu  H��$�   H��$�   I�}譟��A�ƅ�t<��t�����   �   f��$�   ���#  vP����  ��u0�   I�}Ǆ$�   EBDAf��$�   H��t1�H��1��E���A��E������f.�     ��u�   I�}Ǆ$�   CBDAf��$�   �D  �FH���{��� A�   �����D  �   L���;s����$�   ���*���H�eTypeFonI�O@H�%!PS-TruH3QH3H	�u�yttǄ$�      L���ot��D��$�   E�������1�L����p����$�   �������I�( M�g�N  H��$�   L��L������D��$�   H��$8  E�������L��H��L����q����$�   ���k���L��$@  H��$8  �D$|    H��$�   I�H��$�   H��L��$�   Ǆ$�       ��$�   L��$�   M9��F  L�l$(M��H�\$ �xD  </��   I�EI9���   M�uH��L��$�   �ҋ�$�   ����   H��$�   I��M)�A�W���wL9��   H����$�   L��$�   M9���  A�E H��$�   <F�x���I�EI9�v��BH �   L����� ����    H���ҋ�$�   ��t�L�l$(H�\$ �D����A�������     H��$8  L��萾����$�   HǄ$8      �D$|������L��$@  1�����f��   I�}Ǆ$�   1talf��$�   �	���1�I�} Ǆ$�   BODAf��$�   ������H����H����$�   L��$�   M9���   L���3 H����$�   ��$�   ������H����$�   H��$�   L9�s`�8ku�H�PI9�v¿VwH �   H����� ��u�L9�s4H����$�   H��$�   H����$  ��$�   uL��$�   fD  L��$�   �3��� L�l$(H�\$ ��$�   �D$|����������  *�  �D$|   �����A��wH �x1H 1�E��L�d$8M��I��L�t$0M��� ������  M�.I��0M��t�A�E A8D$u�L����_ I9�u�H�|$0L��L���3� ��u�Hc�L�d$8H�IH��H�wH �P���.  �@����  H�D$ H�   H��$�   H�4I��	E1�1�H��H��H�ƀwH ��H��$�   ��  ��$   ��$�   ���	����l���@ H��$8   ��$�  �D$X���  u�D$|   H��$   ��   HǄ$8      H��P  H��$H  H���  H��$P  H���  H��$�  HǄ$�      H��X  H��$�  HǄ$�      H��H���  ������$x  ����  H��8  ��L�l$`E1�H�D$8�D$XI��H�L$ H��@  ���D$\    H�L$(H��$�  H�D$PH�L$0H�\$h� I�GL;|$8��   I��H�D$ E1�fF�xH�D$(J���1H H�D$0N�$�A�G�D$DM��t�D�D$XE��~�E1�L�|$HM��L�t$P�f�I�GM9�twI��K�\� L��H���� ��u�M��H�D$ L�|$HH�߾�1H �   fF�4xH�D$(J����� ���I����D$\�L$DD9�OȉL$\�2���f�L�d$8����fD  L�|$H����fD  ������H�s0������    L�l$`H�\$hǃ,      �D$\��0  ��$P  ��(  �x���I�GL��IL��H��$8  L��$@  Ƅ$H  �j����$�   ���-���L��$@  ������tQ������H�D$ H0  H��$�   �
����D$\    �a�����$(  �#���H��H�|$ �P��$�   ����H�D$ H�  H��$�   �����@ H�H���   �Pt�W�@u��)ЉG1��+w1�9wv�F�f���O�P�   9�s��)�9Gv���щ�fD  1�1��ÐH���   �o@�oHN�oP(V �oX8^0�o`Hf@�ohXnP�ophv`�oxx~p�o��   ��   �o��   ��   �o��   ��   �o��   ��   �o��   1���   �@ U1�SH��H��H�?H���   �/���E\�������UlH�K0)���H�H�C8�Er��H�CHH��1�[]�@ AVAUATUSH��H�6�D$    H����  L���   �   M���H  ;V �?  ���J  ��E�L$I�t$fA�� �h  ��v   A�   H�V�L)�H9���   I�$�   D�@D��D� ��A	�E��D���   fA�� ��   D�h�PA��D	�D��I9���   A�t$lA����H��Ƈ�   A�D$\H�0�wh�����   ��Ǉ�       �G`stibL�H�wL�G H�G    H�G�-����  @ �-  H�EI��$�   H���   ���   D�pA��D���   t���   ��A��L�I;D$vmD  �   H��[]A\A]A^�fD  A�T$v����D  D�h�����    H���#   []A\A]A^�fD  �RA�   �� �   ���� E1�D��L�L$1�����I��H���   �D$���u���A�F�J�+I�D  ���   H�H9�v#L���    �2H��@�1Hc��   H�H9�u�I��L9�u�H��(  �@   �D$�����    ATUSH���   H��tWH���    H��L���   tH���   H���   �g��H���   L���*���H��L��Hǅ�       ����Hǃ�       []A\�@ ��}H ��"��fD  �FL�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H����t?��uI���   �Hl�   H9�t�@ �   �f.�     1��I���f�     I�@@H�@H�� H��H9�t۸   �D  UH��SH��H��H�7H����d����tH��[]�fD  H�S�@~H H���q����u��C���f�� ulH�Sf= tYH��uv\f= uHǃ�       Hǃ�       �CTu:H�3H���Vd����u�H�sH��H���   H��[]�ig��f�     H���   w�H���   []�ff.�     AW��I��AV��AUATU��S��1�)�H��8  L���   D��Hǆ�       H�<$L���   1�L��L����c�������D$0�L$���  ��$�   <�e  ��$�   ����  I���   f�{l ��  I�G�KrM�wH��H��I�Wf9Kp�  �{b tI�Of�{fvI�OH��$�   E1�1�L��    I���   H�D$謉����$�   H��I�G@���!  �Cp�{VA�G8   �H   D�cZD�sXf�E�C`��fClfE��Hc�f�E �H   LD�fE��H�}LD�L�������{lH�� ��H���Hc�H�EH9��q  H�}�H   L�����H�� H���H�EHǄ$      L��$  �{hMuǄ$  nmra�   f��$  1�H��$  1���}H 輏����$�   ��u<�Cu�St8�r%)�H�S��H�I�G H���   H9���  fD  Ǆ$�      I���   L�������I�w@H���:���I�G@    ��$�   A�G8    H��8  []A\A]A^A_ÐH�T$6��H L���nn���������f�|$6MZ�D$0   ��   L���i����D$0����"T$��$�   ��u�����@ H��I�G����� L��H��$�   ��   �su��H��I���   ��$�   ���W���H�4$I�   H�    H�FH���   ������$�   ����������������;���Ǆ$�      �����f�     �t$8L���`���D$0�������H�T$:��H L���em����������D$:�D$0   f=NE�5  f=PE��  I�H����  I9���  �D$0�������Ǆ$�       ���u������� H�}L��H   �?��H��H�E�v��� L�t$H)�L��H�rH��L���6t����$�   H���   �������H��H���   H��H��   �RQ H���   �( L���   L���;R H��M��M��H�H�   L������H��H���   ��$�   �������I�W(I�WI�G0�BH H�у�����   H�ɺDH ��|H HE�I�W0�~����t$8�D$<L���Hc��_���D$0���b����t$>�D$<L��)�Hc���`���D$0���?���L����b��f�D$f��wBD�t$�$��b��f����e  ���@��   H�ID$@L���b��L���f��u��b��Ǆ$�      �����H�������I�G0�|H �����t$8L���c^���D$0����   H��$�   �`H L���"k���D$0����   H��$�   PE  ��   H���  ����H�L  � H#�$�   H9���   f��$�    I�    ��   1�H��$�   D�t$H�D$���'H��$�   H9�$�   ��  ��f;�$�   �}  H�T$�@H L���xj���D$0��t��\$1��)���Ǆ$�      �����L�l$�\$�l$ �   1�� �����L��\$�T$ ��]��I�L$@I+L$HL��H�DH�D$�`���T$ f�������H�|$ ������Hk�vI;T$�m���I����z  I9��j���H�T$0��   L���-q��I���   �D$0������Ik�L��Ht$�\���D$0���w  �   L���^���D$0���^  L���`���L$I���   L����H���L$H��k`���L$I���   L����H��H���   I�D$@�_��I���   L���V����D$0������\$����H��$  L��\$�\���D$0���x���H�T$p� H L����h���D$0���Z���H��$  f�D$&  L�l$H�D$�\$�l$ ��$�   ��$�   �D$&�9��^  H�L$��L��H�H�t�[���D$0���'  H�T$@� H L���Qh���D$0���	  H�D$H�   ������H��������L��H!�H�D$HH�$  H��H�D$(�+[���D$0����  H��$�   � H L����g���D$0����  E1���$�   ��$�   A���9��v  H�L$(��L��H�H�t��Z���D$0���^  H�T$P� H L���g���D$0���@  H�\$X��   �����H��������L��H!�H�\$XH�$  H���fZ���D$0����   H��$�   � H L���%g���D$0����   1�H�������$�   ��$�   ���9���   �4�    L��Hc�H���Y���D$0����   H�T$`� H L���f���D$0��uz�D$[��V���H�|$@u�H�t$L��Ht$h�Y���D$0��uMH��$  ��~H L���tf���D$0��u0M;7tlI��M����D$0��������A���l���f�D$&����L�l$�\$1ҋl$ �����L�l$�\$�l$ ������|$0 �����Ǆ$�       ����H�|$H�T$0��   �Wm��H��I���   �D$0��u�H��$  H��$  L��H�$  H+�$�   H�H���   ������D$0���0���L�l$�\$�l$ �^���D  H��t;USH��H��H���   ����H�s@H������H�C@    �C8    H��[]�@ �f.�     D  H�H��  H��   H�WH�G 1��@ H�G     H�G    �ff.�     @ L�G L�O��1�L9�s?J�H��H��H��L�H92t1w"�5D  H�H��H��H��L�H92tv(H��H9�r�1��D  �B���H��L��f.�     H�xI����    �SH�_L�G 1�D�HM��I��L9�sDJ�H��H��H��L�L;
tnr'�vf.�     H�H��H��H��L�L;
tJs`H��H9�r�H9�s+H�������[L�L��G��I9Һ    DG�D��@ E1�1�[D��fD  �B[D����H��L��fD  H�xI���S���ff.�     �H��P  H�H��X  H�1��f�     �   �f.�     �   �f.�     1��ff.�     f��ff.�     @ USH��H��H�/H���<��H���  H��H�C0H���  H��H��H�C8���  ��H�H�CHH��1�[]�f�USH���FH�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H������   ��u H���  H��  �   H9�tH��[]ÐH���   []�@ H��1�H���s��H���  H��H�E0H���  H��H��H�E8���  ��H�H�EHH��1�[]�f�     H�C@H�@H�� H��H9�t�H���   []�ff.�     @ AVAUATUSL�6M���l  �   A;V ��  A��M���   1����  I�  �   �uD�MD�E �EƇ�   A��0  f���   �   A�D)�D���   �����   �����  ~&����  ����  �P?�������   � ���  �P�����   �U�����   ��D���   A��H�Hc���A��H�G0D��Hc�Mc�H�wHH��H�WPI���  H�0�G`stibI��  L�GH��H�G�J��A��  @ ��   Lc��   ���   H��L��L���p������   H�uL���S������   H���   L��L����T������   I��0  H��H�������   H��H��1��tdH���   ������(  ��uJH���   I��v;I��I��J�t�fD  ��HH���H��H��P��P��H��P�H9�u�@ 1�[]A\A]A^�D  �B�H�,@H�������[�   ]A\A]A^�f��P�������   �i���@ �P��҉��   �R���D  [�#   ]A\A]A^�f�H���   M������J�<&@ �H��������   ��U	щ��������   ��3	ʉ�������	ʈV�H9�u�I��0  H��H������H���   I������I��I��J�t`�     ��HH���H��P�H9�u�1������ H����   SH��H�F 1�H��H;u�2f�H��H�� H9H�t#H��H9�u�   I�    H��[��     H�GH�sH9�wH)�L�$L�D$�Q��L�$��t
�S   � H�SL�D$I�H�SI�H��[ø   I�    �f.�     ���H ���fD  AUATUSH��H��L���   H��   L���]���H��  L��Hǃ       �C���H��   Hǃ      H��t���  ��~b1��fD  H��   H��9��  ~EH�Dm L�$�M��t�I�4$L������A�|$ I�$    t�I�t$L���Ο��I�D$    � L��踟��Hǃ       H��p  L��螟��H�s(L��Hǃp      臟��H�C(    H�s0L���s���H�C0    H�s@L���_���H�C@    H��P  L���H���H��X  L��HǃP      �.���H���   HǃX      H9��   tH��[]A\A]��     �kO��H��H  H���   H��[]A\A]�f�H��t�V���fD  �ff.�     @ ��~aAVA��AUI��ATI��UH��S1�fD  H�} L����� ��tH��A9�u�[1�]A\A]A^�f�     Hc�H�[[]I�D��A\A]A^�1���     SH��H��   H�Ӌ��  H���t���H�¸   H��t�z H�Bt�   H�C1�[��    �C1��   [�ff.�     SH��H���� ���u �����H �`�H HD��:[��H��[�@ H�T$�@�H �![����u��T$�f��T$�f�S�T$�f�S�T$�f�S�T$�f�S1�f�S
H��[�fD  ATH��UH��SH��H�� H��p  H��h  L�L$L�D$������D$��t
H�� []A\ÐH�t$H���Z��H��H�D$�D$��u��� ���uу�H��x  ���H t���H H���MZ���D$��u�H���  H�H1�H)�H=�  ~H�� ��H���  H���  H���  H�H1�H)�H=�  ~H�� ��H���  H���  H�t$H���  H��I��   ����L!��l����D$���&���H�t$H���  H��L!��I����D$������H�t$H��� ���H��   t?H���  �o��  �o��  H���  H���  ��  ��  H���  ����H���  L!�H��������D$�������H�t$H���  H��L!������s���ff.�     f�AWAVAUATI��UH��SH��H��   H���   1�H�D$��K����$�   ��t A�   H�Ĩ   D��[]A\A]A^A_�D  H��`  ���H H���X����$�   ��u�H��`  fcpu�H��h  H��t�H�EH��v�H��H��	wH9�vH��	�	   HF�H��h  H�|$E1�1Ҿ    L��$�   ��q��D��$�   I��H��p  E���D���H��h   ��  E1��$f�     H��h  A�WI�� I��H9���  L�꾠�H H����W����$�   ��t�H��p  H�|$�9�����$�   Hǃp      �D$X�������H�   H�C    M�������H��h  H��p  L�D$`H��L��$�   �   L���   �����D$\���8  L�|$\H��L��L�|$�V���T$\H�D$`���  � ����  ���  H�t$H���rV��H�D$D�|$\E����   H���8��8��H��H��$�   H��H;T$��   H�D$A�   L�L$L��   H=   LF�E1�1�E1�D���  L��L�t$ �-p��D�t$\I��E��uvE1�H�|$ I����  H�\$(L��L�t$ ��    H��I��L9���  L�� �H �D$`t� �H H���V���D$\��t�H�\$(E1���D$\   �E1�E1�L��L������L��L���t����D$\�D$X������H��h  H��p  H��t/H�>   �4  1��H��H��H�<   �  H��H9�u�   H��H�������D$X�������H��h  H��p  E1�L��$�   L�D$`�   H��L���   �����D$\���p���L�t$\H��L��L�t$�T���|$\H�D$`���J���H�� ���� ����6���H����H����  H�t$H����P  �M���ȋt$\������H�|$`H��$�   �� ����  H���������H��H��H��H9������H�������H��   A�   L�L$L��LF�   1�E1�L��  L���	n���T$\I��H��  ���{���K�Dm M�,�f.�     H�t$`L��H��������D$\I�F    ����  A�fA9F|A�FA�V��9�}"1�fA�F1�fA�1�fA�F1�fA�F1�fA�FI��M9�u��D$X    fD  H��h  H��p  L�D$`H��L��$�   �   L���   ������D$\��������   H���H���D$\�������H����J��H��H�D$`���  ��J��H�D$H����I��H�D$`� ����b���H�D$A�   H=   LF�L;�  �@���L�L$E1�L��1Ҿ   L���l��I�ƋD$\������1�H�|$ �u  L�d$ L�d$H�\$(H���D  ��O��I��H��I9��.  L��H���D$`u��R��I����f.�     A�   ����D  L��H���O��H�D$�n��� ����  L��H���eO��H���g���H��  L��辔���D$\Hǃ      �D$X���[����F���fD  H��L��p  I����  �D$    1�M��E1�E1�1�I)��~f.�     H��I�T A�HH��L�JI��H�zH��L�H�pI9�v3�oL�H�r
�oPRL�A�   H�pL��H�xL�HH�zH9���   H)�H9r��   L9�r�E��t�D$�D$L9��V���H�UI�EH9��
  H��H)�I;}��  1��I�MH9���  H��H)�I9}��  �HI�� H��L9�r�I�EH9���  H)�I9UvI�U�D$X    �=����     Ǆ$�   	   �����H���������H��H��H��H9������������L��������H�t$H����O��H�������H��H�D$����H�D$H+D$ H��H�4�H�\$(�C���D$\����
  H�D$����  H�t$H���D$`�6  �0M��D�\$\E1�E������H�|$H��H��$�   H)�H9���  H=  �  L�L$L��HFо   E1�H�T$0H�JI��1��`i��D�T$\I��E�������L��H��H����C���D$\�������L�L$H�L$ E1�1Ҿ   L���i���|$\ �d���H�|$ H��   �  I�H;T$0��  H����  E1�I�OH�l$H��H�\$(L��I���fH����  H;D$0��  H�T$I�t L���"���D�D$\H�EE���w  H��H;\$ ��  I�H��I��H���c  H;T$0�X  I�t H�T$L���Б��D�L$\H�E E���%  A�V��UI�F����b���H�E�D�\$\L�d$ H�\$(E����   �   H�\$ H��H�t$H���D$`�}  �WK��D�T$\E���u
  H��u�1�H�|$ H�\$ H��$�   t2@ I��H��xH9�wL��  H�@HUI��H�QH��I9�w�H�D$`H��0  L��L���S����D$\�D$X�������H���   L�D$`H��H��h  H��p  L��$�   �    H�D$������D$\��������   H���vB���D$\�������H����D��H��H�D$`���  �-D��H�D$0� D��H��D���D��H�D$ �D��H�D$@��C��f��(  H���C��H�D$`� ����#����D$0������D9�����A���   �����t$ ��������|$@9���������   �����D��L�L$E1�)�H�|$)����   ��Hc�H�H��H�T$8H��I��1��f��D�D$\I��H�D$(E�������K�t- H���VA���D$\��u`D�|$GE1�H�\$H�\$ D�|$0���4 �C��f���tL��A�<I��H��L�H�:f�BA��E9���  H���D$`u�� C����H�t$(H�|$�_����D$\�D$X�������E���\  H�CH�ʒ��{   H�St�H�C���  L��   H�C    ��H �D$\    L���   H�D$`    L���H�D$h    H�D$p    H�D$x    ����H��t;�x t5H�P����<It<Ou#H�C   ���|H ���<O��H HE�H�D$p��H L��������H��t&�x t H�@� ���<BuH�KH�D$hDH @ ��H L�������H��t$�x tH�P���t���<NtH�T$x�    ���H L���Q���1�H��t*�x t$H�x�����  ���<N��  H�|$`D  E1�1�HǄ�       H��t��/ H���   M�lH��H��tH�|�`���    L��M��uH�D$`�BH �   HǄ$�      H�T$L���QQ���t$\H�C0���	���E1�J�t�`J���   H��t7H��H9C0t�  H��H��H���\. H��M���  I���  H�H��I��I��u��  �D$\�D$X�������H��   ���  ��H �!���H��t
�x �  H�C(    L�t$XH��  1�M��E1�H�|$�   �    �C8   H��H�C �b���T$XH��H�C@���(���f��A��   @H���  H���  H�2H��H��?H1�H)�H=�  �2��1�A��A)�D���  fD�} ���H L��   D��L���X���H����  H�@H��H��?H��H1�H)�H���� �N  ��  f�E�Z�H L��D������H��t'H�PH�xH��?H1�H)�H��� ��  H�E�  �K�H L��D�������H����  H�@H��H��?H��H1�H)�H���  �
  H�E�� A��� ��H L��D������1�H��t*H�@H��H��?H��H1�H)ʹ�  H���  ��1Љ�)Ѻ$�H L��D��L$�L����L$H���  H�@H��H��?H��H1�H)�H���  ��  M����  L�}��  A��  L�}L���H   D�D$�L$�l����L$D�D$I��H�E�   f���_  ���W  I��H��L���6���D���  L��   H�E�1�H L��D������H��H��t%�B�H L��D���|����} tH��t
�x ��  D�t$XE�����������@ H�������H��H�)�: u�-H��H9�u�������   H��H���z����D$X��������q����D$ �D$ 9D$@�����H��D�|$GH�\$H�<��H�|$L�L$L��L�D$(H�T$8�   �_���|$\H�D$(������L��  H��   �D$X    ����1��o����:E���~�����<��H�D$0��<��H��D���<��H�D$ �<��H�D$@�<��f��(  �n���Hkt$ �H����8���D$\���/����D$\S   E1��M���I�������G���L�t$XH�pH�|$L���U����L$XH�C(��������H���H�gfffffffH�HH��H��?H��H��H��H)Ș�1�)�f�E�����ZD���������1�)�A��A��Mc�L�}�������1�)�A��M����   f��������D���  L��   L�}�����   H��H)���7���������D$\    �;���L�}����M��u�L�}L�}뺺N �  ����D���  L��   H�E����Ǆ$�      �[����D$\   ����L�}L�}f���f���H������I���   �   �+���D���  L��   f�E�o����   A��  ����H�\$ �����L�|$H�pL��L���Ɔ���|$X H��P  �����H�uL��L��襆��H��X  �����H�l$H�\$(�`���H�l$H�\$(�D$\	   �I���H�l$H�\$(�D$\    �2���H�U�4��� AVAULc�ATL��I��UL��SH��H�� � �����tWH����  H��L���   �����L��L����2 <��  ����  L��H  L��H��L��L���   ��������  1����  t	f����   H��X  L��P  H���	  M���   ���߀�I��   �P��߀�S��   �P��߀�O��   H���S�H �   H����� ��td�Y�H �   H����� ��u�4hH �   L����� ��t2H�ƿ^�H �	   ��� ��uj�g�H �   L����� ��uRf�H�cinu  H�\$H�D$�Hf.�     �   H��tH�߉D$�����D$H�� []A\A]A^�f�     H�\$H�D$    H�T$1�1�� �H ��a��H�� []A\A]A^�f�L��L���9 <t���`���H��t?H���,���H�� �   []A\A]A^�f.�     L���   A��   �1 <�����   �U���f.�     �H����   �1�����   E1ɀ�-��   I����������H�ʃ�������`�H 1���r�<D  L9�KH������H H��H�P���H�ʃ�@������`�H ��r�H��H��M��HE�� 1��D  H��������H��H��M��HE���     �WA�   H���O���ff.�     f�H���   �1���txE1���-��   ��H�ʃ�������`�H 1���r�9 f=�J����H H�����B���H�ʃ�@������`�H ��rʉ���fE��E��fD  1��D  ��  ����fE��E���    �WA�   H���c���D  �����H�VH9W|�����f.�     H�H��  H��  H�RXH�G 1�H�W�H�G     H�G    �ff.�     @ L�G L�O��1�L9�s?J�H��H��H��L�H92t1w"�8D  H�H��H��H��L�H92tv(H��H9�r�1��D  �B�����H��L���    H�xI����    �SH�_L�G 1�D�HM��I��L9�sDJ�H��H��H��L�L;
tnr'�yf.�     H�H��H��H��L�L;
tJs`H��H9�r�H9�s+H�������[L�L��G��I9Һ    DG���D�ÐE1�1�[D��fD  �B[D������H��L�� H�xI���S���ff.�     �H���   H�H��   H�1��f�     USH��H��H�?H��  �X���H�E@H��H�C0H�EHH��H��H�C8�E��H�CHH��1�[]�f�     AW�   AVAUATUSH��L�6A;V �  �B����E  I��  H��    H��H)�H��H�Q`D��� H���PD�hD�`�hH�p H�H(�@���   ���   ���   ����fA����   ��   fA����   fA��u�   ƃ�   f���   �    ��A��I��H�{0���   ��A����? H����   ��H�CH���   Hc�ǃ�   stib��L�kPH�C0���   H�S@��H�C8I��  �p
��Hc��e���1�H��[]A\A]A^A_�@ fA���m���ƃ�   �a���f�     A��0  ����@ ƃ�   �<���@ ƃ�   �,���@ U1�SH��H�W�D$    H9�sRH��H��H�l�@   H�����t9H9�wAH��H�����w5H��H�L�L$�   L���T��H��D$��uH�kH��[]�fD  ���������ff.�     �H�GH��tSH�7H��H���X}��f��C[� ��    AUI���   ATUH��SH��L�eH��H���   H���� L���   L�L$�D$    J�"�T��H��H���   �D$��u$H��   H��L��H���� �(
�D$L��   H��[]A\A]��     ���H ����fD  I����������ʉ���������`�H ��1���r�L@ L9�w;Hc�H��H������H ���H�P��@��������`�H ��r���    H���������    ��ʉ���������`�H ��1���r�DfD  f=�w2Hc�H��������H ��΍B��@��������`�H ��r�ø������f�     �FL�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H����t?��uI��  H�HHHH@�   H9�tø   �f.�     1��I���f�     I�@@H�@H�� H��H9�t۸   �D  AUATUH��SH��H���� H�7H����z��H���   H�E     H��t"H�������H���   H����z��Hǅ�       H���   H���z��H���    Hǅ�       H���   tPE1�� I��L;��   s;O�,dI��J�.�xu�H�pH��I���Yz��H���   J�D.    L;��   r�H��E1��5z��H�}X L�e`Hǅ�       t@�    I�4$H��I��I��8�z��I�t$�H��I�D$�    ��y��I�D$�    L;mXr�E1�H�}p L�ext:�I�4$H��I��I��8�y��I�t$�H��I�D$�    �y��I�D$�    L;mpr�H�u`H��E1��y��H�E`    H�uxH���ty��H���    H�Ex    L���   tF I�4$H��I��I��8�Dy��I�t$�H��I�D$�    �.y��I�D$�    L;��   r�L���   L��H���
y��H��� H��Hǅ�       ����H���  L�� � t^E1��f.�     I��I��L;�� s7I�4$H���x��A�|$I�$    u�I�t$H���x��I�D$    � L�� � L��H���vx��Hǅ �     H��[]A\A]�H����   USH��H��H���   H��  H��t�&���H��  H���'x��H���   H��Hǃ      �x��H��   H��Hǃ�       ��w��H�s(H��Hǃ       ��w��H�C(    H�s0H����w��H�C0    H�s@H���w��H�C@    H��  H���w��Hǃ      H��[]� ��    AWAVI��AUATI��UH��SH��(L�oH�G    M��t*H�H�  �H H�@ �H H�@ �H H�@ �H H�@  �H 1�M���S  �U ���G  ��   ���7  f��E1��   )$)D$��ȉ��������H��t���t��+u܀~ u�A�   H��u�I�1�A� �H L9��#  fD  ����  �Ѓ�H���������s�  @ �����������rH�����u�I9��P  H9�IC�I�$H�FI�D$H�,�E����   �; ujE1�I;D$�V  H�pL��������u<I�t$I�$H��    H�M���,  H��I�t$H�  �H H�DH�     1�H��([]A\A]A^A_Ð� H�kI�t$H9���   1ɀ}  ��M�l$I9��&  �U �������H�1I��I9D$�o����U���������   �������4�у�����   H���fD  ����������o����E  H���E ��u�I�t$H9��_���1��a��� H��L�������������I�t$A� �H ����@ H��I9�tн �H �}���H��H�     H��(1�[]A\A]A^A_�I9�vHH��1����� M�l$I9�v1H��H�������M��tI�$붾   �V���H��H��I��H������1���f�     SH��H��H���   �����H��tH� H�@H���   [H���@ 1�[�ff.�     �H��  H����   H���    ��   H����   �> ��   SH������H��H��t1�H��tO��t2�   ��t[�fD  H�B�   H�C1�[ø   [��    H�@�   �C1�[��    H�@�   �C1�[��    �   �f.�     AWAVAUATI��UH��SH��H��(H���   L���� H���D$    ����H��tFH� H�@H���   H�ЋC����  ����  ���F  �D$H��([]A\A]A^A_� L��� H��L���^���I��H����  L���   L;��   �^  I�H�IH��H�� �H H��RvH�� � H��8���H���   K�RL�4�H�I��PA�V�P�@A�V���  ����  ���n  �P�H �   H����� ����  �E< ��  H�&     H����  I���X�H �   H��L���   ��� ����  �E< ��  H�&     H����  I�FH�C8�D$�����f�H�sL���q��H�C    M�������A�<$ �����H�T$L��L���r���fD  1�M��tA�<$ tL������H�C�[����M���_  L���   I�JL�L$L�Ҿ   L���7H��H��H���   �D$������H���   f��H�@H�� H�@    L���   H���   �1����    I�F    M�������A�<$ �v���H�T$L��L���<q��I�F�D$�������L���   �J���1�M��tA�<$ tL�������I�F�+����H���   I�>L��L���;R���D$���]���L���   �9��� L�������I�F������    �e�H �   H����� ��u0�E< w(H�&     H��sI�FH�C@�D$������    �q�H �   H����� ����   �~�H �   H����� ��������E< �����H�&     H�������I�FH����  ��D$��߀�P��  �C0   �j���@ L�������H�C�D$H��([]A\A]A^A_�f�     L��H��L���� �D$    ����H��ty�D$�D$������L��H������I���,���fD  L�L$E1��   1�����@ �E< � ���H�&     H�������I�FH�CH�D$�����    H��� L�� � L�L$L���   H�J�E��H��H�� � �D$���l���H��� f��H��H�@L��I�B    AL�$�Q L��L�L$E1�L�X1Ҿ   L��L�\$� E��L�$H��I��D$������L�\$H��L��� L�$L��L��H��� I�B   I�:H�pS�O���D$�������H��� �D$    ������Mu�C0   ������C������C0    �����   ����@ AWAVI��AUATUSH��H���   L���   1�H�|$�T$�D$x    L�<$����D$x��tH���   []A\A]A^A_�@ L��H�T$|�x@ L��H�      �D$|    H��$�   H�       H��$�   �1��I�ǋD$|����  H��$�   f��E1��   I�G@��  I��H@ �   fA�GI�FIǇX@     I��p@ H��$�   I��h@ I��I��`@ A�H@ I�~8H�T$@1�H�|$ Ǆ$�       H�D$8�NC��I�Ë�$�   ����   H�\$PE1�E1�   HǄ$�   �pC H�D$   A� H�D$(   L�|$HM��H�T$H�|$K�4/L)����H�D$0I�M9���  H�|$0 tSM����	  H�|$��  ��  L�l$L�L$8M���   H�|$ K�\- L��H���B��D��$�   I��E����  M��H�\$PL�|$HH�|$ L���Fk����$�   I�o8�D$|���   I�H��H����  �}0t�Mf�M4H�uXH�MpH�<I9tA�   fD���� I�@D�'E����   H	���   E�GA�wD����D)�D�ED9�t)�A�   f�}fD���� f;MtA�   f�MfD���� A�wf9utA�   f�ufD���� A� f9}t��A�   f�}��fD���� f�MD����D�D�E
D9�t�f�u
H���	  H���   H���1  H���� L���   �   H�JL�L$|�A���t$|H���   ����  I�G8H���   H���   � I�o8��  fD  O�'I�D$E�D��A9���  A��
��	  A����	  M���fD  ��
tI��I�vI9������C�\7M�7��u�A� A�D��<#��<����tI9�|uM�fH�D$(�   A�A��
�e���A���
   �   E��O��� M����  �D$x<������H�������   �����f�     H�\$�����fD  L)�L�T$hL��L�D$HD�L$`H��H��$�   H�T$(L�\$X��$�   L�\$XD�L$`�����$�   L�T$hu:L�T$`L�D$HH��L��D�L$XH��$�   H�T$(��$�   L�T$`D�L$X��$�   ������������D  H��u�D$|   �Af�     � �����   �D$|H��tH�������I�o8H�<$H��1���g��I�G8    H�|$@�n���L�4$I�w(L����g��I�G(    L��L���g���D$|�D$x<��������������D$H��  ��~	f���S  H�   H�C    H�K�   H����  H���    ��  �~�H H��� ���H��t
�x��  H���    �  ��H H�������H����  H�pH����  H�<$H�T$x�g��H�C(�D$x�������L��  �D$|    L���   HǄ$�       HǄ$�       HǄ$�       HǄ$�       H�C    M����   I��$�    ��   ��H L���/���H��t
�x�H  I��$�    tj��H L������H��t
�x��  I��$�    tC��H L�������H��t
�x�J  I��$�    t��H L������H��t
�x�  1�E1�E1�JǄ�       H��t�	 J���   M�tI��I��tJ���   ��@ L��M��uHǄ$�   �BH �   HǄ$�      L��H�T$|�f*��H��H�C0�D$|���U���E1�L��$�   K�4�N���   H��t5H��H9{0t� H��H��L���g H��M����  I����  J�<0I��I��u�� �D$|�D$x�������H�EP�C8   E1�1�H�<$L�L$x�   �    H��H�C ��;��I��H�C@�D$x�������f��A$AD$H�E@H���  ��H����  ��  H�EHH���  H����  �  ���H���    fA�<$��  ���H H������H����  H�@H���� H����	 ��  ��  fA�L$H���    �#  �Z�H H�������H���  H�xH��� H=�	
 ��  I�D$�  H���   H����  �K�H H������H��t!H�@H���  H����  �S  I�D$�� H���   H����  ��H H���=���H���t  H�PH���   E1�H��t#H���  A��  H����  w����1�A��A)�H���%  �$�H H�������H���  H�@I�|$H���m  H��u
I�|$I�|$I�|$H�MPH�<$1�L�L$xE1��   L�e`�	:��H��H��  �D$x�������ǃ0      H�}PH���\  H��L�M8I�L$1�A������fD  H��H��8H��H9��+  H�1f�PH�0L9�w�L9�u׉�0  ���    H��M���:���H��J�<1D  �8 u� -H��H9�u�����f.�     L��  H�C(    �1���@ I�Ľ   �G��� L��K�4'L��L)�E1�H��I���r �����     H�xH������������������<N�����H��$�   ����H��H��?H��?H% ����H�  f���H�E@������     H�H��?H% ����H�  f���H�EH�����D  H�@H���
���� ���<Mt<C�����H�K������    H�@H����������߀�Ot	��I�����H�K� ��|H ���<O��H HE�H��$�   �o����    H�@H�����������������߀�N�����H��$�   �����    H�@H���J���� ���<B�<���H�KHǄ$�   DH �&����    I���7���H���    t=�1�H H�������H���    I��t#�B�H H�������M��tH��tA�|$�f  H�BODA   H��$�   1�1����H H��$�   H��$�   �	>���SH�D$x�������H�SPH�H���   �����    A� I��M���p����H���  H����  �T  H���  I�|$��  A��  I�|$�H   �4���H��I�D$�   fE���O������G���I��I������I�D$�5���fD  H��������   ����fD  H�E(������    H���   H�U ����H�EH����   H��H��H=�  ��  HF�I�D$����� A�<$H���   �   �x���fA�D$�|���D  E1��w���H�gfffffffH�HH��H��H��H��?H��H)���1�)�fA�T$�9���f.�     �1�)���H�I�D$����@ ������1�)�A��H����  f��������fD  A�D$��H�I�D$���� I�o8������    H���N �  H��?H1�H)�蜾��I�D$�����f�M��H�\$PL�|$HǄ$�      �`����x�����I�|$ �����H�pH���w���L�4$H�T$xL���^��H���   �D$x���N���I�t$H�T$xL����]��H��H��   �D$x���&����E ���<I��   �E���<S��   �E���<O��   H���S�H H����� ��tL�Y�H H���� ��uH���   �4hH �Γ ��t&�^�H H��轓 ��uvH���   �g�H 訓 ��uaH�cinu  H��$�   H��$�   1�H��$�   1����H �:���c�����   A��  �	���I�|$I�|$���P���H�������H��$�   HǄ$�       �I��H@ 1�H�D$@�D���ff.�     �H�    L�WM��toH�1�E1�H� D  M9�sJH�N��A���t!I)�f�     H���L�A���u�L�WI��M9�v�� L�WH��M9�r�H= �H t� H��1��ff.�      H�OH��t0H��v1H�H�t��f�     H�PH��H�P�H9�u�H��H�O�fD  H�G    ��    AWAVI�ι   AUM��ATI�����H UH��L��SH��   ��À� �ۅ���   A�D$< ��   H�&     H����   I�x8H���t  H���    �f  �e�H �l���I�}8H���O  H��H����   H���    H����   �q�H �8���H����   �����I!E I��yC H�Ĉ   ��[]A\A]A^A_� ���H �   L����À� �ۅ�tl�P�H �   L����� ���  A�D$< ��   H�&     H����   I�T$��tA�D$ I�T$I�}8L���������h����    A�D$< w�H�&     H���C����q���D  I�E8H�H���H H��H�HHH��1��s� I�}8H��q�H �(������P  �������f�     H�G���H H�G@H��H��1��/� I�}8H��e�H �������u�I�}8�   f���� �x��� A�$M�}8�����  L���	u��  f�     <	�H  H�����u����  ����   I��� L���^���H����   A�����H�H�RH��H�� �H H��RvI�� � H��8���A���tD�3H��tr�ytlM��H@ H��L�⾮�H L��������Å������I��H@ L��L�����H������I�}8H��L�������������I�E8�   f���� ���� �I�4,����   H9�s4�F�<	t< u �     H��� H9�t�F�< t�<	t�<"��   I�}8H��L���a������;���f.�     � A�<$ A�	   tI��� L���!���H�������D�3I�4,H���  �@H����u�a���f.�     H������H���< t�<	t�<"����H��0���f�     �F� �W�����L���0���D  H���A�$ A�	   �{���� A�<$ D���Q����d���ff.�     �AWH��H��AVAUM��ATI��U1�SH��8  M�@8�D$    M��tI���� �P�H �   H����À� �ۅ�u]�H�� wTH�&     H��sDI�u@�v��tM��t����  H��H�pL���������H��8  ��[]A\A]A^A_�fD  M�M A����   ���H �	   H�ƻ�   ��� ��u��@	< w�H�&     H��s�M��h@ H�T$�8� I�E    I�E8    L������\$���m���I��h@ I�E8L��� L��L��H���� Iǅh@     �U���ÉD$���0�����H A� �H 1�� H��I��H��S��  I�<$L��L��H���$7���ÉD$��t������D  �   ���H H������� ����   �H�� ��  H�&     H����  A����   �����H��I��H@ H�¾��H �<����ÉD$���t���I��H@ I�]8H�xH����  �? ��  �����I��p@ H���   H��I�EH9���  Hǃ�       �   ����@ �   �˃H H������� ����   �H�� ��   H�&     H����   A����   �����H��I��H@ H�¾��H �l����ÉD$�������M��H@ M�M81�I�{H��t
�? t����I�{fA�AE1�H��t�? t����A��fE�Q
I�{����fA�AI�{ ����fA�AA���fE�QfA�AI�M �,���fD  �   ��H H������� ����  �H�� �v  H�&     H���b  M��H@ H�Ѿ��H H��L�������ÉD$�������L���b���H�t$�����I��H���  I�E8H��H�0��R��I�]8H�D$1�L�L$E1��   H��H�    H�H��)��H��\$���Y���I�E8L��H�8H�D$H�P�� I�m8H���{  H�] H���n  �; �e  I�E@f��H��H�D$     )D$H���� �@H�T$(�E0�V� L�`I���   �$  H��L��H�|$0�2� L��H�T$0�ۃH H�|$�p����Å���  H�|$ �=  H�|$�`���I�M ����fD  H�pH���o��� �   �n�H H������� ����   �H�� ��   H�&     H����   A����   �)���H��I��H@ H�¾��H ������ÉD$������M��H@ M�M81�I�zH��t
�? t�~���I�zI�A1�H��t
�? t�e���I�zI�A 1�H��t
�? t�L���I��X@ I�A(��  �   fA��� I�M ���� �݃H �   H����� ����   �@< ��   H�&     H����   A����   �:���I�P���H H�|$01�I�P@���A� I�}8H�T$0�e�H ������ÉD$�������I�U8���H H�|$01�H�JH�JH����� I�}8H�T$0�q�H �����Å������I�E8�   �����f���� I�$�yC ����fD  �   ����fD  Hǃ�       1�I�E    L�L$E1�1Ҿ   H���&��H���   �\$��tI�E8Hǀ�       �7����I�M I�$�lC �$���fD  I�]8H�T$�(   L���"��H���   �\$�������I�E8L��H���   �N���ÉD$�������I�U@I�E8�RH�@8�����P0�����   ����I�z �`���f��vfAǁ�  �����H������f���   �   �   E�F�fA��� �����H�D$H�@X���C��-�����H�        �   H��H��u.H�      H��u+H�      H���r����E0    �f����E0   �Z����E0   �N���H�|$���������f�     AW�   AVI��AUATUL��SH���P�H H��H��(M�h8��D$    M���� �� ��u �C���r  �P����&  <�  H�E � ��   �݃H �   H����� ����  �S�� ��  H�&     H����  H��H@ L��H�ھ��H ������D$����  H��H@ H�xH����  �? ��  ����H���������I�EPH��H�EH��H��p@ H��H9���  I�UPH�UH���Z  H���� ��  H�U �D$   ��@�[@ ��H �   H����� ����   �S�� �  H�&     H���  ��  ��  �D$�   ��@H��H����   �\$�0f.�     I�V�H�s����   L��������D$�Å���  H��(��[]A\A]A^A_�f�     ��H �   H����� ��uw�S�� wnH�&     H��s^%?���H�E0    H�E 1��f�     ��@�D$�   H��H���I���H�u(L���K��H�E(    �0���H�sI�V��C��� H��@tH�}0��}  �	   ��H H������� ��u4�K	�� w+H�&     H��s��  ��  �D$�   ���� �   �J�H H������� ����   H�}0���  I�uXH��    H)�I�u`L�|��I��A��   ��  H�uA�WH9���  �   ������H���   1�H�E fA���� �l���fD  H�E    I�EP@   �@   L�L$E1�1Ҿ8   L���!��D�T$I�E`E��tVH�U ��@�����f.�     �K�� �0���H�&     H������H����  �D$�   ����f�     H�M  1������@ H�M@D�IE���r���1������     I�uXI�}`� FC �8   ��� ������\$H!E �u����    H�u(L��L��H@ �I��L��H�ھ��H H�E(    L��������D$������L�������H�t$�4���H��H���(  H�D$E1�L�L$1Ҿ   L��H�H�H ��D�D$H�E(E�������H�L$H��H��H�Q�-� �\$H�M @��������C���@ �   ���H H��L�D$����� ����  �K�� �9  H�&     H���%  ���  H��H@ L��H�ھ��H ����L�D$���D$����H��H@ H�xH��t�? t����I��fE�G1�H�M    ����@ H��H��H@ L�񾮃H �����ÉD$�������L��H@ I�z����H�E0H����  �  H=�� ��  H��x4H��H����H�L� H�QHH���"  �   H�E0����fA���� H�E@�@����  I�UpM�ExI;Uh��  H��    H�M(H)�I��H�H�JI�MpH�PH����?����H#E H�E(    ��\$H�E ����f.�     I�upH��    H)�I�uxL�|���C���M�G(L��I��Iw H��'  �A�ɉ�A����A��E��@�H A����  E1��8�A��t�F H���I��A�ʉ�A����A��E��@�H A����  �Hc�I�Q�����H �H9�u�H��A�Of����  B�C��������@�H ��sH�E �   @uH   @H�E fAǅ��  H�E�\$�����   ��H H������� ����   �K�� ��   H�&     H��s{��tiH��H@ L��H�ھ��H �`���L�D$���D$�y���H��H@ H�xH��t�? t����I��fE�GH�E    �	  H�M    �\$�\����D$�   ������   ��H H������� ����  �K�� ��  H�&     H����  ��t�H��H@ L��H�ھ��H �����D$�������H��H@ H�{H����  �? ��  �����A��H�{fE�_H���o  �? �f  ����A��fE�OH�{�E���H�{ fA�GA���4���fA�GA���fD9MfE�OfDMMfA�Gf9E fME fD�Mf�E C�f9Ef�E"fMEfD9Uf�ED��fNEfD9UfDMUf�EfD�UH�E    ufE�_H�E@�8 ��  H�M    �\$�����H�U �D$   ��@����H������H�E �   @uH   @�   H�E fA���� A�Of�������H�E8��� ����H���0�H  H9��l����,����   ��H H������� ���A  �K�� �4  H�&     H���   ���k  A��� A�G��A�O����Hc�I�w(H��=��  ��   H����  ��   fA�O0E1�1�L�L$�   L���)���|$ I�G �����H�E    1�H�M    ���� H�E0����H��X@ w	H�E0�����I�z�\���H�����  H�E0���������H��M�E`H�QHI�UXI;UPt]H�JI�MXH��    H)�I��H�M(H�BH����?����H#E �H�
H�E(    H�E �"����D$   ������D$�   �����H�J@L�L$�8   L���<���|$ I��I�E`�����I�EP@I�UXH�E0�i����D$�   ����1������1��Q���H�JL�L$�8   L�������|$ I��I�Ex�_���I�EhI�Up����H�u(L���A���'���I�UI�U A���@ �?���fA�G�����E1�����E1��o���I�UI�U �@ A�����fA9G����H�}0�fA�GtII�G�   H�ƃ�H����H��I	���   H�M    fAǅ��  �����I�MP�{���H�E0�����I�EpH�P�����H�����   H��I	���@ ��    ���   ���$� �H fD  H���  �1�H���   t^H���  �@ H��0  �H���  ��     f��h  �t.H��h  �fD  H���  �1����   tH���  �D  1��D  1���w�����   ��������H ��!��ff.�      �Wи   ��	v���1���A�����@ D��0  ����������E��tWH��H  1�I�������  �f���H�� D9�t4f9pu�f�x t�f�8tAL�M!�I��uՉ9��H�� D9�u��    ��   ��x�@ �������     f�xw�f�x	u��:�ff.�     f�H�H��   H�RH9Qw���     H�w1��f�     1����   wH�W�F��f.�     D�A�PH��HW��BH����u��A�ȁ��   v�1�E1�D��ff.�     f�H�OH�F    �A�����A	���H�1��ff.�     �1�����  wU��H�WH��  ��u�H���N��f	�HD��D  �H�������B�    	�%��  H�H9�HD��H�A������H��1�H��t|�JE�������J	��2�ɉ��r��	���A)��r���r��	���D9�v9��t5B�A�rD�JH�|
����W��f	�tA����	����� 1��ff.�     f��I��L�OD�@A����  wGD��L�������H��tV�P�����Pf	�upA��   tA���   vE0�A��   A����  v�1�1�A�2� A��L��D������H��u�A���   v�A��   u��   L���e���H��u���fD  ��pA������	���9�v~E0�1�A�4D�@D��D�@��A	�H�LE��D9�s^A�A)��x�����x	���@ H���A������A�f	�t������6�����D9�u��D����     )�D�ƍz�A���*���ff.�      H�OH�F   �A�����A	���H�1��ff.�     �H�w�F�����F	�f�����G0�����H�G(1���     D�G0L�OA9��  G�\ AUE�P�L��AT��USH���  ��  �fD  f�����   ��A9���   �6I�D������PL�	��҉W<������PH�	��҉W8������PH�	��҉W@������P	�D9�r�H9_8u�f��t7L�'��L�l(I��$8  I�$0  I9��[����G@   1��
�     1�[]H�GH1�A\A]�w4�fD  [�����]A\A]�f��t���H��Ѹ�����f�     AWI��AVAUATUS�_(����  ��   L�7��A�   9_8C_8M��0  I��8  ��A�G4L���p������x}A�G89�B�A�w<9�w�I�WHA�@H��tw��A+G8�H�I�,H9�w��f�     ��9�r�H���B������B�f	�t������t�A�_([A�G,]A\A]A^A_��    �����[]I�G(A\A]A^A_�@ A�N D�>�2fD  ��xL=��  �9���A����  �,���D��)���9������;��9�vʅ�t�A�_([A�W,]A\A]A^A_� E�������������f�     AWA��AVAUATUSL�w�ӉT$�A�VH�t$���A�V��	���  �����|  ����������  �w  H����D$�H��8  H�0  H�\$�H�t$���1�I�|6H�D$�L�wH�H�|$�H�t$�fD  A�|VH�D$�E�DV��A	��<P�DPE����	���9�vE����   ��A9���   H�\$�A�z�4SD�LS��A	�A�2E����	���D��I�\:D��H�\$�!�9T$���   f�����   f���
  H�\$�H9\$��J  �   D  D�A��E��t\L�l$�A;E ��   ���Ä��9  ����  w/��A9�s��    H�BI��H9T$��  H�������D  1�H�T$��
[]A\A]A^A_�@ [1�]A\A]A^A_� f���t�E��t]��D��)��A�DL�H9D$�s��u�D�(D�@1�A��fE	��Y���E�A��L�D$�A;@ sV��A��D!��9����     D�������     E��xsA����  �.���A�=��  �����   )������ 1������f�     f����I���H�BI��H9T$������ 1��|$� ����������fD  D����������������@ AWAVAUATUSH��PH�OD�aD��D�a��A	�A����  �F  D���T$ ���H�t$H�|$�D$����   �D$���  A�T$D�L$1�� A9��  �nD9�sHB�t ��6H�D�8D�@H���D	�D� D��E��D�@A��E	�E��A9�v�A��D9�r�1�|$  ��   A9�s��9t$��   H�|$�������^  H�D$�X(��tV�h,H�D$��hfD  �����<���1�1�A���  말A��f�����  �|$  t4H�|$1��@�����u&H�D$�X(H�\$H���W����k,����  @ 1�H��P��[]A\A]A^A_�D  L�t$M�>M��8  L�|$8M�0  E��L�M��L�L$0�(D�HN�48A�L�t$(��A	���A��E�N�l$D	�L�L$��l$$�l$E�I ��D�L$@A��9�w]D!�f���uTf����  ��I�|>I9�s>E����  �FA��   E1�D$HA���  �D$@��  �A ����������� E��������~�|$Hf����F  D�T$@�|$A��E��D�d$$���  ������H�lD�E �EA��D	�A��D��A9���  D�T$DD�\$L�4f�     G�T �J�lD�m D�UA��E	�E��A9��	  E��H�D A��D�D��D�XL���A	��8E����A���xL�D	�D���A��D��D�PA	�fA���E��EE�E���t���D�\$@D�T$DD�\$LD�t$DD;L$H�  E9���  C�	H�DD�D��D�XH�D���A	�D��D�PL�E����A	��E�҉��P��	��ʉL$J�8�H�L$(�����A	����D$$�L$$��tf��D)ЍAHD$(H9D$0sD��1��D$ �������@��f	��X  fD$D����H�D$8;h �    C��j���A��A���  fD  �L$�|$  ��������H�T$8D��;j �@���1���  =��  �+����L$�   A�)ȁ���  O�����D�L$H�|$E��D�T$@A���  ����E���t����FA��|$E1�D$HA���  �D$@��  ����D�\$@D�T$DD�\$LD�t$DD;L$H�[���D9��X  H�D$(D�\$DA���|$D�T$@D�d$$D9L$��  C�	I��H�D�(�xH���	��(���|$D�x��	���A��9��_  A�|$E��H�L$D�t$DH�lL�l9D�ωt$$E��H�A��H�T$(�<f��u A�E�I���UA�M�����	�	�H��H������9�wCA��A��E��L�E�P�8���xL����H	������	�f���D��EE�D9T$u�H�L$�t$$D�\$@D�t$DH�T$(D9��&���D��D�\$D1��W���D�\$DD�T$@H�D$(�|$D�d$$�q���A������D���(���E1�D;L$Ht9H�D$(D�l$D�������D�������������A���D$   A���  �����|$E��D�T$@D�d$$�Z���A�y�D�d$$E��D�\$DA��D�T$@�|$�@���A�A��|$E��D�d$$A��D�\$DH�D$(D�T$@����H�D$�X(����H��1��t$����  w1�H�t$�G t����H����    �{���H���fD  H�OH�F   �A�����A	���H�1��ff.�     �H�O�A�����A	��Q��)Ɖ��Q	��	�1���9�v�H�L1
������A	�����    ��P1�����  ��   L�OA�yE�A��A	�A��E�AD��E�A	��A	�9�B�E��A��A)�C�M�T	
E9�vcE�
I�JE�RA��fE	�uP����  t8A���H���A��y���f	�u$����  t��A9�u�1�1҉�D  1��D  ����1���A�����     H�OH�F   �A�����A	���H�1��ff.�     �H�O��   H��   ʅ�t6��H�RL���   ��     9�sI9�t��HH���x���9�v�1��)�ω����9��    C��ff.�     L�G�1�A��   �����   Ƀ�M��   ����   �A�AVH�@ATUI���   SL�'������    A�9E�QI��E�A��9�A�B�A�A9�r_��I��E��)���I)�M9�wK��D�u<���t(����A9�r4��I��I)�M9�w'A�)�u�����u�1�[]�A\A^�@ A;D$ r�L9��w���1�1�[]�A\A^�f.�     �1҉�f.�     H�GH�F   �@ȉ�H�1���    H�O1��Q�9�w#)֋Q�9�v�H�L1������A	����ff.�     f�H�G�D�@L�HD��D�@1��Aȃ��tq��9�C�A��A)�C�I�E9�vgE�I�IE�IA��fE	�uU���t;A��@ H���A��y���f	�u$���t��A9�u�1�D��f�     1��D  A����D��A����A��A����H�GH�F
   �@ȉ�H�1���    H�w�F�G( ȉ�H�GH1��f.�     H�G0�����H9���   AUL�_@H��ATUSH�_HL9���   H�OK�[H�/A�����L�L�D  A�1A�IA�Q�A��ɉ�L9��A��IB�H9�r[O�,I)�M9�wO)�A�Չ�A�ukL9�tOH�PD�,H��H9�r.L��H)�L�L9�r E��uCA�   L9�t!H��H��H9�s�@ I��I��L9��o���[]�G( A\A]�@ �G( � D;m s�[]D�o8A\A]H�G0L�_@��    AU1�ATUSH�_D�cA�E����   D�����   I��H��E��E1�� E9���   D�QE9�s)C���I��H�t�D�F�A�A9�s�A��E9�r�1���t6E9�v��A9�t)D���E(H�E0��H�E@H���Q����}( usD�]01�E�] []A\A]�f.�     A���t�A���X����D�ߋv)ǉ�����9��    BƄ�t�D��H�U �E(H�}0��H�}@;B s���t��E8��    �E8D�]0�ff.�     @ H��1҉t$H�t$����H����    H�GH�F   �@ȉ�H�1���    H�w�F�G( ȉ�H�GH1��f.�     H�w0�����H9�wrL�O@L�WHH��M9�saH�WK�IL�H�L���    I��H��M9�t;��QD�Aȉ��H9�A�HB���H9�r�E��t�E;C s�H�w0D�G8L�O@� �G( �ff.�     AU1�ATUSH�_D�cA�E����   D�����   I��H��E��E1�� E9���   D�QE9�s)C���I��H�t�D�F�A�A9�s�A��E9�r�1���t6E9�v��A9�t)D���E(H�E0��H�E@H��������}( u[D�]01�E�] []A\A]�f.�     A���t�A���X�����FȄ�t�D��H�U �E(H�}0��H�}@;B s���t��E8�@ �E8D�]0��    H��1҉t$H�t$�����H����    H�GH�F   �@ȉ�H�1���    H�w�F�G0    ȉ�H�G8    H�G(1��ff.�     @ 1��ff.�     f��    1���    �����H�F   H�1��ff.�     f�D�E1�A��A�E9�v{G�A��B��    H�T��J����	��J	��JD��9�rB�Lf�     C����    H�L�D�Y��A��D	�D�Y�ID	�9�vA��E9�r�1�ÐE��H�L9�s	D�R�h����   �fD  D�E1�A�E9�sfG�A��C��H�L��Q����	��Q	�9�r8�>�    C�
���H�L�D�A��A��D	�D�AD	�9�vA��E9�r�1��D��E�� 9�vD�RE���y����A�����A	����ff.�     f�D�E1�A�E9�vqG�A��C��A�AH�D��HH������	��H�	�D��9�r8�K@ C�
����AH�D�D�@��A��D	�D�@D	�9�vA��E9�r�1��fD  H��E��9�v�D�Q�m���@ AUATI���U��SH��H�_H�{�B���H��t�D�h�Aͅ�uE��u9H��1�[]A\A]�@ �׉�H�������t�I�D$L��H�@H��[]A\A]��H��E���J�<+[]A\A]�(����     ATU����SH�_H�{���������H��t�D�`�A̅�u2�����E��u[��]A\ÐE���J�<#�����1�[]��A\���ډ��f��҉�H�<�����   ��t����     L�H��E1��pD I��x  I�Q I���   H�@��f.�     H�H��x  �` H�H��x  �` H�GH�@`H��t�����   �f.�     AWH��  AVAUATUH��  S��  HŅ���  H�HH��
H9���  A���D��  E1�I��A�   I	�f.�     D�AD��D�A��A	�E��I�L9�LF�E����   �QH�qM��I)���Q��	��ҍR�H�I9�}H��������*I��I��?D)�D�y�AA��A	�fA�� �uRD��   uy��tE�Aȉ�I9���   �B�H�@H�TA��    �ȉ�I9���   H��H9�u��     Eۃ�tI�@L��H9�����[D��]A\A]A^A_�f.�     E1�D9�v�F�2A��C�I�H��ɉ�I9�t=v)�kf�     C���I�H��ʉ�I9�twUA��E9�r��x����     �P�@��	ИA�A��DE��R���f��F�����F	И��D��A���     D�qD���W���E1�[]D��A\A]A^A_� H�L�HI9���   D�L�GfE�D�PfE�PfD�PfE�PfD�PfE�PD�PfE�P��t6L�HI9�wMf�PfA�P
f�PfA�P�@fA�@1��G L��fD  1�A�@
    fA�@1��G L���    �   �f.�     L�WH�GE�ZD�H����  AWAVAUATUSA�	D9���   E����   D��   C�A;��   �_"A�ٍ{��A��Hc�H�H9���   IcjA��A��D��E�Mc�MJ��A����   E��tl�S�Lc�A� �  ����A����I���,�f�     J�<L�ȃ��P  H���V�H��H9�u�K���H����tD��H����"M�A��u�1�[]A\A]A^A_�D  [�   ]A\A]A^A_��     E��tэS�A� �  1�����A���؍�I��L�ʉD$�N�&����    H���F�D��	�������@:H����L9�uދD$�K�!D�:��tf��I�rE��E�A��D��D�E!�D	�A��A��E	�D�:��~��D����@zI�A���&���N�&L��1����v�����I��D�:��u����D��L����D	�����    �   �f���L��H������ AWAVAUATUSL�OH��H�GE�QH�T$��P���  D�
E9��	  E���   D�8�   G�E;��  D�w"D��D��A�փ���Hc�H�H9��  E���t  E���k  IcAA�˺   ��A��)�D��A��D����   H�D$�E��D�|$�E��E�Mc�MYD9�N�1�E1��ى\$����)�����D��)ى|$��L$��   )ىL$�f�E����   D9l$��L  D9D$��1  H9t$��F  DD$���D��I�[�����L$�"T$�AA�ʃ��)  A��H��D��D����A��I��N�&H���~�H��	�������@z�L9�u���A��L�E��L��E��~F� �  D���;��E9�}kL��L;L$�s
A�	H��	�D��D����A��D!�	׺   @�;D)�A�L\$�A������1�[]A\A]A^A_� E��L��I��A���:���� D����E)���!�L��	�@�;�f�     [�   ]A\A]A^A_�f��D+D$������f��E��H���������H��	�����I������f.�     � �H �f���fD  AWH��AVAUATUH���nrekSH��H��(H�L$��@  A�����  H�t$A��   H����  H��  H�������A������  H��  H�|$A�    H��  �AH�L�A�����A	�f�� DF�E��f���k  H�A
H9��^  �A�Q�q�I	����	�	�D��f���6  A�   E1�1�1�I��������*A�   �S�    ��A9��  E��H�FA��H9��  �F�VD�F��	��V��D	�I��D��f����   ��L�H9�HF�A��u���f��u�M�pL9�r�A�@����A�@	�H��L)���I�֍@�Hc�I9�}L��I��?I���D)�D	���K���A�PM�pʉT$�P���t5E�@A�D��D9D$r� ���E�A�E��I9�����L��I��H��u�E	������f�     E1�1�1�f�     ��  ��  D��   H��(D��[]A\A]A^A_�ff.�     SH���  H��H���   �I���Hǃ�      Hǃ�      [ÐD��   H��(  I��I�L9�r�3 H�� I9�v'H;0u�L�HM��t�H��tL�	H�pH���%���D  ��   �f.�     AWAVAUI��ATI��UH��SH��8L���   �    ��L   ��  ��H  H��(  ��    �t$H�L$M����   H����   H���F� A�   I��H����   �t$����   H�L$�A
D�AH�\H�Q��A�����AE��D�A		�A�E	���fD9�t[��H�t��,��
H�����J���	��B���A���B�D	���f9�t%���H�H9�u�A�   H��8D��[]A\A]A^A_Å�t��H�D�L�<C�CD�K��A	�A��D�L$tv�3M��@  Ή�L9�sdL��L�T$H)�L9�vTI��8  H��H�H�D$�M A����u6�CD�L$ȉ�D�ȃ�f���*  L�T$��  f����  D  H��
L9��c���A�   �6����     L��(  f��H�L$(H���   �(  � FDBI�F     AFH�T$�������4  H�t$(H���%  H�|$L���������  I��(  H�T$(H�I��0  �1D�I�A���qA����A	��A	�ȉ�f����   H����   H�p�A��H��H9���   H�pH9�r|A��H)�L�I��@  ��    H�QA��H  H�<M��8  fE��t4�F�L�L��    �BH����A���B�D	������H�L9�u�I9�rAƅL  �����H�|$L������f��A�(  I�F     AFA�   �����    A�$   A�T$����fD  ��D�D$I9��0���HD$1�L��H��H�D$�L D�D$H������H�D$A�$   I�D$�B���@ A�$   A�T$�,���ff.�      ATI���1�H UH��SH��H�� H�T$�������tH�� []A\� H��B�H H���������u��|$u�<$tH�� �   []A\ÐH�T$I�$H�T$H�U �ff.�     �AUH��ATUH��SH����tLL��X  L���  �xtmvH�L$H��H����@  �Å�uH�D$H��I�E ����I�$H����[]A\A]�L��P  L���  �xtmh�ff.�     AWA��A��AVAUI��ATM��USH��H���  H��8L���  H��P  H��X  H���  H���  E��uH���  H��H���@&f��t.��H���   H�D9���   B��    H�H�FH9��P  1�1�fA�E fA�$M��tTA�$�D$(A�E �D$,E��uVI�H��tH�T$(D��H����I�FH��tH�T$,D��H���ЋD$(fA�$�D$,fA�E H��8[]A\A]A^A_�f.�     I�FH��tH�T$(D��H����I�F H��u���    D������H�$Mc�I�I�@H9��9���L��H��D�L$L�D$H�L$����D�L$���D$$����H�L$H�t$$H�������t$$D�L$fA�$�������D��L�D$H�$)�H�L$�t L�H�FH9���   1�fA�M ����� H��D�$H�L$�/���D�$���D$$�����H�L$H�t$$H���-���D�D$$D�$fA�$E���f���H�L$H�t$$H�������|$$D�$fA�E ���M����:���f.�     H��D�L$H�$����H�$D�L$���D$$����H�t$$H��D�$����D�$fA�E �����ff.�     UH��1�E1�S�   H���_H�oH��L�L$�K������T$��u]��ti�U H�u��t]�{�H�HA�?   L�L=�f�     H���V�H����t�z���`H��ACЈQ�I9�u�� H��[]ÐH��1�[]��    H����ff.�     ATH��1�E1�U�   SH���_H�oH��L�L$f��D��A�L$�����T$����   f����   �u H�M���u��	���f��trA�t$�H�xA�?   L�Tu�#@ H���q�H�����q���	���f��t�r�I����`ACшW�L9�u�A�  H��[]A\��    H��1�[]A\�D  I���� USH���G0�D$    9�r1�H��[]�f�H��I��L�G8��H�S@L�L$�¾   L��H���)���H�C8�D$��uĉk0��     AUATI��USH���Ʌ���   D�i�H��H�F1�J�|�D  �0H���L1H9�u��qL��H�]�Q�����uYI�D$8J�|�H����sH������	��s�	��s�H�t�fD  �
H����H9�u�H9�u��    H��[]A\A]�H��1�[]A\A]þ   �������u�I�t$8H����ff.�     @ ATI��UH��S�ˍs������uVI�D$8��t]�S�H�MI��H�t�	H� ��yH��I������	��y�	�A�P�H9�uډ�H���    []A\Ð[1�]A\�f�     H����ff.�     AWI��I����AVAUATUSH��L�wI�~�=���H����  D�(�@A�D��ȉ�	���  I�4>L��E����  E��M����q  I�A�m I�EA��˅��S  �U�I��I�t�1��    �H���T
H9�u����+  ���X  �tL��L���q������)  A�UM�UI�G8E1�A�MA�vI�~	A�   ������	�A�ME�m	�A�NF�*��	�A�vA�   	� Ic�A9�rFH��L�<09�vA�A��L�|0A��D9���   ��wH������	��w�	�Ic�A9�s�H�4��@ D���D�zH��A9�u�A��C�tE�A9��?  A�E�BA��I��E�j�A����D	�E�B�D	�F�*�Q�����u5H��L��L��L��[]A\A]A^A_�����H��1�[]A\A]A^A_��    L��L��H��L��[]A\A]A^A_�L���@ A9���   Ic�H���fD  ���rH��A9�u�C�TA��Hc�L�<�A9�sdE)�O�\�@ A�2A�RI������	�A�R�E�J�	�Ic�H���VB�<
�
�    ���1��H��9�u�G�DM9�u�Mc�N�<�A�    H��[]A\A]A^A_�Hc�L�<�A9�w�A��A�A9�sNIc�H�4��S�D)�L�D�I�D  ��OH��H������	��O�	ʉV�I9�u�D)�A�Ic�L�<��Mc�N�<��x���AWH��AVA��H��AUATI��USH��L�o(H�oA�u��������   M�|$8E����   A�E�H�]
M��H��H�DPH��fD  ��utH9�tP�CH���S��ʅ�t��D��I|$�T$�"����T$��t��C��S�I������	��S�	�A�E�H9�u�A�E     H��L��[]A\A]A^A_�D  ��D��I|$�y������u�����    E1��� M���ff.�     ATH��I��USH�o(H�_�u������ubI�D$8��ti�U�H�K
H��L�D�f.�     ��yH��H������	��y�	��V�I9�uۉ�H���    []A\�f.�     [1�]A\�f�     H����ff.�     AVH��1�AUATUH��SH��H��L�f8�psag��@  �D$��tH��[]A\A]A^�D  �   H��賹���D$��u�H��胻��H��f���  �t���H��f���  ����f���  v1�f���  H���   []A\A]A^�D���  E1�1�L��L�L$�   L�������H���  �D$���Y���J�4�    H�������D$���=���H���  E��t4A�E�L�d�f.�     H��H���ĺ��H��f�E�踺��f�E�L9�u�H���G����D$�����ff.�      AWAVAUATUH��SH��(D��0  L���   �D$    L��H  fE���  I������L��1�E1�Ic�Mc�D�D$A�   �D  ��H�� fA9��   f9pu�f�x t��f���  f����   f����   f��u����t�Hf���f��	u��Hf��
w�M��I��A��  t��HHc�f���f��	A���v���fD  A�����   ���t
E��x<E��u7I��L��A��C L�����t7H�{ ��   L��H��A��H�D$� H��L��Cf��vf��
t1�1�H�U H��([]A\A]A^A_�f�A���C ��     Lc�������     f�x u9Lc����������uC�|$���   A���t�I��L��A���C L����N���f��L$f�x DʉL$�{��� Lc\$E�������E����KL��`  1�E1�L�L$�   L���3����T$H�C��uH�sL��苴���D$��t(H�CH��L������1�H�C    1�f�C�D$������SH�sL��苵���D$��������Lc\$�|��� AUATUSH��H�����   t"H���  L���   H=   t$H= P ��   ƃ�   H��[]A\A]�fD  H��  L���A��1�f��   Hǃ      f��   H��  t71�f.�     D��L���J�4�����H��  J��    f9�  w�L������1�Hǃ      f��  �\���@ H��  L�����1�Hǃ      f��   �0����     AUATI��USH��H���   H��H  H�hH��tXD��<  I��I�L9�s.f�     H�sH��H�� �@��H�C�    I9�w�I��$H  H��H��� ��IǄ$H      I��$X  H��tSA��$P  H�@L�,�L9�s'f�H�sH��H������H�C�    I9�w�I��$X  H��H������IǄ$X      AǄ$P      1�fA��$8  IǄ$<      H��[]A\A]�fD  H���g  ATUSL��p  H��H���   M��t!I��$�   H��t��I��$�   H��tH���Ѐ�L   H���   ��  H��  �l���H��  H��Hǃ      Hǃ      ǃ       �� ��H��(  H��Hǃ      Hǃ      �� ��1�Hǃ(      H���   f��   H��0  �������   Hǃ8      Hǃ�      Hǃ�      �  H���  H���d ��1�Hǃ�      f���  M��tH��A�T$hH�s(H���7 ��H�C(    H�s0H���# ��H�C0    H�s@H��� ��H�C@    H��   H��������C8    H��`  H��Hǃ       �����H���  H��Hǃ`      ����Hǃ�      Hǃp      []A\�f�H��(   tH��(  �ڱ��H���   Hǃ0      Hǃ8      Hǃ@      �5���D  H��   H���I���H��(  H��Hǃ       �/���ƃ�   Hǃ(      �����     �ff.�     @ SH��H�8H�3�����H�    H�C    H�C0    [��    H�G@�G0    H��t H�w8H��tSH��H������H�C8    [Ð�ff.�     @ SH�H��H�w H���   �y���H�C     �C    [��     AWI��AVE1�AUATI��UH��SH��H��(�rH�T$D�D$f���D$    ����������T$����   I�wH��I��蔮���D$����   A�wH���k����D$��usA�GH�]@f������   �B�M��L�|C �; u�{A�ԅ�u�|$ t�CI��A�E�H��L9�u�A�E  H��臱��H��(L��[]A\A]A^A_�D  L��H��E1��b���1�I�wH��fA�GI�G    �G���I�G    �D  M��� AWE��AVAUI��ATI��UH��SH��H��(�BH�T$�D$    H�p������T$H�D$����   I�t$L���k����D$����   A�t$L���A����D$��uqA�D$I�]@����   ��L�t$L�df.�     �;�Յ�uE��t�I��A�F�H��L9�u�A� L���b���H�D$H��([]A\A]A^A_�fD  H�t$H���;���1�I�t$H��I�D$    fA�D$����I�D$    H�D$    �f�     H�D$    �D  L�t$�x���fD  I��H��H��tE��   H��(  H��H�H9�r��   �D  L�HM��uWH�� H9�v�H;0u����    H���   L�HM��t9I�H��tH���   L��鹬��f�     M�1��f.�     LPM��u�H���   L��L��酬��D  AWAVAUATUH��SH��H��H��   H���t  HcW8A�   H9�vu�4����  ���D  ��vw���6  H���  A�   �t�΍FH;�h  w7L���   ��H�`  L���7���A�ą�u�   L������A�ą���  H��D��[]A\A]A^A_�fD  H���  H�vH��H�T�B,f�E H���B-f�ED�JA��A��Ic�H�u�J��Hc�H�E D�R����   E����   H��H)�H��H����   H�E(�J�B�  @ E1��R����R  ��H�H�E0�Z����R  �}�  @ H�E�vZ��H�E�%���D  A�   ����D  ���  A�   H9�����������fD  A	��]����B��D��8  ��A��Hc�Ic�H�uH�E �4���fD  I��A���?  L)�L�E(H�u �)���D  H��H�H��H�M ����fD  L���`���L��A���U���L��E������D��R  fD�} I��fD�}H���  L��L���Y��H���  L��L��H�E�iY�����  L��L��H�E ���  )����  �Hc��>Y�����  L��L��H�E(�(Y����R  �} �  @ H�E0�Y����R  �}�  @ H�E��X��H�E����D  L��H�E     H�����?  H�uH��������    H��1���n��fD  AWH��AVAUATUH���CLBCSH��H��(HǇ�      HǇ�      H�L$HǇ�      ��@  ���`  ǃ�     H�|$wN�   H���   tL���  L��H��D$蹩���D$Hǃ�      ǃ�      H��([]A\A]A^A_ÐH���x���I�ŋ��  ���g  ���n  ���U  �   H��舩�����w���H���X���H��A���M���H��A���ҫ��H��I���ת��fE����  A���fA���0���I����  �#���H�D$J��   H9�vL�p�I��H���ϧ��H��H�p������������B�4�   H���  H��H���  �����������D���  ���  �>   H�L$H��CLBEH����@  ��uǃ�     H�|$���������� H�L$H��colbH����@  ��t�H�L$H��xibsH����@  ���G���ǃ�     H�|$�,����u���D  L���  H�t$H��L���Y���������H���  H�L$H���  ��RȉƁ�  ���H��   t%��  =   t�   �����fD  ����  �,  ��H�@H��H��H9�sH���������H��H��H��H�����  ���  Hǃ`      Hǃh      ��u@H�D$L��`  H��h  H����   1��w����    Hǃ`      Hǃh      ��t^H�L$H��TDBCH����@  ��t\H�L$H��TDBEH����@  ��tBH�L$H��tadbH����@  ��t(H��h  �u���@ ǃ�      1�������    H���h���H��`  H�D$H��h  �9����   ����fD  �   �m���fD  U1�H��H��S�TLCPH��H����@  ��tH��[]�f�     H��H���  H��@�H []����fD  AWH��AVI��AUATUSH��H��(L�f8H��`  �emanH�L$��@  �D$��tH��([]A\A]A^A_��    H��舤��I��8  � �H H��H��衰���D$��u�A��<  �I��L�lH�D$H�H��H�D$��   I9�w�fA��8  �6  L�L$E1�1Ҿ    L�������I��H  �D$���^���A��<  H�ߍ4@���/����D$���=���E��<  M��H  E���:  @ L����H H��D�$����D�$���D$uHA�Wf��t>A��@  H�IGI�GL9�r'H�H;D$wfA��8  ��  I�� f.�     A��u�M��H  E��<  M)�I��D��D��D�ʾ    L�L$L���
���A��<  H��I��H  �ԥ��A��<  fA��0  �D$�V���@ L��H���=����D$���;���H�t$H���D���D���D$L��E��P  ������L�L$E1�1Ҿ   L������I��X  �D$�������A��P  H�ߍ4�    躣���D$�������B��   M��X  I�A��P  H�@I��H�$I9�sM@ L����H H���`����D$A��@  H�IGI�GL9�rA�H�H;D$v1�fA�I��L9<$w�H��诤��H�uH���3���A��<  �D$���� A�Gf���T���- �  A;�P  �P���I��X  H�@H��f�8 �)����2���1�M��1��G���fD  U1�H��H��S�tsopH��H����@  ��tH��[]�f�     H��H���  H����H []�f���fD  AUH��1�ATI���pxamUSH��H����@  �Ņ�tH����[]A\A]�D  L���  ���H L��L�������Ņ�u�Hǃ�      1�H���  ��  Hǃ�      Hǃ�      f���  ~�L��`�H L���Ĭ����u@f���  ?w�@   f���  f���  ��b��������1�f���  �O���f�     ���?���f�     U1�H��SH��H����H��@  H��tD�aehvH���  �Ѕ�u$H�ھ �H H���2�����uH�C(    H�C0    H��[]��    �aehh�Ѕ�u�H�Ð  �ff.�     �L�W8LWHA��d��  AWAVA��AUA��ATE��UH��S��H��HH�w@H���E  I�BL�PH�D$(E�D��E�Z��A	�I�BH�D$(A�BE������A�B	���9�L��wD9�sHf�     H��H����   D�D��D�X��A	��PE�ۉ��P��	���9�r�A9�w�H�PH�T$(�@L��L)�ȉ�H9���   L�H�HL9���   H�PH�T$(����P��	�H�pH�t$(�xD�PH�L$(@�|$D�@f��wE���$�8�H D)ۍ�    H�H�AL9�w%H�QH�T$(�H�D$(�Iʉ�ɉ�H9��,  �A���%�   ��H��H[]A\A]A^A_� H��H�   []A\A]A^A_�@ �   �H�PD�L$D�T$D�D$I9�r�H�P�   H��D�XH�T$(H�t$(L��������u�H�T$(H�BH�D$(I)ǋ2L���H����H9��^���H���U���H�BD��D�D$D�T$H�D$(�Bɉ�D�L$�����B1�	���9�u6�L  �     L�\$(I�CH�D$(A�����A�C	���9��O  H��H9�u������f�     H�PL9������H�HH�T$(L9������L���pH)�H��Ή�H��H9������H�������H�xH�|$(�x�@��	���9���  1��4D  H�zH�|$(�z��A���zD	�L�ZH����9��Z  L��H��H9�u��#���D)ۍH�H�qL9�����H�AH�D$(����QH�t$(��	��A�I����	���H9������H9������H��D�L$�   D�T$H)������A�D��H�H;M0�����L�}HU(H�L�������������H�T$8H��L���3������y���D�T$�D$D�L$A��A	�H�D$8E��H�fA��H�D$0w!�   D��H��� ��  � ��  fA����  B�$�ؑH H�PD�L$D�T$D�D$I9������H�P�@�   H�t$(H�T$(H��L���D$�������������D$��D�D$D)�D�T$D�L$ȉ�H��H�������   H�t$8L���D$�Л���D$����H�D$0H��H9��  H�D$0A�p�C �}! �
  E����   E��E��D��H��H�t$0H��A���A���C ��H�UA���C �
�B�P�����у���9�s�H��H+D$09¸��C LD��A���C �I��1�H��L�\$(�Q���Q��	�H�yH�|$(�y���I��	���H9����������@ H��H�����D�L$1�H��H�t$0H������D�L$���M��������D�L$�   �Ҹ   ����1������}  t3H�MH�U�1�A�2H��B�}"�w�@����   @���$�x�H �   �r������B�Bf�B HcrH��H�������L�T$E��u�H�E H���   �X������/����E!L�T$�k����B�Bf�B 밃��B��f�B �B뜃��B��f�B �B뇃��B��f�B �B�o����   ������     AWL�~�   AVAUATUSH��I9��  D�6E��D�FA��E	�E��F��    M�L9���   H�WA��H���Bf�D$�Bf�D$�Bf�D$�B
f�D$
�Bf�D$�Bf�D$fE����   A�@�A�iL�t��	@ M9�t9A�7A�WI��E1�A��H�߉�A�w�A�O�D���	�D����������t�H�Sf�L$fD�|$f�J�L$fD�zf�Jf�L$
f�J
f�L$f�J�L$f�JH�K�q�	f�rf�
H��[]A\A]A^A_�1��D  H���   H��0  H��8  H�D$H�H�D$8H�D$8H�4$H���|  H�D$8H��H9��j  H�D$8H��H�D$8H�D$8H�T$8�@��R���f	��>  H�D$8H��H�D$8H�D$8H�L$8�@������A�	����D$,�D$,����  H�D$8H��H9$��  H�|$�4f.�     �D$,���D$,�D$,����  H�D$8H��H9$��  H�D$8H�|$H��H�D$8H�D$8H�L$8�@������A�	�f�D$lH�D$8H��H�D$8H�D$8H�L$8�@������A�H�|$`�D$h    	�f�D$nH�D$8H��H�D$8H�D$8H�T$8H�L$8�@�H�t$8�R�����	��V�	��Q���	��%���H��8  ��H�V�H�t$H9��
���HD$H�D$@H�D$@H�L$@� �����A	����D$0H�D$H@�H H�D$HH�8 u&�   �     H�D$HH��H�D$HH�D$HH�8 tdH�D$HH� H�D$PH�T$P�D$09BPu��D$4    H�$H�|$p1�H�t$@��Q��H�D$H�|$p���  ��$�   �� ��t>��$�   ��tSH�D$H�9���f�     1�H���   �fD  �   H���   � H�D$PH�t$pH�|$@�PX�D$4��     H�t$@H�|$PH�L$XH�T$`�'�����u��T$4H�D$X�P �D  AWAVAUI��ATUH��SH��   H��p  ���~	  �A�E1�E1�   H��I�T ��H=spgiDD�I��L9�tI� H=fpgiu�I��A�   L9�u�I���   H�xh �)  1�H��xibsL��A��@  A�   ���  H���   H����  H��L���Ѕ��D$<�$��  �D$ E����  A��R  �P�   f���?�=  H��L���SHH��L��D$<�S@H��L��D$<�S`H��L��D$<�SX�<$ A�ǉD$<�  H���   H��tH��L���ЉD$<H��L�����   H��L��D$<�SxH��L��I�m(�D$<�SpI�E(    fA��h  ��D$<A���  I�E0    I�E �D  A���  �6  E���}  H��   L��������D$<���X  E���	  I�}0 �(	  I�EA���  H���W���@��HB�H��H���|$HD�H��H��E��uI���     t	H  H��I��   tH��A���   tH�� A��  ��tH��@A���  �z  A��   I��(  H��H�H9��[  H��� H�� H9���  H�:fylgu�H�z t�H���fD  H�� H9���  H�:ravgu�H�z t�H��   �  I�U�D$<���,  H��I�UI��x  A���  I�UhI��z  fA���   I�UpI��|  I�UxI��~  I���   A��R  fA���   A���  fA���   fA��  )�fA���   H�  ����  I���   uJfA��h  �t?I���  ��  A���  A���  fA���   fA��  )�fA���   fA���   A���  A���   fA���   ��  A���   A��  fA���   A��   ��fA���   f���f��)�fA���   H�Ĉ   []A\A]A^A_��    1�H��L���S8�D$<���  1�H��L�����   �D$<<��R  ��u��   H��L���S8�D$<���@  �   H��L�����   �D$<���#  Aƅ�  H��L���SP�D$<���b���A�����fE��h  �O���@ H��   L��������D$<���+���I�E(E��u	H���  H����  I�m0�   L��H�������D$<�������A��I�E0u	H���3  H�������H��   L���U����D$<���t�������@ �$ �D$ H��L���S0�D$<���9�������D  A��   I��(  H��H�H9���  H���@ H�� H9�vH�8fylgu�H�x �����H�� H9�w�H���D  H�� H9�v=H�8 FFCu�H�x t��a���f��$ �D$�[���H�y �F���H�� H9��@  H�92FFCu����    H�x ��   H�� H9�vH�82FFCu���<������I��  eurt��  I���   �D$<�   H�Ph��   H���~���H�H�z �p���E1��D$<    fE���  ����<�������K���H��   �|$I�u��  A���  H�Ѓ�H�H��H����HE�I	EL�������A�MH����  M�MP1�E1�fD  I�<�   �`�H D�G�O��    H��H=�H �(  �9�u�P���tA9�u݋@�G=cinut=bmysuA�   H��A9uH�E���3  E���  E���)���I���   A��R  H�@8H�$f����  fA��h  ��   A��D�fEE�j  E��H�<$E1�L�L$<L��1Ҿ    L�|$ ����I�E@�D$<�������H�<$L�L$<E1�L��1Ҿ   �ű��H�D$(�D$<���������A��f�l$L�|$@f���D$    ���t$�D$A�F�E1�H�D$    H���f�     I��M�e@L��L��L�����   �D$<��uzH�L$�t$@�|$H��H��I�H�D$hH��fA�$�D$��D$�����fA�D$��I�D$�D$B��Hc�I�T$I�T$t��t�D$H�t$(�D$D�4�H�D$ I�FI9��[���H�T$ L�D$(L�L$<�   H�L$H�<$詰���T$���v���I�UI��   �D$H��I�UA�E8�Z���D  �G    �����E1�E1�����fA��h  ��<���A���  1�f����H��H���� HE��6���L�|$@1�1����H H�cinu  L��L�l$@H�D$H������t<������D$<    ������� ��������@ H��   L���x����D$<�������I�}( �x����W���@ A�   �   ����A��  �u���H��   L���+����D$<�������I�E0����H��   L�������D$<���Y����d���I���   �D$<�   H�Ph��   H��������>���I�U0�   L�������D$<�����������I�U0�B���H��   L�������D$<�������I�E(������D$<    �D$ �*���A���  A���  ��fA���   ���fA���   fA���   �N���1�H��xibsL��A��@  ��A�������ff.�     AWH�GAVI��AUI��ATUSH��(H�VHH9��-  A�E����A�E	�I�VHD��K�L% H�L$H9�w^f=vXI�]E1�I��  �D  ����A9�DB�L9�tAH���C������C�	�A�vP���vШt̾   L���'E��뽾   L���E���F�,�   J�+H��H�D$I�FHH9���  E1��A��L���C�sL�k��f	���   ���CA�vPD�[D�C�D$�C�$��vE�3���s��	�f��� w����   v#�   L��D�D$D�\$�tD��D�D$D�\$D����fD	�t2��I�t5�H9t$w�|- H�H9t$s�	   L���2D��A�vP��uA�GE9��-���H��(1�[]A\A]A^A_�D�D- M�M9�s��l$�$��	�L�����f�     I9�vCH���E������E�f	�t����A9FXwھ   L��L�$�T$�C��L�$�T$I9�w�H������H)�I�I��O�lE�T����   L���qC��������   L���_C���e���f.�     AWH�GI��AVI��AUATUSH��xH�VHH9��#  A�_I�VH��A�_��	�����L�H9�sA�FP����  I�^HD)����|  A�G����A�G	�A�VP��A��A���v���  B��   9���  A�FP��v^A�GE�oE�O
E�G����A�G		�D��E�o����A	�D	���  ����D9�w���D9��  �   L���JB����%��  I�TH�T$H�H�,H�T$H�H�D$XA�FP��v'A��$����I�L������A	�f����m  E���,  A�D$�E1�E1�E1ۉD$dI��L��H�D$0���D$`    H�D$hL�|$��   fD  E��E9�w(E��t#�rP����  E9��  D9��v  �L$`����@  ����  �4  �JP��LÅ��k  H9\$Xw��H�t$Ht$hD)�L	H�H9�vH�׾   �D$@H�T$8�#A��H�T$8�D$@�JP���_  I�L$E��A��I��L9d$0�>  I��H�D$H�|$I�h�]��M�F�4`F�|`H�D$B�4g��A��	�E	�F�|`B�D`��@�t$ B�tgE��A��A	�@�t$(A��A9������H�׾   D�T$TL�D$HD�\$P�L$D�D$@H�T$8�\@��D�T$TL�D$HD�\$P�L$D�D$@H�T$8���� f��������JP��wD;L$d�+  H�׾   �D$(H�T$ �@���D$(H�T$ ������    D;L$d�E  H9\$X�������H�rHD)�L	H�H9�������JP�������fD  A9�������H�D�|$ �D$ D)�L�tK�L$(A��H�l$(L��H��I��A	�E��D��I���	@ M9�t;I��A�F�����A�F�f	�t����9EXwپ   H���4?��M9�u��    H��D$ H�l$(�����    �L$`����fD  H�׾   L�D$H�L$D�D$@H�T$8D�d$P��>��H�T$8�D$@�L$DD�L$PL�D$H�@����D$`    �D$`H��x[]A\A]A^A_�D  E!�fA����x�������D  �   L���{>������fD  �   L���c>��A�G����A�G	�A�VP��A��A���v �t�   L���/>���i���f.�     �   L���>���]���fD  �   L����=�������fD  E!�fA�������������D  E��A��A�D D9��l���D��A����	��   ��9��Q����Y��� �   L���L$D�D$D�L$�=���L$D�D$D�L$����D9��������� �   L���S=��I�^HD)��R����    AVAUATI��UH��SH�FHH�_
H9���   A�D$E�l$H�MH����A�D$	�D��E�l$	��A	���L�E��H9�rfC�T6
��9�wZ�EP��tEfE��t?A�F�M�dD�f�L9�t-H���C������C�	���9EXw�   H���<��L9�u�[1�]A\A]A^� �   H���s<��뗐�   H���c<���=���ff.�      AWL��   AVAUI��ATUSH��H��H�FHL9��H  I�UH�CH)��9��<  =   �1  I�UH��   �����H�kL)�ȉǉD$������9��  �T$���$  �$    1�A��   �A�A�GI��E�O���A��9��"  �$��t9�w�   L��D�L$�;��D�L$A�UP����   D��A�UX)�9�r�A�D)�D9�w�   L��L$�I;���L$����  ����   ��u*�p�ډ��������  �t D������tz�SA9�tJ�Ӊډ������t ��D������u��   L����:���fD  �   L����:������fD  �$D��$9D$�����H��1�[]A\A]A^A_� �   L���:���t���fD  �   L��T$D�L$�j:���T$D�L$����@ A��  ��uO��u�f�     �SA9��t����Ӊډ��������  �t D������tԾ   L���:����D  �   L��L$��9���L$�f�     �   L����9������fD  �   L���9�������fD  AVAUI��ATI��USH�FHH�_H9���   A�EI�T$HE�u�L)��A�D��H9�rH��vH��H��H9�s�   L���S9��A�D$P��tE��u([1�]A\A]A^�f.�     �   L���#9��H��t�H���C������C�	���A9D$Xw���fD  �   L����8���U���fD  AWAVI��AUATL�gUH��SH��(H�FHL9��3  �E�]I�VH�ˉ���H)�H�$H9�r H��vH���������H��H��H��H9�s�   L���p8������   1�E1��l�M��t$I9�w�   L��L�D$�D$�@8��L�D$�D$A�VP��t-��A�VX)�9�r
��)�9�r�   L��L�D$�8��L�D$I��L��L9,$tUA�$A�l$I��A�D$���A��A��M9��p����   L��H�T$L�D$�D$�7��H�T$L�D$�D$�B���f�H��(1�[]A\A]A^A_��    �   L���{7������fD  AWI��AVAUL�oATUH��SH��H�FHL9���   �E�]I�WH�ˉ���H)�H�$H9�r H��vH���������H��H��H��H9�s�   L��� 7������   1�E1��8�M��tH9�w�   L����6��A�WP��tD���A;GXsFI��H��L94$tSA�m A�]I��E�e��ˉ��H9�v��   L��H�T$�6��H�T$� �   L��I���o6��H��L94$u�H��1�[]A\A]A^A_�D  �   L���C6�������ff.�      AWL�
AVAUATUSH��H��HH�FHH�|$(L9���  H�|$(H�CHD�w�oH)�A�D���A��H�t$H9�r"H��	vH�V�H���.�袋.H��H��H��L9�s�   H���5�����  H�D$   K��I�DD
HD$(H�D$ �*@ I�D$H�D$E����   ���`  L9|$ ��  E�'A�GI��H�L$��A��A	�A�G�A	�A�G�A�o���A�ŉ�M��H�D$L9��,  H9��#  L;d$s��   H����4��I�D$H�D$E���w���Ll$(H�CHM�uI9���  H�CHE�e L)�A�D��H��H�<$H9��T  H�<$ �4���E1�L�|$0E1��l$<M��L���f�M9�rRM�}I��L94$v_F�d�B�D�A����A	�B�D�A	�B�D�N�, I���� v��   H���>4��M9�s��   H��M�}I���$4��L94$w��l$<L�|$0�������L�l$H�CHLl$(M�eI9��z  H�SHA�m H���������L)�͉�H��H�4$H��H9��5  H�<$ �M���E1�L�|$0E1�M���Ef.�     L9���   �CPL�z��tA��@��A	�E��D;kX��   I��L94$��   A�$A�T$I������	�A�T$�E�l$�A�l$�	Љ�=�� v��   H��H�T$�3��H�T$L9��z����   H��H�T$��2��H�T$�^���D  �   H����2�������fD  �   H��I����2��L94$�X���D  L�|$0L9|$ �F���H��H1�[]A\A]A^A_��    �   H���2�������fD  �   H���k2���t���fD  �   H���S2������fD  �   H���;2���`���fD  �   H���#2������ff.�      H��tKM��tF��   H��t,D�ȸ�   A9�v1��H��H�(  H�H�H�FH�H�FI� 1���     �   �f.�     �=��  w'�G u;G(t$�   ���f��   �։��fD  1��D  UH��SH���[����C,��t�S(�U []�ff.�     �( t�H9G0t�   �H����     UH��S�&���1��( t
H�W0�G8�U []Ð�( t�H9G0t�   �(����     UH��S膚��1��( t
H�W0�G8�U []ÐUH��H��H��8  S�pamcH��H����@  ��tH��[]�@ H��8  H��0  H���u����t�Hǃ8      H��[]�@ AW�tsopAVAUATUSH��H��XH���   H�L$HH����@  A�ǅ�tH��XD��[]A\A]A^A_�@ H����r���    H��L�l$HI��L���  �Tr��A�ǅ�u�I��   t$A�   I�� P �a  ƃ�  ��     H�t$DH��L�u8��v��D�|$Df�D$E��u�A�   f;��  w�D��E1�L�L$D1�L���   L������D�D$DH�D$E����  K�4?H���Ts��A�ǉD$D����  �D$f���6  H�t$��L�d$ H�\$0H�DFH�t$(H��H�D$I��H��H����t��f�C�L9�u�H�T$(H��L�d$ H�\$0H�T$ �_t��H�T$ H�|$1� �
�ȁ�  ~D�Ɓ�  f-D9�O�H��H9�u�f�t$��L��L�L$DE1�1Ҿ   �'����|$DH�D$ ���  f�|$ ��  K�,D�|$<E1�I��H�\$0H���   fD  H��D$(��p��H��L)�H9���   D�l$(A�ML�L$DE1�1Ҿ   L��謖���L$DK�����  E��H��H��L���;q���D$D����  K��I��B�( fD9d$��  H��E���{p��H9��2  H�t$DH���Ut���t$D���V  D��L9��D���H��A���Ap��A)Ÿ    DH��I���H�t$DH��L�m8�t��D�|$DA��E���}���A�   f;��  �j���D��A�F�=  �W���E��L�L$DE1�1�L�Ѿ   L��L�T$襕��H���D$D��utL�T$H��H��H�L$L��L�T$�-p��H�L$��A�ǉD$DuGE���0  H�L�T$I9�|(H��x#�   @ A9��  H�H�H��I9�s��D$D   H��L�������D�|$D�����H�D$     H�t$ L���ڽ��H�t$L���ͽ��D�|$D�r���H�\$0�D$H�T$ ��H����L�d�fD  H�u L��H��落��H�E�    L9�u��H���yq��E1�1�1�L�L$D�   L��耔���|$D H�D$ �i���f�D$  �D$f��   �D$f��  H�D$H��  H�D$ H��  �����fD��   H��  ����H�D$0L��D�d$D�|$<H�D$(A��1�L�L$DE1��   �   L��H�\� �����T$DH���u1A���  fE9�r�H�l$ H�\$(fD�d$�M���D�|$<H�\$0�>���H�l$ H�\$(fD�d$����f�AUATUSH��L��x  M���  H��H��A��1�A�T$ H�E H���  H=   tkH=   tH= P �   H��1�[]A\A]�f����   ��   ��   A9�s�H��  D���<pf��vlH��  H�������H�E �D  A��  w�D��A�T$ H�E H��1�[]A\A]�fD  ���   tg��   A9��h���H��  D���<D�A�T$ H�E H��1�[]A\A]�H���x������M����,��� H���   []A\A]��     H���H�����t�� ���ff.�     @ H��t���  9�v���� �   �f��#   �f.�     AUATUSH��H�G H��xT�����H9�~cA�����I��H��1�D  ���  9�v$H�T$��H���&�����uH�t$L���s� ��t
��D9�r�1�H����[]A\A]�f.�     A��H��u���fD  H��H��t���  9�s
H�T$�����H�D$H����     ATUSH��H��tS���  A�   9�sH��H�T$������A�ą�tH��D��[]A\�H�t$��H��豺��H��D��[]A\�D  H��A�#   D��[]A\�ff.�      AWAVAUI��H��ATUSH��H��hL�v8��j��H�t$H��H�D$0��s��H�D$ �D$��tH��h[]A\A]A^A_�f�H�T$ � �H H���v���D$��u�H�D$ H=OTTO�]  �L$(I��fE��   E1�1�L��I��  L�L$�    ����I��(  �D$��u�H�D$0H��H�p�gi���D$���j����t$(H��H���:k���D$���M����l$(f����  1�E1��3f�     I��xtmh�s  I��xtmv�f  A��fD9|$(�f  H���Nm��H��I���Cm��H��H�$�7m��H��I���,m��H�SI9�w�L)�H9�w�I��(  f��t-L;7t��M�H����H��H���     H�� L;2t�H9�u���H�$��H��H�L�7H�OL�gH�G�W���D  H�D$0H��H��H��H�$�@h���D$���C���f�|$( �x  E1��D$    1�E1��D$    �4fD  H��GNIS��   H��ATEM�   DD� ��f;l$(��   H�T$@� �H H���t���D$����   H�t$PH�CH9�w�H�L$XH)�H�T$@H9�vH��xtmht	H��xtmvu�A��H��daehtH��dehb�h���H��5��   H��H���Zg���D$���]���H�t$H���Aq���D$���D�����H�߃���Hc�H4$�g���D$��� ����D$   ����@ �D$   ���� ��f�l$(fE��t2�D$��u��   D�|$������D$    H�D$ A������@ �   ����fD  H�Ѓ�������D  fA��   H����i���D$������   �|���ff.�     f�UH��1�H��SH��H��H����@  ��t
H��[]� H��H��0  H�ﾠ�H []��r��ff.�      �dehb�f�     �daeh�f�     AUH��1�ATI���2/SOUSH��H����@  �Ņ�tH����[]A\A]�D  L��h  � �H L��L���r���Ņ�uѸ����f��h   Hǃ�      Hǃ�      Hǃ�      ǃ�      f���  t�L����H L���*r����uNf��h  �n���L����H L���r����u,f��h  �L���H��L��L�羰�H []A\A]��q��@ ���'����AWI��AVAUI��ATUSH���   H���   L��p  �T$@H�_M����  �   ��BH �B��I���   I��x  �f  I���   �0  I�G8L�t$Iǅ�       H�D$Iǅ       Iǅ      f�     L����d��H�t$PL��H���8n��H�D$P����  H��FFOw�d  H��L���d���D$P����  H�T$`� �H L��I�_8�D$T    ��p���D$T����  H�D$hH=FFOw�j  H=fctt�^  H�D$pI;G�O  �t$xf���A  H��H��,   H9��,  H��H��$�   H��H9��  ��H�l$�  H��$�    H��$�   �  H�$�   ��   H��$�    uH��$�    ��   H�T$TH���iw��H�ŋD$T����   H�$    E1�E1�L��H���a���H�4$H���U���D�\$TE����  �D$P    �    M���   �l���@ L�t$H��   �  Iǅ�   fcttH��fctt�I  I���   �@�H L���Zo���D$P��uI��  H���R  f��   H���   []A\A]A^A_�f�     H�������H��$�    �������fD  H�T$T�P   H���^v��I�ƋD$T���  �T$x�Ѕ���  1��@ ����qu��   ����A��A����H�t$h��)�H��f��@�u H�t$hH��@�uH�t$hH��@�uH�t$h@�u�t$y@�u�t$xD�ML�L$T@�u�0   D�EE1�@�}H��f�U
1҈M	�L$x����H�$    I�ËD$T���?����L$xE1�1�L�L$T�   H��L�\$ 誇��D�d$TL�\$ H�$E�������D$xL��H�4�H����b��L�\$ ���D$T�����1�f�|$x M����  H�\$ H�\$H�l$(H�,$L�l$0I��L�\$�(f.�     H���D$xN�d� I��I��0D9��B  L����d��L��I�$��d��L��I�D$��d��L��I�D$�d��L��I�D$�d��I�D$ I�$H9�w�L��H�\$ H�l$(L�l$0�c���D$T   L�\$����H��H���u���L����_��L��H���b����D$T�D$P����������D  ��1H H���=��I��H���o  I��p  H� I���   I��@  �����f�H��fctt�����H��OTTOt:H��eurtt1H��1pytt(�dbk�H9�tH H9�t�   H��   ������Iǅ�   fcttH�|$H�T$P�   Iǅ      Iǅ     �ks��H��I��  �D$P�������H��D$X    f.�     �\$@I��  ��A����A1�A)�A�ǅ��[  Hcи   H9��_���H��    I��  I���   H�4H���^���D$X���1���H��L��A���   �D$X������A��H�L$`H��L��M���   D�<$�ravfA��@  ��uH�|$`�  1�A���  E1�E1�f�|$1ɨ�?  E1�E1�1�L��L���|���L��L���q���1�H�ھfylgL��A��@  ��t91�H�ھ2FFCL��A��@  ��t!1�H�ھ FFCL��A��@  ���]  D  ��9$��   �D$@1���6  I��  I�mI�E HcD$@I�E�D$X����D  ��H�H9���	  1����� ��.H H���:��1Ҿ�1H H���L;��I���  ������.H H���:��1Ҿ�1H H���$;��I���  �r����     ��H���^���@ H�$    E1������A��1�D$H�D$XH�D$�D$H�T$L��E1�D�L$(��H�L$ H�H��H�D$0��p���t$XI�ǅ��{���H�T$H�t$0L����p���L$XD�L$(I�ƅ�H�L$ �P���H��D�L$ H�L$�]��H�L$�T$D�L$ Hȅ�H�D$L�X�t|�D$M��A��f�l$ fD�L$FH�̓�L�|$(I�D�L�d$8M��L�l$HI��M��fD  L��L��   H���\��I��I�D$XM9�u��l$ L�|$(L�d$8D�L$FL�l$HE��D�L$H�L$E1�Ic�L�L��ŉD$�D$H�D$f����  f�l$H�l$0L�d$ M��L�l$(E��� Ld$A��D9l$�n  L��L��H��H���\��H��L��L���D$X�� ��u��l$L�d$ L�l$(����f�     I�GH��H9��  H�|$L�L$PE1�1Ҿ   �v���I��  �D$P���x���I��  L��H�4�    �\���D$P���U���1�I��   ~(@ I��  L��H�,�H����^��H�E I9�  �L����]���D$P�D$X���t��������    1�1������    �����A�   E1ɸ   ���b���fD  H�D$XH��H��H�D$�d��D�T$XI��E�������H�t$H���_��D�L$X��E��������   H��H�L$�"Z��H�L$���D$X�����H�t$H��H�L$��^��D�D$XH�L$A��E���\���H�t$H��H�L$�^���|$X H�L$A���7���H�t$H��D�L$H�L$�}^���|$X H�L$��D�L$�	���H�t$H��D�L$ H�L$�O^���|$X H�L$f�D$D�L$ A���  tf�D$  E1�E1�1������fD  I��   �����fA�������A�V�f���?weA���t$��   �|$9�t��9������f���~w;�|$��������Hc�H�Hc�H�H;T$`w��A�   A���  ���� A�   �>���D  �   �����fD  �   �����fD  H�\$ H�l$(L�\$L�l$0L��L�\$ �[���t$xH�<$���C �   �S �L$xL�\$ I��H��H�L$(H��H��fE��H��,   H�L$��  H�<$H�7H�~H9���   H�FL�d$pL9���   L��H)�H9���   H�VL��$�   L9���   L�$A��L�|$ I�HO�L�M��I��H�L$�QD  H9�r[H��H��H�N(������H�H�M9�toI�0H9~u5H�FI9�r,L��H)�H9�w!H�VI��L9�wM��I)�I9�s�f�     �D$T   ����� �
   �����l$L�d$ L�l$(������H�L$L�|$ H��$�   H��tH9�u�H�$�   H;|$pw�H��$�   H��t"H�W���H9�u�H�$�   H��H;D$p�u���H�D$H9�$�   �b���H9|$p�W���H�T$(H�L$I��H��L�L$T�   L�\$ H��H���|���|$T L�\$ H������f�|$x L�`�D$(    ��  L�\$L�l$ M��M��I�$I��L��H��A�E�I�$H��A�E�I�$H��A�E�I�$A�E�I�D$ H��A�E�I�D$ H��A�E�I�D$ H��A�E�I�D$ A�E�I�D$(H��A�E�I�D$(H��A�E�I�D$(H��A�E�I�D$(A�E�I�D$H��A�E�I�D$H��A�E�I�D$H��A�E�I�D$A�E�I�t$�#U���D$T���(  I�t$L����V���D$T���  I�|$(M�D$I�D$I�O@H�I9���   H��H�T$XH��H�D$X��T �D$T����   H�D$XI9D$��   L���X��I�D$ID$(�t�     �D  H���u�D$(�D$xI��0�L$(9��y���L�\$L�l$ H��$�   H��L��L�\$��S��I�G8I�uI�F0��C I���   I�F8H��
���@��M���   L�\$I�e��������L��H���E �I���H���*���L�\$L�l$ �����L�\$L�l$ �����H�������     ATH�GI��UH��SH�VHH9���   A�D$H�MH����A�D$	���L�H9�rSf=vM�EP��t:I�\$I��  ��     L9�tH���C�;EXr�   H���A��L9�u�[1�]A\�D  �   H���#��뤾   H������j���ff.�     @ AWAVAUATUSH��x���  ����  H��A�Ճ���  ����  H��   ��H��$�   �     H���  D�t�A�D;o �s  H��h  E��L9��`  B��   L)�H9��L  �D$   M��H��`  A��L��I�tL��NR���Ņ��)  �   L���'T���Ņ��  L���V��L��I���zV��L��H���U��A9���  ��   A��E)�A����   H��h  ��L)�H9���   H��`  E��L��L�L���Q���Ņ���   D��L���S���Ņ���   L���lU��L���dU��L����U��= gpj�1  w=epud��   �l$�1  L���1U��L��D����T��D;k �#  H��h  L9�vL)�B��   H9������ �   ���   H��x��[]A\A]A^A_�f.�     =lbgr��  =ffit��  �   L���MT���� H��h   ��   t�H��   L���   A��M�ϋ�H��`  L��D$�P���Ņ��z���H���   L�d$D�d$H�\$H���   H��$�   H�D$ 1�f�D$0H��`  H�L$(H���  H�D$8H��h  H�L$XH�D$@H���  H�H�T$`K�dH��H�r7H9������H�t�ʉ�H�T$H�Nɉ�H�L$P�v.@�t$2H9������H)�H��H9������E��E1�1�1�A��D��H�|$A��詰���Ņ������A��  P �����A��|���H���   H�|$L� � �   H�T$L��L���� �Ņ�tPH�t$L���K �;���fD  L��   �R���#���fD  �   �I���fD  �   ����fD  �D$*H�t$ A�G�D$H���   A�G�D$(fA�G����H���   H��(  �H����D  AWAVAUATUSH��HL��`  M��tH��HL��[]A\A]A^A_�@ H���   H��tH�G  �uq�G�ukH�L$0H�T$(�   H����]����t�HcD$(H��H  H��`  H���   �����  H��A�   ���C H��>���I��L��`  �i����    H���   L���   H���  ��  H�T$L�D$ 1�H��H�t$�S@H�EH�T$ �  ��I  �E��?  H��L��p  %�  H�X�H�BI��$�   H��H؋pH�D$(    �� ������~  ��  ����  H�T$0H���p��H�|$0H�T$ H����   ��? ���  L����H�tH�T$�a���L$I�ą������H���  H���o� ���  L�� -H�L$0H�p���t/fD  �Ѓ�0��	v��߃�A��w�H��H�����u�� H�^H�t$0L��M���(����x   HcD$0A�   ���C H��H��Ԟ��I���a���@ �D$L�bL�������tH�T$��  �`���T$���-���H���  H���� ���  I��HËD$����  H�D$1�H�t$0�����I�T$H9��  �_H�D$H��Ѕ���   L�Sy
�C-L�S��D����A����  H��f.�     D��H���������A)�D��A�Ӄ�0�C���u�H9���  M��H��� �B�I��H��A�C�H9�u�H)�L�E��tP�.C��L�S�D L�[��M�J��A�Ճ�0A�Q�%��  �  ���M9��!  M����@ �C0H��I�D$ H��H���� t*D��A��0A��	vA��A���A��AA��w�I�D$ H��H��H���� t*D��A��0A��	vA��A���A��AA��w�I�D$ H��H��H���� t*D��A��0A��	vA��A���A��AA��w�I�D$ H��A��< t�Ѓ�0��	�;  ��߃�A<�-  H�D$H����I��0H�D$;L$����M��L)�H�������ۍCI���A����A����Mc�M���  ��    ��Hc�A��[H�Hcɿ�[��[H��I��A��[M�L @ i��#H��iQ��J�8��i������iғ��1�iA����D1����������VD�i��J�81�iA������D�D���5͖�����G��i���#D1����D���;�2I9��v���H�؃��$�x�H f�     D�H��H�D$������    M��I)�I��t,��0��  L���	fD  H��H�C��@ �{�0t�����f�=�B ̀�1�p  = � �U  ��t�A�U/�S��    ��H�T$(H����L�|$(M����  L��M���(; I�\�E���1�A�@1�i������i���#A1�A�P����A�P
��1�A�@	��1�A�@1�i��J�8��i����A1�A�P����A�P��1�A�@��1�A�@1�i������i��J�81�A�P����A�P��1�A�@��1�A� 1�i���#��i����1�1�1�A1�D1ۍ>D���Aʉ�ˉ�����1�1�i�k��i�k�녉ȉ�����1�1�i�5���D����i�5���A1�Ai�k�녉ȉ�����A��1�A��D1�i�5�����1׉���1��>1��i�k��A��A��D1�i�5���A��A��D1�L�D$0�ƉD$0���t$4���  I�x�D$8L�T$<H���F�-�F	... H�F�     ��H����������H �HH9�u�H��L9��}���H�����1�����1�����1�����1��`���1��c���1�A�@��1������1��U���1�����1������1������A�P����fD  L��M��H)�H���!�����1��   ��0����A�U/A�S�����fD  L������H�L$H�T$�   H���yU������   HcD$H��H  H��`  H���   �����   H��E1����C H�躖��I��L���=8 ��[vA�D$[ �[   L���  ���  ���� L���H���=� �A����T���A�C�0�S���fD  H�L$H�T$�   H����T�����P���H�L$H�T$�   H���T����������,���HcD$E1����C H��H��4���I���E���A��[A��[��[��[����H�D$ I��$�   HXH���?����     AWAVAUATUS�H�|$����Y  �{  �C�L�~I��H�@M��L��L�\�0�    H�M H�E�H��� H��H9~0�o H�zH��L�J BL�PL�R(H�xH�x�H�L�HH9�u�H��I9�u�L�&D�k�1�   ��    D9���   D��D9�v��D�OH�@H��L)�L9�~�9���   A��K�RH�Ɖ����L�H�@I��1� HH�    H��H9�u��H�H��K�RH��D9�s�D��D��D��H�@L�$�D9�w� �    I�8 t���Ao��H�RH��
I�HH�JI��M9�u�H�\$��[]A\A]A^A_�f��GD��A��9��F���1�A���w����   ��ff.�      H��t
H��(:  H�H��t
H���  H�Ð��AWHi��	  AVAUHi�88  ATL�4USIcFXH�<M�N`LcPH��H�P�����L�|$�I�����fHH�\$�����I��H�H�� �  �    H��H�H�� HN�H�T$�I9��  ���  H��   H�t$��D$���H��H��    H)�L�$֐�T$�H�D$�E1�L�l$�����   �    �P0I������   ��A�I��A;Nh��8�tzI�1H�H�hH��I��H)�I)�H��L��H��?H��?I��I1�I)�H��L1�H)�I9�~
L�XL��H��H)�H��HH�Hc�H�T$�H��H��?H��
 �  H��Hc�L9�}I��M��H��8I9��U���M��tM�y(I��XL9L$�����[]A\A]A^A_�f�H�FP�N4H��   �V0H�GH�FXD�B�A�щ�  H�GH���8  H�GH���8  H�G 1�A����A���A���uE��A��uBA��A����AD�H�V@H���  �ʃ��~  t���ʉ�  1���  �@ A��t̃��ff.�     f���t\�F�L�GA�b   H�@L�T� H�� I�0H��H��H)�H)�HH�L9�}H��I��I��M9�u�H�H H���H9�~H��/H9�HO��H�J H��H���H��/H9�HL��f�     �F4H��   ��  H�FH�GH�FH�GH�F H�GH�F(H�G 1��ff.�     f�����ff.�     ����ff.�     H��t
H���I  H�H��t
H���  H�Ð��AWHi��	  AVAUE1�ATH�USL�@PHc@HL��I��M�t�F�H�@L�,�H��   �hH�   I��I��LD�Hi�p  H��M9��/  Hi��	  L��I��)g>îH��D  H��PI9���   D�^D;[hu�H�~L���fD  H��PI9�v��QH�AD�u�H9�}�D�I�QfD9NfDNNf9VfMVM��H��I)�M9��H)�I��M��t<H��
A� }  H�I��H-   H='  E1�H��~H��I��H��I��f�     H��H�I��L�H9F0~H�F0H�N H9A0�M���H�A0H�q �@���I�@ H��tL9@ tI�@     H�@ I�@(I��PM9�w�[]A\A]A^A_�ff.�     f�H�VPL�VH��   �F4�N0H�WH�VXD�A�A�ɉ�  H�WH��H  H�WH�� H  H�W 1�A����A���A���uI��A��t`����tFA��t
A�Bt ��H�N@H���  �y  u����  1���  �f�A��t҃���u���A�Bt��fD  ��u�����fD  H�S      H�G<	  H�G�   f�G H��  �  H�G$H��    H�G,H�  H�G41���     �ff.�     @ AWAVAUATUSH��   H�D$�L��   �     H��I9�u�L�_0H�_ I)�L�W(H�GN�,L��L)�M9�L�_8A��HL�K�,M��M)�L9�MO�)�A)�D9�A��A��@A��E��  ���  �L$�)���$�   A�݉L$�A)ͅ��  H��$�   Mc�Lc�Hc�H��$�   H�h��$�   ��H��H��L�tRD  H�E D�]H�T$�I��H��H��?L�� �  �EI��I�A)�H��M�I)��    I� ��?���H A��T��H��A9�}�H��PH�T$�I9�u�HcD$�D+d$�E�H)��f�     tCH��A9�|(�D��A�9Gh}�GhH�H���OlH�wXH�G`A9�}�H�İ   []A\A]A^A_�9Ol~���Hc��ff.�     @ AWAVI��AUATUSH��H��XH�GL�g�G,    L�o�D$L    H�D$H�G H�/�G<    H�D$��GH    �GX    Ǉ0
      Ǉ@
      ���?  H�@ ��  A�F�P����`��  H�{0 ��  �C,A�L���Ch   �C<ǃP
  �����?5����u�Ch����ǃP
     H�D$L�cL�kH�CH�D$Hǃ(      H�C HcC,Hǃ0      ���u  L�{0H��M�FH��M�^M�NI�H��   M�H�$H�@K�<�L�\$H�����   L�����	�D$4I9��  1ɉ�L�D$ L��L�D$L�|$(Mc�Mc�L�t$H��A��L�t$H�\$8�y��������f��N�P�^)�Hc�H��H��?H1�H)��H)�Hc�H��H��?H1�H)�H�H9�}f� H�pHH�F@H��H9���  H��PI��I��H9$��  �@�@I�I�Sf�HHc�I��f�PHc�I��H��H��?H�� �  H��Hc�L�H�H H�HH��H��?H��
 �  H��Hc�L�H�P(H�PL��H��HT$H�
H�Rf�Of�WA���������   f�������W89������L�G@H��8  I9��c  ��L�L$L�   H������I���^��H�C@�D$L����   A�FD�{8�P����`�|����s(9��|���L�C0H��x  I9��  ����L�L$L�P   ���H��A���^��H�C0�D$L��u-D�{(A�F�1���H�S@HcC<�l$4H��I��H��H9�ww�D$LH��X[]A\A]A^A_�H�\$A��H���D9��O���H�\$ Ic�L�SK�<�H��H|$(H���-���H�\$8L�D$ L�|$(H�S@HcC<H��I��H��H9��A  1�H��@ H��H��I��H��H��L�H�B�A�@���H9�r؋D$4L�|$I���������I��D�d �Mc�f�I�H�KHD�A�yH9���   �sD�K��)�H�H�H1�H)�D��D)�Hc�I��I��?L1�L)�H�I9�J�\  D  D�N��D�VD)�H�H�H1�H)�D��D)�Hc�I��I��?L1�L)�H�L9�}H��E��D��H�qHH9�u�H�A0    H��H��1�H�A8    E1�A����    f�
H9���   D�BD�RH�R@�zD)�Hc�I��zD)�M��Hc�I��?H�L��I��L1�I��?L)�M��I1�M)�N�I9�|�I��I)�I��M��L�P0I��L�R8M��I��I9���  A�   L9�}L��L��A�����L��    �   I)�L��H�H9�DM�D�HH�@@D��H9�tfD  @�p@�pH�@@H9�u�@�rH��E1�H)�H��I��H�p0H��H�q81�H9�����I��M9�����L�|$L;<$�H���L��H�4$I����������D  H��PH9���   ���u�f�xu�H�x8H�H0�XH�<�H��H��H����L�8L�E�CD)�E�BA)�D1�x��XE�C��D)�E�BA)�D1�x���H)�H��Pf�P�H��H��I��I�S0H��I�R8H9��m���H���������H�$�%A�WA�O8�t[�tfD  I��PL9��[���A��u�tσ�fA���fD  L9�}H��A������Z���D  L��L��A�   �D�����u�I�G0A�wL�$�I�G8I��L��O�,'A�GI��A�MA�UO�4L�$A�~)�)�Hc�Hc�)�A�~Hc�)�Hc��o���L�$���C���L��L)�H��H��I�F0H��I�E8A��:���H��E�ȉ������H��8  �G8   H�G@A�F�P����`������]���H�G@    E1�����H�C0    E1������H��x  �C(`   H�S0�1��� AW��$I�f��AVAUATUSH��  H�)�$�   H��$�   H�G@)�$�   H��H��$�   HcG<)�$�   H��)�$�   H��$�   H��   )�$�   HǄ$�    }  �PH���������H�D$h��H��$�   Hi��	  H��Ph�Hh�@H    H�G0��1�)�HcW,�L$PH��H��H���  H9�vf�H�HH��PH�H�H�H�H�H�H9�r�H��$�   H9�$�   ��  Hi�$�   �	  H�|$XE1�H�|pH�D$`H�|$x�|$P�|$H��$�   H� H�PHH�D$�B����1�)�;D$P��  E1��D$ 1�1�H�D$H ���H�\$H�� ���E1�H�D$@ }  E1�1�A� }  H�D$8 ���H��� }  H�D$0 }  H�D$( ���H�D$  }  fD�L$f�L$V� }  f�t$TH��D  H9\$t<��uLD�cE��E��A��E��E1�E)�D;L$P�:  H9[H�0  H�[@H9\$uĀ|$ ��  �D$��t�H�[@L�K0D�L9�IO�L9�IL�L�K8L9�~E��L��L9�}	fD�T$L��A��uM9�MO�L9�IL�D�KD;L$u�   H9\$�B���M��tM�OHM9K@�w  L�I�[HI��fE�KI��I)�I��fE�KD�L$E	�A��tI��M)�L;L$h}A�D�|$A��fA�K1�A)�fA�sfE�K
fD�|$VM��E1�H�|$HL�D$@fD�t$TH�t$8H�L$0H�T$(H�D$ �����    Ǆ$�       H�L$XHL$`HcAH����   H�QPH����  �pL���qHI��I�fo�$�   I�C�M��fo�$�   fo�$�   LE�I�[@fo�$�   AE�kD�3ASH�C0H�K8A[ H�SHAc0I�[HA����   H9���  fD�t$H��H��H�� ���D�d$A� }  ����@ HcQL9���   ������`  ����D�TD9��m  Ic�A������]  L�t$XLt$`D�T$L��$�   M�FPL;D$x�  H��$�   �P   �eT����$�   I�FP���   IcFHD�T$�PL��E�VLI��A�VHM^P����D  H9��O  H��I��fD�t$H��H��D�d$�B��� H�D$x�AL   H�APHcAH�PL��I���QHLYP�e���D  L�T$ L9�M��L�T$(LN�L9�LM�O�d L�T$pM)�L��I��D�SH��E8Q��   L�T$8L+T$0M��I��?M1�M)�I��I)�L�T$ M��I��?M1�M)�L9L$ �6  L�\$pI�_HfE�gfA�oL�\$(L�l$ L�\$XL�T$`1�C�lHE1������    A�H�� ���A� }  fA�C1�fA�KH��fA�S
H��fA�KE1�fD�t$D�d$������     fA�CH��I���� H�D$0H9�~	D�t$TH��H�D$8H9�}�t$Vf�t$H��H�D$@�T$I�_HfE�gI9�fA�oLO�H�D$HH9�HL�D	�A�����   H��L)�H;T$h��   ��A���H�T$p)�fA�OfA�G
L��fA�w�����@ �D$I�[HfE�cD	�fA�k�tH��L)�H;D$h}A���fA�KH�T$p)�fA�sfA�C
�Ao+�D$H�|$HA/�Aosf�D$VL��Aw�Ao{ L�D$@A �Aok0fD�t$TAo0�Aos@H�t$8Aw@H�L$0H�T$(L�l$ �9���f�����!����     �@   H��  []A\A]A^A_�f�     ����A��������H��$�   H��$�   H9�$�   �M���Hi�$�   �	  HD$XH�PPHc@HL��I��I�L9�r7�~    H9�~
H)�H��fJ
H�O@H�I8H9�~
H)�H��fJ
H��PL9�sLH�r@H�zHH�N8H�G8H�vHH�v8H9�|�H9�}
H)�H��fr
H�O@H�I8H9�}�H)�H��fB
H��PL9�r�1�����fD  H��$�   E1�1ҾP   �AP����$�   I�FP��t�������H�t$xH�xH���H�H�H���  H���  H)�H)��  �����H�IcFHD�T$��$�   �PL��E�VLI��A�VHM^P���X������f����H�D$�@����1�)�;D$P����H�t$�|$P H9������H�RH�B����1�)�9�t�H�B@H�D$�����H9��^��� H�HH��PH�H�H�H�H�H�H9�r��;���AWAVM��AUA��ATI��U��S��H��(�G�D$    ����   L�GE1�M���Q  Hc�H��H�JI��L9�w_�v 9�@��@��uc9���   �oB��oJ�H��X�oR �oZ0�ob@H�JPBXJhRx��   ��   H���   L9�v�r�@��u�9�@��@��t�A�D$��A�D$D��I�H��([]A\A]A^A_��     E9l$ �p����� HcW9�}L�GE1��+���@ ��]t��   ��L����D�|D9�}Ic�A��]tqM�T$I��$�  I9�toL�L$M�оX   ��M��D�L$1�I��I�D$D��E���U���E�|$A�D$����L���  �G   L�G�����@   1��#����]tA�]t����1�L�L$E1��X   L�T$�dM��1�H��I�D$�D$�������L�T$H�yH���I�L��H�I��$�	  H��  H)�H)΁�   ���H�M�D$D�L$�I����     ��AWHi��	  AVAUATUH�SH��(H�h`Hc@XH��H�PH����E�L�D A���A��L9��%  HcG,H�_0L�<�I��I�L9��	  H���.�袋.H��A��H��H��f��3��D����   ���   A���   H�CL�cH�u L9���   I�x�I9���   H���  ��   H����  L9���  �X   1�� L�HXI9�~L��H��L�T H�t H9��I9���  L�\�I�C A�;M�KH���  A)�H�Mc�I��H��H��?H��0 �  H��L�E��u&H�C fD	+H��PI9�����H��([]A\A]A^A_�f�H�C(��f.�     HEH+E�fD  H�CL�c�����f�I+@�I@��fD  I��1�L9�}KJ�4H��H��H�FL�T� M�
M9�|)�B�    H�7H��L��N�HN�T� M�
M9�}+H��H9�|�H��H�GH��L�T �����H��L���    M9�~cH�xI���|����    A�2H�L$H�T$)�I�zL�\$Hc�L�$L)�����L�\$H�L$H�T$L�$M�KA�;I�C ����@ I�B����I��1��]���ff.�     f�AWAVAUATUSH���҉�L�~L�n LD~LDnHi�88  H�L9�x8  �m  Hi�88  L�4A���  M��x8  M���8  M�~PM�nX���J  Ic�H��   E1��D  A��H��8E9��  �   H��c0�Hc�H��H��H��?H��
 �  H�KH��Hc�)�Hc�H��H�L�H��H�{H�{H��H��?H��2 �  H��Hc�L�H�S H�S(H�H�� �  H��H�H��0H��`�j���H�� L��H���H�{����H�SH��H)�xBHc�H��H�H�� �  H��Hc�1�H��~H�B H���H�s�K0H)�H�s(����fD  H)�Hc�H��H��H��?H�� �  H��H�H��+1���    L9��8  �����H��[]A\A]A^A_�@ H�� H���H���ff.�     U1�H��SH��H���oG�oNO�oV W(�����H��H��H�ߺ   []�����ff.�     f��ff.�      AW��I��AVAUATUSH��XH��   H�$Hi��	  H�U �RH�\HH�L�`PH�\$H�� �H HcPHH��@X    L�,�H�GI��H�\$ M����  H�_H�ƿ@   � ����D$ I��H�޿    �����Hc�   H�D$Hi$�G  H�t$(Hc��  H��H��H�H�� �  H��H�H��HN�����H��M9��5  Hi$�	  L�T$K�4vL��M��D$L�d$M��I��D$4L��M��I���f�H��PI9��3  H�S
H��L9�|�H�SL9��D�KA��t�H�{( t	�H�L9�|�A�GX�s��~C��I�W`H��H�HL�D�X����)�Hc�H��H�߅�HH�H9�}
D:J�  H��XI9�u�L�D$ �L$4A��L�L$HH�|$L�T$8L�\$�����L�\$L�T$8����  H�D$HH�xH�     H���H�@P    H)��HX1����H�H�T$HH�ZHH�ZP�C�BH�Cf�H�D$(H��H��?H�� �  H��H�BH�BH�[H��PI9������f�Hi$�	  L�d$M�I�s`McSX�D  I��PM9�vA�|$u�E��~�A�B�E�D$H��H��H�HL�L�X�fD  H��XI9�t��D��)�Hc�H��H�߅�HH�H9�}�H�BHI�D$H�BPL�`L�bPI��PMcSXI�s`M9�w�D  K��H��I�BH�,�H9�r�x  �    H��XH9�v/H�JHH��t�H�� H�PH�@H9�u�H��XH9�w�f.�     L�^H1�E1�L���   �    H�x(A��H�H H����   H�WH9�A��H����A!�H���6  H�y �+  H�V0E1�E���$  H��t:D��>D)�Lc�M��I�م��yMH�D�HA)�Ic�I��I��E��IH�I9�~H�QE����   H�V8�JH�@I9�t>� �M���H�x(��H�H H���N���H��t�H�y t�H�V0E1��n���f�     E����   A9���   �FH�~8 tH�~0 tH�F8    H��XH9������1�H��X[]A\A]A^A_�fD  H�BHH�CH�BPH�XH�ZP�W����    H�V0�@����    E���0���H�V8H��A�   �����D  �F �m����YE1��\$H���l���Hi$�	  M�McSXI�s`�����ff.�     AWAVAUA��ATUSH����L�~L�f LD~LDfIi��G  H�L9�H  ��  Ii��G  A��H��Ic�H�L��H  L��H  ���I  ��t/��J  H��PJ  ��t��   f��
H��H����   ��9�u�Ii��G  H�L�xPL�`XE���'  L�{L�c(Ii��G  1�H�3H��hH�ǋ@`��t=@ �Ѓ�H�@H��H�HcH��I��I��?J��  �  H��H�H�AH�A9W`w�Mi��G  I�Ic��  H��H�H�� �  H����'A���  A����   H��[]A\A]A^A_�1�fD  H��H�K@Hc���I  �IH��H�H�� �  H�CH��H���   Hc��@9�@�ƃ���@��t	�4   ��u�(   H�H���H9������A����  L�{PL�cXL�{L�c ����� L9�H  �G����O���fD  ���I  ���;�����H���I  A�@   A�    L��I������I������I��J��J  �>@ E1�H��~H��/M��MO�H�� ��H����r@H�BL)�H�B(H��HH9���   H�
L�rHc�D)�H��Hc�H��H��H��?H��0 �  Ic�I��H��I��?H��J��1 �  H�H��L�I��Hc�H�BI��?L�q0H�BJ��> �  H��Hc�L�H�r H�r(�r@����r@I��`�f���H���0���H����~   E1��2���fD  L���I  J�� J  L���@ H��HH9�������y0������u�L���f�     H��HH9�tϋP0��u��t�H�YH9�H�H9X|؃���y0�H���M��ML�����H��L���������I  �sH��t9��H���I  H��L���@J  f�H�QH�9H��H9�HL�H9�HL�H��HI9�u߉�Hc�D)�Hc�H��H��H��?H�� �  H����Hc��ޅ�Hc�HI�H�ƀ���uHc�I��L��H  L�� H  �\���ff.�     U1�H��SH��H���F(�G0H�H�G�F,�G4�z���H��H��H�ߺ   []�d���@ USH��H�/H���	  H�wPH�GpH��H�GH    H9�tH����f��H�CP    H�s`H��  H�CX    H9�tH���f��H�C`    H��8
  H��X
  Hǃ0
      H9�tH���xf��Hǃ8
      H��H
  H���  Hǃ@
      H9�tH���Gf��HǃH
      H�s@H��8  H9�tH���$f��H�C@    H�s0H��x  H�C8    H9�tH����e��H�C0    H�C(    H�    H��[]�ff.�      H��twATUH��SH�1�L���   �     H�t H��t6H��`�H �@H�� �H H�@ H��t
H����H�t L���ye��H�D     H��H���  u�[H��L��]A\�Te��� ���H �F���fD  @����   SE1ۉ�H��xk��tt��Hi�88  D�D`����   E��t"��Hi�88  H�DpH��H)�H��'H��N�8  H��5��   �6   H)�H��H�H��[H��E��HE�ÐH��A�   ��u�����   ���8  H���8  H�ʉ�����H��?��   �@   뱐H�|hH��D���p�����H��tX�@   H��?~�H�B H�������H���@ H��H���   �h���H�ʃ�?H��	�X���H���H����   H�A
�A����H��/:H�B@H���.���fD  D���8  E��� �������� H��H������� H���i���H�BH��������f�     H��0�0   HL������fD  H��*H��6H��HB����� AWI��AVI��AUI��ATUS�@   H����  ���T$u+�F�q  A�G�f  A���7   �1   HE�@ M�gI�mD��H��   ��L��H)������H��I�,H��H��?H�H��H��?H��H�L�H��H)�H�4
H��H����?��?�\  H���S  A�@   M��I)�H9���   H��?'H9��/  L9��&  I)�L9��  H9��  H�Ѓ� �  A�@   I)�L��I��I��H��L)�M)�H)�M)�I)�I9�IN�I)�L9�IM�H��H��?I��I��I��?I1�I)�L��H1�L)�I9�HOƋt$��u|H��~gH���   H�4
fD  I9�~jI�MI�wH��[]A\A]A^A_�@ 1�A����H�\;����D  1�H9�~�L9�}tD�D$H��H��E��utH���H������HL�H�H�4
I9��I�uI�OH��[]A\A]A^A_�f�1��q���f�     I��A��?M9��X���L9�������J���f�L�������     H)�H�4
�,���@ Hc�H�<�H��H�H9�w�; � H��PH��H��H9�v$H�F H�H�F(H�B��u֨�������f��ff.�     @ @����   ��A��Hi��G  ��>�   ��   U1�SH��H��yH�۽   ����   Hi��G  D�T`A����   A���O  H��O�@   HN�E����   Hi��G  H��H�DpH��H)�H)�HH�H��'��  H���   �v  H����  M����  H�FH���   �@��	�  ����   H�K H���H��[H�؅�]HE�H���fD  H���@ H�|hH��D������A����   �@   H��?~�H�H H����f�     A��u2�D$uD��(H  ������    H���   �H���w����    ��(H  H��0H  H�ډ��1����@   H��?�J���H�HH����=���D  H��8�8   HL�����fD  H��/~BH���U���H�HH��H���H��H)�H)�HH�H�������H�K@H��H��0HM������f�H�H@H�������@ H��H�ك�?H��	�����H��H����� ��   H�J
����@ H��0�0   HM�����fD  H���o���M���f���H�FH���   �@��	v;���I���H�gfffffff�   )�I��H��H��H��H��?H��H)�I��H���}*L������   )�I��I���������H��I��H��I��L)������H��6H��6HL������@ UH��A��D�ESH�ZH�BH��   H�I��  API��D�JH)�D��I)�����ZH�H�][]��    UH��SH��H��H��H���������tH��[]�fD  H�MH�U�D$H�s0�{,� ����D$H��[]�D  AW��I��AVAUATI��UD��SH��XH�D$Hi��	  H�H�XP�hH���������  Hc�H�4�H��H�H9�sV��H�S@L�KH����
�L9�t4H�R@�:A��	�A����u��H�R@�
��A	�tA��I9�u���H��PH9�w�E����  I�wHiD$�	  ��   L�H�XPHcPHD�hhI��   H�,�D�pHH���ɽ��H�D��H��H�T$H��H9�r�  D  H��PH9���   D�ZE9�u�H��fD  H9���   �qD���   D�A�rA)���   �q�yf9rfNrf9zfMzH��H��H)�H9t$lL�R0Mc�J�<�    N��    O�4L9�}M)�L9�|H;r8~L�B0H�r8H�J L�Q0N��    O�4L9�}M)�L9�|H;q8~L�A0H�q8H�Q  H��PH9��3���H��PH9�����H���f�     H��PH9��+  L�A M��t�I9H u�E�PD�IfE9�~�L�i0L9�~�N�4�    H���fD  H��PH9�v��rfA9�|�H9�t�H�z H��t�H9W u�fD;W�ufA9�t�H�r0I9�}�L9�}�H�r8H�4vH9q8��  H���D  L9���  H��PH9�v�L�^ I9�u�H�F     L�F(���    E����  E9���  �@H�x8 tH�x0 tH�@8    H��XH9���  1�H��X[]A\A]A^A_�fD  I�w�q����    H�S H��t)H9Z t#H�J0H�C     H9�
H��H9K0}H�R H�S(H��PH9�w�HiD$�	  I��   I�\HL�H�\$(HcPHI��@X    H��H�\$0H�XPH��H�<H�|$ E����  I�wHiD$88  L���  Hc�H��H�D$8Ic�H��H�H�� �  H�����i  1�H;\$ ����HiD$�	  H�D$fD  D�k���s  H�D$���  I�t`�A�H��H�PL�FX1�I��H�D$�*�     H��H��f.�     L��L;D$��   I��XD8nu���C)�Hc�I��I�م�L��IH�L9�HN�H9�~�L�[ M��t�L�VH1�M��M���f.�     A)�Ic�L9�}�M�IM9�t$M�Q M��t�A�BE�SfA9C�D)�H��� L9�HL�HL�L��L;D$�]����    H���o  H�BHH�CH�BPH�XH�ZPH�D$H��PIcLXH9\$ �����HiD$�	  H��H�QI�D`H�,�H��H9�r���� H��XH9�v/H�rHH��t�H�� H�QH�IH9�u�H��XH9�w�f.�     H�XHE1�E1�H���t�H�q(A��H��txH9FtrH�P8A�   H��t3D�
�8D)�Lc�M��I�څ��~MH�D�QfA9�~VA)�Ic�I9�~H�VE��tbH�P8�JH�IH9�������u�H�q(A��H��u�H�q H��t�H�P0E1��f�     D)�Hc���     �@ �e����    H�P0�f.�     �sL�D$01�A��H�|$(L�L$H�"������M���H�L$H1�H�yH�    H���H�AP    H)���X���H�H�T$HH�ZHH�ZP�C�BH�Cf�H�D$8H��H��?H�� �  H��H�BH�BH�[����f.�     H�F     H�N(�`����    I�w�d����    �   �.���I��HiD$�	  IcLXH;\$ �~��������D  I�@     H�A     �S��� AWAVAUATI��USH��H��L�j8H�i8I9�H��L��I��H��H��H��L�q0H�z0M��H��I)�L)�I9�tL9�uWI9�s�<�     L�H��PH�C�L9�w$H�C8H9�~�H�L9�H��IL�H��PH�C�L9�v�H��[]A\A]A^A_�D  L��L)�H�L$H)��5���I9�r�H�H�L$��    L�H�S0H��PI9�r�H�S8H9�~�L9�|
H���D  )�Hc�H��H��H��?H��2 �  H��Hc�L��@ AWAVAUATUSH��8HcG,L�G0L�O@�t$$L��HcG<I��M�M�<�����   L��M9���   H�P(H��PH�P�H�P�H�P�I9�w�A�   M9�s4M�1M�fHM9���   @ I��M9�wo�D$$����   M9�sfD  I�@0I��PI�@�M9�w�H��8[]A\A]A^A_�M9��s  L��@ H�P H��PH�P�H�P�H�P�I9�w�A�   M9�sL@ M�1M�fHM9��x���A�L��D��t�Jf.�     �D��u8H��PI9�s��J���M9��r����I�@0I��PI�@�M9�w��[���f.�     H��H�xPL9�s�PPD���'  H��H�xPL9�r�I9��  �PPD����   H����VPD����   H��H�nPI9�s�H9���   L9�s6H��H��L��L�D$(L�L$L�T$H�D$�����L�D$(L�L$L�T$H�D$I9��z���H�s�L9��m���H��H��L��L�D$L�L$L�T$����L�L$L�D$L�T$I��M9�������8���H��H��f�     H9���   H��H��L�D$L�L$L�T$�]���H��L�T$L�L$L�D$�����fD  I9������H9��K���fD  H�C0H+C8u����f�     I�V8I��PH�I�V�I9�r�H��PI9�������    H�S8H��PH�H�S�I9�s�I��M9�������k���f�H���;���A�   M9�������u���A�   M9�������a���AW��AVAUATI��USH��(H���  �  ��Z�W���I��1�I���  �/  �E$D�E(D�}<M���1  A��Ic;   Mc�L��L��H��?I�� �  H��Hc�A���Ƀ�)Ή����   ��   B����)����-�V  D�����ǉ���H9���   D�M,�U0�M4D�u8E�ʉT$�m@A��L9��[  ����H9���   D����H9��&  A)�H���s���E���  D)�A)�Ic�A��Hc�Ic��r���D��H��H���D���H�| �D  A��H��D���)���H��L������ �  ��H��([]A\A]A^A_��    �   A�  K �  K ����� ��L��H�މL$D)ʉT$�а���L$HcT$�������<���D�|$A)�Ic�E)�A��Ic������D��H��H��蒰��H�| �b����     Hc�H��H��H��?H��1 �  H��Hc�����fD  ��H�މ��K���H������ D��H��L�T$)L$D�D$D�L$�T$����HcT$D�L$D�D$�L$��L�T$����D�|$A)�D�D$Ic�E)�Ic�����D�D$H��H��A��D���ʯ��H�| ����AWAVAUATI��UH��SH��8H�G H���   H�4$H�T$(H�� �  ����I�ǋD$(��t H�$L�9H��8[]A\A]A^A_�f.�     H�U H���   1�I�/I���  M���  I�WI�_fA���  IǇ�      IǇ�      IǇ�      IǇ�      IǇ�      H�D$��t$��H��I��W�  @ ��?  H��f�H�H9�u�cinuH����������  E1�A��H ���H H�D$��H A�p�H �7f.�     I��M���c  A�EH�� �H H�D$L�pL��N�,�h�H M��t΃x
u�E�E��twL��H��L�D$����L�D$���D$,t3����    A�VI9�w:I;GsH�C�f%�?f=�?ufD�"@ L��H�T$,H��� ���I���D$,��u�I��E�E��u�H�D$L�@E�0E���4���@ L��H��L�D$����L�D$���D$,t;����    A�PI9�wLI;Gs!H�C��Ɓ��?  D9�u��@f��    L��H�T$,H��L�D$�c���L�D$I�ƋD$,��u�I��E�0E���s���I��M�������fD  A�0   f.�     L��H���������t��I;Gsf�C �I��I��:u�I���  �p���?  t:I�GH��~1H�<Cf.�     ���f���?f���?u	f% �	�f�H��H9�u�H�t$H������A�G    1������AWf��AVAUATUSH���3  H�GH�nL��$@  H�|$H��$1���  L���H��   H��$�   H��$@  �H�D��L��$�   H���   H���   ����H��(  H�|$H�7H�AP)�$�   )�$�   H�t$)�$�   H�pH��t9Pt*�oQ�oY(�P�oa8H�IHPH�pH�H@X `0H�@ L���   H��$�   H��$�   H��$�   ��$�   H��$�   L��$�   M���!	  �D$p    �$A�   I;E��  I�U�Bf%�?����I�L� L�y M����  I��@L��$�   L�,� �H I�EH���  D�D$ H��$�   L����D�D$ I�E0H��tD�D$ L��L����D�D$ ��A����  A����4$H��D��(  �J���A�ƅ���  ��$�   L�\$p�<  H�D$�P��$�   ����  H�l$H�����   ltuo�y  A�   IcwH�CXH+C@H�K`H�H+KHH��Hc�H��H��?H��0 �  H��H�H�D$`IcGH��H��H��?H�� �  H��H�H�D$h���$  H��$  H����  L��H���H���H�T$pH�t$xH��$�   H���H���H�H?H��$�   H�T$pH���H�t$xH��?H��$�   H)�H���H��$�   H�K0H��H�S@HT$`H)�H�CHHD$hH���H�����$�   H�K8H�C`H�CPH�SX��  H�S�B��  IcWH�Hǃ      Hǃ      H��H�H�� �  H��H�IcOHcShH�� ǃ�   ltuoH���H��H�CPH��H��?H��
 �  H��H�H�� H���H�ChHǄ$�       L��HǄ$�       HǄ$�       �����H���3  D��[]A\A]A^A_�D  fo�$�   fo�$�   fo�$�   AoAwA(�i����L��`�H L�\$pD�D$8L��H�L$0A�BL�T$(L�� �H I�E I�qH���   L�L$ H�|$@�G��D�t$pH��E���0���L�T$(L�L$ L�h@H�L$0D�D$8L�I�AH���^  H��H�T$(I�u ��H�T$(H�L$0��D�D$8L�L$ �D$p�0  I�A H��tD�D$(H��H�T$ ��D�D$(H�T$ H�|$@H��D�D$ ��E��D�t$pD�D$ E���7�������@ H���   �xp t�����H�D$�x! �����H���   �  �L��$�   H�D$X    H�D$@H���   L�D$0H�@PH�D$`    H�D$�@f�D$ A���  f�D$(���   ��H��H�D$H�����f���    L�D$0H�D$p   H�D$8H�D$x    HǄ$�       HǄ$�      ��  I��@H�� �H H�@(H����  L�D$0L��H�T$XH�t$`���|$(f9|$ H�L$XL�D$0uH���A  I;��  �4  H���   ���   L�D$0H��$�   ����H�|$H�t$8��HcWH�H��H�H�� �  H��Hc��ץ��L�D$0H�T$XH�|$ �  I���  ���WH���|$(I���  fA���  f9|$ ��  H�L$`H���   ���   L�D$ H��$�   �����H�t$8��Hc�H�D$H��Hc@ ��H��   H��H�H�� �  H��Hc��3���L�D$ H�T$`H�|$ �  H�t$HI���  ���WH��H��L�D$I���  H)�fA���  ����L�D$I���  H�l$@I���  L�D$I���  H���   H������L�D$L�\$pH��L��L�\$I���  H��$�   �=���L�\$����� H�D$L��L�\$�oH�o@ �oh0�$�   �$�   �$  )L$p)�$�   ����L�\$����  H�l$��$�   H�����   ltuo�������t&H��$  H��$  L�\$H���   �w���L�\$HcSPHc�$H  H��$P  H��$`  H��H��$  H��$   H��H��$0  H��?H�� �  H��H�H�f���    H��$(  �  M�E8M��t!L�\$L��H��L��<$A��H��$(  L�\$��$�   ��  Hc�$�  ���  ��$X  ��  H��$�  H�4�H�rL�iL�AH�TѨL�JH+BL��L)�J�4I��H�W�HL�H��H�VHL�H�O H�V H���H���H��$  H��$(  I9�M��~H��@H��$  I9�|H��~H��@H��$(  H)�H)�H��  ��$�   H��  �����H�Q I���B���@ H���N���H��$(  H+�$  �9���f�H�T$H��$�   H��D�D$ �f���A�ƅ��U���L��$�   D�D$ Hǅ�   �aD L���   �����    H��1�H��L�$�o���L�$�����fD  L��$�   H��L�$L���i���L��H�|$`�<���L�$���� H��$  H�P H�N H���H��$  H���H)�H��$(  H)�H��  H��  ��$�   �����    L��H��$  �����L�\$�	���fD  H��$  H��$h  H��$p  H�H�� H�H���H�� H��$  �u���f�     H�L$`H������I;��  �H��������L�\$p�:���fD  H��t[UH��SH��H��H���   H�D$H��tH�E 1�H��[]ÐH�t$�������u�Hǃ�   �aD H�D$H���   ��f�     �#   �f.�     SI���   �ȟH I��H��H����� ����   �ܟH �   L����� ������   ��H �   L����� ������   ���H �   L����� ����   ��H �   L����� ������   ��.H �   L����� ������   ��.H �   L����� ������   A�Q!��f�     A�QH��`�H �R�H��[�f�     H�;L��H�t$�p�����u�H�T$H�RH�SH��[�f�     A�Q�H��[�@ A�Q ���    H�;L��H�t$� �����u�H�T$�R�S��    A�Q$�A�Q(�SA�Q,�SA�Q0�SA�Q4�SA�Q8�SA�Q<�SA�Q@�S�=���@ �   �/���ff.�      AVH��AUATI�ԉʹ   UH���ܟH SH��0��À� �ۅ�u@��u\A�4$1�1ɸ��H �D  H��H��`�H H��t7�H9�u�x
u�U�*D  ��H �   H����À� �ۅ�u��t`�   H��0��[]A\A]A^�@ �   ���H H������� ��tO��H �   H����À� �ۅ�us����  A�$�E 릐A�$�EH��0��[]A\A]A^�f.�     �   ���x���I�<$H��H�t$�����Å��]���A�T$H�D$�P�K���fD  ��.H �   H����À� �ۅ��8  ����  L�l$M�u�
   H�t$L���"� A�E H�D$�8,�����L9������I��L�`M9�u�L��
   H�t$��� �ǉD$,H�D$� ������I9������L�d$A�$A�D$��������������A�L$A�t$���v������n���9��f���9��^���E�T$A���  �L���9��D���E�L$E�D$A���  A��A���  A��E��������  �����U$D�U(�E,D�M0�M4D�E8�u<�}@������    ��.H �   H����À� �ۅ�u8��uQA�$�E!�����1��
   L����� H��t'H��������E �����   ����A�|$������E  �|���1��
   L���� H���E!�a���ff.�     �AWAVAUATUSH�Ӻ   �H��HL�fH�FH�WhH�VPD�vHH�L$L�gXD�N,H�G`H�$H�V0D�t$L�#H�E����  �JA����  A��L�Bh��O��I��N��
�   �A�9�O�9�L�I��PM9�u�9���  Hc�Mc�Lc�H�T$I��M��L�T$ I��I��?N��
 �  M��I��I��?J�O�� �  M��I��I��I��H�L�I���I���L�OL�H?M�{ I���H�GL�OI��I���L9�L�_ LL�L9�M�Q LO�M)�L�W8M)�L�(L�O0L�G@I��@�0  H�W(M��A�   H�G0L�GHL�WPM��M)�M9���  L�HO�M9���  L�OPO�@M��M�SMI�I��M9�~L�WHM��O��M��M�SMI�I��M9�}L�WPM��L�\$Mc�H�\$0H��H�t$(L�\$8M9���   )�Hc�H�|$�    H�K I��H9�~I��I)�H��M�, �։�)�)�H9�L�I9��   D)�D�4H�t$I������H��G��M��I�4E�H��Hc�H�D$H��H��?H�� �  H��H��H)D$P�t$����XZL9{P|?H�H�CL�C@L��H��L)�H)�M9��O���H�s(I��H9��X���H)�I)�H���J����H�KXH�s`H�\$(��D)�Hc�H�D$H��H�H�� �  H�D$ H��H��H�H��(  H�H�� �  H��H�H��0  H�D$0H�H�D$8H�0H��H[]A\A]A^A_�f.�     D��)�D�4
�����f�L�OP�$����    L�H�����    L+O(L�WPL�OHI���   ~A�   �����E1�I��`A��N��   �����     AWI��H��AVL��AUATUSH���   H�T$H�L$�W����D$���U  A��  ��4  ��T  E1�I�XM��E��H�|$ E��tA����  H�D$ �	  A��E��u�u�H�|$��G0�  H�D$ �D$0    H�XHc H��H�\$8H�PH��H�,H�D$XH9��#  E1�D�d$(M���:�     L�i���CL�kH��tH�z( ��  M��LD�H��XH9���   �C�u�H�K(H�S0H��u�H��t�H�B(H��t�L�h�JI��L�jI��   A��  I�L$H+J�T$0�,���A�L$I�M�l$�@ 1�L���>�����tJ�D$�D$H���   []A\A]A^A_þ   L��������u�H�t$�   L��轡��A��  �}����H�t$1�L��衡��A��  ��^����D�d$(E1�E1�L�|$@H�\$8E1�D�L$4M��D��D�d$TI��D��H�D$H    ���D$P�AI��   A��  A���T$0H�KI+M�=���IED�sH�CL�T$(H��XL9���   D�sA��u�L�k0M����  @��tI�B?H;C��  I;E�z  I�}( L�T$(�z���I9���  �D$P��  H�|$@ ��  E1�1�L��H��L���g���H�D$H�K�   M�UH�\$@H��XA�ML9��_���fD  L��D�d$TD�L$4M��E����  H�D$XH=  ��H=   ���Ƅ���  ����  E���=  H�D$8�     �P��u#H�p8H��tH�H��H+NA��HN�PH�HH��XH9�w�E����  L�l$8M��L���D  H��XH9��c  H���Cu�H��XI9�w��@u	H��XI9�v�H���
@ �Au2H��XH9�w�I9�w�H�SH+PHPH�S�f��D$4�:���fD  I9���  H�CH+AHAH�C�r���f����   H�D$ �D$0   H�XHc H��H�\$8H�PH��H�,H�D$XH9��<����A��  ���H9�sl�    H�CHH�K����   H+K@ H�P@L�@H�fD  ��HJ f�2L9�tH�R@�2E��t��HJ(f�2L9�u�H�@H;CHu�H��XH9�r�L��D��L�\$(�Ӻ��L�\$(D��L���s���A��L�\$(��   H�D$I�s0A�{,H�HH�P�Z����/���D  H�@H;CHt�H�KH�P@L�@H��     ��H�J f�2L9�t�H�R@H�K�2E��t��H�J(f�2��D  L��H�T$`H�|$pL�\$(H�L$h�t���L�\$(L�D$hHc|$`IcC,I�S0H�4�H��H�H9�s1D  H�BH��PH��H��H��?H�� �  H��L�H�B�H9�w�A��  �=���M��H�D$ H�XHc H��H�PH�,�E���<���A��  ���9���D  D�D$0H�L$HL��H��L��������i��� I��   A��  A���   �T$0H�KI+M�����IED�sI��H�C����@ E�������H�D$ H�XHc H��H�PH�,�����H=  ��H=   @�Ƅ�u	@���F���H�\$8E1�f.�     H�D$8H�HX��u[H�D$8H���  L��  H���   H�GM�PI)�H��H+QM��I)�L)�IH�H9Y0��   E��t+H;l$8��������� H��H���   H��L��`  �f�H�D$ H�XHc H��H�PH�,����� ��0f9�u%H�@H�C������     I��H���Y���D  �;L�p��H�q)�)�Hc�L)�Hc�耎��I�L�s����@ H�GXH9G0�B���I�@0I�XXH9��1���H���'���H�WH�H+QH��I�PI�HH)�H��t*H)P@��tH�|$8H)��  H)��  A�H�H�����@��tH�D$8H)��  H)��  A�H����ff.�     f��;���ff.�     AWI��H��AVAUATUS��L��H���   H�T$8H�L$腢���D$����  A��  ���  ���  E1�M��tA����  A���J  I��M��u�A��  H�|$��W0��  �u�IcGXI�`�D$O E1��D$    H��I��H�|$@H�PH��I�H�D$PI9��R  �D$H    H�\$@L�t$XL�l$ M��M��D  D�cA����   H�k0H���4  H�}( �i  �EH��L�sE1�L�UI��   E�̈D$8A��  PM)�T$L��L�T$8�����M��ZYL�T$(D�\$0��  A���+  H�uH)�H�sA��D�c�MH;\$@vM�|$O H�CH�S��  H9�����t0H�C0H��t'H�@H)�H��H��?H1�H)�H����
  f�     H��XH;\$ ����M���D$HL�t$XM��M��L�l$ ����	�M���  ���o
  �T$Hi��	  L�H�BPHcRHH��H��H�H9�sKf�     H�xH��t0H�P@H�pHH�f�
H�z(H9�tfD  H�R@H�z(f�
H9�u�H��PH9�r��\$L����耴����L���&���A�������H�D$8I�w0A�,H�HH�P�����D$H���   []A\A]A^A_�@ H�D$1�L���h`�&������>  �D$���     H�D$�   L����(H  �������u�L�t$��L���   I��0H  蹚���   L���̸����u�I�F@H�@�DX@�����Ic�@
  I��H
  H�t$H��H�PH��H  H��H�D$H9�������FH�����Hc�������H��H�H�� �  H��Hcظ    H�� HN�H�D$(���I  �D$ ��H��H���J  �    �t$ ���N	  H�D$L�\$(E1�E1�H���I  � H��HH9��	  �A@�t��WA��A��A;�P
  ��D8�uE��t�H�7L�H��M��I)�L)�IH�Hc�H��I��I��?J��2 �  H��Hc�L9�}	I��E��I���G�{���H���r������j���L9���A8��[���H�AH��H)�H)�HH�Hc�H��H��H��?H�� �  H��H�L9��%���L�aI��E������fD  A��  �����Ii��	  E1��D$   M��I�t`IcDXH��I��H�t$@H��H�PH��H�D$PI�I��   H� �@H�� �H �@�D$OI9�w~����D  H���  H�}( t(�M����  ���H�E(    �MH�S(H��t3�C��H�R�CH�SH��H��   L���o����M M��LD�H��XL9���  �C�u�H�S(H�k0H���s���H��t�H�E(H��t�H�S(H�@�MH�EH��u�H��H���H�D$1ɉ�L��H�Ph諗��1�L��������������A��  ����������D  �t$H��H��L�������K�E���D  L��M+wMwH��L�H��_�  H�J �    �&   A�   H���H��AHL�LL�H��H)�H��I��H��I)�H)�IH�L�I��I)�H)�IH�H9�H��HM�H��?H�H��H��H��H��H�H)�H�KH�E�H����     �D$H����fD  H��@��  H��_��  I�� I���L�sA���t$H��H��D�cL��I��������N���fD  ��  H�R���CH�S�5���D  H9��������D  M�F H��H��I��H��I���I�4H)�H)�HH�K�| H���I��I)�L�I)�H)�IH�H9�}I�< M��L�KH�}�a����M��   �     H�D$PH=  ��  H=   ��  ���k  L;l$@��  L�d$@�l$OL�� �rH�ZX@���  H�K�H���)  H�{�H�AI��I)�H)�IH�H��O�
  LAL�C�I�Ѓ�@�s�M9�sKH�C�H��`���@����  H9�����t-H�C�H��t$H�@H)�H��H��?H1�H)�H��~
H�S�fD  I9��  �T$Hi��	  L�H�BPHcRHH��H��H�M�������H9��F���@ H�xH��t0H�P@H�pHH�f�
H�z H9�tfD  H�R@H�z f�
H9�u�H��PH9�r������f�     I9��p���H�������    M����   H�C�I��L�C�H�� H���H�C������ L�C�I9��"  I9��  I9��  I9��  H�QH�xL�HH9���  L�K���@�s�M9�������    �C�g���H�C�H�S@���M  H9������H���H�C�H���;���H�@H+�`���H��H��?H1�H)�H������H�S������    H9����4���D  H��P���I9�w#��h���t�f�     �@u	H��XI9�v�I9�v'H���Ct�����fD  �A�����H��XI9�w�L�C�H�C�I+CH��H���ICH�C�����@ �    �    L��H��I�I�N H���H��H)�H��I��L��M)�H)�IH�H�H��L)�I)�LH�L9�HM�H��H��?H�H��H)�H�H�SH�E�����D  H9�������D  M�������     IcWHI�GPH��H��H��k����     H�|$P  �1  H�D$@H�xXL���  H��  I�HH�^H)�H��H+GI��I)�H)�IH�H������I�@H�NH�H+G�~H)�H�FH�F0��H����  H)HH�|$P   uH�\$@H)��  H)��  @�~�H������     L;l$@���������H�S�7����    ���H�C(    �CH�E(�W���f�     H�C�H�qH)�L�\$0L�D$(H)�L)�L�L$ H���Ȁ��L�L$ �s�L�D$(L�\$0I�L�K��
���f�     H�|$@L���   H��`  ������     M��tL�g(E��t�OH��XH9|$����������f.�     H�T$`L��H�|$pH�L$h�����IcG,I�W0L�D$hHc|$`H�4�H��H�H9������ H�BH��PH��H��H��?H�� �  H��L�H�B�H9�w�����H�|$P   uH�D$@H)��  H)��  @�~�E����T$Hi��	  L�H�BPHcRHH��H��H������   �&   ����� 1��ff.�     f�H��H���   �   H�T$�v���H��ÐH���   ���@ ATI��UH��S�< u�    H���< t���H�_H��v"H���   ��   �W��H�_H����?H	�E1��f�     H�{D����x4H�����u�M����   H�E     H��[A�$    ]A\�f�     I���   vWI���   I����   A��A�   E��H��I�H��L��D�A�H��A��?I	�L9�u�A�B�H�\�y���f.�     D���H��H��A��?I	��T���D  H���   H��vs��A�   D��H�D  �GH��H����?H	�H9�u�A�@�H�\����� H�F@H��H�8�y�����H�E H��[A�$   ]A\� A��A�   �$�����A�   �fD  AW1���  AVI��AUATUH��SH��X�  L���   �E`    �   L�l$H��$�2  ǅ�8      L���H�H�E L��L�D$�@H�� �H H�X �B���I���    �����  < uf�     H���; t�H��H��$�2  L��H��������$�2  H��w�M�<$M��t�I���   L�������   D��L���,������l  I���   f���    �W  1�H��$�2  ��p  蠽 �EHL��H���   HǄ$�2     ��$�2  H��$�2  HǄ$�2     L��$�2  H��$0  Ǆ$(      ��������   L�uhM��1ۉ�L���D$    �d�������   1�L���1��.���IcT$HI�D$PH�<�H��H�H9�sGLc�D�D$E1�Mi�88  f�H�P H��tH9B @��H9���@ ��+  H��PH9�w�E��tD�D$���QL��H�|$I��88  ����$�2  I���	  ��聆���D$A��������t�   �1���I���   L���x���U`����   �EHH��H��H��
H��H���  H�gfffffffH��H��ƅ�   H��?H��H)��8  H���  ��ud�EHH��H��H��
H��H��(:  L��H�gfffffffH��H��ƅ0:   H��?H��H)�H�� :  �ٲ��H��X�  []A\A]A^A_�H�Mh�`���H���8  ��R�p)�Hc�I��I�ۅ�IH�A�������D��A��A��H�4vI�4�H�T5h����fD  AWAVI��AUATUSH��x  H�H���   L��$�  H�t$�   �XL������I�ǋ݀�H H�,݀�H =)  ��  �     H��@�H �EI�FP�D$    I���8  �D$    A�   HD�H�D$ ���u�d  @ H���< t�<|��  H��H�L$,L��L���"����|$,H��w�I�7H��t�H�|$�   �����H�|$H���   f���   ~���u����   f����  H���   ��D�d$1�L���   �����L�FI�<@1�I��D  �6�~9�}JD�UE��A��A����   Hc�H��L�fE��t8�     L���xL9�}��L�у�H��9�u�Hc�L��M9�t0I��� L���xL9�~��L�у�H��9�u�Hc�L��M9�u�D�d$E���p  �D$H�L�0�@�D$���������    �|$��D$��   H���E =)  �6���H�D$L��H���   �2��H��x  []A\A]A^A_�H��E1��<���@ fE��t:f.�     H��H��I�|9��xH9�}��H��H��9�}ލ~����fD  H��H��I�|9��xH9�~��H��H��9�}ލ~�������v]�D$H�|$0A�   E1�I��D�X�I��@ L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��M9�u�H�D$�|$D���  A�[�'  �D$M��   E1�D�P�I��f�H��I�HL��L)���H��H�H9�~H��H�P�H�L9�u�H��I��I��I9�u�H�D$���  �D$�L$J��    L)�H�|$��H����  ����   H��H��H���  H���  �U��H9�t?@��@��f9�t2H�H�|$H��H��?H�J��    L)�H��H��H���  H���  J��    H�|$L)�f��uoǄ��      ������D$H����  �@�D$�*���H�|$�t$���  ���"����D$��H�L�0J��    L)�H��H���  H���  H���1���Ǆ��     �S���H�4׋T$H���  ��H�L�0H���  �����1������f�AWH��AVE1�AUE1�ATUH��SH��Hfo: H�8H�t$H�T$�   H�\$ H�D$    )D$ �D$08 9 ����I��f�     �; t\H��H�L$L��H�������|$H��w�H�E@M�<$H�L$�  H�8D���!���M��t�H�D$E��tI9�u5�; I��A�   u��   H�D$L��H�8����]8H��H[]A\A]A^A_�1���@ ATUH��S���   H��L���   �cinu�GHH���������tL��H���y���[1�]A\�f�H��H���u���H��H�������H���   H��������f�     ATUH��S���   H��L���   �cinu�GHH��舔����t$Hǃ�       L��H�������[1�]A\��    H��H�������H���   H���6�����@ AW1���  AVI��AUATUH��SH��x�  L���   �E`    �   L�l$H��$�2  ǅ(H      L���H�H�E L��L�D$�@H�� �H H�X �"���I���    �����  < uf�     H���; t�H��H��$�2  L��H��������$�2  H��w�M�<$M��t�I���   L�������   D��L���������l  I���   f���    �W  1�H��$�2  ���  耳 �EHL��H���   HǄ$�2     ��$�2  H��$�2  HǄ$�2     L��$�2  H��$0  Ǆ$(      ���������   L�uhM��1ۉ�L���D$    �D�������   1�L���1�����IcT$HI�D$PH�<�H��H�H9�sGLc�D�D$E1�Mi��G  f�H�P H��tH9B @��H9���@ ��+  H��PH9�w�E��tD�D$���QL��H�|$I���G  ����$�2  I���	  ���a|���D$A��0�����t�   �1���I���   L���X���U`����   �EHH��H��H��
H��H���  H�gfffffffH��H��ƅ�   H��?H��H)�(H  H���  ��ud�EHH��H��H��
H��H���I  L��H�gfffffffH��H��ƅ�I   H��?H��H)�H���I  蹨��H��x�  []A\A]A^A_�H�Mh�`���H��0H  ��R�p)�Hc�I��I�ۅ�IH�A�������D��A��A��H�4vI�4�H�T5h����fD  AW��$I�AVAUATUSH��8  H�H�|$ �XH�t$H�݀�H H�D$(�GHH���   �   �$���������H��$�  H�D$x�����H�$�݀�H =)  ��  fD  �D$p    H��@�H 1�E1��D$T    I��I��L�� A����|  < u�     I��A�; t�H�$H�t$ L��H��$�   �������$�   I�Å�t�H�D$(�D$S L�\$8�@f�D$��f��H�E1�H�D$�D$H�D$H�D$   ���A��D9�$�   ��  H�$H�0H��t�L�t$�   L���0���I���   f���   ~���u�H�D$(���   �pf�t$Pf����  H���   ����E1��D$    L���   1�A������D$    L�HH�l$0M�4Q���    �0D9�~]Ic�D��f��ty� H9�|"I9�LO�H��9�|(H��A��H��I�T��y�H9�H��D��HL�H��9�}�D9�t�t$A��D�\$D�^L��M9�tGI��뉐H9�"H9�HL�H��9�|�H��A��H��I�T��y�I9�H��D��LO���f.�     H�l$01�E����  �D$P��  H;|$�z����D$SA��H�|$D9�$�   �q����    H�|$L�\$8H��   ������H�����������|$S ��  �D$pH��Đ  �@�D$pA��������f.�     I�܋D$p�\$TL��	��  H�D$(H�D$(� =)  �"���H�D$H�4$H���   ����H�D$ ���I  ���?  H�D$ D�e�L��$�   I��L��H�I  K�LH�H��H��HH9�u�L��A�   E1�����  H�KM��E��H��M)�D�I@A���+�     H�:E��t-H�1H9�~.J��H�P�H�I9�tH��H��B@u�H�zE��u�H�qH9��A��D9��H  I��I��H����    H;|$������V���Ic¹����H�\$HD��L���   H��L�l$@H��D�d$X�l$A�I�D�|$��H�T$0I��<ADʉ�A���fD  A9�tq��9��N�AM�Lc�L��H��L�H�BH)�I��I��?L1�L)�H��~$H�H��H��L)�I��I��?L1�L)�H9��  C���<u���E��y�A��A9�u�L�l$@�\$@H�\$HD�d$HD�d$XL�l$`E��D�l$�L$hD�|$D�d$t�L$@H�\$XD�d$H��    A9�tpA��E9�A�sAN�Hc�I��I��M�I�AH)�H�H1�H)�H��~&I�H+T$0H��H��H��H��?H1�H)�H9��7  A���<u�A���y���A9�u�H�\$XL�l$`�L$@D�d$HHcL$hD�d$t�D$Pt_H�D$ ���QD�XHD����Hc�H��I� ��A��Hc�H��L�|$XI+H�H1�H)�I9�~���T$+T$)ȃ�9��5  �    HcD$@��x+HcT$H��x"H��H��I�I+ H��H�H1�H)�H;D$xBA���<t'�   �D$P������k���H��8  []A\A]A^A_�Hc�A�6��<u�1������D$TH�L$H����   �@�D$T�����L$@H�\$XD��L�l$`HcL$hD�d$HD�d$t�����L�l$@��\$@H�\$HD�d$HD�d$X�����1�1��I�����vh�D$pL��$�  �   E1�D�P�I���     H��I�HL��L)���H��H�H9�~H��$�  H��H�P�H�H9�u�H��I��I��I9�u�H�D$ �|$TD���I  E�k�V  �D$TH��$�   A�   E1�I���X�H��f�L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��L9�u�H�D$ D���I  �D$T�L$pH�\$ ��H����   K�ۅ��  H��H��H���I  H���I  H�D$(�@H9�t:@�Ǩ@��@8�t+H�H�\$ H��H��?H�K��H��H��H���I  H���I  1�H�\$ �K����H���L���I  H�� J  ��J  �tK�ۃ��J  �tH�\$ K�ۃ��J  ��'���H�\$ K�ۃ��J  ����H�\$ �t$TD���I  ��������D$p��H��Đ  K��H��H���I  H��H���I  ����H�4ËD$pH���I  ��H��Đ  H���I  �����D�Ћl$L�|$0�L$`�L$�	A9��s����P�9���M�Hc�H��I�L9�t�HcL$`A9��K���H;T$0��L��$�   �D$tA��A��D�؉�$�   �t$H�D$h1�D��$�   D�d$�D$`    �D$0    L��$�   H��$�   �   Lc�M��I��M�I�BI�L)�I��I��?L1�L)�L�H��L)�I��I��?L1�L)�H��~L��I��I9���   G�>A��A����   L9�A��D:T$tuH9T$X�  �   9�tgIcՄ�u&Hc�A���<��   �D$`����A���D$0����A9�EN�H��L�L�J��H��L)�I��I��?L1�L)�H;D$h����1�9�u�H��$�   L��$�   ��$�   D��$�   ����D�T$0�l$`E���A����l$0�8����l$`A��l$0�w���M��"H�HH�PI�@�@@t2H�@H9�~H�I��M9�����I� �@@u�H��H�I�@�@@u�H� ��L�L$XH��L��$�   D�T$`�T$0D�l$hH�<�    H��$�   L��$�   D��$�   9l$�END$Hc�H��H��H��I�D H+D$XI��I��?L1�L)�H��~I�L)�I��I��?L1�L)�H9�~1A�6��<u��H�A��9�u��L$H��H�|$X�T$@HcL$h������T$@D�T$H9t$}�v�HcL$hH�|$X������t$HcL$hH�|$X����ff.�     f�AWAVAUATUH��SH��H��HH���   H�D$���   �cinu�GHH���ك����t%H�t$H���X���H��H1�[]A\A]A^A_��    H��H��L�|$ E1��]���H��H������H�T$�   fo�' H���   �D$08 9 H�D$    )D$ ����H�$    I�� A�? t_L��H�L$L��H���'����|$I��w�H�E@M�4$H�L$�  H�8D�������M��t�H�D$E��tH9$u3A�? H�$A�   u�A�   H���   L���F��D�m8�����D  E1��� USL��H��H�.H��tH�G@�  ��H�8�L���H��tH�    H��H��[]�fD  D�A9�vx��H�vH��HG�P��ubD�G��USH�_�PH�@     E��t,D�D�PA�P�H�l�H��E�H�2�D9�-NA9�%H�p E9�vA�P�WJ��[]�fD  ��    H��H9�u���ff.�     f���Hi��  H�7�B����   L�D7Lc��  IcI��H��H��?H��
 �  H��Hc�H�Q I�HH���I�PI�P��tg��H�@M�T�0��     I�HHcH��I��H��H��?H��0 �  H��H�H��H)�H)�HH�H��HN�H��H�B�H�� H���H�B�L9�u��ff.�      AWI��AVAUATUL��SH��H9��  u	H9��  tI���  L��1�I���  �����I9�(  uI9�0  ��  I��(  L�߾   I��0  �����I��8  H���I��  H��H��H)�H��I��X  H��H9���A��`  A��l  ��~PLc�Hc�I��H��H��?H�� �  H���� ~.L)�L���! H��I��H)�H��?I�� �  H���� ~��u�A��d  1�Hc�M��@  M��P  M��H	  @ �H�G����   ��H�RH��H�|8f.�     HcPH��0H��I��I��?J��" �  H��Hc�H�H�P�HcP�H��I��I��?J��" �  Lc`�H��Hc�L��H�H�P�HcP�M��H��I��?I��I��?J��2 �  H��Hc�H�P�K��, �  H��Hc�H�T H���H�P�H9��\�������tlL�׃�� �����L��ID�����f�     []A\A]A^A_�D  I��X  H���S㥛� H��    H��H��?H��H��H)�H9����<��� 1�Hc�M��P  M��H	  D�P����   A��@  L��I��H  ����   D���H�_H�t@A�@�H��H�@H�H��H�l8f�     E��tD�	D��+GH�I��I��?L1�L)�H�H��I��I��?J��0 �  I��H����?=�   D  D��A+H�I��I��?L1�L)�H�H��I��I��?J��8 �  H����?~MI��0I9�u�H��0H9��o���A�������D��D�P������A��8  L��I��@  �������� I�F(H��0H�A�I�F H�A�I�FH�A�I�FH�A�H9������f�     H���   ��     H���   ��     H���   ��     �G    �G   �G    �G(    �G8    �GH    �GX    �Gh    ��    �G    �G   �G    �G(    �G8    �GH    �GX    �Gh    ��    L�GH�G     H��H�wHǇ�       H�(��H���)����   1����H�L�BHǂ�   ��D Hǂ�   @�D Hǂ�   @�D Hǂ�   @�D Hǂ�   0�D Hǂ�    �D Hǂ�   ��D Hǂ�   P�D Hǂ�   ��D H���   Hǂ�   ��D Hǂ�   0�D Hǂ�   `�D Hǂ   @E Hǂ  �E Hǂ  ��D H���   �UH��SH��H��H�w(H�������H�C(    H�sH���C     H�C0    �����H�C    H�sH�������H�    H�C    H�C    H��[]� AUI��ATUH��SH���GH�_��tK��H�D@L�$�f�     H�sH��H���`���H�C�    �C�    �C�    �C�    L9�u�I�]H��H���/���I�E     I�E    H��[]A\A]�@ D�H�GE��t(A�K�H�LIH��H�@ �`�H��0�@�����H9�u����   �F�UE1�1�SH�\@H�O1�H��1��H�    A����E��t.L�WI�E�BA��uA��E�BA9�vA���N��fD  H��0H9�t��u�D�
�@   H��A��   �fD  �o��~pI�ɍ]�I������E1��     I�qI��>;:/J��    O��D  H�T�H��9:|H�TI�t H��u�I�BI��I��I9�tI���fD  []��G    �ff.�     f����`  A�   AWA��Mc�AV��   AUE��ATUSD��D�AD�A�݉D$��A�H�D�	�\$�L�$G�L�T��WfD  E9���  D�Z!E9�tTE��t	E9��o  ��@t"�L$���   �L$���   H�z( ��   H��HL9�t`�J��u�D�Z H�B0E9�u�I���u���     I��M9�t�I�+I��Hc] I)�M9�}�H)�L9�}݁�  H�j(H��H�J�L9�u�[]A\A]A^A_�@ ��t�I��I�+I��Hc] I)�M9�}H)�L9��  I��M9�u�H�z( �N���I���f�     I��M9��3���I�Hc+H��H9�|�KHc�H9��H�Z(�����������I��D  I�+I��Hc] I)�Hc]M��I)�M9�}L)�L9���   I��M9�u�H�z( ������q����    �������I��� I��M9������I�+I��Hc] I)�Hc]M��I)�M9�}�L)�L9�}ρ�  H�j(�J�e���D  ��  H�j(�J�N���fD  ��������;��� ��    ��  H�j(�J����ff.�      AWI��1�AVI�΍6AUI��ATM��E1�U���   SH��L��H��(L�L$����H�C�D$��tH��([]A\A]A^A_�@ ��L�L$E1�1�H���0   L��H�$�����H�C�D$��u��    A�ML�L$1�E1�L�������t$H�C(����u�H�SH�<$�+�C    I�H���C     H�SH�SH�C0    ���  �E�H�t@H��H�D  �H��0H���BЋA��BԋA��B�H9�u�M����   A�M�~L�s8����   ��H�D@I��H�D$D  E�7M�o1�E1�1�E��u�I ������u$A��E9�t5��u�A�U ��   I���@   ��t�D��H��A���$�����$E9�u�I��L;|$u��+;kt8��tE1�D��H��A���q���A9�u�D$H��([]A\A]A^A_�f�     �t$���J���D  M���<���A�M�~L�s8���������"���ff.�     f�AUI��ATUSH��H����WL�G�i9�r0��H�@I�T��1��    �B    �+I�U H��[]A\A]�D  D�aH��L�L$�   A����D$    D������1�I��H�C�D$��u�D�c�@ D�GE����   ATU��SH��H���t�   �CH��[]A\��    �G(L�'��tH�O0H�@H���p�H�{(H�T$L��������u��CX��tH�S`H�@H�h�H�{XH�T$L���������u�H��[]A\�fD  �ff.�     @ AT��U��SH����D$    D�@1�A��A9�r	H��[]A\ÍZH��D��L����I��H���   ��L�L$H������I�$�D$��u����] H��[]A\�ff.�     �ATUH��S��97v#�؉ٺ�   ����HE��1�[]A\�D  D�fH��H�wD��H��9�����u�D�e �ff.�     @ AWI��E1�AVM��AUI��ATA��U��SH��8����   M��tA�����A�M M�E���N  L��1��fD  ��H��9�tE9*u�D9bu�A�E��tdH�@I�EH�|��L�ډ�������uM��tA�H��8[]A\A]A^A_Ð��A�ED�yA9�sqD��E�} H�@I�D��(D�`D�PA�E��u�I�}L��H�T$(L�\$�����H�|$(L�\$��t�H��8[]A\A]A^A_�@ ���tsA�   E1�����D  �D$(    v�����L�L$(�   ���L��D�T$�L$L�\$����I��I�E�D$(���+����L$D�T$L�\$A�M�3���@ ��A�   E1�����1��
����     AU�   ATI��U�j�SH��H����E�H��H����H�H�vH��L�lf�     I�$�SE1�L��3������uH��H9�u�H��[]A\A]�@ A�D$H��[]A\A]�ATA��UH��SH��H��H�:�'O��H�{H��H�$�O��H��H�D$�E��uH��   D��H���3���H��[]A\�f.�     AWAVAUATUSH��  H�<$�t$����   A��H��E1�fD  A��A�   EN�E1�C�\6��\$�@ I��N|� L���N��H��J�D�I�D$L9�u�D�d$H�D$A��I��J�L$(�    H�P�H)H��H9�u�H�$�P��u�t$H�L$D��H���a���E)�E���e���H��  []A\A]A^A_� H��H��tHH�?�F    ǆ�      ǆ8      ǆ@      ǆH	      ǆP      �7����    �ff.�     @ �D�P�E���o  AWIc�AVI��AUATL�$@UI����   S��   H��8H�t$fD  M�^E�j�D��K�#I��L�HD� K�#f�D9D��F
H�B����  A�1@�0uiL���@ D�>D�8uW��H��H����w��t�6@"0@�Ɖ������х�u-��H�����u�E��E���m���1�H��8[]A\A]A^A_�@ D��A��9�wsӉ�E���    E9>v�D��H�RM��E�E��tKH�@M��E�E9���   I�SA��I�pA��t%A�y�1��f.�     H���H�HH9�u�A�     A�@    A�����D)�A����~[��E�HI�HI�pH�@L��Mc�H��D�L$H�L$��� D�L$H�L$I��K�I���     D�HH�H�@    A���A�E��E���R��������D  L������H�L$I�sI�{D��D�T$,L�D$ L�\$D�L$�7����������L�\$L�D$ D�L$D�T$,I�S�    E9vD�щ�D�Ѓ��������� I�SA��E9�u�����1��ff.�     @ �G��t	��     ATUS�G(L�'��tH�O0H�@H���p���H��H�8L���2�����u.�CX��tH�S`H�@H�h�H�{hL��[]A\�����     []A\�ff.�     AVAUATU�)SA�����   ��A�����L�t��   fD  D�D�
D�Z��   D��I�p��E1�D)߅�u�   fD  ��   H��0��tZD9~�D�H�M��O�II��I���     A�����AoI��0H�@H��H� �AoI@H�AoQPP D��E��u�D��~E��tL��H��1�I9��J����)A�[]A\A]A^�@ D��H�qD)υ�t@��E��A�   �Y���E�XA�xf���� �F��x9�}��~��     9�~���D�I�y념AVM��AUA��ATUS�D$0D�˅���  L��  H��	  A�$    L��I��1��E     �i���D��L��   �Y���E�$�u I�L$E��tME��H���D�XԉP�D�H�A����xH��0A��vD�E��A)�A9�|�D�:��fD  �P���P�E��t�H�}��tJA��H���# E��D+A9�~D�X�D��D�D�@؉P�A��D� �PH��0A��w�D�D�@؉P�E��t�A�   E��uA��H��A����   A�   E��t�)Y�QA����   A�B�L�T@I��I����H��0�A�A؋QL9�t2D�I<E��A)�D����D���9�|ӍA)�H��0�A�D�I�QL9�u΍H��A�BA��A���u���[]A\A]A^�f.�     I��H��  �\����I����ff.�     AWAVAUI��ATUH���p  SH��H��(H�T$蚫��I�ċD$���A  ���   M�,$I��$�  A��$�  ���   H���   ��t!�O�H��M�    �H��H���J�H9�u����   ��I�T$(A��$�  A�D$���   H���   ��t"�O�H��M�   @ �H��H���J�H9�u�H����L�UD�M|A�|$L�}(�M	L��j �uM��L�mXI��$8  L�u<H��L�T$H�D$����H�D$M��L���M�u
�$   D�M|H�������D�EXH�MZ1Ҿ   L�T$E��t����fA+zf9�L���H��A9�w�D�E	E��t&H�M*1�@ ���fA+f9�L���H��A9�w�D�E
E��t&H�M>1�@ ���fA+~f9�L���H��A9�w�D�EE��t'H�MZ1�@ ���fA+D} f9�L���H��A9�w�H����  �eF��H9EpHNEpI��$X  �ExA��$`  �E|IǄ$�      IǄ$�      IǄ$(      IǄ$0      A��$h  �D$L�#H��([]A\A]A^A_��     �G��  AWAVAUI��ATI��USH��H��8HcHc�Hi��  H�|$I��L�Lc��  I��H��H��?H��9 �  H��Hc�H��  H�L$HcK�L$(I��H��H��?H��1 �  H��Hc����  A���    ��  A���    �k  H�k�D$   H�D$     L�{ M��t\A�G��  �T$(��A�A�W��AA)�I�WMc�M��H��IWH��L��H��?I��6 �  H��Hc�H�H��H��H)�H�T$A���    twH��@�M  HiT$�  H��I�TH��H)�H)�HH�H��'�6   H��/~>H��H���   ��  H���?H��	~"H��H���@�� ��  H��5H�i6�    L�\$H�kI�K I�T+ H���H���H��L)�L)�H)�H��I��H��?I��?H1�H)�L��H1�L�L)�H9�HO�E1�H�K�T$��tYH�SH�KH��?�B  H�� H��H���A����  A��t,A����  H�sH��H��@�9  H�� H���H)�H�K���CH��8[]A\A]A^A_�fD  ����  A���    ��  A���    ��  H�k�D$   �|$(E��$8  I��$@  A�8A��$l  �|$,E��tpE��$h  ��A+�$L  E��A��A9�SE��$H  E�D9��,  A�y�H�<H��M��<p  � fD  ��+~D9�|D�NE�D9���  H��0L9�u�H�D$     E1�A��$@  I��H�IH��I��  E��tlE��$h  �OE��D)�A��A9�S�wD)�A9���  A��I��J��    I)�I��I��D  �OD)�A9��wD)�A9���  H��0L9�u�1�A���	  A����   H�T$ H�sH)�H�S�����f.�     ��    H�k�D$    �����    H�T$��H�k�CH�SH��8[]A\A]A^A_�fD  A����   A�������A����   H�C@   �    H�� H���H�� �����@ H�k�D$    � ����    L��L��L���B����CD��D$(�C����A�������H�T$ H)�H�S����D  H�s�����    �@   H�T$ H�sH)�H�S�C���fD  �@   H�s�/���f�D�L$,E��uA9�$d  �����H�~A�   H�|$ �����@ �t$,��u1�A9�$d  �e���A��H�w�X��� H��~"H�T$H��H�@   H���H�T$�����@ L�t$I�V H���H��~@I�4.M��H��H�N I)�H���L)�IH�I��I��I)�I)�L��IH�H9�HN�H�L$����H�T$����H�� H�������H�i
����ff.�      AW1�I��E1�AVAUATUSH���  H�H�|$8H��$�   L�L$p�L$@�   �H�H�NH�T$ �H   1�H��H�\$0H��$  ����H��$�   �D$p�D$��tlH��$  H��$h  H������H��$   H���t���H��$�   H���t���H��$   H��HǄ$�       �X����D$H���  []A\A]A^A_�f�I�H��L�L$pE1�1Ҿ   �E����|$pH��$   �|$���a���E�GA�?L��$�   D��$�   ��$�   ����   I�W�O�L�JI�I1��f�H��L�ʉ�L9�t|I���2����)�H��M�̉PL�tԉ�I�BH��I�L̸I�
���`  ��H�T�	M��L��f.�     H�JHH�I�H�RHH��H�AL9�u�M�SH��L�ʉ�L9�u�I�GL��1�E���I  L�d$I����   �    D�[D�߃��|$H��Hc�L�H��L�iL�L�1L��H+rL��H+:I��H��I��?H��?L��I��H1�I1�L)�I)�L�II��M9��\  ���D�BH�D�C H��L�H�H�HL)�L)�H��I��H��?I��?I��I1�I)�L��H1�L)�L�@I��M9���   H����  �D$�C!����   A����   �    ��$�   ��H��H9���   H�|$H���H�9��8��8�H�CH)�H)�H��H��H��H��I�w�������C   A�   �D$   �����@ D�l$�C!E��u"A���x����D�����k���D�[�    A��D�[�S��� O�II��L9�~�H����  D�t$�C!E��u�A���"�����K�@A�   H��H9������A��E�B�����@ H�D$ L��$  I�W��$�   H��$  H��$�   ��t?�q�H��H��H�fD  H�
H��H��H�@�    H�@�    H�H�H�J�H�H�H9�u��D$    ��u�  @ �D$�D$;�$�   �r  �D$H��H�$   �xv�L�L��fD  H�[I9�t�H�k0I+i0L�s8H��M+q8L	�t�H�l$L��H�\$L���D  L��L�e L9�t�L�m0M+l$0L�}8L��M+|$8L	�t�H�|$L��L��L����B����t�M��M��H�\$�D$(H�l$HL��H�l$L�l$f.�     E1�H�C0H�K8I��I��E���f.�     H�U0H�E8H��I��H��I�n�   H9l$DD�H�U0I��I)�H�E8L��H��H)�H	�t�H�t$H��L��L���>B����t��|$(M��E��I��L��1���
  H�\$HL��H��L�d$�D$(E���U����x���H�D$8L�D$0H��$   �pH�H(H�P ������D$�D$p���R���H�D$8L�D$0H��$h  �pHH�HXH�PP�����D$���$���H��$  H�D$ H��(  Hc�@  L���  Hc�H�|$`H��L�t$XH�H�� �  H��Hc�H�u H���I���s  H9��j  H���*8��L��H��L9���  H��H��$  E1�1�������D$WH��$  �|$@A�  �D$    fD��$�  �G�����$�  ���H��$   H�D$H�D$ ��$�  ����$�  HH  H�D$hH��$  D��$�   L��$�   D��$�   H�PE����
  A�y�L��D�\$H��H��H���    H��H�H0H��HH�p�H9�t0H�rH�
�@    H�@(    E��t�H��H�p0H��HH�H�H9�u�E��t#H��$   E1ۋ}����  A��H��E9�r�E1�E9�s$D��H��I�z@��@�   A��E9�r�H�|$�H�o��t?��D�l$L�d@I��I�@ H��D��H��H��0H��$�   �f���L9�u�H��$  H�D$�    H�@8L�`D�8HcD$H�D$(D�hHi��  H���  �7���   D��$�   H��$�   ��OǉD$0A���y  E����  A�G�E9t$D��AFL$H�@D�l$8I�l$L�|$I�D�0��I����    H��D��L9��4  D9uE��DFeA9�v�E��u L��A)�H��H��H�U����I�wA�D��D�L$8D�D$0H�������D��$�   H��$�   � H�U H����    H�r0H9p0uH� H9�u��q����L�`L��H��fD  H�RI9��#���H�r0H�O0H9�t�H;H0~H9�|H�H���� H9�~� �O@H�H9�t��O@H�H9�u���@ �D$W �����fD  H��� H�p8H�J8H9��  H� H9�u������f��  E���  A�F�I��H�D�	H��H��fD  H�x( t�P��u���PH��HH9�u�HiD$(�  H�$  �|$L���  ��  K�D�	Mc�H�,��$f�     LiL�k@�� �CH��HH9���   H�K(H��t�CL�i��u���u�HcH�{0H)�H����  HcQH�qH9���  )�L�Hc�I��H��H��?H��
 �  H��Hc�H�H�S@�L��H��?L�t$XH�ףp=
ףH��L�H��H)�L��F����H��$  H��$�   HiD$(�  L���  ��$�   H��L�$�L9���  H��1�f��P�������H��HI9�w����  L��$  H�l$p���=  H��E1��D  H��HI9�vM�At�D��H�D� H9�s*H�P�H�q0H9r0�@ H�P�H;r0}H�H��H9�r�H�H��HA��I9�w�A�F�I��H�D� H�D$0�<�    �S ��t:S!uH�   @   H�{��  fD  H��HI9���   D�CD����u�C�u�L�M H�{0I�A0E���,  H9��#  H�E�@ H�0H��H9~0
�эQD9�u�H�D$0H�0D��L�V0I9�}�N  �p�H��H�t� L�V0I9��1  �Ѕ�u��H�L� H�A0H9��F  I�Q0I�q@H9��>  H�s@��  @ H�D$pH9�tH��L������HiD$(�  H��$  L���  HiD$(�  L��$   L���  ��$�   ��t~D�P�Mc�I��I��M�@ A�GI�H��H�4�H9�sKH��1�1�D  �@ t
H��HD؃�H��HH9�w�I�܃�w��  f��A ��   I��I�L$H9�u�I��M9�u�H��$  ��$�   H��$�   D�\$L�HL�P1���u0�  �L���tL׹    �7	�H��H��;�$�   ��  �ǋJL�B@H��H����L�E��t�L�F��t�L׹@   �7�fD  H��D  H�m�E t�I�t$0L�E0L�]@I�|$@L9���   L)�L)�I��H��H��L��L�T$HL�L$@L�\$8L�D$0H�T$(�0��L�\$8L�D$0I�L$L�T$HL�L$@H�T$(L��L��H�L�:�<�    L9�|{D)�Hc�I��I��I��?J�� �  H��Hc�L�H�Q@H�IH9�t9H�Q0H)�H���Hc�I��I��I��?J�� �  H��Hc�H�H�Q@H�IH9�u�I��H9��S����X����Hc�H����    L��H)�I)�M����  �   �E���@ u.HcC0L�K@I��H��H��?H�� �  H��H�I)�f.�     H9�t$HcB0I��H��H��?H�� �  H��H�L�H�B@H��HH9�w������f�     �|$W ��   H�D$H�|$�����H��$  �D$   �����    L�t$H A�NM�vL9�u�K����f�     Hc�I��H��H��?H�� �  H��Hc�I�L�k@�����)�Ic�Hc�H��H��H��?H�� �  H��H�IA@H�C@A�� D�C�i��������C�}���H�T$`H�t$XE1�1�H��$  �I�������D�l$8L�|$I�G8L��H�@H�P�0����I�wA�D��D�D$0H��E�������D��$�   H��$�   �����/-��IŋCL�k@����H���	 H;H8uH�@H9�u��D���H9�}H;H8�5���@�π�z�)���M�����������H;H8������   �z����E������������D  I��   E1�1�L��������t$pH�Ņ����������A9�u7D)�Ic�Hc�H��H�H�� �  H��H�HF@H�C@����H�A@H�C@����L�L� ����D��H��L�D$ L�L$hH�D�	H�,��fD  H��HH9�������G ����t�G!����u��Gu�A��8  H�w0I��@  ����   Ic�L  I��E��h  I)�L��E��A��Mc�L9�|`��H�RH��M��p  � HcPH��H)�L9�|9�PD�Hc�H9�"A��l   uIc�d  H9�|H�P �O0H�W@H��0L9�u�A��@  I��H�@H��I�T�E������E��h  HcJE��H)�A��Mc�I9������A��I��J��    I)�I��I��@ HcJH)�L9�������BD)�H�H9�|"A��l   uIc�d  H9�~H�B(�O0H�G@H��0L9�u�����H�D$ L��$  H��$  ����D�L$�C!�E������A����u�������D�T$�C!�E�������A����T��������H�I@H)�H)�D�\$@H)�H�L$8�3*��H�L$8D�CD�\$@H�H�K@�[���I��I���'���ff.�      f�~ tf�> u1������ff.�     �G����  AWAVAUATUSH��H��8���  ���   L�/I��E�H�l$$��H�vH��H�D$L�tI��H)��I�?I���=)��L��I��L��H��H��L��H����������.  H��H�D$0I��H9�u�H�D$D�t$,D�d$(�l$$H�H�z@�B8H�|$����   ��   ��A��E����A��A��D��A��D���A����A��H�D@Mc�A��D����Mc���Hc�L�<����    �9�vH�OB�	D����   D9�vH�OB�D����   D9�vH�G�0���|   H��H�|$L9�u�H�D$H�T$L��H�|8������u0��xH�|$L����H�����uE��y_E��xH�|$�9 �   �CH��8[]A\A]A^A_�f�     ��    ��y�E��y$E��x�L��D���������t��f�     H�|$L��D���������t��f.�     USH��H�PH��H�GX    H�o�HǇ�       H���4���H�{@H���(���H�s8H������H�C0    H���   H��H�C8    �����H�{pH�������H�shH������H�C`    H�Ch    �C     H�C    H��[]�ff.�     @ AWAVM��AUI��ATA��UH��S��H���G��tH�WH�@H��D�@�L�}H�T$L��L���	�����tH��[]A\A]A^A_�fD  �E����   H�@H�EH�l��H�uH�}L���������u�D��D�῀   �] ����H�u��Iչ�   ��t�@ �E�M A��A��A!�	�A��AD����u	I����   ��u	H����   ��u�H��[]A\A]A^A_�fD  H�T$L��L���8���H�l$���S���H��[]A\A]A^A_�ff.�     ��G��u)AVAUATUSD�gD�oHC�,9�t[]A\A]A^��     ��    L�7H��H��E1�1�H�D��H��M���h�����uE1�H�{HM��D��D��H���L�����t��C[]A\A]A^�ff.�     ��G��u)AVAUATUS�GD�gHF� D9�t[]A\A]A^��     ��    L�7I�͉�H��A��H���D��M��L���������u1�H�{HM��A��D��L��������t��C[]A\A]A^�f.�     �H���    H�O8��   H9O0��   H���   H�@(    H�@     H�HH�@    H�@8    ��8  ��u=A��A����E��AE�f�HH���    t6�   ���   f���   1��f�     ��tT��(H���    ��f�Hu�H���   ���    �G@b   �   � H���   H���   H��@H�O8�/���D  ����f�H�q���f�     H�G8H���   H��H+Jx|tRH��H�J @��t�rA����A�� ����AD�f�JH�H@H���   H�O8H�@     H�HH�B8H��f���   H9G0vƇ�    1���     �G@b   �   � �G@c   �   � HcGDL�_(I��M��H��D��I)���x/I�S�Lc�L9�~OA�B�H���    H��I�T�L9�~2����y�H�G0H��H�G0H;G8vjA�BA��Hc�Mc҉GD1�K�4�� 1�L9�}ALc���I��H��K�O�D�I)�Hc��	 H�Hc�H�H����L9�u��f.�     ��    �G@b   �   �ff.�     H�W H�OH�W@H�HH��H��?H�H��H��H�G0H��H��?H�H�OH��H�GH�H��H��?H�H�W(H��H�WHH�HOH�G H��H��?H�H��H��H�G8H��H��?H�H��H�GH�H��H��?H�H��H�G(��     H�OH�H�W H�w0H�H�w`H�LH�tH��H��H��H��H�GH�TH�DH�OH�wPH��H��H�w8H�G@H�DH��H�W H�W(H�G0H�GH�whH�tH�H�LH��H��H��H�wXH��H�TH�GH�DH��H��H�GHH�DH��H�W(H�G8�ff.�     �AWI��AVAULc�ATI��USH��H��(L�gHH�w8M�t$O�,I�QI9��  L9���   �H��H�����Hc�I!�M9�MN�H9��  ���    t�H���   H��H�B(ƃ�    L9���   �L��L��H)�H��L��H�D�H��H9C0wT�>  fD  J�/L�RL)�I��HcCI9���   H�L$H�t$H�T$A��H�T$H�t$H�L$H��L9�r8L9�3ƃ�    H�GH9�|�uƃ�   H�H��H�F�HcCH�H�L9�s�L�cH�fD  L��H��I�H�s81�L�cHH��([]A\A]A^A_�fD  Lcǃ�I�D�H!�H��f����������    ��   H��H��I�I�, H����    ���������fD  L�H�H��H�L)�H��L)�H��H�I��L�H�F�HcCH�����fD  H�s8�   �C@b   H��([]A\A]A^A_ÐH�N�ƃ�    �v���ATH��UH��SH�_HH�[H�[H�[(��uH�[8L��H��D���   H��H��I������E��t���    uH���   H�Z(H�[[]A\�ff.�     @ AUI��ATL��@  UL��SH��H��H�GhL�gHH��P  H��`  H�GpH��X  H��h  L��H��@  L��H  �> H9���   H9���   H9���   H�� H�{HI9���   H�G(H�WH�oL�/H9�}�H9���   H9���   ���   ��tX�sA�   �V�Hc�H!�HcSH9�A��E�Ʌ�tD��H����������   D��D��H����������   A����   H�KxL���   �PE H�߾   �f�������   H�{HI9��E���L�kh1�H�kpH��[]A\A]�@ ����H�CHH�x H�{H����f����   �4�����t/HcsA�   H��H�t0���Hc�H!�H)�HcCH9�A���$���f�H�KxL���   �PE H�߾   �������]���H���   []A\A]�ff.�     AUATM��UH��@  SH��H��H�GhH�oHL�l$0H��`  H��p  H�GpH��h  H��x  H��P  L��X  L��@  L��H  H����   �     H��L��L9�~	I��L��M��H9���   L9���   I9��  ���   �  ���,  HcsA�   H��H�t0���Hc�H!�H)�HcCH9�A��E�Ʌ�tD��H���������  D��D��H����������   A����   H�KxL���   ��E H�߾   �l�������   H�{HH9�wAH�G8H�W(L�GL�oL�'I9�����L��H���
���@ �K���H�CHH�x0H�{HH9�v�L�ch1�L�kpH��[]A\A]�D  H��0H�{H�fD  ���^����sA�   �V�Hc�H!�HcSH9�A������D  H�KxL���   ��E H�߾   �������7���H���   []A\A]�ff.�     H�H����   H�АH�pH�H��H��f��H�H�h H���H�LH�HH�@H��u�H�BH��H��u�G�    H�JH�RH��t;H�BH��t&H�0H92~�H�H�HH�JH��H�PH�H�BH��u�� ��    �ff.�     @ Hc��   H����f��  ���H�H��H��   H��~���   ��H��H�H��   �ff.�      LcOE�@I�ʋL��A����Hc�I�D�H!�H��fA����   M��I)�H��M)�LcOM9���   H����   D�GPL��I9���   H���    HI�I9���Hc�I�ɾ�   ��H�����Ѻ   H����I���A����H��   D)ȉ�L�HOX�����~ZA	�D���t+��H��H�|H��f�     H��� �H9�u�Hc�H�L@q��    L!�H��H��H���@����D  D!�	�@�1�ff.�     @ AUATUSHc_H��L�T���H�I��I!�I!�M9�D���I��L��M��x'�GPL9�~L�Ѓ���   H��H�   HGX��[]A\A]��    L�L9�u�A�h���f��tf����   f��t#f��u�M9H8��   M9A8��   L��f��tH�T
�H��H��?H�HcWH��H�H!ƋH��x��H��H��H���WPH9�|_L��M��I�҉�I��M���&����WPL9�����L��A��H��HWXH�   D���2��   ������������� L��� L9�t�M��I��� I�x  �<���@�������I��LcgI)�M9���������� H��I9p(������ �����I��HcwI)�I9����������f�     H��  H�   ��ff.�     @ LcGI��I)�L��M9�}��I�T�H�H!�H!�H9�t
�f�     �H��H��x싇�   I��H9�v�Lc��   ��   f����I������H��H)�HGXE��~A�P�L��L��ff.�     f�AVAUATUSHc_H��L�T���H�I��I!�I!�M9�j���I��L��M��xK���   H��L9�v=Lc��   ��f��A��   H����I��A��H)�H�GXH�E��~
��L��L�D []A\A]A^��    L�L9�u�E�`H��D���f��tf����   f��t#f��u�M9H8��   M9A8�  M��f��tH�T
�I��I��?I�HcWI��I�I!��M��x L�É����   H��H9���   L��M��I��Lc��   ����I��f��M��H��M��L)�HWXE��~���   ��L��L�M����������   L9��������A��   ��A��D������������M���c����     M9��y���M��M���n���@ I�x  �	���A�������I��LcoI)�M9���������� I9h(�����A�� �����I��LcGI)�M9�������l���ff.�     ��ff.�     @ �ff.�     @ 1��ff.�     f�H��H��1�H�hH�@1�H�@p�P1�H���ff.�     @ H��H�hH�@H�@p�`ff.�      H��H�?�%���D  AWM��AVI)�AUATUSH��8M9�A��H;T$p��A���  M���{  I��M��M��I��H��I��I��I)�L9���  �H��H��H��I�ŋG��!�L;t$p�Q  H�|$pH��1�I�����X  E9�L�T$ L�D$�L$D�L$�  A�t$L��L��L�\$(A��)�Hc����L�\$(D�L$HŋL$I�D$8L�D$L�T$ ��A��$�   A��$�    tI��$�   Ic�H�J(AƄ$�    E)�E��E�MIc�H��I9D$0�(  Ic|$D�L$M���5  L��L��L�\$����L�\$D�L$H��IcD$I��H�I���   L)�M�D$8H��E���1  K�t�@ I��I�h�H�H�xL)�H�L9�u�I�t$8H��81�[]A\A]A^A_��    A�t$L��H���N�I��D!�������A��$�    I�D$8�����H��I�D$8�����f.�     H�t$L��L��H)�L��H�L$L�\$���L�D$A�$L�\$L�T$I�, I��1������    A�D$@b   H��8�   []A\A]A^A_� M)�L��L��L�D$���L�D$D�L$H��H��IcD$I��H�I��H���������� L�������AUATI��UH��SH��H�����   ���N  ����   ��u^H�WpH9�|pH�CxH��H�shI��L���   H��L��I��H��D���   H��PI�������ZYE��t���    uH���   H�Z(��uKL�ch1�H�kpH��[]A\A]�fD  HcO1�H��H�L
���H�H!�H)�HcWH9�@���������0  H���   []A\A]��     H�GpH9���   ~��O�Q�Hc�H!�HcS�   H��H9������K�����u����   ����   H�SpH�����   H��I��H�shL��L�Kx�����^_���'����m���D  H�WpH9�~ËG1���H�H!�HcGH9�@����������:����G��H�H#Gp�\����HcOH��H�L���Hc�H!�H)�HcGH9��¾   H�����������@��������f��������H�Sp�6���fD  HcWH�OpH��H�T���H�H!�HcWH)�H9��D  AWAVI��AUATUSH��X���  @�t$@ ����  H�IcNI�^(E1�I��E1�H��R  H��I���   H��P  H�S�Iǆ�       H��fE���   fA���    I�V0I�F@    I�FxI�F I�F8I���   H�@fE���   �  H�D$    1�f�     H�|$I���   ��Aǆ�       A�NMcFIǆ�       H�?�<zH��H�D$(I���   H��I��I��I�H�H�M�MH��H�PH��I��I�U L)�I��H��L��M)�H��H��L)�L)|$ tH��L��I��H��H��H��M���   L����t��A��8  ������T  ��u9A�8�����_  H�I�H��L��H��?H��?H�I�H��I��H��H��I�nhM�fpI9��Z  H�l$L�d$ �SL�xH�k���W  ��uZH�PH�@A�NIc~H��H��H��H��H)�H)��|$ t	H��H��H��L���������  H��M9���   L����    H�P I9��{  �S�����k  H�PL�@L�x0L�H(A�NH��L��L�@ Ic~H��H��M��M��H)�H)�I��I��I)�I)��|$ tM��M��M��I��H��L��M9��!
  L�X0M��L�X8I��L��I)�H��H)��|$ t	L��I��H��H��L��L��P����AXAY���3  H��M9��"���H�l$L�d$ L��H��L����������  �  �H�PH�@A�NIc~H��H��H��H��H)�H)��|$ t	H��H��H��M9��5	  M��I���WD  ���@  H�D L��I��I��?I�H�3H��I��H��?H�H����������}   M9��4  A�NIc~H��H��I��M�I��A�E L��M�G��H��L��H)�H��H)��|$ t	H��H��H��<�m���I��H��L��L��M��M���n����������fD  A�~@b��  Ic��  A�F@    I��H����R  ��P  A��։׉����������  f9���  f��T  ����fD��V  f��R  A���  ���\���H��X1�[]A\A]A^A_� A�F@   �   H��X[]A\A]A^A_�@ I��I��H�������I��L�d$ H�l$M��H��L��H��L������������I���   H�\$(I�VpI�v8�A�FM���   �H���Hc�H!�u6I;Vx|0I;��   'I���   H��t�fA3y��uH��I�v8D  Ic~I9q��   A�A��   H9�@��@��L���t������|���I���   H��tI�A8H�D$A���   H�|$9������E���   I���   fA��@��H����@ �uA�  f�     D�l���L���������	���A�u�����������H�[fA��tmH�C 1�fA��tH�SH��H�SH�S(�Cu��rA��)�H������HCHc�H�K(�D  Hc���H�L
�H�H!�H)�H9�@�������f.�     I�F0I9F8�r���I���   H����   A�I�FxE1�E1�H�D$8    H�D$@    H��A��f�D$6I���   H�D$H    H��A��f�D$41� H�r(�J H�z��fD9�}A��A��fD9�~A��A��H�    H����  H�8 ~�  @ H�8 H�HH�@H��u�H�BH�H��tIH�D$8H����    I�V0I�F8Iǆ�       H9������A���  ��A���  �>���fD  E��tfD�D$6E��tfD�L$4A�ND����  H�T$6H�t$4L��A��  H�D$8H���  �L$4��D  �P()ʉP0H�@H��u�A�ND����  ��I�v(H����H�H9�u��A�ND1�f�T$f�     ����  H�D$8D�l$H��u�    H��H����   D)h0H�pu�H�T$8H��t%H9�u��  fD  H9��7  H��H�JH��u�H��@�.  H�T$@H���`  H9
~�V  fD  H9
H�zH�RH��u�H�PH�H��H���w���H�|$@����H�|$H�w���A�FDI�V(�H���H�A�NDL�$�D��)�f�D$fA9���   A�\$�D��)�A�o�ۍ+�D$H�\$@L�l$H1�H����   �l$ ���     H�I�M H9�~	H��H��H��McFH��H)�L��I9�|9��N�L�Hc�H��L!�H!�H9�t!H9�tH9���  L�H9���  �    M��I��D��L��A��   H�[M�mH��u���l$ f���I  L��A��A��0  9l$�  A�NDD��H�T$@H��u�W�    H��H��tHH�z  H�zu�H�D$@H��t�H9�u�  f�     H��H�pH��t�H9�u�H��H�8H��H��u�H�T$HH��u�����H��H�������H�z  H�zu�H�D$HH��t�H9�u�  D  H��H�pH��t�H9�u�H��H�8�fD  H�T$HH���J  H;
}�@  �     H9
�����H�zH�RH��u�H�PH������fD  H�|$@���K���H�|$H�A����	���@ H�\$@L�l$HH�������D  �C0��t!�C0    M��I��H�I�M D��L��A��(  H�[M�mH��u��e���fD  �s��f���2���H���I�M �C0   ����f�     H��H�2�����@ H�L$8�i���fD  f;l$6�����D  L����A��0  f9l$6}��s����    H�|$@H�PH������    H�|$HH�PH������    H�T$8�z���fD  H�D$H�k���fD  H�D$@�����fD  H�l$L�d$ I��H���H��� A�F@   H��X�   []A\A]A^A_�@ L�d$ H�l$L��L��H��ATI������^_���0������� Aǆ�      �   A�F@   ���� �l$4������   ����@ H�VH���  H����   H�zf����   H�f����   L�BM����   H�JH����   E�D@�D�ϸ   A��E9���   �   �F��   L�M����   E�HE����   A�0��tzI�x tkH��H�9H9�svH�1H��   H��   wKH�qH��   H��   w7�    H��H9�v?H�1H��   H��   wH�yH��   H��   vи   �f�1��D  �`   �f�H��G  �o�AoH��$�G  �$�   �oJ�$�   H�B )�$�   �AoXH��$�   )�$�   I�P H�L$(H��$�   H��$�  H�T$ ���u  �$   �   �   H�      H�L$�   �t$�L$�T$�T$��  Ƅ$8  ��	1�1�H���HǄ$   E ��HǄ$   PE ��$9  ��$�   HǄ$(  �E ��f��$P  f��$R  ��$�   HǄ$0  @E f�D$PH��$�   Ǆ$�      H�D$X�:�����uy��$9   tw��$8  tm1�H��   HǄ$  PE f��$P  ��$�   HǄ$   `E HǄ$(  �E ��HǄ$0  E Ǆ$�      f��$R  ����H�ĨG  �1��������� �JDш�$8  ������$   1Ҿ@   H�       H�L$�    ����ff.�      UH��SH��H��H�    �   H�T$�Na���T$��uH�(H�H����[]��    f��B�G 9��   t
�f�     H���   H���1A���AWAVL���   AUATUSH��H��   L��G �D$    9��   tF�D$   1�E1�E1�H��(  �@�e  H���  �D$H�Ĉ   []A\A]A^A_�fD  �   ��u�H��(  H��I���@�W  L�Ҿ   H��L�T$�b�����   E1�1�Hc��   L�L$L���sr��H���   �D$���Z���D���   H��(  D���   L�T$A��D+��   �HA��A��Mc�Mc�M��tM"MjL��L	�unH���   H�L$H�}hH�t$ H�D$ L�t$(�D$0    �UpH�L$���D$�����ǃ�   stibH�������L��L��L��H��H����?��������    L��L��L��H�L$�?��H�L$�u��� H���   L��H�L$�T���H��(  H�L$Hǃ�       �`��g���@ H���   L��H�L$����H��(  L�T$Hǃ�       �`��u���ff.�     �ATA�   US�G 9��   u6H��H��H��tH���   H���A��E1�H��tH�UH�u H���   ��>��D��[]A\�f.�      �ff.�     @ 1��ff.�     f�H��H��1�H�hH�@1�H�@p�P1�H���ff.�     @ H��H�hH�@H�@p�`ff.�      H��H�?����D  A����H��A��A��	A1����   tSD�Ⱥ�  %�  )�A��   L���   E�M��tJH���   �D$H�T$
D��f�t$
�   fD�D$A��H��ÐA���   ��   AN�L���   ��M��u�D���   Hc�Mc�L)�H��   H��A��wYE��B�$���H fD  �H���H�G�H�x�H�W�
H�B�H�x�H���D  H���� H���� H���� Ic�����9 �R����     f��B�G 9��   t
�f�     H���   H����<����GDH�Wh+GP�O@H�H��H�H��t;|�tNH�PH�@H��t9~�H���   H;wx}=L�FH�4vL���   L�GpI�4���OX�N�O\H�F�NH�2� �WXP�W\P�AQ�   ��: �    SH�� H�|$�D$    �: ��t�D$@   �D$H�� [� H�\$���H H���   H����*���D$�C`��u�H�|$�����D$H�� [��     AWAVAUATUSH��@  �WP�GT�OH�D$)ЉL$�OLHc��T$�L$H��Uv(H���������H�VTH��H��H��1�H��H�D�H��H��L�$�   H���������I�T$�H��H��H��$�   H�OhH��H�RH��H�Gp��  H)ЋT$H�Gx9T$��  I�D$�t$I��L�l$ H�$H�ϋD$�L$L��t$D�d$A�GP�D�t$9ƉD$N�D�d$$D�t$ A�GTD��E��A���8@ ��@�G  ���?  D�D�uH���] L9��  D�e D�uI�hH�$1�D��D)��P7 A�G`   L��IǇ�       E�wHE�gL������u�E�gPE;gT��   D�� D��I�Wh)�Hc�H��H��tm�E1�fD  �S��	A�D��+KtA9GH~aH�[�pH��t%�E��t�9�}�)�D��D��L��A�������� E��tE�GLD��D��L��A)�����A��E;gT}$A�GP�k��� ��A�   D��L���u����눐H��L9�������|$9|$~ I�h�k����   H�Ę@  []A\A]A^A_�1���D  H���7  �V�   ����  H�~H����  �Gf���l  H�f���_  L�GM���Z  H� �O  A�LH���9��>  USH��  �o��H�.�$�   �oO�$�   H�G H��$�   �  H�FH���  H��$�   H�F8H��$�   H��H���8��H�$H��   ���   H�D$H=   ��   H�t$H��   ���   H�T$H��   ��   H��?H��?�{H��H��H��H�$H��H�t$H�D$H�T$@���  D�MD�E 1�E1�L9�IL�H9�HL�L9�IO�L9L$hIOЉt$p�D$l�T$t9�}A9�}=H�|$ ������D  1��D  �   �f��   H��  []ÐH��t�E��u$H��  1�[]��     �   ��f�     �E ��t�H�UH��t��M��x	����H�H��$�   ��$�   HǄ$�       HǄ$�       ����@ �   �f.�     ��tL�S@H�{HL�KPL�CX�����H�� ���A��  A��  I�������ff.�     SH��H���GH�H�9��G`O��uH�X uGH�CX    �   �s@�SD9ST~9SP~�C`H��[�f�     1�9sL���C`H��[��    �T$�t$�{����T$�t$뢐AWAVAUI��ATUSH��XH���   H�t$H��H�T$H��H��H�ՉT$ 9�N�9WT�4  �WPA��9���  9��  H���   H�L$I��H��I��H��H)�H��I��H�|$I��A��Hc�D�T$0H��H)�H)�Hc�H��I)�D��H���R  M����  M��H�؋L$0H�D$@    M��H��I)�A9�tH�������� H�I��H�D$@H�D$8    9�tH�������� H�H��H�D$8H��I��H�l$HL��H�|$(L�|$M��I��L��E��E���     L����H+T$�C\�sXM����  H�L$(L�H����  )�M���<  H�T$8A��C\A���D$4   �   H��I��L|$H��8I�I��D��D)ƉsXD��D��H������D;d$0�t���D;l$ �i���I��I�݋L$4L��H�l$H�RD  H���   L�\$I��H��H��I��H��D�\$0Lc�A��I��L)�Lc�I��M)�D��D9���  9���  Lc�H�T$A�E\I��L)��L)�)�H�L$A�E\HcD$0H��H)�H���A]XH�D$I���   H�D$I���   H��X[]A\A]A^A_� A��H�\$H����  A��H�l$ D��E�̐A�E\��D��L���   D)�A�E\�   L)����AEX����E1�A9�u�H�\$H�l$ 1��3���fD  H��~CH�T$@)�A��I��L+|$(H��8ЉT$4�C\H��H)�H�Չ�A��A�   ΉsX�^��� H�L$(L�M��~JL�T$   A���D$4    )�M)�L�T$8�C\I�׸   H)�1�I��8K�M����ΉsX�����)�H�|$(L������H�T$@I��   A��I��E1�H��H��8ЉT$4�C\H��H)�H����ΉsX���� ��t$0L��L$ L�\$�i���L�\$�L$ M�������     H�|$M��L�|$H)�I)��]����     D��E��A���    E)]\I�ۃ�D��E�މ�L��E�E]X�����A�   A9�u�H�\$�   A�   ����ff.�      H��H��H�OH�7H��H��    H���.���1�H����    ATI��USH�H�_L��H�,�    H��H��H��H��H���p���I��$�   1�I��$�   []A\�f�     UH��SH��H��H�    �   H�T$�P���T$��uH�(H�H����[]��    AWI��AVAUL���   ATUSH��H���   H�G� �D$\    H�$H��(  �@��9��   t2�D$\   E1�E1�1��u:M��ua�D$\H���   []A\A]A^A_� A��D9�t`�D$\   E1�E1�1��t�H���   H�<$����H��(  Hǃ�       �`�M��t��L��H��L��H��H���0���f.�     I�υ��-  L��D��H��L�T$�������   E1�1�Hc��   H�<$L�L$\��a���L$\H���   H��(  ����   ���   ���   ���   �H����L�T$����Lc�Hc���I̀��   Hc�u��VUUU����)�Lc�I�M��tI/MgI��M	��  H���   L�l$hM�BpH�D$`I�zh�D$p   A����   A���z  H�t$`A�ЉD$\����   ǃ�   stib�a����    �@E1�E1�1���C���D  H���   H�<$L�T$蓉��H��(  L�T$Hǃ�       �`����� ���   �����L�T$H�t$`D���   �D$ ���   �D$$�����ȉL$H��   H�D$A�ЋL$L�T$���D$\t:H��(  �@�������     L��H��L��L�T$�.��L�T$����� 1�H������L��L$L�T$��-��L�T$H�D$H�t$`H��   I�zhA�RpL�T$�L$���D$\��   H��(  H��M��I	�@�������    �����L�T$H�t$`Lc��   L��   C�6�D$D����   �����   �ꉓ�   A��L�T$���D$\����1��   L��L�T$�:-��L�T$H�t$`L��   I�zhA�RpL�T$���D$\��  H��(  I��I��M	�@���Z���@ 1Ҿ*   L��L�T$(�L$H��M����,���L$L�T$(I	�H�t$`�	I�zhH)��   H�D$A�Rp�L$���D$\�O���Ic�H�<$H�T$\�L$(H��H�D$�,L���T$\�L$(I�ƅ������D$ 1�1�����   A�   A�   L�l$0A��E)�E)�H�l$8L�d$@D��A��L�|$HE��H�\$(H���    H�D$(H���   H߃|$$vGH�D$H�L$L��L�L�1� ��
A�4A�A�4A�4�L H��H��A�4A9�w�H�T$L��A���( H\$D9d$ u�L�l$0H�l$8L�d$@L�|$HH�\$(H�<$L���I����D$\�b���H������1�L��I��L�T$�V+��L�T$Lc|$H�t$`L)��   I��I�zhM	�A�Rp�D$\����������   �VUUU�����ꋃ�   �@)򉃘   ���   ������     ���    D�E1������ff.�     f�A�   �����D  A�   �����D  AWH��I��AVH��H��AUATN�$�    USH��8  L���   L���   H��$p  L�d$ H�L$0H�,�    �GTL�D$8I��H�l$(I��H�t$@H�T$HL�t$PL�T$XA9�|M��I��D9���  �GPH�|$A9�}-M��I��D9�~!I��I��D9�~M��I��D9���  D  H�\$ H�\$fD  M��L��M)�H)�L��H��?I��M1�I)�H��H��?I��I1�I)�M9��  K�<[H��L�H���  ��   I��L��M��M)�N��I)�L��L�l$M��M�H��L)�I��I��?L1�L)�I9���   H��L)�I��H��H)�I��L��L)�I��I��?L1�L)�I9�|H��L)�L��L��L)�H�D$I�M��aH��L)�L��H��L)�H��L�H��EH�|$H��L���u���H;\$�x  H�K�L�C�I��M��H�s�H�S�H��0H�kL�#�����@ I�M�6H�L�L��L��H��I�H��?H��?L�s`H��?L�L�L�ShH��H�H��M�H��H�CL��L�$0H�H��?H�{PL��H��L�H��?H��?L�H�L��H��H��H�C H�H��?I��L�H�K@I��?H��I�H��H�sXH��?I��H�L�c0H��H��H��0H�,H�H�C�I��H��H��?I��?H�I�H��H��H��I��H�C�L�H��L�CH��?H�H��H�k�����D  K�|m H��L�������    I��I��D9��N���M��I��D9��>���L���   H���   H��8  []A\A]A^A_�H���rH��L�
L�FH�H�WH�7H���m���1�H���fD  AUI��H��    H��    ATM��UI��SH��  L���   �_TL���   H�L$H��    H�$L�D$H�L$L�\$ L�L$(A9�|H��H��9�L��H��9���   �_PA9�}H��9�~L��H��9��`  �L�H��A�   H)�H��H��H��?H1�H)�H��K�H)�H�H1�H)�H9�HM�H��@~H��E�H��@�H��H��D  A����   L�C L�[�   H�{(L�S�
�    L��K�L�L�C@H��L��H�{HL�k H��?H��?H�L�H��H��H�sH�I��H��H�C0H��?H�J�LSI��H��I��?H�s I�L��H��?I��L�L�K8H��H�SL�I��I��?L�M��H��H�S(D���e���H�������A���+���H��  []A\A]�D  H�SH�3H��H�� ����A���������H���   L���   H��  []A\A]�D  H��H��L�FH�WH�H�7H�������1�H���ff.�     �ATA�   US�G 9��   u6H��H��H��tH���   H���&��E1�H��tH�UH�u H���   �u$��D��[]A\�f.�      AWH��AVAUATUSH���   H�L$�L��$(  H�D$�    H�D$�    H�D$�    H�D$�    H�D$�    H�$    H�D$    H�D$    �T$�H��$  L�D$�A��L�L$�N�� H���H��D��L9�u�D�T$�A9��i  ��D$��   fD  �l�؉�����   H��H��u��D$�   �   �   D�L$�D9�v	�L$�D�L$�L�\$�   �A���uYI����u����    D)Ӊ\$���  �D$�E1Ƀ���D$    �D$�    �D$�    �   @ �D$��   ��� �t$�;t$�s�t$�A��\$��9��  ��+D���m  D�Q���J�T��I�J�L���fD  +H�����B  �H9�u���+\�؉\$��)  �D�؃��D$    ��1�1��f�     H��T��H�H�T� H9�u�L��$0  1�f�����t�L��qA���t�H��L9�u�HcD$�E��H�D$X    A��H�ËD��D$    ;\$��  E1�H��$0  �D$�    H������A�   H��1�H�D$�HcD$�H�D��H�D$��D$����D$�1�H�|$����|$��|$��O�D����|$ċL$�����  �|$��l$�G�D)�D)��J�D��L�\�XL��B�\�A��L)�A��H��D��A��I��A)�@�2D�|$�D�JD�zE��D)�D)�Ic�E�D;D$���   D����D�R����9D$�s�t$�9�A����DG�A9�wEE�u A����  ��   L��$   A�M O�4�Mc�N�t�XE���P���H�t$�L�6�fD  �wA9�v/L�|$�+D$��A�9�w�@ I��A��9�s
��)�A9�w��D��E�u ��A����  �}���fD  �����H���   []A\A]A^A_ÐD�D$������H�|$�E)�H;�$0  v4H��$0  H��$0  �?�|$�;|$���   ��   �`   �    E��L$�D��A�ڋl$�D)���D��A��D��D9�vfD  A���O��A�2E�BA�j9�w�|$ĉ���tfD  1����u�1�D��D��Hc������!�;L�t+��D��Hc�D  D)�D��Hc�H�����!�;|�u�A�˃l$�����f�     H�D$�H�     1��    ������    H�|$��L$�+L$��<��|$��|$��wPH�|$��<��|$������D$��|$�H�D$�;|$��-����t$Ѕ�t�|$�u1��q���������g������+\�؉\$��P����D���D$    ���G�������ff.�      UH��SH��H��H��tH�GhH���P���wH�sH�}P�UH���uH�sH�}P�UHH�C@�    �C,    H�CXH�CPH�C`H�C0    H��t1�1�1���H�ChH�E`H��[]�H��tGH�W8H��t>H���zH��H�G(    �H�G    ��H�G0    H�z ���1��;���1�H��ø�����ff.�      H��tsH�w8H��tjH�GHH��taUSH��H��H�n H��t51�H��H�������H�u@H�{P�SHH�u8H�{P�SHH��H�{P�SHH�CHH�s8H�{P��H�C8    H��1�[]� ������f�AWD��H��AV��AUATUSH�D$�H����  ����  I��f����  ��  ��F�)ǉ|$����  ���D$����D$�H��H��L�H�D$� A�E�rI��E�j�E�b�L�A�j�A�Z�I�E�Z�E�J�M�L�E�B�A�z�M�L�A�R�E�z�L�L�H�H�I�4E�Z�H�H�t$�H\$�I�A�r�L��E�Z�H�L$�H\$�I�A�J�M�I�M�M�L�M�H�L�H�H�H�H�I�H�L�HT$�L;T$��.����D$��|$���)ǉ���   H���/�  H�|$�I��L��H)�H��H�H���/�  H��Hi���  I)�H��H��H)�H��H�H��Hi���  H)׋T$�H�|$����u���H�D$�[]A\H��A]A^L	�A_�fD  L�T$�H�|$��H�L$�H��H�tH�� H���x�I�L�H9�u�H�|$�Hc�H�L$�L�T�5���[�   ]A\A]A^A_�ff.�      ATUH��SH�_L�g8H��tiH�{�#���H�CX    H��L��H�C`    H�Ch    H�C    H�C0    �C     �C8    H�C    H�    H�C    �Ku��H�E    H�}( t[]A\��    H�u L���$u��[H�E     ]A\��    �u��ff.�     ��t��ff.�     �҉�H��H��H�T$�9��H���D  �҉�H��H��H�T$�9��H���D  U1�SH��H���0%���D$��tH��[]Ð�   H�t$H���N&���D$��uހ|$�   uҀ|$�uˀ|$u��D$�u��   H���(%���D$�D$�uj�t%H�l$f�H��H���U)���D$��u���u��D$�t0H�l$f�     H��H���%)���D$���O�����u��D$�uF�D$�9���H�l$H��H���1-�����D$������H���$���D$�������D$�Y����   H���g$�������f�AWAVAUATUH��SH��H��L�PH�GXL�fL9�sH�GH�M L)�9�F���thE1���u`)�A��Lu(�M H�K`H��tH�{h��L����H�ChH�E`L��L��L��M��2 M�L9sHt&L�eD��L�sPH��[]A\A]A^A_�@ A��� H�SXH�K@�E I9�txH)�9�G�A��)�O�<N�4��tA����    DD�E H�C`LE(H��t#L�D$H��H�{hH�$��L�D$H�$H�ChH�E`L��L��H��M��� �[���f�     H�KXI��M��E1�1��ff.�     @ H����  AVAUATU��SH�G@H��H�G0    H���%  H�PH�{H �  �(   �   ��I��H�C8H���r  H�@     ����   �@    �E����7  A�D$��H�{PA�l$A�   A��OE �p   �   A����    LE��S@H��H����   H�{P��  �   �S@H�{PH�E8H����   D��   �S@H�E@H����   L�L�u`1�H��H�EHH���E     ����I�l$ H���.���1�[]A\A]A^� ���@   �/���f�H�CH�RE ����� H�G@�RE ��RE H�GP    1������@ H���SHI�D$     H���)���������f�H�u8H�{P�SHH�{PH���SHI�D$     ��H�������������b��������ø�����R���ff.�      H���w  H�O8H���j  AWAVAUATUSH��hH�/H���L  E1�������A�ă9G�d����   �H���$� �H �    ����������   H��W�H�C�SH�pH�3� �   H��H�AD������   H���H�C�SH�pH�3� �   H��HAD����t\H���H�C�SH�pH�3� �   H��HAD����t/H���H�C�SH�PH�� HAH�AH�C`�   �   H��h[]A\A]A^A_��    �GA���������  ��H�C�CH�H�PH�� HAH�AH;A�  �   H�C0�H �A   H��h�����[]A\A]A^A_�@ �W����  H�E��H�GH��W�u ���q��<��  �   H�G0�H �A   렋W��������*���H��z��q�{H�PH�C��H�� ��B�A�������)����������)�9��R  �   H�C0=�H �A   �0����W��������� �   �����H�G0T�H �A    H��h[]A\A]A^A_��    �W��������z���H���H�C�SH�pH�3� �
   H��HAD�����I����B�H�H�C�CH�rH�3��   H��HQ�=���@ �W������fD  �W������l��� �W��������� ������S�������H���H�C�SH�pH�3� �	   H��H�AD���*����   @ �   ����fD  A�� �[  �   H�+D��L�Q D�sM�ZXM�BPM�z0E�j,M9�s%M)�A��A�D�$$M��A�҃�	�_  �$Ő�H �E�BHE)���M��L��M�|$0H��H+�����E�l$,H��L��HCD�sH�+M�\$X�������m  I�t$H�{P�SHM�\$XM�D$PH�+D�sM�|$0E�l$,M9��+  M)�A��A�T$(����  A�$    E1�A���#  E���6  �E D��A��L�MA��E1�H��I	�D����A�D$(D��������l  ����  ���i  A��A�$   I��L��D���I��A)�A��w@E����  D���f�     E����  H���E�A��H����I	ǃ�v�A��E1�L��H��H��L1�f����  E��E�l$E����  A�t$(����  D��M��E1�D�$$A�   �[  M��D�$$M�z0H��H+E�j,HCD�sH�+M�ZX�����H��L������D  �����
  ���o
  D���A���E�L$A�T$���������э�  D9���  A�t$D9�v>E����  D����     E����
  H���E�A��H����I	�9�w�A��E1�I�D$ D��#���H H�ȋxD�@���  I�D$A�QD��E)�A�T$I��B�<�E�L$�M���A�D$A�t$D����
��9���   H���w!E���   �E A��H�UE1�H����I	Ǎ~I�D$�4�@�H ��A�|$D��I�����<�A�D$A�t$��
��9���  H��H���v��f��VI�D$A�T$��@�H ��    A�t$��v�M�D$8I�D$M�L$ I�L$D�T$<H�{P�   �   L�\$0A�D$   L�D$(L�L$ H�L$H�D$�D$X    �S@H�L$L�L$ H��H�D$L�D$(L�\$0D�T$<�0  D�T$ �   �   L�\$�t$H�D$`PAPE1�QH�|$01�� ���H�� L�\$D�T$ ����  H�SHH�{P�����  A�|$ ��  �D$ H�t$D�T$L�\$�ҋD$ L�\$D�T$����  A�D$    E1�A�$   �v���M��D�$$M�z0H��H+�   E�j,H��L��HCD�sH�+M�ZX�$������������������D$�t$(L�\$0A� I H�|$ �t$��I ��H�<�H�T$TR1��t$(H�D$`PL�L$x�!���H�� L�\$0���(  �|$H H�SHH�{PD�T$<u�|$  �P  D�T$0H�t$L�\$(��H�L$PH�{P�0   D�D$HD�L$D�   H�D$XH�L$ D�D$D�L$H�D$�S@D�L$D�D$H��H�L$ L�\$(D�T$0�s  H�|$D�HD�@I�t$H�x(H�{PD�T$L�\$�     H�H I�D$�SHA�$   D�T$L�\$I�t$PH��M�D$M�|$0E�l$,H+D�sHCH�+M�\$XL9��m  L)ރ�L��A� I��M��I����	��
  �$���H A�$   I��A��L��A��w:E���p  D��� E���  H���E�A��H����I	ǃ�v�A��E1�D��D��%�?  ��A�D$����  ��������  D�T$��  H�{P�   L�\$�S@L�\$D�T$H��I�D$�   A��I��1�A�D$    A�$   D������A�$   E1�E1�E����  E��uRM9\$H��	  M�\$XD��H��L������M�\$XI�L$PI9���
  I��I�T$HM)�A��I9��e  E����  A�L$H��L��D�D$D9�AG�D9�AG�A�ɉL$L��L�L$�� �L$L�L$D�D$I��L�A)�M�A)�A)L$�����A�$E1������D��M��D�$$M�ZXL��H��L�$�����L�$M�ZXM;ZP��  A�   �\���E1�D��#���H H��I�D$H���B��A)�I���
�ȅ��O  �BA�$   L��A�D$��u_M9XH�g  I�HXD��L��L��L�L$L�D$�>���L�D$L�L$I�HXI�PPH9��+  H��I�xHH)΃�H9���  ���  A�D$L�Y��E1҈A�T$I�D$ A�$   A�T$I�D$D9��$���E��u�
  @ E���$  H���E�D��A��A��H��I	�A9�r������A�T$A9�s4E��u�	  E����  H���E�D��A��A��H��I	�A9�r�E1�D��#���H H��I�D$H���B��A)��I���	  ��A�D$�BA�$   A�D$A�T$D9�v9E��u�:	  D  E���\  H���E�D��A��A��H��I	�D9�w�E1҉Љ�A)�A�$   �<���H D!�I���AD$A�D$�A�D$L��I�P@H)�H9�sI�@HH)�f�     H�H9�r�A�L$����   �r���fD  M;XH�&  M�XXL��D��L��L�L$L�D$�:���L�D$L�L$I�xXI�PPH9���  H��I�HHH)���H9���  ����  �L�_��H���I;XH�U  A�l$A�    ��������m���L����A�T$�����M��L��M�|$0H��H+�   E�l$,H��L��HCD�sH�+M�\$X���������L��L��M��I��A��vA��A��H��M�\$XD��H��L��L�D$�M���M�\$XM;\$PL�D$��  A�    �t������  ��A�D$�BA�$   A�D$A�T$D9�v<E��u�5  �     E���T  H���E�D��A��A��H��I	�D9�w�E1҉Љ�A)�A�T$�<���H I�D$(A�$   A�T$D!�I�D$I��A|$�����L������ �������H�K8H�މ$H�y H�Q����H�K8�A��t]�   �$�����    H�C8�    �@    �����f.�     ����;qvu�   H�G0)�H �A   ���� �   D���_���f.�     M��D�$$A��1�M�z0H��H+H��E�j,L��HC�C    H�+M�ZX��������@ �   D������I�X@����M��H��H+�����M�z0H��L��D�$$E�j,HCD�sH�+M�ZX�U����P���������A�t$HD)�����E�D$HE)������I�@PI�x@H9��������  H)��p����
���I������A��D��M��D�$$����I�|$8I�t$  L�\$0D�T$<�   H�|$H�{PH�t$ �   �L$(I�D$     �D$D	   �D$H   �D$�D$L    �S@L�\$0H��H�D$��  PA� I ��I H�T$TR�  �t$(H�D$\P�t$0H�|$@L�L$p����H�� L�\$0���}  �|$D ����M��D�$$H�C0��H �����H�{PH�t$�D$L�\$L�$�SHL�$L�\$�D$����D$�!  I�rH�{PL�\$L�$�SHL�$L�\$�D$A�	   M�z0H��H+H��E�j,L��HS��D�sH�+M�ZX��������M��L��E1�M�|$0H��H+D��E�l$,H��L��HC�C    H�+M�\$X�Y����������������I�HH��)��+�������  �G��D$   �D$�D$A�4 D9�v@E������D���f.�     E������H���E�A��H����I	�9�r�A��E1�D��L��D�D$A)�H��I�t$I��D��I��D��#���H �L$�D�9��3  ��u	E���%  1҃�uA�A����I�t$A��A�AB��9�u�A�L$A���}���M��1�D�$$A�   �l���D��)��-���I�x@H9��h  ��  H)��r�����������r���M�x0H��I+�����E�h,L��L��M��IAL��E�qI�)M�XX������?���I�T$PI�D$@H9��8����  H)�D�B�I��E���f��������    A�$    E1��Y����D$   �D$   �^���L�L$H�{P�0   �   L�\$D�T$�S@L�\$L�L$H����  �	  I��A��L���     D�T$f�xH�@  �H H�@( �H I�D$A�$   �%���M��I��A��L��D�$$H+A�	   H�C0d�H M�z0E�j,D�sHCL������   D���]���I�T$HA��E)��U���A��H���*���L�d$H�t$D�$$H�C0��H L�$��L�$L�T$I�rH�{PL�\$L�$�SHL�$�����L�\$A�	   ������)��E���M�|$0H��H+H��E�l$,L��HS��D�sH�+M�\$X�!����{���I��������@��  A�D$�BH��I�D$A�$�P���M�\$@L9���  I��L)�M)�A��L9�DF��t���H������M��L���.���E��A)������H�{PH�t$L�d$H�C0X�H D�$$L�$�SHL�$L�T$�����M�x0H��I+L��E�h,M��L��IQ��E�qI�)I�xXL���N��������@u3A�L$�BH��I�D$A�$����M���H��D�$$L����������L��L��M��I��� ��  �   �|���I�PPI�@@H9������H��I)�H��H)ƃ�H9�AF��������e���M��H��H+D�$$M�z0E�j,HCD�sH�+M�ZX�����H��L����������M��D�$$A�	   H�C00�H �9���L�d$H�{PD�$$L�$�SHL�T$H��L�$H+A�	   H�C0��H M�z0E�j,D�sHCH�+����I�������I�x@H9�������  H)�H���r������I�xH��)������M��D�$$A�	   H�C0w�H ����M��D�$$����������M��D�$$���uH�C0��H �������������n���M��D�$$���tc���uOH�C0��H H�{P��H�SH�D$H�t$L�\$L�$��L�$L�\$�D$�W���M��D�$$H�C0��H �������H�{PH�SH���t���H�{PH�SHH�C0��H ��	   I�A0��H �3�����H��)������M�x0H��I+L��E�h,L��M��L��IQ��E�qI�)I�HX������"���M��L��D�$$H+I�B    M�z0E�j,D�sHCL������M��D�$$�����L��L��M��� 	   I�A0 �H ����ff.�      AUH���  L�oATL���   USH��H��H���   H�G0�G8   �JD  �   L��H����H����   ��HEL�c�S 1�L���+�������   ��uv�C8����   �S ��u�H�+H�E(H�uH��u�H�EH)�H=   ��   H��t<��Hu ����sW���   ��t��>A�<$���{����t�fA�t��k��� H���   H���   �U   H��[]A\A]�f.�     H�I�$��H�|�I�|�H���   L��H���H)�H)�����H�����@ H�C0H���   H;��   t#H��1�[]A\A]��    �   �   �/����U   �r����>A�<$�t�A�t����� AVAUI��ATI��UH��SH���   H��H9���   H9���   M����   E1��    H���   H���   H)�L9�r*M�L��L����  L��   L��L��   []A\A]A^�f�L��H��I�I����  H��   H��I)�H��   ������t�[L��]A\A]A^�fD  H���   H�?�������   E1�[]L��A\A]A^�f.�     H)�D  H���   H���   H��H)�H9�rH�H�H���   H���   ����fD  H�H���   H���   H)������H��������u�H���   뙐H�{�����H���   �C     H�CH���  H�C0H���   H���   H���   1��C8    Hǃ�       �p���ff.�     �H��7����    H���  H���v  AWAVAUATUH��SH��H��H��L�n8�����D$���5  f��H�T$��   L��C0L�k8CC C@��'���L$I�ą���   H�XH��H�(H�C8IǄ$�       I�D$I��$�   I��$�   I��$�   �
������*  H������I�|$�����I�D$X�RE I��$�   H�E8I�D$`�RE I�D$hI��$�  A�D$     I�D$�2������:  I�|$ �.  �D$    L�cH�EH��L�uH�p������tJ�D$A����L�{H�C    H�    H�C(@uE H�C0 RE H��[]A\A]A^A_�fD  �(   �f�H�t$H�������T$L��H��I�ǅ�uR�M��I�G�H=��  �5  H�T$L��L���}��H�ŋD$��t:1��k��� �D$L��L���yP���D$�s����� ��A�����D$�<���@ L��H��1�L������I��L9�t*1�1�1�L�������H��L���'P��1�� ����D$   �I�|$����I�$    L��L��I�D$X    I�D$`    I�D$h    I�D$    I�D$0    A�D$     A�D$8    I�D$    I�D$    �O��L�s�D$H�C    H�C    H�+H�C(    H�C0 RE �{����D$M���K���A�����@���H��A��H����A���   H����   USH��H��xH�H�t$�   H�|$PH��H�$D�D$�D$ H�D$@�RE H�D$H�RE �������uC�   H�������Ń�tOH���_�����t3���tf���t)1������H��x��[]��    �   H��x[]�@ H��x�
   []�@ H�D$(H��H��������@ �   �f.�     �@   �f�     S1�H��H���������tH��[��    �   H�t$H���������u݀|$tH���   [��     �|$��   E�H��[�ff.�     f�USH��H���G �o<�W@�wD���
  �9{�&  9�w5f����k<���G  9k0�0  �   ��H���   �SD����   �C���  �S<H���   H�s�O����S<HC(�C    H9�H�����҉S��    9���   )ʃ��SH����   ��   �   1�1��K�D���H����M�L�B��vL�B�R��   )���M�	Ѕ�t�������A���!ʉ���	�H��[]�D  9�� ����C<	   �	   �CD   �C  ����@ 9���������L= �   ����)�H�P�Z���@ �s8�V������S������ H���   �Ox1�H9�rUH��SH��H�lH���   H��L�GpL���   I9�t_H��H��   vH��   tl�   �   H��L�L$�   L���#��H�Cp�D$��uAH���   1�H��[]��    ��    H��   �   H�Gp    HG�1�E1�H��랸������ff.�     @ H�G    �G  H�G(    �Gx    �G<	   H�    �fD  H�    H��H�1�HǇ�       H��H���H)����   ���H�H���   H�F8H�BX    H�B`    H���   H���   �Bh    H�BpHǂ�   @   H�B    �B  H�B(    �Bx    �B<	   H�    �fD  H����   H����   AVAUATUH��SH��H��H�� L�f8�0����D$��u_f��H�T$�  L��C0L�c8CC C@�;��I�ŋD$��t@H�C���H�C    H�    H�C( �E H�C0�~E H�� []A\A]A^�@ �(   �f�H�C8I�]H��M�uI�m I�EI���  I��   I���  Iǅ�      �t�����tL��L��D$��I���D$� H��L���D$�I���L�k�D$�L���ff.�     �UH���   SH��H��H�wp�G  H���   H�G    H�G(    �Gx    �G<	   H�    H9�tH���?I��H�Cp    H�sXH���+I��H�{H�    1�Hǃ�       H���H)����   ���H�H��[]�f�     ATUSH�_H��t:L�g8H��H�{�C���H�C    H��H�    L��H�C    �H��H�E    []A\�@ AWAVAUATU1�SH��H��(�GPD�wLD�oH�$H��t�I��I�ԃ�t\����   ����   �$D�kHD�sL�CPH��(H��[]A\A]A^A_�@ =   �}  �K4����  �C@    E1�E1��C H��������y��   �D  ���CxM��tH�Sp�A�/H��I9��x����Cx��uՋC@;C8s"D�[hD9���  H�SXfD�,BH�S`D�4�C@�   D�,$��    H���   �   ��������   H���   �   H�t$�A���H��H����   �D$����������щC4�S0H��H�⍲ ����s8��wg���C<	   H�������   ��
���C@�   CЉSD�	���=�   w*M��tA�I���!  �   A��A���$    �����$    �1��   �W��� ��=�   �@  �$�KxH��H;��   �}  H�sp��A�։Cx��   ����f��C@�   �$   ���  H�{X uD�H���D  H�{`��   ��H�sp�CxH���H�CX�P���   �w���H���	����KxH��H;��   r�H�߉T$������������Kx�T$H����    H���   E����   D����B��L$L�CXL��L�L$�   L�\$����T$H�CX��������T$L�\$H�<PJ�4XL��H�{`���  �L$�C@�Kh������ ���;K@��   �$�F����SxH��H;��   seH�Kp���CxD�4D��A���   ������y���f�     H�߉T$�����T$��x�KxH���d����   �D$   �%���A�������H���o�����������SxH���A��A���$    �Q����$�L���D  AWAVAUI��ATI��UH��SH��H�_H���  H9���   H���  H��H���   H)�H��H)�H9�wvH��H���  H)�H�H���  M���\  H��   H���  E1�L���   H)�K�|= L9��=  L��M��-�  L��  L��  H��L��[]A\A]A^A_�f�H�;1��f�������   H�C0    H���  �C8 H�C@    ǃ�       �CT	   H�C    Hǃ�      H��   H���  1��    H9��0���H���  H��   H)�H)�H9�HF�H�H�H���  H���  H)������I��L�{A���  �6�    1��   L���q���H=�  v/H���     H��   �����I9�u�1�L��L���?���L9�sZE1������f�H��I�I)����  H��  L��H�{L���  �   ����H���  H�,H��   H���j������� L��  �5���@ ��G�H��H	��FH��H	�H9��H9Ѻ   G���    L�E1�I9�sUH�B�I��H��"wHAUATUSA��Cը�ugM�HL9�tQA�H�Aը�tE��-������H�I��L9�wOD  L�� L���@ E�����L�LE�L��H�؄�LE�[L��]A\A]� ������M��1�H�I���� ��   ����   ����   E1�E1�H� 6     �=f�A�   I��L9�v�A�	I��A�    I��A����!ECń��f���E���]������I ���N���L��M9��A���I9��u8��M��M��D  A�6  E1�E1�I���l��������L�E1�����f.�     AT�
   I��USH��H�H�|$H�\$�n���H�L$H9�t9H9�rI�$H��[]A\�f��9#u�H�YH��H�|$H�\$�5���H�L$H9�u�H��1�[]A\�H�H9�sWH�6     �@ H��sAH��H9�s8��� v��%u+H9�w��D  ���tր�
t�H��H9�u�H��H9�r�H��ff.�     f�H�H9���   �E1��@ <(��   <)��   H9�sC�H��H�Q<\u�H9�t0�AD�@�A��Lw2E��B�$� I fD  H�QH9�r��    �   H���    H9�v�HЀ�w�1ɐ��H����w�H9�������D�@�A��v��y���f�     A���_����    A���N���1��H�ʸ   ��     H��H�I��I�� H��H�T$L9�s7L��H�|$�u���H�T$L9�s �
�ȃ�߃�A<v̍A�<	vŸ   ��>uH��1�I�H���ff.�     f�SH��H��H�H�T$H9��  I��E1��<�    <%��   <(uLL��H�|$�_���H�T$����H��H�T$L9�sA��t=�<<tLv�<{��   <}uA����   @ H�T$�   1�H��H�T$L9�r�E�۹   E�H�H��[�f�L��H�|$�����H�T$������    I9�w� f�     �<t<
tH��I9�u�L�ҹ   1��H���D  A���o���H��1�H�H��[�1��ff.�     �UH��SH��H�_H�H�|$H��H�D$�����H�T$1�H9���   �
�q����   ��   ��{��  ��(��  ��<�  ��>��   ��/�?  �� wH�6     H����   H�     � PH�rI�6     �ȃ�߃�[������>wH��H���	Є���   H��H�t$H9��H  �H���� w�I��H�rs�1��fD  H��H�T$H9�vH9U �   D�H9�sH�] �EH��[]� H�\$�EH�] H��[]�D  H�JH�L$H9���   �z>t/H�ʸ   �fD  H�T$1���    H�JH9�v�z<uH��H�T$�l��� H��H�|$����H�T$�R����H�rH�t$H9�si�JH������fD  H��H�|$�����H�T$����f�     H��H�|$�s���H�T$�����f�     H�ʸ   ����� 1������H��������H�w������    AUATUH��SH��H���F    H�    H�F    H�w����H�L�gH�D$L9�sX���[��   ��{��   ��(tNH�E �8/�����D@�E�M����SH����?  H�EH���     H��t@H�H��[]A\A]�D  �E   L��H�|$H�E �p�����uHH�T$H�UH��H��u�H�E     �E    �f.�     �E   L��H�|$H�E ������t�H�UH�D$�v���fD  H�PH�E L���E   H�H�T$����H�H�D$L9�st�wA�   ��t7�eD  ��]t;H�H���P���H�sH���D���H�H�D$L9�s7�K��u0���[u�A����f�A��u�H�PH�UH�������f.�     H�U������    AWAVI��AUATI��UH��S��H��X�����H�t$�����|$ tH��X[]A\A]A^A_ÐI�D$M�,$H�D$H�[M�<�H�D$H�PH�D$I�$H��I�D$H9�swL���0D  M��tI9�vH�D$@foD$0H�CH��I�D$I9$sH�t$0L���x����D$@��u�L)�H��ië����E H�D$M�,$I�D$H��X[]A\A]A^A_�1���ff.�     @ H�w�����H�w�n���ff.�      AVI��AUATUH��SH�wH������1�L�H�OI9�s/I��E��t0A�:<�  I��L9���   H�    I�z1�I�9[]A\A]A^�H�D)�H9�HG�H����   1�E1�   1�I�6     1��I��s�}H��H9�sOL�I���7@�� v�@��x>�����I ��w/��	���t�A��A��}�   D��H��I��H9�r�@ L׃�t��E�eA�L�#E��u5I�91�[]A\A]A^��    H�D)�H9�HG�H���@���H�    ��I��M9Q����A�:>�����[�   ]A\A]A^�H�    L���ff.�     @ �G    H�wH�WH�7H�O H�G(�E H�G0��E H�G8��E H�G@`�E H�GHp�E H�GP�E H�GX��E H�G`��E H�Gh��E H�Gp��E H�Gxp�E HǇ�   ШE HǇ�   @�E �ff.�     �ff.�     @ H�GH��t&H�W �o��   �oJ��   H�R H���   �H�G(H��t7H�D�@f��~0H�pH���LN���A��9���   fA���? ��    1�f��u�fA��~�M��H�xHc�M��H��I��H�J�|�L�L9t$f��~��p�~���9�t9H�@f�|P���    H�H9~u�H�pB�|�u�A��fD�@��    ��f�xf��D  ��f�ÐH�GH��t&H�W �o��   �oJ��   H�R H���   �L�G(���    I�@t-H��
H��H��
I@H��Ix��H�W��H�7�A�@��fA�@��     H�G(H��tfH�f��~]H�pH���|V��P��f��~/L��L�@Hc�M��H��I��L�O�D�M�L9t-f��~�P�r���9�t:H�@f�tH���P1�f�����f�M�XL9^u�H�pB�|�u���f�P봐��f�pf��D  H�GH��t&H�W �o��   �oJ��   H�R H���   �H�7H9�sF��H9�HF�H��t8��E1�1ɐH�A���A��A1��i�m�  D�A�II���X  ��H9�r�É���1ǉ���1�����1��f.�     �G(    H�G0    H�G     H�G    �H�H��  ���  H���  �O(H�G0H�B(H�G H�B0H�G1��ff.�     @ H�H��  ���  H���  �O(H�G0H�B(H�G H�B8H�G1��ff.�     @ H���,  ��0  H��8  )щWH�G 1��O�ff.�     H�G    H�G     �ff.�     @ �W1�9�wW9�v
H�G ���p�D  �D�O�PD9�AB�DOD9�sEH� ���G��u*��H��H�<W�D  D�H��E��u����A9�w�1҉�@ D����1�1���ff.�     �H���  ��H���f�L�H��E1���E I��  A���  I���   H�@���    H�H��  �` H�H��  �` ��L���   H���  Ǉ�       H�L���  H��x
  H���  H���  H���  H9�vwM��A������L�^<��   <s[<vc<��   <u_L�¸�   L)�H���B  Ǉ�      I�@�HG@I�@�H�GX    H�GP1��D  <s�H��w��   �fD  <s�<t�<v���<���   ��u���L�����- <v�<�u�H�NH9�r��Fȍ� }  �� �  w���H��L��L)�H���  �I��H�I�@�L���  H9������t����     L9��c����~�Y���L�¸�   L)�H��U� L�^L9��7����v<�w���   ���DlL���F���fD  ���   ���1D��)Ɖ�L���%���D  �Ǉ�      I�@�HG@I�@�HGHI�@�H�GPI�@�H�GX1��f.�     D�G E����   � ��   �G$A����PH��H��9t8��D9�r��tC��H��H��D�D8D9���   ��H��H��H�L8�D  H�� D�A A9�~{���Ѕ�u�O8���W<�G$    )�H�9�K1�H��Hct@H��H��H��?H�� �  H����fD  HcGHc�H��H��H��?H�� �  H��ÐHcw�f.�     �щG$H��D)�H���T<Hc���     ATI��USH�����t�I�����   1��fD  I��1�E�Q E��E���g  A�y8A�s9���   I�IX1�� H�� �y�9���   ��D9�u�I�y� t
A���   A�B�H��A�D<A9C|[A�q A9��  E��L��H��A�D<����  A9C1�~����   w&��A��D)���   �     �   �F9B�<���H��[]A\�1�@ 9�t��t9z}��H��H��A�D	u�I�y� tlA�ufA���O  rH�T$�����������H�T$�J��A+s�����Icq��Hc�H��H��H��?H��1 �  ��H���)�A�s�BD�Ѕ��-  E�A D��E1�A9�������~�A���tA������   �%���D��E��D)�t=��)�)� ���>��H��H��H��H��L�L��oA@�oIH9�u�I���AoI��K�P�Ao[XA�D$A�A �������A�B�o"A��H��H��L�`�ojhE�a H��[]A\� �~�9B�6����h���H�T$�]���H�T$A�CD�������I�y1�� �����E�A�������A�s�h���A������ff.�      L�SD����)�)�L�T$A��4   ��   A��A)�D��A��E)�E��A�    A�    ���H   t~����L�_��������)�AC ��xwE���  C� 9���   �Hc�I  D9���   Hi�3�  H�H�� �  H��A�Hc�I  Hi��L  H�H�� �  H��A�[��    A�����X���fD  ��E��xiC� 9���   �Hc�I  D9�|jHi�3�  H�H�� �  H��A�Hc�I  Hi�3� H�H�� �  H��A�[�fD  A�    A�    [�A��C� 9�|M�Hc�I  A9�~W��A���I  A�[��    A��C� 9�|��Hc�I  A9��Hi��L������� A�    ��I  �A�[�@ Hi��L���<���@ �ﾭ�H9Gt�@ USH��H��H�o8H�7H���h)��H�    H�s(H���U)��H�C(    H�s0H���A)��H�C0    H�C    H��[]�f.�     USH��H�GH�/H��t&H�W �o��   �oJ��   H�R H���   H���  H��t&H��H���  ��H���  H����(��Hǃ�      H��[]�ff.�     @ SH��H�wH�?�(��H�C    [�fD  SH�H��H�w H���   �i(��H�C     �C    [��     ATUSH��L�'M��t#H�o8H�wH��H�T$H�������T$H���tH��[]A\�@ H�SL��H���,�  H�C(HcS H�3H��L)�H9�s!f.�     H�H��tH�H�H��H9�w�H�CL��H��H�C�'��H��[]A\�ff.�     f�AUI��ATI��UH���    SH��H��H��H�T$�X���H�D$��u)L�bL�"L�j�B   H�+H�SH�C    H�C    H��[]A\A]�f�     AUE1�ATLc�   UH��L��SH��H��H�W81�H��L�L$�����T$H�C(��t#H��H����&��H�C(    �D$H��[]A\A]ÐL�L$E1�L��1Ҿ   H�������H�C0�D$��uZ�ﾭ�D�c H�K�C$    H�    H�C    H�C    H�C@��E H�CHp�E H�CP��E H�CX0�E H��[]A\A]�@ H�C(�T����    H��������AT1�USH��H��H�O�D$    H��H9�s%H�S1�H��t�
��u�@   H��[]A\�D  H��H�W0L�G8I��H�?L�L$�   H��������|$H�C8��u�L�c�   H�k0L9c(v�H�CH��t�0��u� �   L�c(H��1�[]A\�f�     UH��SH��H��H�(H;{t*H�SH��H��H{8��  H�C(H��[]�f.�     H�s H�H���������t�H�{(��    AVAUATUSH�o(���    H�Eu��f�E[]A\A]A^�fD  H��I��HEA��I��H��I��Lm�P���L��H��I�E �@���H��E��I�E������E��f�E[]A\A]A^�f�     AWAVAUATUSH��8H�/H�l$(H9��Q  �E I��I��I���PՁ��   �  E1�<.�
  L��H�|$(L�D$�h���H�L$(H��H9��  H=�  A�   L�D$�8  L9�s	�9.�g  A�   1�H�QL9�s����<E�#  H��1�H	�I�H����   E���f  @����   M���^  H������G  H�gfffffff�8 I���.  L��I��?H��H��L)�I��I����  H������  H��H�H��H������H�l� H���fD  H�MH�L$(H9�t�U�rՁ��   u 1�H��8H��[]A\A]A^A_�@ <-A�ǀ�.�f  L9���   E1�1�A�   1������fD  ��E1�L9�����������@ L��H�|$(H�T$(H�T$L�D$D�L$�����H�L$(H�T$H9��l���H��D�L$L�D$H	�H=�  �o  I�H���C��� ����H��H��E��HE��+���H��fD  E1�1�H�MH�L$(L9��'����U�� �o  �B�<�B�@��<��@�� ����������H�EA�   1��P@ I��H��H�D$(I9��������� �  �r�H��@���r�@��@��@��@�������������H���I ��	��   I������H������H�L� H�,JH��u	M���z���O�$�M��r���ttH�����������     O�$�M�H	�����I��tJH��H��H��H��H��I�����~�H��H��H��H����f��   H=�������I�1��
���D  H���|���L��H���l���H��i���H�L$(�����H��1�H	������H��A�   1�1������H���X���H���A���ff.�     AWAVAUATUSH��8L�?D�D$E1�H�|$�T$L�|$ I9���   A�H��I��<[��   �}   <{��   I��L�|$ I9���   E1��nf.�     A8/��   M��tD9t$~rM��O�D� H�D$(H��HcT$IE�H�|$ I���E���H�T$ I�$I9���   D�D$A��@��t]I��H9�sTH��H�|$ D�t$E���7���L�|$ I9��y���H�D$L�8H��8D��[]A\A]A^A_��    �]   �-���fD  I���� 1��*���f�     I���f.�     A������E1�� H��A��H�wI��A������H�wL��D��H���w����    AWAVAUA��ATUSH��H��   H�t$H�t$pH�|$0H�T$������$�   ����   H�T$p�KL�t$xH�T$h�L$ ���R  �D$    �D$$   ����  B��    D�d$H�D$8C�D- �D$@D�D$XA�E��D$D�    H�t$H�L$D��H�|$h�YH�L��������D$ ��w�$�h
I �    �   H�ĸ   []A\A]A^A_�f�     H�D$0H�L$8E1�1�L�L$d�   H�@ H��H�D$H�����H�ŋD$d��u�1�A�   ��E1�D��L��H�L� H�|$h��������  D9���  L��H�|$hD�����A��u��D$DE1�H�D$(E����   L�t$PL�t$D�d$\M��D�|$X�@ I��J�|� K���}��H�C�D% H�|� �}��H�C�D$@D�H�|� �}��H�CC�'H�|� �v}��H�CI�D$L;d$(u�L�t$PD�d$\H�|$HH�������mD  E1��   H�|$hH��$�   �.����������H��$�   �}��H�H��$�   �}��H�CH��$�   ��|��H�CH��$�   ��|��H�Cf��D$$A��D$A9�����1��9���@ H�|$h�f���H�t$�V��tc���O  ���6  H�뱐H�T$hH�BI9�v	�:t��  H�J1�I9�v�:fu�za�-  �    H�t$H�T$h�V��u�f��]���D  �   H�|$h�����n���@ H�D$hL9��2���H�T$0��$�   H�J L��H)�A�׃���   ���W���H���j�D�z�H�D$hH�3H��tH��H�L$(�B��H�    H�L$(H��D��H�T$d����H���D$d������H�t$hH��H���2�  �( H����� 1�H�|$h�\��������    ��y���f�     ��i���f�     E�������H��D�l$$I�^�H�T$hI���D$   ����D  H���j�H�D$h�(����    1��zr������zu������ze�����H���   �r���f.�     L�|$0H��I�^�H��$�   M�'I�oI�L��I�_�������$�   M�'I�o�D$    �D$$   �w���E�������H�D$h�D$    �/���@ H�|$HH���D$d   ����D$d�����zl������zs������ze�����H������ff.�     AWI��AVAUATA��UH��SH��H��H  �o�oN�oV �F)D$)L$ )T$0�D$   ��
��   ����   H�L$�    H�t$@L��������D$����   �S 9���   �{M�7M�ot�S$����   H�\$@��&�   D  �D$,D$(H���D$���D$��~tH�E1�D��H��H�t$L��I�H�CI�G������t�M�7M�oH��H  []A\A]A^A_� �ЉT$�j���D  H�M ��D$�m����D$   ���� 1��@ ��   묐AWE1�AVI��AUATI��USH��(�t$H�w����H�L�oH�\$I9���   �<[��   <{��   �D$}H��H�\$I9���   L��E1��^D  �D$8��   M��tD9|$~W1�L��H�|$����H�T$H��M��HE�f�H�D$H9�t{A���|$ tHH��I9�v?L��H�|$�����H�\$I9�w�I�H��(D��[]A\A]A^A_� �D$]�O���fD  H���� �D$ �I���fD  H���f.�     A�������     E1��ff.�     H��A��H�w�p���H�wIc�H���0���H�    I��H�1�H�G`    L��H���L�V0H)�L�N8��p���H�H�~@H�NPH�F`L�M�L�^M�XL�^M�XL�^M�XL�^ M�X L�^(M�P0M�X(M�H8I�x@I�HHI�@P��t;A�@X ���   A�@Y���   A�@Z���   A�@[A�P\I�@` �E I�@h�E ����   A�@X���   A�@Y���   A�@Z���   A�@[�f�ATf��UH��SH��H��))BH�H���   H�xh t5H�L$H����x  ��uH�$H�L$H�H�SH�KH�SH��[]A\�f�L��  I��$    tG���   w?I��$h  ���A�L$$��t*I��$   1�H�Wf;u� @ H��f;B�t��9�u�   땅�x�H�}�^��� f��SH�Ћ\$))GH;V(rL�V1�M��tE�E����   H�FHF8D�XD�PD��D)ց�  ����   ��  ��tM����   ����   �   E�ھ   ��0  D�OH�WE�HE�D�G�8 t/�@���G[�7�@ ����   DG�    D�GD�OH�WMc�Mc�[M��L��H��?I��  �  H���G��     ��t��   �   E�D�OD�GH�W�8 t��@��     A��   ����@ �   E�Ӿ   ��   �   �)�����t�   �   ��    �   �   �����     H�|$�H�zH��1�H���H�T$�H)�H�    ���  Hǂ�      ���H�H��P  ��HǂH      Hǂ      H���)���   ���H��~@��H  ��t�     H�LFH���P  H��9�w��~	1�@��I  ��tf�     H�LF(H����  H��9�w��~
1�@��J  ��tf�     H�LF<H���  H��9�w��~1�@��K  ��tf�     H�LFXH��  H��9�w�H�FpH���  HcFxH���  HcF|H���  ���   H���  ���   H���  ���   1�@���  ��t"f�     H��F�   H���   H��9�w����   1�@���  ��t H��F�   H���h  H��9�w����   H�L$����  �F���  H���   ���  H���   H��  H���  H�D$�H���   �Vt���t.���  ��t.@ ����1Љ���1Љ���1�x�Vt�D  ���  ��u1H�T$�H�D$�1�H�T$�1Љ���
1�����1�9¸�s  EƉ��  �ff.�     �U1�SH��H��H�G�    H��HǇ�      H���H)����  ���H�����   H���������H���  H��(  H���
  H���  ���
  ��h  H���
  H��`  ��h  ��l  H��`  H���  ���
  ��@  H���
  H��P  H���
  H���  H���
  H���  H���  H���  ���  ���  ���
  ���  []�f.�     H��1��&���H���   H��  H�  H��(  H���  H��   ���  ��D  H���  H��X  ���  ��L  ���  ��@  H���  H��P  ���  ��H  H���  H��0  ���  ��8  ���  ��l  H���  H��x  H���  H���  []�ff.�     SH�_(H��tn���    t=H��W�G`�D;Gw8H�f��~�sH�K�V�f�TA����f�1�[�f�f�1�[��     1��   �������t�[�fD  �   [ÐS���    H�_(tbH��W�G`�D;Gw-H�f��~�sH�K�V�f�TA����f�1�[��    1��   �d�����u�H�f�����D  f�1�[��     AUATUSH��H��Ƈ�   H���   Ǉ�       H�wH�OH�H��t\H��(  I��H��E��H�8H�GH�{H�C H�G`H�C(�x��I�EPH� Hǃ�       H���   E��tH��(  H�@@H���   H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    Hǃ�   ��E Hǃ�   ��E Hǃ�   ��E Hǃ�   ��E Hǃ�   ��E Hǃ�   ��E Hǃ�   @�E Hǃ�   ��E H��[]A\A]�ff.�     �AU�   ATUSH��H��f���   H���   H�wH�OH�H��tuH��(  E��I��H��H�8H�GH�{H�C H�G`H�C(�Tw��Hǃ�       Hǃ�       E��t.M��t)I�D$PH� H��tH� H���   H��(  H�@@H���   H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    Hǃ�   кE Hǃ�   ��E Hǃ�   `�E Hǃ�   �E Hǃ�   ��E Hǃ�    �E Hǃ�   ��E Hǃ�   @�E H��[]A\A]��     H���  ���   ��   AUHc�ATUSH��H��H�P0�<r�P(I�ŋ�h  ��tUH��`  D�`�1��fD  H�CI9�t7H��H�|� H��t�A�E 8u�L���'B ��u�H����[]A\A]��     H�������[]A\A]ø�����f.�     AW1�AVI��AUI��ATM��UL��SH��H��H��H��H�T$D�|$P�   H�G�    HǇ�      H���H)����  ���H�H���   ��BH �4���H����   H���
  L��L��H��H�T$E���M���I�E L���
  H��`  ���
  �D$XHǃx  ��E ��h  H�D$`Hǃ�  ��E H��p  1�Hǃ�  p�E Hǃ�  `!F H��[]A\A]A^A_�f�H���   []A\A]A^A_�ff.�     �AV�A   1�AUI��ATI��US�/�0I ������IKHc�H�<��I ��XHc�@8�u��    L��L��D�s��A ��t�؃�I�H�<��I H��@:/t�A�K   [D��]A\A]A^�ff.�     H�OH�f�     H9�w������G   �fD  H��H��B��� t؃�	tӃ�t��
u	�G   Ð��;u�G   Ã�t��ff.�     f��W��YH�������G��JH�H�H�B�H9�w
�F   �f�H�JH���� t��	t��t��
t��;t��t�H���� 1��D  �F   ��F   ��     �WH���������W1���?H�H�~H�B�@ H9�w�F   � H��H��J���t��
t��u���@ ��    �F   ��     AWAVI��AUA��ATU1�SH�^H��(L�g�K�L�����   �_���H�D$H��t?M�<$I)ǃ{�I�O�wT�S��$հ
I f.�     1�H����   ���H��A9�u�H��(��[]A\A]A^A_�D  H�4H�|$�������H��A9�t΋K�L����r����Q���H�D$�m����    M�FM����   I�V H��H��A�Љ�f�H�41�H�|$�`���H�� I�>H�T$L��H�L$������T$H�L$H����o���H�t$H��H���ڨ  H�B�D8� �Q����H�ƿ9I ��� �������D  �    �%���D  H��t;H�D�Gf��~4H�OH���TQ���A��9���   fA���C�    ��    1�f��u�fA��~�M��H�wHc�M��H��I��H�J�t�L�L9t$f��~��O�q���9�t9H�Wf�tB���    H�vH9qu�H�OB�|	�u�A��fD�G��    ��f�wf��D  ��f�ÐSH�_8H�{(�����CX [�ff.�     �ATUH��SH�GH��P  ��0  ����   H��h  H���  H���   ���  H���  1����  ���  t�k   ���  v��l�  �%k��� �  ���  H��   H���  H��  H���  H���  1�[]A\�fD  H��h  I���H��8  �P�и   ;�0  s�Hc�H���    H���8  �@���M���7���I�L$PH�	H�D�H���   �����    I��UMc�H��Ic��H  I��Ic�SIc��H  H��D��L��H��L��H��H��?I��  �  H��?H��H��
 �  H��H�������Hc�I�H�HcqDHcQLH��H��H��H��?I��H��> �  A���H  I��?H���J�� �  HcQHHcIPH��H���H��Hc�H�u H��H��?H��H�� �  A���H  H��?[H��]�H��1 �  H���H�I��f.�     AWAVAUATUH��SH��H��   L�?H�4$H�L$D�D$ D�L$$E��uH�� �@  H�$L�p(H�D$�x ��  H�D$H�C     �oh �o�oX)�$�   )�$�   )l$)�$�   L9p�  A��A   ��  M���`  A�����1�L��$�   �,fD  H��A���H��u
I��A�����H��L9���   E�e t�H��D�KL��H��jD�D$0H�t$H�|$P�H���D�D$0H�t$L��D�KH�|$p�$    �&���D�\$PAYAZA��u�D$`�D$����  H�T$`H�t$@H������D����A E �L���@ H��H� H��t�(��u�    �y �����A� t
�     �C H�ĸ   []A\A]A^A_�@ �|$$ ��   A�����1�L��$�   �) H��A���H��u
I��A�����H��L9��r  E�e t�H��D�KH��L��jD�D$0H�t$H�|$P�(���D�D$0H�t$L��D�KH�|$p�$    ����H�T$pH�t$PH������XZ�u���D  �K ���]  �{8���R  �A�H���t8���?  H�CH�@(     1�fD  L�mI��L��H���D;A��A��tM��H�� L�m��Z  H��   �    A�    H��D�L<L��H��E��D�T<D)�E��E�A�º   )�AD�9�N�A9�AN���A��A��I9��F  L��A�� �  H��9L3<�-  H��tH�M�� ���)�H��D�9t<�L  E��9�}�D;(�K  D��H��D�H���t<E���@  L��H��D|<H����  L��I��H��I��H�I܋p8A�T$89�t)֋x<A+|$<Hc�Hc��a��A�D$@�C L��H��L9������L�kM�](M����   M�eI�{�I�m8L��I��H��    H��H��I9�w$I�EH��H��tD�0E��u� �   f.�     H�
D�BH��H�AH��H��H�H�D�J<E�E�� �  D9P<|D�J<�@tH��H��DD<L)�H��u��|$$ ��  H�D$�C�@	 �����@ �Cf��H�T$`H��H�t$@D$DH�D$T    �D$\    �D$X�D$@1   )D$`)D$p������K H�CH�@(    ���t����f�H��t6H�M�H��H��H�L�<�u8A�G89�t)Ƌ}<A+<Hc�Hc��_��A�G@E���A����w����    D��H��tHH�M�� ���I��)�I��D�B9|<~,H��A�H��D�L<E��t�L��H��T<�q����     9�AO�A������f�H�������G���f�A��<  A��L  �������D�T$pD�L$PD��L�l$(D�D$D�\$4I���  ��D�T$<E��E��D�L$8A��
�=fD  ��t$D�A)�E9�D�HF�E9���  �     ��H��9���  �x u�E��t�D�E��A)�E9��D�PA�E9��A��@   L�l$(D�\$4�L$t��  ��H��A����  ��)�E����  �D$t�D$���D$`�]����H�M(L�H��`�o���H�D$H�qA�  H��H�HH�pfD�XH��t;H�D$H�� H�0H��t�     � �H��H9�u��ٸ��������H�L$ D1H�$L�p(�����f��K H�CH�@(    ������f�     D�S E������H�S(1�H�<$��    D�@� �C H�� H9�������2H��@�� u�H�BH;G(r#L�G1�M��tE�E��uA� �   �2�    H�GHG8��
D�Bu�D�@��     L�l$(����fD  f��I��x  H�T$`H��)D$`)D$p����I��X  H�t$`H�������,���D  H�f��A�   H��$�   �$�   H��$�   H���$�   HǄ$�       �?����z���f.�     E1�E1��D;(�����H�{D)�H�t$`L�d$`�T$h�����H��H���t<����D  �|$$ �K �]����`���A��@   L�l$(D�\$4�L$Tt=��H��A����  D�D$��A���D$T)�D�\$@E��������L$t�
�w���@ �� �  D+L$8f1�E;�H  |���H��A����  ��   9�O�럋t$<�� �  f1�D)�A;�H  ������H��A����  ��   9�L������A��T$TD�\$@�u���f�     H�H��t���u� U   1��f�     H�GH��t���u� �   �f.�     �O H�WH�GH��H9�t�0H���@�   H�G�f.�     �ff.�      �O H�WH�GH��H9�t�0H���@�    H�G�f.�     �k���ff.�     H�GH;GtFH�P�H�W�P��@���t������D���    ��x    ��� �    )�����ÐH�W1�H��t�
��u���   ��     H�WH�GH)�H��9�s-��H��P� ��t������D�Ð��x,    ��� H�W1�H��t�
��u���   ��     �    )�����ÐH�WH��H+GH��9�w��H��H)�H�W��    H�GH��t���u�� �   �f�H��tKUSH��H��H�/H�wxH���c���H�Cx    H���   H���L���Hǃ�       H��[]�f.�     �ff.�     @ AWAVAUATLc�USH��8E����  H���   D9g �J  H�A��H�]I��L�u J�/H9��  M��M)��9  L9�H������LF� H��H��H��   H�� ���H9�w�H�E8H�T$,H�މL$L�L$H��H�D$�[���L�L$�L$H��H�E �D$,����   M����   H�UL���L$L�L$�l�  H�E(HcU H�} L�L$H�4ЋL$L)�H9�sH�H��tH�H�H��H9�w�H�|$L���L$L�L$�����L�u L�L$�L$K�I���H�]H�}LE�H�E(I�L��L��N�4�H�E0H} B���ۗ  Lm1�H��8[]A\A]A^A_� I��� I�����������@ H��8�   []A\A]A^A_�@ L�u H��8[]A\A]A^A_�D  AWM��I��AVAUI��ATI��USH��(L�JL+JI���l$`D�˃�@��u��uwI���8   uS��E��A9�v>��L��������s��ŉl$����H��L���$ H�D$    ŉl$�G���A9�w�I�D$I�D$A�H��([]A\A]A^A_�D  A�? u�H��1��`���I�H��   H��  ���A��^���f�AWL���I  AVAUI��ATL���I  USH��H��xD��|I  H�t$H�L$L�D$D�$A��tL���I  L���I  I�I�M I�WI�}H9�uH9�t{I�,$M�T$D�D$D�L$)�D)�A)�A)�������A��A����A��A��H�Hc�Mc�Mc�I��I��H��I��H��?I��?H��0 �  J��2 �  H��H��)���  E1�1��o�XI  )D$ A���0  E1�A����   H�D$ �<$ M�MH�L$8M�E H�T$0H�$��  H��H��8  �����H�$H��XI  H9|$0��  �o�XI  H�S�D$`   H��)L$ H���RfoT$0�XI  E����   H��x[]A\A]A^A_�f�A�   E1�L�t$D���I  H�L$8H�T$0D���I  H��D�\$L���D$`   �2���H�L$HL��H��D���I  D���I  H�T$@����H�L$XL��H��D���I  D���I  H�T$P�����H�CH�t$ H���Pfod$PD�\$�XI  E�������I�m M�eH��x[]A\A]A^A_�f.�     )�D)�Hc���������Hc�Hc�L��L��L��L��H��?H��?I�� �  I�� �  H��H��)�Hc��NS��I�7M�$H�M�L$��D)�Hc�H��H��H��?H��
 �  I�WH����B�,D)�Hc�Hc�H��H��H��?H�� �  H��F�$Mc�I9�u����1�)�9�$I  HO�I9�u����1�)�9�$I  LO�I�E H9D$u���)�)�H�9�$I  HO�I�MH9L$uD��A��E)�)�AH�9�$I  LO��H��D��|I  �������Hc�)�H)�H�H��HH�Hc� I  H9������L��������Hc�D)�H)�Hc�H��HH�H9������I�/M�g�o�XI  )\$ A���>  A��A�   D�$���������@ A�   E1�H�D$ �<$ �D$`   H�L$8L���I  D�\$H�T$0L���I  H�D$��   H�t$H������D�\$H�D$H�|$0H9|$ ��   H�SD�\$H��H���Rfol$0D�\$�XI  ����@ H�t$H���;���H�$H��XI  H9|$0�l���H��`I  H9t$8�Z�������fD  H��H��8  �����H�D$D�\$H�|$0H9|$ �h���H�t$8H9t$(�X��������f�     D�$A�   �����SH��H��H���   H�@hH��t8H�xH� H�����u!H�$HcT$H�    H�CH�CH�H�C1�H��[ÐH���  H���  ��H��Hc���fD  S��pI  H��Ƈ�H  ��hI  �  ��xI   u1�ƃ�H  f���H  ƃxI   [�f�H��8I  L��@I  H�sH��H��(I  A�   �������    ATA��U��S���H   H��u{Ic�HcՀ{( ƃ�H  H��hI  H�� I  H��HI  H��pI  H��PI  t
�y	 H�kt$H�kH���H  E1�H���H  D��I  H���W���H��8  H��  �H�[]A\�������{���fD  ATI��UH��SH��H��P�o�XI  �( �D$@   )$tUH�L$H�T$A��E��H�sH�������H�CH��H���foL$L��(I  H��0I  �XI  H��P[]A\�f�     ��pI  ��hI  ������ff.�     f�AWAVLc�AULc�ATM��UL��SH��(H�� I  H��PI  H��HI  �x	 ��   ���H   ��   A�   H�D$D��A��H��PL�L$�+����L$�D$��HI  ��PI  �A��΀��H   Mc�Hc�Hc�Hc�H�t$H�T$ X��   ��xI   ��   foD$ƃxI  ǃ|I     )��I  L���I  H���I  E��u<L��HI  L��PI  H��([]A\A]A^A_��    E1�I9��8���L9��/����ӐH�� I  H�{E1�H���H  H���H  D��I  �H����fD  H�sE1�L��I��H�T$H�������D���������ƃ�H   ƃ�H  L��8I  H��@I  ����f.�     AWA��AVMc�AUA��ATA�̉�UD��A��SH��H��H��PI  ��HI  H�D$$PL�L$(诿��H�D$4��D��PD��$�   D��L�L$8菿����D��D��D)���H�OD�\$8������D��E�E�D)�Mc�Mc����֋�HI  )Ћ�PI  A �D$4�L$0�AǋD$<�F�)Hc�Hc�Mc���$�   ���H   Mc�H�t$@Hc�H�H�T$HYAX��   ��xI   ��   foD$0H�� I  ƃxI  ǃ|I     )��I  L���I  L���I  L���I  H���I  L���I  H���I  �y	 ��   Lc�$�   L��HI  L��PI  H��H[]A\A]A^A_�H�D$L�\$L�T$�,���L�T$��xI   ƃ�H   ƃ�H  H�D$L��8I  L�\$L��@I  �6���L��H�sE1�M��H�T$0H��H�D$L�\$L�T$�����H�D$L�\$L�T$������    H���H  H���H  H�{E1�D��I  �����%���f.�     AWE1�AVAUI��ATUH��SH��H��XE�`	D��H�$E��D�\$A�ǉD$E1�1�A���D  I�BM9�t4D�\�I��C�< F�\�t�H��D�v�o���D��A�I�BF�\�M9�u�E���  D�t$<E����   A�E D�|$8E��H�߉�E��D)�A)��E DHʉ�D)�A)�DH�����E9�}A�M F�$0�L$H���D$4PD�L$8D�D$4�L$0�T$,�t$(H�|$����D�L$E��D���T$D�t$@D�$$H�|$����H�CH�C�D$A�E D�e H��h[]A\A]A^A_�@ D�D�e �D$����A�x
 u9A�E A�x �D$@uL�D$@D�e D�|$8�D$�S���@ D�u ������    D�T$8H��D�N�/���D�A�x D�ΉD$@t�H������D�|$8E�$�D$@�D$�����H��G�Wb��;Gw1���     1��)���f�     ��t��f.�     1��ff.�     f�ATI��UH���   SH��H��������tH��[]A\��     L��H��H�߹   �D$�y����D$H��[]A\�ff.�     ����   u1��@ ATI��UH��SH��Ǉ�      �4�����t[]A\� L��H��H��[]A\�V���fD  H�?�G�Wb��;Gw1��f�     1��)���f�     H�O(�Y H�At%H��
H��H��
HAH��HyH�7H�W� �A��f�A�@ AUATUSH��H�o(�GXH����   �Y I��I��H��tvH��W�G`�D;GwqH�E f��~�uH�M�V�f�TA��E ��f�E H�{�   ������uL��L��H�߉D$�8����D$H��[]A\A]�f�     f�E �f�     1��   �$������{�����f.�     H���   []A\A]�ATI��UH��SH�_8�{X uH�VH�6H�����������   H�{�   �w�������   H�C(�{Y H�Pu ��f�PH��f�Bf�@[]A\��    H�uH�}H��H��HPHHH��
H��
H�9H�q��KYH�S(f�@����   H�BH�u(H�} H��H��
HBH��H��
HJH�9H�q� �KYH�C(f�B���n���H�PH�u8H�}0H��H��
HPH��H��
HHH�9H�q��;���@ I�T$0�
���-����[]A\�H������f.�     H��G�Wb��;Gw1���     1�鉻��f�     ��t��f.�     1��ff.�     f�ATI��UH���   SH��������uDA��$�    I�t$(H�Vt(H�NH��
H��H��
H��H~H�H�/H�_��V��f�V[]A\�ff.�     ����    t1��@ ATI��UH��SH��Ƈ�   ������t[]A\�fD  L��H��H��[]A\�F���fD  AWI��AVAUATE��USH��(H�D$`E��u*�E��A��E�A��A�E�H��([]A\A]A^A_�fD  D�Hc�Hc��Hc����0D�@H�у�D�HH��H��?L��
 �  �   I��A��)�A�̓�A)�D��-��   D�ɉ�����9���   D�P�PD�pD�$A��D�P�@A���D$D9��V  D����9���   D��Ic�H��D�L$)�D�T$�D$�C��D�T$HcT$D�L$D��������   A)�D+4$Ic�Ic��B���<$H��I����Hc���B��A�| A�?�    �4Hc�Hc��B������D  IcՉ�H����H��H��?H��
 �  H��9�����A��H��Ic��zB����A�� D����9�}VE)�Hc�H��D�$�TB��D�$E��t;�t$A)�Ic�Ic�D)�A��Hc��OA��Ic�H��I���!B��A�| A�?�L���@ �|$H����Hc���A����A��,���@ ��Hc�D�\$)�H��D�L$D�T$D�D$�T$�L$��A���L$�T$D�D$D�T$��D�L$D�\$�i����4$A)�Hc�D�$Ic�D)�Hc��@��D�$H��I��A��Ic��pA��A�| A�?���� AV��AUATUSH�GH���<p�S �k(��t<L�c0I��D�m�1��f�H�CI9�t7H��I�<܉�H��t�A�8u�L���W ��u�[��]A\A]A^�f.�     1�[��]A\A]A^� ���   w�s��� 1��ff.�     f�ATI��US��X���   w4H����    ����   t��H���+�����t�A�$[]A\�fD  1�1�A�$[]A\�ff.�     L�GI��A�xL���J���A�@    L������H��u%A�xt�M��u	��     1�I��f.�     M��t�H��H��II��ff.�      AWAVAUATUSH��   H�oH����  H�t$(H��L�/A�   �\���H����   H�|$(��   H�ƿ>I �   ��� ����   A��   H�t$(H������H��tYH�t$(H���������1w܉��$��
I �     H�C�   H�t$@H���D$@   H�D$�������,  @ A��   H�u8L���n���H�E8    H�uHL���E@    �S���H�EH    �EP    �E  H�Ę   D��[]A\A]A^A_� E1��� �   H�t$@H���D$@   ������u�H�D$HH�E0���� �   H�t$@H���D$@   ��������S���H�D$HH�E(������    I�      � A�   H�t$0H�������H������H�t$0H����������7������$�pI f��   H�t$@H���D$@   �f����������D�T$H�fD  1�H���v���A��H��t>E����%fD  H�t$@H���3������*  ���!  H�t$@H���4���H��u�A��   ����@ �   H�t$@H���D$@   ��������C����D$H�E ������   H�t$@H���D$@   �D$P   �D$`   �D$p   �����������H�D$HH�EH�D$XH�EH�D$hH�EH�D$xH�E �g���@ �   H�t$@H���D$@   �>�����������D$H�����2���A�   ����@ H�C�   H�t$@H���D$@   H�D$��������\����D$H���P���H�T$�BP��  E1��;D  H�t$8H��������H�A����7����L��H�� @ ��  L���^  H�t$8H������H��u������ A�   ����D  �D$H�������H�T$�B@�  A�����H�t$8H���k���H�������H�t$8H���5�����tv��8t9��Kt����������s���H�D$A��D�`@�9����E1�������     H�L$A��D;a@�=���Ic�H�t$@H��H��H�A8�D$@   �D$P   H�к   �D$`   H�L$�D$p   Ǆ$�      �|�����������D$HH�L$�H�D$XH�AH�D$hH�AH�D$xH�AH��$�   H�A �����H�;1҉�L�L$@E1��(   �3���H�T$D�d$@H�B8E��������}���H�;1҉�L�L$@E1��   �����H�T$D�d$@H�BHE�������H���H�D$D�D$D9`P�.���L��   H�t$@H��H��HHH�D$@   H�L$�D$P   �D$`   �D$p   �|�����������T$HH�L$D�D$��T$X�Q�T$hA��%tN�QA��"uA��u<�D$x�AI������������H�D$Ic��P�E �   D�`PH�xH�=�  �P���1����A    �Q��     ATI��1�E��UH��P  E��SH��H��H�G�    H��HǇ�      H���H)����  ���H�L��H������H��@  ���   H���   H���  1����  ���  t�k   ���  v��l�  �%k��� �  ���  H�D$ D���  H���  H�D$(H���  []A\�f�     H��`wjH�B�  H�WH��f�OH�GH��tGH��tBI��1��H�PH�V� A�D H��I;Hs!H�FH;Fr�H���T���A�D H��I;Hr��@ H�H��t�0��u��    �ff.�     AUATI��UH��SH��H�_8�{X uH�VH�6H��������uH�{�   L�mH�m������tI�T$0�
��u�H��[]A\A]ÐH��L��H��H��[]A\A]�����     H�GH;Gt6�x�t H�W1�H��t �
��u��   ��     H�P��@�H�W�@ H�W1�H��t��2��u���   ��     AWf��AVI��AUATUSH��H�wI��H��hd  H���   L�'�8H�T$`H��$�  L��$�  H�D$HH��   H�L$h�   D��$�d  �|$\H��  H��1��H�D��$�   L�ߺ�I  D��$�   H�t$x)�$�   H��$8  HǄ$�       Ǆ$�       HǄ$�       L��$0  HǄ$@      HǄ$H      HǄ$P  
   HǄ$X      HǄ$`      HǄ$h      H��$x  H��$�  H��$�   1�L��$p  HǄ$�     HǄ$�      HǄ$�  
   HǄ$�      HǄ$�      HǄ$�      L��$�  HǄ$�     HǄ$�      HǄ$�  
   HǄ$�      HǄ$�      HǄ$�      �$�   �$�   HǄ$�       �u  H�T$`�|$\H��$�  H���H  A��   L��$�  H��$�  H��$ K  H��$K  H��$�2  H��$�  A�F,H��$K  H��$�2  H��$�  H�T$h��$hc  A�F4fo
��$K  H��$p  ��$lc  I��8  ��$�2  ��$�  L��$(c  L��$0c  HǄ$8c     HǄ$Hc  
   ��$K  L��$ K  ��$�2  L��$�2  ��$�  L��$�  ��$pc  )$�$xc  H��$�c  A��  H��$�c  H��$�  ��$�c  A��0  H��$�c  H��$�   ��H��$�c  A��,  ����$�c  1ȉ�$�c  )ȉ�Ƅ$�c  ��D��$�c  Ǆ$�c  �  1�)�H�L$H9�L�H��$�d  �A�~ ��$�c  H��   ��$�   H��   ���A�~ ��  H��  D���  D�l$p�(   L��H��$p  Ǆ$p      �|�����$p  I�ǅ�uL� H�D$xI�GL��L��$p  E1�1Ҿ   L��腨����$p  I�G���  �L$pI�GH��$H  A�O �?  HǄ$X     H��$h  foA�VfocH�$)d$`���i  ���D$@    E�f���D$W H�x�D$( -1�D$8    �D$0 Ǆ$�       L�t$��$�   H�H H9���   �|$@ۃ���E��t_�|$W u�؃��<t�C�<�R  f.�     �L$8��t�C�<v���    G��D$8�|$0 t��������!ȃ��D$0����   �l$(�   ���J  ���$�0I E����  �    I�GH�$H�II�GH9��@���H�$H�AH�C���t	���0���H�D$�x �    E�����@ �D$@���$  L�t$A�   E�nH��$`c  H��$(c  HǄ$@c      HǄ$Pc      HǄ$Xc      �\���H��$�  H��$�  HǄ$`c      HǄ$�      HǄ$�      HǄ$�      ����H��$�  H��$p  HǄ$�      HǄ$�      HǄ$�      HǄ$�      �����H��$h  H��$0  HǄ$�      HǄ$H      HǄ$X      HǄ$`      ����HǄ$h      M��t"I�I�wH���m���I�G    L��H���Z���H��hd  []A\A]A^A_��     A�0   �D$p0   �q���D  �������I�GI�GH�$H�H�Z���f.�     H�$H�QH9��  H�$H��������H�yH�AH9��  H�$H�PH�Q� ��L��	��������'  @ I�GI�oH)�H������)�9���   I�GH�$H�H�����f�     ��L���6����$�d  A��A�ƍED��A��L���������$�   D��A�������uF�������u��A������H��E��D��ATF�,D��D��E��H��$�  ����D��$�   D��$�d  ^_9��R  ��D��$�d  D�M)�E����o����J���f.�     I�GI�oH)�H������)�9�������D�M)���   f�D��$�   E��L�����;����$�d  D��A���)����uA������u��F�����H��E��D��F�, D��D��AUH��$�  �����D��$�   D��$�d  AXAY9���  ��D�M)��p�����L�������$�   A��A�ÍED��A���V��� I�oI+oH��A�����  E1�D  D��L��A�]�i���A�u�$�   �Y�����$�   �$�d  H��$�  ��$�d  �u���A�EA��D9�r�9���
  �L���������s�$�   A�������s�$�d  A��������sF�4������sF�������s��F�,0�����H��E��D��B�, D��D��UH��$�  ����D��$�   ��$�d  AZA[D9��m����+
  �     I�GI+GH����v��$�    ��  H�D$HƄ$�   ��8   �_  L��������$�   ��$�   �Ƌ�$�d  H��$�  ����I�GH�T$H�$D�b�RH�yH�I�5���f�     I�GI+GH�����  H�\$HƄ$�   ��8   ��  L���I����$�d  �=������  �$�   �Ɖ�$�   ���t����[���f.�     I�GI�OH)�H����v��$�    �����H�D$H��D��L��j L��$�d  H���   L��$�   H��$�  �	���]A\H�D$H��8   �,  H��$�  H�$�  ����  H�\$1��  L�4$H��$p  f��HǄ$(      �H���   L��H��$   �$  ��$�  �D$\�$  ��$�  H��$ K  H��$x  H��$(c  H��$�  H�D$xH��$p  H��$   ����H��$   E1�E1�H��$�  H��$p  H��$p  ����I�GD�c�SI�~I�N�Z���fD  H�D$�x �9���H�D$H�xh �����H�X`H���   ���   ���   H���  H���P��t-H�D$H��H���   ���   ���   H���  �P ����  L���������9D$p��  L�t$A�   A�F����������@ H�D$�x �����H�\$�{a �����L���z������u  H�T$���   I�G����fD  �|$W �  E���  ��$�d  ��$�   H��$�  �����H�D$x�\$@f���$�   HǄ$�      HǄ$�      �$�   HǄ$�       H��$�   Ƅ$�   ��ttH��$@  Hc�D�S�H��$h  H�A�L��$X  H��L��$8  H��L)�H��H��     I��I9�wI��M��tE�E��uA� �   �H��H)�H9�u�L�$H�$H�T$�D$@    I�G�D$WH�KH�{H�KD�b�R�9���D  I�OI�GH)�H�������Å���   E1��8@ �$�   ��$�d  ��$�   ��H��$�  A���������A9���   D��L��������u��$�d  ��$�   ��$�d  �@ I�OI�GH)�H���Å�th1�f�     ��L���F����u�$�   ���4�����$�   �$�d  H��$�  ��$�d  �P���9�r�H�D$I�OD�`�PH�$H�xH�$I�OH�H�b���f�I�GI+GH����v��$�    �-  H�D$HƄ$�   ��8   ��  L���/����$�d  ��$�   ��$�d  �[��� E���  ��$�    �����1�H�\$H��L��D��PL��$�d  H���   L��$�   H��$�  �NfD  E����  ��$�    �I���1�H�\$H��L��D��PL��$�d  H���   L��$�   H��$�  �����AYAZH�D$H��8   ��
  H�$I�GD�c�SH�yH�I�����I�GM�WI)�I����D��A�ƃ��A)ʉL$XA9���   �%����    D��L��E1��j������$�   D��$�d  A���Q���B�D�ƉL$t�A�����F�(�6����L$tB� ��A����  H��D��A��D��SH��$�  �������$�   E�≜$�d  ZYD9d$X��  D�L$XA�jE�BA�ZE�bE)�E���P���D��L��D��$�   A�   �������$�d  A������B�D�ƉL$t������F�(�����L$tD�Í,A���M���D���g����L$tB� E�b�4���fD  HcD$@�������H��H;�$X  r$H��$8  1�H��tD�*E��u��   �    H��$@  L��H�$h  H�$�#���H�T$�z t(H�T$HH���  H��t����/��H�¸����H��t��f�����c  L�$H�\$HAAC�H  ;�@  �����H��P  ��H��I�K�{\ ��  H���  H����  �<�H�I�{�  D  E���w���H�D$HH�x(�����Ƅ$�   ����@ I�GI+GH��A�Ń��!  �   �\$X�D  ��L���u�������u��$�   A��������u��$�d  A��������u�F�4������u�F������u�F�$0����H��D��E��B� D��D��SH��$�  �i����ED��$�   ��$�d  A^ZD9��k����\$X���  I�GI�GH�D$D�`�PH�$H�xH�H�����    H�$H�AH9��7  H�<$�������A���Q����#  �$�0I D  I�GH�T$H�$D�b�RH�yI�GH�$H�H�N���fD  �   H��$0  覙�������������f�     �À����  H�4$H�V�����  ��	�����H9���  H�<$�8����tlL���l��������    ���D$@H�H;�$X  r-H��$8  1�H��t�)��uH�T$��   D�b�RD  H��$@  H�$h  H�xH�HH�$�n���fD  H�PH�Q�A�������D  ��$�    �����1�L������H��$�d  �$�   ������f�H�BH�A�2H9������H�<$�S��������fD  H�D$HH�@@�@�P����    H�D$HH�@@� �����H�$H�T$HC�L  ;�D  �����H��X  ����H��H�KH�KH�<�H�{H�D$�D$@D�`�P�w����    ��u���L�����������D  L���`���H�\$HH�H�SHH�H�B    �E���H�K@��Hc�H��{[ Ƅ$�   ��  H�L$�|$W �Q��  �$�   H�L$I�GD�aH�$H�yH�I����@ H�L$I�GD�a�QH�$H�yI�GH�$H�H����fD  D��� ����L$tE�b�,�����L��L��E1�A�@   �,����r����    ����2  �������H9���  H�$H�BH�C�������L��)�������[�����H�<�H�$H�xH�$H�H����1�L������H��$�d  �$�   �����1�L���j���H��$�d  �$�   ������E1�A�@I H��$�  H��$�d  L��H��$�   �K��������A�   A�I ��E1�A� I ��E1�A�0I H��$�  L��H��$�d  H��$�   ���������H�BH�F��g���D�aH�$I�GH�yH�I�����H9��O  H�$H�BH�A�
H�$H�SH�CH9��  H�zH�{�2H9���  H�$H�WH�SD�H9���  H�$H�BH�C�����H�\$	�A��D	�	ƀ{ �  �� }  �   L��=�  �D$0CD$0����H�$D�c�SH�xH�H�o���1�����1�����H�D$�x �����A��%�����H�T$D�bE���]  �\$8����  A����  H�$I�G�D$8    �RH�yH�I�����    H�$H��$�   H������H�T$I�GH�{H�KD�b�R����L�����<����u�$�   �-�����$�   �$�d  H��$�  ��$�d  �I�������H�D$M�_A�   M+_D���   I��D��E)�B�,A�����   �\$XL�t$�    I���   D��L��H�X����A���   A��vKD��E��A)�@ L��H��D�V����HcS�H�D��H��H�H�� �  H��A�C�A;��   r�E��I�WI�GH)�H��A9�w>D��H��D� �@    A��A9��`����\$XD��L��)�����H�D$�@a�����L��������H�<$轿���"���L�t$E1��V���H�\$H�    D���  E��I��  H�$��Hc�H�H�KH�<�H�{����H�<$�i����H���H�$H���X���H�SA��H�C����H�$H���<���H�{��H�C�����H�<$�$���������L���u���I�WI+WH�������������  1�9�s��)�L��������L���Z�������I�GI+GH��L�t$�����u��$�    �  H�D$HE1�Ƅ$�   ��8   �<�����$�c   ��  E1�fA�~ ����I�GI+GH�����
�����$�    A�   �����L������A���������������$�d  ����H�|$HH��$p  D�Ɖ�$�   蜡��A�Ņ������L��$   A�   L��AT��$�d  PD��$�   H�L$xH�T$pH��$�  H��$�  ����L�l$XH��$�  H��H+�$�  I�}A���  ��L��H��$�  ����Y^A�Ņ��(���ATE1�A�   L��j H�L$xH�T$pH��$�  ����H�D$XH��$�  H��H+�$�  H�x���  XZ�����D  ��w	���$� I H�$H�T$I�GH�y�RH�I�i�������$�   H�D$�PH�$H�xH�H������!w����$�I H��$�  �����7���A��L�t$�X���1�L���ӽ����$�   �H��$�d  �(�����E���h���L��1�訽���   A��蛽���   A��莽���   A��聽��I�OI�WH)�H������   A�D���A    D)؉A�   L���I���I�OI�WH)�H������   E)��A$    A)�D�I H�D$HA��H�@@ty�@H��$p  H�\$�SH���   �T$XL��ASPL��$�d  �|$hL��$�   ������|$W �}���L���O�����$�d  �C�����$�   H�D$Hǀ�      �}���� H��$�  ��w����b����m����"���E���L�����$�   ���3����|$8 ������l$8HcD$8����   �-���E������L���^���A���V���Lc�I�GA���q  D���$�(I E���r���H�D$HH��   ���  ����1��҉���1�����1��r���  L������H�D$�D$8    Ǆ$�      D�`�PH�$H�xH�H����A�����������A������A��������� ���E9�LƉ��H�\$HH���   �����A��������t����������9��  �����H�T$HH�H���  H�4��J���H�\$HH���   �v���A���l����'���Hc����\���9��  �P����k���H�T$HH�H���  H��H�D$�D$8    Ǆ$�       D�`�PH�$H�xH�H����A�����������Hc������������Hc��A��������A�����������Hc�����H�H��H�H�� �  H���k���A�������軹����费��)����L���A�������蜹����蕹����/���H�\$HA��L���  �X���M���O����
������B���A��;��  �0���H�L$HH�I��  H��H���  H�<���S  �����H�T$HH���  H�������1�A����E�L�A��A9������M�WI)�I��E)�G�$
D��D��L��D�u��C���A�   A���4H��  D��L��H�,��"���H�Hc�A��H��H�H�� �  H��A�C�4D9w�I�WI�GH)�H��A9���  D��H��D�(�@    A����E9��q���D��L��D)��%���H�D$�D$8    D��$�   D�`�PH�$H�xH�H����I�G����E��������|$W �����H�T$H���   ��������  �C���  �C����t���H�D$H�   H�x�*�������������~�D��P���$�   ��Hc�H�����   ��$�d  ����   ��t	������S��$�   P��$�   ��$�   D��$�   D��$�   ��$�   H��$�  ����H�D$ D�`�PH�D$]A]H�xH�H�D$8    Ǆ$�       �����E��������|$W �����H�\$H�   H�{�J������Z���Hǃ�     �i���A��������|$W �V���H��$�   1��
   HǄ$�      HǄ$�      H���H�D$xƄ$�   H��$�   ����A���=����|$W tH�D$H���   �$������  ������$�   L��������$�d  �ܵ��H�D$�D$8    Ǆ$�      D�`�PH�$H�xH�H�����H�D$HH��   ���  ����1��҉���1�����1��r���  ����L��諵��A��裵��A��蛵����蔵��E9�LƉ������L�������������H�����  �����L��� ���Hc��X������j�������  �^���E���`���L���2���H�\$HH�H�SHH�B����H�SHH�H��������	���H�S@�
�Hc�H�
�JƄ$�   �Hc�H�J�{[ �e���H�L$�|$W �Q�k����$�   �$�d  ����E�������H�D$HL��L�t$L�@�8���A���0�����艴���$聴��Hc��y�����$�    �D$�L���H�D$H�x[ �=���H��`   ��  H�D$HH�@@HI���   H�xh �S  ���	���E��� ���H�D$H�xZ �z  H�H�   H��(  H�L$0H�H��H�T$(臈��H�T$(H�L$0��A�������H���   HcD$H�L$8H�T$0�.H)�f�FH��H�F    D�f0f�F4 H�t$(���H�t$(Hc<$H���F8H�t$���H�T$0H�t$H��H�L$8�F<H�BXǁ�      H���   ǁ�   pmocǂ�      ����E������E������A���   �   IN��D$8L����   I��;t$8�$  L������A� ����L���>����w���L�l$H��L��躟��D��L���譟��A������I���   H�xh �����H�D$HH�@@H�f���L�l$HI�}�d��I�}��L�l$HH��$p  �����A�Ņ��L���H��$�   A�   L��E1�Uj H�T$pH�L$xH��$�  �3���L�l$XH��$�  H��$�  I�}H��$  H)�H���   ��$  ^AXH�@hH��tH�xH� H��$   �PI�}H�T$HD��H�B@H�RHH�H�L$(H�HH�L$@H�
H�RH�     H�@    H�T$8H��$p  H�L$0�!���A�Ņ��q���U�D$A��A�   L��PH�L$xH�T$pD+L$ H��$�  �X���H�D$XH��$�  H�PH��$�  H��$  H)�H���   ��$  ZH�@hYH��tH�xH� H��$   �PH�T$HH�L$(E1�H�B@H�H�L$@H�HH�BHH�T$0H�H�T$8H�P����Ǆ$�       H�D$D�`�PH�$H�xH�H����L��衰��Hc�虰��H�H��H�H�� �  H�������L���x������q���9�@��@�������x���L���U����k���L���H���1��������Hc�H���	~
��Hc��H��H��H���^
��H�DH��H9�u���h���L������=   �th�؉��P���L������������)����8���L��E��t�D$0uB�Ư��L��A��軯��Ic�Hc���	��������L��衯����蚯������������������$���A�������D$0 �L���m���=   �tә1�)Љ�����L���R�������������L���>������7���A������D������L������1���@��蒮���(���L�������������	�@��@���o�������L���������ۮ��������@��@��!��E���������r�����L���P���A���H����ƃ������H�$M�_H�xH�HI�GL)�H��9���   D��E��xw���H�D$D�`����   ���A�   E1�E1�A���&)�Lc�A��O��A�(A�XE�E�PA��A��D9�tWA9�uA�ELc�A��O��E�E�P�9�~���y����ؙ�����I�GH��t�8 u� �   H�D$D�`�P����H�D$��D  AWI��AVI��AUATUH��SH��   D�g\�D$<    E��tH��    �F  M��(  I�] H���	  I�L���   f��L���   H���   H���   H��$�   H��$�   L�D�BpI�WHǄ$�       D�H<)D$`��0   H��$�   H�D$p    ��1  ��  �D$`   �D$l   E����	  �C D�c�C    ��tE��ty	E��u�K�P@���   ��  �PD��  �PH��  �PL��  �PP��  �PT��  �PX�@\���   ��  ��   ��tR�l$`����  D�d$lE����  ���  ��
  ���  �Hc��l��A9��{
  9��s
  L���   I�H�D$X    D���   E1��D$@    D���   H�D$P    M��   �D$D    H�D$H    �C    L;��   tL���   A�   �{ uI��  D���  E���;	  H���   �@��;C\t	�C\A�   �CH�L$h1�H3K����   H�T$`H3SH	щ���  @�ƃ�����  foD$`H�t$pH�       H�C$    H�CD   CC,H�s<H�{L9�t	����  D���   E���0  �  ��A��H�H�$=�  I��A��I��   �{\   �   Mk\H���  ����$  ����
  H��  E��D�\$H��,  H�D$��  D��  ��$  ǃ,      E��tE��uH��E1���D���t$�f���XZI��   H�4$H���  ������~��9�$  �J
  �  n �P����(  ��D��  E��ǃ0      ��E������u%E��u H��H��0  E����t$D������AZA[D��,  �   E��uD��0  E����H��@  ��  ��H���   H����  �Hǃ8      )�ƃ4   ���  1�Hǃ�      ���H��C8��8  H��   H���  �{��H��   ��D  ���  ����H  ���  ����L  ���  D��H  D��I  D��J  D��K  ��  E1�1�M��uH��   @ ��0  ƀ�   ���  򉐜  ���  ���  ����<  H��I9���   ��<  ���X  ���P  ��H��H��H����A�҉��  ���  A)�x�E9�EL�H���x������  ƀ�  ���  � L��8  A�s_A�� AI����t$`H��@  �V_�� I����T$lE���  �C D�c�C   ����f�M��tsI��H���  I��I��N���  ���<  �H��H����H���F���  �����  )�x#A9�Ƃ�  DL����  �����  ��<  H��I9�u�Hc�8  �   �����<  H���  E1�H�<$��tz�    �~ ���  I��vS��0  A����A�   D�	B���  ����D�A��A)�)�AH�D9�E��DN�A9�~	���tA��I��M9�w�I��H��L;$u�Hc�D  E����  Hc�8  9��  ��   t
ǃP      D��<  M��tsLc�8  ��P  H���  1��!�    )�H��H�� �  f1��B�L9�t:HcI��H��H��?H��8 �  H���z uƍ� �  H��H��f1��B�L9�uƋ{����  ƃ4   ��  L�d$@L���   H���   ǃ�       H�x�5	��ATL��E1�j E1�H��H��$�   H�L$`�����sZY����  @��t���   ����  H���   H�}(賗��H�}��
���C�T$@���[  H���   �y\ u�� �  H��0  ��H��H�H�Ĩ   []A\A]A^A_�D  ����M��tBE1� B��͈  A����A��A)�A)�EH�9�A��DN�E9�~
�>E��tXD��I��M9�w�I��������  ��A��A)�)�AH�9�N�9�������>I��H��L;$�l���������    1��@ 9������E���k�������f.�     I�I�E@�E H�T$<��  H��H�$��a��D�L$<I�E �@   E�������I��(  H�$H�H�E��uI��  H��h  H���  f��H�CHǃ�   0�E ��   ��   ��   H���   H���   Hǃ�   @�E Hǃ�   ��E �J���@ E1�H�$   A�   A��  �����@ A��Hc�H�L$(Mc�H��H�T$ L��L�D$����Hct$L�D$H�T$ H�L$(H9�I����  ǃ,      ��$  A���  �����H����E1�E���t$D���?���Y^������     ��x  �C �C    �S�'���fD  ��x  �C �S�����D  ƃ4  1������f.�     Mc�   L�������H9��G  ��D  Hc�8  9������ƃ@  Hcտ��  ��������  )Ё��  ��  O�P  ����@ H���  D�$E1�1�H���  H�L$HH�t$D�P@�C���  I��   A��  H�L$H�T$D�UD�$��t I��  �T$DL��A�   H�L$H�UD�$I��(  �Ca I�H�ChA��  ���   �D$D���   H�D$HH���   ����@ ��   �W���fD  H��L��H�L$�������$  H�L$ǃ,      ��A���$������� L��   �����ŉ�D  ����fD  �   �����fD  M��tcE1�1�I���������P  ��=  ���w�����X  ��=  ���c�����`  ��=  p�O�����h  ��=  p�;���@ Hc�8  ǃ�  ����ǃx  1   H��H�򉳐  H����p  H)�ƃA  ǃX  2   H��H)�H��H��?H�� �  H�� �  f1�- �  ���  ��0  ��  pHc�h  H��H�H�� �  H�� �  f1� �  ��l  ����fD  �   ����fD  H�4$�  K D�D$D�\$�(���D�D$D�\$��$  �5��� �  K ������(  ����f�     �$   �_���fD  ���ωЁ����%���9�t�   w���    9��9Ѻ   G��f�     H�W �GH��H������H�rpH��H�<9�t^E1��,fD  H9�t;9�v.H�WH9�r.H��H)�H��H�<9�t-%���9�u�H9�tI��H�O�H9�s�1�M��u	��     L�ǋG�1��fD  S�_�����   ��L�_ D�@���M��A�
A9�txA��1�1��*�    v^�zD9�s0D��)���:M��H��A�
D9�tE�����A9�u�A��A�BD9�rЅ�u.E1�9�s'I��[D��BA�����D��D  A��� A�BD�[�1�E1�����   ��  w��H��?��I H�J Ð���  w��H��?��I H�J �fD  1��ff.�     f���I �f��fD  SD��4   E1�B����	H����I f����D���I L���I D����A9�tP~E�@  f�     A�	���H����I f����D���I L���I D����A9�tc��A9�|�1�[�H��H9�s/D��E�B�I�BE��A��E�ل�yID9�u�I��H��H9�u�1�E��x�A�z y�A�B[f�����@ ��D�JA9�����1��D  I��E��IH�H�PE���t���D�@fA��E��M���I E���I E��A��D9��z���E�C�N�L@�'�f����D���I L���I D����9��H���H��I9�u�1��������\���f��<utQ����   �WH����     ��.uH9�r�VH����u�H9�sv�0�����    �#���   ��D  �W��nt_L�GA�Ҿ   1�E��A�IЃ�	vA�I���w/A�IɃ�w&��I��E�ȃ�u�E��t�A��.�d����1�Ã��V����᐀iu�H�OL�O1�D�A�pЃ�	vA�p����w���A�pɃ��j�����H���L9�u��O��t��.�K����2����@ AWf��AVAUM��ATA��USH��H��   �F    H�F     L�L$,H�t$�   H�$�J
1�L�D$E1�H�|$)D$0)D$@H�D$P    �fj��H��H�C �D$,���  E����  1��     ��L��H�$��I��H��t[E1�1��fD  Jc<� I H��@I L����� ����   I��I��
u�L�������������   H�D$H��tL��L���Ѓ�A9�u�H�D$�L$0H�x 1��f�     �L0��u���I �L`H���E��M�H��H��(u�H)�H������   D������9���   ��/F �   H���y>  �D$,H�L$�iH�Ę   []A\A]A^A_� J��    H�D$0HЋ���'����    L���\`�������������1Ҿ�  ��    �4��I 9�tH��H��
u�E H���]������@ �E H���]��D�0   �����1�H��������    H��H�|$�s���H�D$��   H�@     �D$,��D����� I��H�|$D��L�L$,H�پ   �Sh���D$,    H��H�D$H�x �����f.�     SH��H��U�  H�C    H�C    H�    [�f.�     H��uH9wrEATUH��SH��L�gH9wu!L��H��H��[�   ]A\��  f.�     1�L���i�  ��@ �   �f.�     H���C  �     H���B  �     H��H���D  D  H����   USH��H��H��H�s �PJ H�C    H�    H�C    H�C(    H�C0    ��  H�Ÿ   H��tB�   1�H����  H���'�  H�CH��t)1�1�H����  H�k1�H�C(�6F H�C0�6F H��[]�H�����  H���Q   []�@ �(   �f�H���    �B  H��tH�     H�@@7F H�@`7F H�@P7F H���f�     �sA  f.�     �H��tH�G     f��G��    ��ff.�      AWAVAUATUSH���D$    H����  H���h  H���_  H9��  �^�BA��A��A��A��A��A��H�~ ��   H�Չ�D�.I����L�EH�?1�)�Hc�L��M���6  ����1ȉE )�Hc�H��I9���   �Ao$E �AoL$MI�D$ L�EH�E E9��  �E I��M�d$I�ݍx�H��H��I���u	�"@ ��L��L��H��I��/0  I��M��u�D$H��[]A\A]A^A_��    �o�o^ZH�F H�B E9�t�ۉZ1�H��[]A\A]A^A_�D  L�L$L��   ��c��H�E�D$��u�L�E�����H���   []A\A]A^A_�@ H���!   []A\A]A^A_�@ H�T$L���3c��H�E�D  I�t$L��L���S/  �D$�c���ff.�     @ AVAUATUSH���D$    H����  H���z  H���q  H���VH��D�mL�EH�Ѓ���vL�D$   �SL�c��y�����Hc�I)�E��y�M ��D��Mc�M)�<�  �$�XJ �    D��D��H�?�E���61�)C�U �u �ED�KA��E�ͅ�~D�ș������   ��D�Ҿ   A��L�L$�Qb��I��H�E�D$����   D�ME���1  D�m�C�8���@ �;�   f�U��tq��C������  �r�1�L�N��     H��A�������A�@A�T@H�PH9�uދCK�K�H�t����HcCI�HcEI���u�@ �D$H��[]A\A]A^��    ��)�E�,E�������     D��   f�EE��t��    �C1�D�H���u�qf�     H��E�\�1�D��E��tEA��A�D�A�T�H��H��H��Hi�|  Hi��  Hi�m6  H�H�1�H��A��)ǉ�A�0H�FI9�u��SHc�I�HcEI�A���i�������@ D��   f�ME������ �C�����2  D�R�L��L��I��O���H��H���Ɖ�����@�r����������J����B�@�r�L9�uʋCM���s  HcCI�HcEI�A��u�����f�D�+�   D�sf�uE���g����    L��L��L����+  I��HcCI�HcEI�A��u��6���fD  D��   f�}E������ �S�����:  D�P�L��L��I��O��     �H��H���ǉ�����@�z������J���@�z�������@�z�������@�z�������@�z������������B�@�z�L9�u��SK�Ѓ�u/HcCI�HcEI�A���O����b���f�A��������     ��A�	H�t@ ��H������P�H9�u�� ��A�I�L��I������A�A�I9�u��g���f�H���   []A\A]A^�fD  H���!   []A\A]A^�fD  L��M���A���D  M��M������D  L��L������D  1�H��t���   stibt�@ H��(  �Bu�SH���   H��f��H��0H�?H��)$)D$H�D$     ������u0H�T$ fo$foT$H���   H��(  ��   ��   �JH��0[ÐH��t;H��t.SH��H�?H�v�f���f��H�C     1�C[��    �   �f��!   �f.�     H����  H����  H�~ ��  L�B �   I��I�����nL�A I��I�����]�� AW�� 1�AV��AUATUS������H��x	ʉ\$�L$��   ����  ���}  �VH��H�����#  ���$ŘJ �fD  A��D�A��H��A����G  D�t$H�t$(�L$�   HcSD�T$0L�D5 ��tEf.�     ����Hc�E��t&H��M��H)�I)��    �2
H��I9�u�HcS��D9�u�HՃ$��<$9���  T$�T$�D$C�D$�1�H��x[]A\A]A^A_�f���   H�T$@H�D$`    )D$@)D$P������u�H��H������H�D$`foT$PfoL$@H�C S�S�D$�sD�k�D$��H�E ��H�D$A�̋A1�A��A)̀���  �$��J �   ø!   ø   �K����|$F�t/A��E��A�   D�L$E���c  E9��Z  �|$B��    H�kB�/A��9��P  A��A� �  N�t% ��A��A��I���-  H�$D�ŉ��M�M���  L����tE /I�L9�s�L��1�H)��a&  �ϋ|$F�t/A��E��A�   �O����|$�   D�n��NǉD$�D$�D$H�E H�D$��vA������A��A1�A)ԋ|$F�t/A��E��A�   ������D$�@�D$�D$�sD�k�D$��H�E ��H�D$A�ԋA1�A��A)ԋ|$A�   F�</�����D$�@�D$�1�������   ������|$L�L$@E1�1ҍD��H�|$H���Y��H�ŋD$@�������D��E��{D�3A��L�kK�D5 E��H�$�D$��E)���A��H�D$ ����  L;,$�;  ��Mc�H�D$(D��I��H�D$0L�H�D$8H�T$(L��L��M��!%  H�T$0K�<&1���$  Lt$8L;,$r�H�T$ 1�L���$  H�sH�|$E��軂���sH�k���=  D�{�E���  �T$A��Hc�HՅ������A�~��t$�$    A�   ��Hcǉ|$ ��H�zH�D$�D$�t$0H�|$(��H�|$�t$ H�A����������D�t$D�t$ �   D�'E��uZ����D  D��)������Hc��D�[D�| ��E��D�A9��Z���D���K�҃�9��J�����9��?����{u�D�����
�E��t�D�O�D��)�A��D	ʈ��H�$H�k��sA�������A�ލP�A��H������A�ދD�s����H��H��1��L$(�5#  �|$(H�D$ Mc�H�|$ K�<4H�H�|$(L;,$�]���H�\$0H��H�T$ L��H��M��9#  J�<#L��1���"  H\$(L;,$r�H�\$0����I������ H��H��E1�E1�H�t$1ɿ   H�D$    ��  H�D$H���f.�     D  H��H��E1�E1�H�T$1ɿ   �  �D$H���f�     Hc�E1�E1�1�1ҿ   �  f�     H��H��H��Hc�L�D$H��E1ɿ   �k  �D$H���D  H��H��H��Hc�L�D$H��E1ɿ   �;  �D$H���D  H��H��Hc�Hc�L�D$H��E1ɿ   �  H�D$H���@ H��H��E1�Hc�L�D$�!   ��  �D$H���f.�     �L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A���	  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�H��H	�t�l   �AUI��ATA��UL)�H��SI��H��H��H���  M��uH��[]A\A]�f.�     J�<#J�t% A��s1A��uvE��t���A��t�E��B�D.�fB�D/��f.�     H�H�OH���H�D��H�T�H�T�H)�H)�D������{������1���L�L�9�r��`����E��B�D.�B�D/��J���ff.�     @ SH���(   �f0  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     US�D$L�T$ ��y�1���y�1�E����E��M�ZA��A��A	�E	�A��   ���~OA;r}I��l��t�D  A�BA��D�ȅ�~9�~���
���A9B~A�E��9�u�9�t	��A9Z�[]�ff.�     D��SE������AQ��A��P�D���XZ[�H��I��H��A��H�� ��H�� ������� AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   �CA9���   D��D��D�\$�NfD  ��L�[�D��    G�L��L�KD��x��E�9E� H�{D�D9�t=�C����9�~0��D�BD�L= �zI�H�A��u��?u�A�8u�D9�u�D  D�\$E)�9t$t��9s�F���H��[]A\A]A^A_��    AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�w���XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_ÐH��H��A��H��APH�� A��H�� ����m���H����     AVA��H�� AUATUS�F��~u�G)Ѕ�~l��I��I��1��D  A�E)�9�~QA�D$A�M�<+B�40��D)�9�N����Ń���D�Hcҍ4�    ��Hc�Hc�It$I}�����A9l$�[]A\A]A^�ff.�     ��NA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      H��H��E1�E1�H�T$1ɿ   �_  H�D$H����     L�D$(H�L$ H��E1�H�T$�   �.  �H���   HD��)  ff.�     @ ��(  ff.�     ��'  ff.�     �����ff.�     ��'  ff.�     �'  f.�     �UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo% SF f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo% SF f��fs�f��f H����H��]Ð�����������                AW�B��A��AVAUE��ATU��SH��H�� �K �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�����_AXA��@�w���A��AV�   ��RD�L$A��   D�D$����Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�s���XZA���%���A��AVA��   RD�L$�   ��D�D$�@���A[XA�������A��AVA��   RD�L$�   ��D�D$����AYAZA�������A��AVA��   RD�L$�   ��D�D$�����_AXA�������A��AV�   ��RD�L$A��   D�D$����A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃��i���XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_�UH��SH�}�H�u�H�U�H�M�L�E�L�M�H�E�L�E�H�M�H�U�H�u�H�}�L���i�[]�UH��H���}��E�H�A�    A�    �    �    H�ƿ   �������UH��H��H�}�H�u�H�E�%�  H��tH��� �   H�5�� H�=�� �
  H�E�H�U�H���  H��H��A�    A�    �    H�¿   ����H�E�H� H��u�������    ��UH��H�}�H�u�    ]�UH��H��H�}�H�E�A�    A�    �    �    H�ƿ    �������UH��H�=� ����UH��H��H�E�A�    A�    �    �    H�ƿ   �w���H�E��E��E���UH��H��0�}�H�u�H�U�H�U�H�E�A�    A�    �    H�ƿ   �2���H�E�H��H�E�H�H�E�Hi�@B H��H�E�H��    ��UH��H���   H��X���H��P�����L���H��@���H��`���H��Q�K H��H���  H��`���H�5%� H���  H��H��@���H��H���  H�5� H���  H��H��P���H��H���  H�5� H���p  H��L�����H���  H�5Ҹ H���N  H�5Ÿ H���?  H��H��X���H��H���*  H�5�� H���  H���e  H��`���H����  ���UH��    ]�UH��]�UH��H�}�H�u�H�E�]ÐUH��H��H�}�H�E��     H�E��@    H�E�H��H����   H�E��@ H�E��@ H�E��@ H�E��@ H�E��@ ���UH��H��H�}�H�u�H�E��H�E��H�E��PH�E��PH�E�H��H�U�H��H��H���   H�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��PH�E��P��ÐUH��H��H�}�H�E�H��H���(   ��ÐUH��H��H�}�H�E�H���2  H�E��@ ��ÐUH��H��H�}�H�E�H���  ��ÐUH��H��H�}�H�u�H�E�H����   H�E��PH�E��PH�E��@��tH�E�H�ƿ   �U���H��H�E�� ����UH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H��H�}��u�H�U�H�E�H��H����   H�E���UH��H��H�}�H�E�H� H�U�H��H��H����   H�E���UH��H�}��]ÐUH��H�}��]ÐUH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H���>���H�E�H� H�U�H�M�H��H���x   H�E�H���������UH��H��0H�}�H�u�H�E�H�������H�E؋ H�U�H�M�H�Ή��_   H�E�H����������UH��H��H�}�H�u�H�E�H�U�H��H����  ���UH��H�� H�}�H�u�H�U�H�U�H�E�H��H���M   ���UH��H��@�}�H�u�H�U�H�U�H�E�H��H������H�U�H�M��E�H�Ή���   H�E�H���+������UH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=e� �Ȣ��H�E�H���   H��u)H�E�H� H�U�H��H��H�������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=³ �͡���u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�7� H�E��E�    �E���~H��    H��uH�=�� ������M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=|� 菠���E��P�U�H��D�-H�U�H�E�H��H���   � 9E�����tE�E�    H�U�H�E�H��H���   � �U�)�9E�����t�U�H�E���H���   �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���b   �E��ڋE����E�}� x!�E�H��D���H�E���H���2   �m��ِ��UH��H�}�H�u�H�E��H�E�� 9�}H�E��H�E�]ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=�� �L���H�E�H���   H��u)H�E�H� H�U�H��H��H���u���H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ��ÐUH��H��H�}�H�u�H�E�H���������ÐUH��H��H�}�H�u�H�E�H�����������UH��H���   H��X���H��P�����L���H��@���H��`���H��Q�K H��H��� ���H��`���H�5� H���@���H��H��@���H��H���+���H�5�� H������H��H��P���H��H������H�5ޱ H�������H��L�����H������H�5�� H�������H�5�� H�������H��H��X���H��H������H�5�� H������H�������H��`���H���������UH��H���   H��X���H��P�����L���H��@���H��`���H��P�K H��H����   H��`���H�5� H����   H��H��@���H��H����   H�5� H����   H��H��P���H��H���   H�5Ұ H���   H��L�����H���   H�5�� H���   H�5�� H���u   H��H��X���H��H���`   H�5�� H���Q   H���   H��`���H���.   ��ÐUH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H�}��]ÐUH��H��H�}�H�u�H�U�H�E�H��H���   H�E��ÐUH��H��H�}��u�H�U�H�E�H��H���   H�E���UH��H��H�}�H�E�H� H�U�H��H��H����   H�E���UH��H�}�H�u�H�E�H�U�H�H�E�Hǀ�       H�E�ƀ�    �]�UH��H��0H�}�H�u�H�E�H������H�E�H� H�U�H�M�H��H���x   H�E�H���f������UH��H��0H�}�H�u�H�E�H���W���H�E؋ H�U�H�M�H�Ή��_   H�E�H���#������UH��H��H�}�H�u�H�E�H�U�H��H���������UH��H�� H�}�H�u�H�U�H�U�H�E�H��H���M   ���UH��H��@�}�H�u�H�U�H�U�H�E�H��H������H�U�H�M��E�H�Ή���   H�E�H���������UH��H��H�}�H�u�H�E�� ����   H�E�H���   H��vH��    H��uH�=#� �&���H�E�H���   H��u)H�E�H� H�U�H��H��H�������H�E�Hǀ�       H�E�H�PH�U��H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D �B������UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=�� �+����u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�=� H�E��E�    �E���~H��    H��uH�=T� �W����M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=:� �헹��E��P�U�H��D�-H�U�H�E�H��H������� 9E�����tE�E�    H�U�H�E�H��H�������� �U�)�9E�����t�U�H�E���H���q   �E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���:   �E��ڋE����E�}� x!�E�H��D���H�E���H���
   �m��ِ�ÐUH��H��H�}����E�H�E�H���   H��vH��    H��uH�=o� �Җ��H�E�H���   H��u)H�E�H� H�U�H��H��H������H�E�Hǀ�       �M�H�E�H���   H�pH�U�H���   H�U��LH�E�H���   H�U��D ���UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�sH�U�H�E�HЋU�H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�H;E�s"H�U�H�E�H�H�M�H�U�H�� �H�E���H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H;E�s4H�E�    H�E�H;E�sgH�U�H�E�H�H�M�H�U�H�� �H�E���H�E�    H�E�H;E�s3H�E�H+E�H�P�H�E�H�H�E�H+E�H�P�H�E�H���H�E���H�E�]�UH��H�}�H�E�    H�E�    H�U�H�E�H�� ��tH�E�H�E���H�E�]�H�H�oL�gL�oL�w L�(H�D$H�G0H�$H�G8H��    �H�H�oL�gL�oL�w L�(H��H�g0�g8UH��H��H�}�H�E��    H���|   fH~�H�E��E���UH��H��H�}�H�E��
   �    H����   ��UH��H��H�}�H�E��
   �    H���   ��UH��H��H�}�H�E��
   �    H����  ��UH��H�� H�}�H�u�H�U�H�E�H��H����  fH~�H�E��E���UH��H��H�}�H�u�H�U�H�E�H��H���  ��UH��H�� H�}�H�u�H�U�H�E�H��H���8  �}�H�E��U�H�E��U��m���UH��H��0H�}�H�u��U�H�E�� ��t"H�E�� �����Wa  ������uH�E��ԐH�E�� <+uH�Q� �:   H�5]� H�=� �^����E� H�E�� <-u	�E�H�E��}�
t@�}� tH�� �B   H�5� H�=K� �����U�H�M�H�E�H��H���   �   H�E�    H�E�� ��tGH�E�� </~<H�E�� <91H�U�H��H��H�H�H��H�E�� ����0H�H�H�E�H�E��H�}� tH�E�H�U�H��}� t	H�E�H���H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H��`H�}�H�u��U�H�E�����H�E�H�E��E�    H�E�H�PH�U�� ���E�E����_  ������t�փ}�-u�E�   H�E�H�PH�U�� ���E���}�+uH�E�H�PH�U�� ���E�}� t�}�u9�}�0u3H�E�� <xtH�E�� <XuH�E�H��� ���E�H�E��E�   �}� u�}�0u�   ��
   �E��E�Hc�H�������    H��H�E؋E�Hc�H�������    H��H�ЉE�H�E�    �E�    �E����\  ������t�m�0�4�E���^\  ��������   �E���_  ��t�7   ��W   )E�E�;E�}r�}� xH�E�H9E�rH�E�H9E�u�E�;E�~	�E������*�E�   �E�Hc�H�E�H��H�EȋE�Hc�H�E�H�H�E�H�E�H�PH�U�� ���E��<�������}� y
H�E�������}� tH�E�H��H�E�H�}� t�}� t
H�E�H���H�E�H�U�H�H�E���UH��H�� H�}�H�u��U�U�H�M�H�E�H��H��������UH��H��`�K H����  %���]�UH��H��H�}�H��� ��   H�5�� H�=֥ ����UH��H���}��E���H��`�K H����  ���UH��H��   ��\���H��`���H��P�K H��H���i���H��`���H�5�� H������H�������H��`���H���f������UH��H�� H�}�H�u�H�U�H�M�H�E�H��H����
  �E��}� tdH�%    H������H�E���    �H�E���UH��H�� H�}�H�u�H�E�H�E�H���!	  H�E�H�}� u�    �!H�E�H�E�H��H�E��    H������H�E���UH��H�S� ��   H�5Q� H�=�� �R���UH��H��H�}�H�E��    �    H��������    ��UH��H��H�}�H�	� ��   H�5�� H�=8� �����UH��H���}������E�������UH��H���}��E�������UH��H���}�H��� ��   H�5�� H�=ߣ ����UH��H��H�}�H��� ��   H�5y� H�=�� �z���UH��H��H�}�H�|� ��   H�5N� H�=�� �O���UH��H��`H�}�H�u�H�U�H�M�L�E�H�E�    H�E�H�E�H�E�H;E�s|H�E�H+E�H��H�E�H�U�H�E�H�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���ЉE܃}� yH�U�H�E�H�H�E�뛃}� ~H�U�H�E�H�H��H�E��H�E��.H�E�H;E�tH��� ��   H�5s� H�=ݢ �t����    ��UH��H��`H�}�H�u�H�U�H�M�H�E�    H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�E�H��H�E�H�E�H;E���   H�E�H�E�H��H�E�H�H�E�H�M�H�U�H�E�H��H���Ѕ�����ufH�E�H�E�H�E�H�E�H�E�    H�E�H;E�sEH�U�H�E�H�� �E�H�U�H�E�H�H�M�H�U�H�� �H�U�H�E�H��EǈH�E�벐H�E��M���H�E��������UH��H���}�H�u� �  H�51� H�=l� �2���UH��H��H�}�H�N� �  H�5� H�=A� ����UH��H��H�}�H�(� �  H�5۠ H�=� �����UH��}�u�E��}�E��E��}�ЉE�H�E�]�UH��H��H�}�H�u�H�ٶ �'  H�5�� H�=�� ����UH��H��H�}�H�u�H��� �+  H�5W� H�=�� �X���UH��SH��HH�}�H�u���� H�E�H�E�H�E�H�U�H�E�H�H�E�H�E�H�E�H�E�H��H�E�H�}� uOdH�%    H������f�   dH�%    H������f�@  dH�%    H�������@    H�E��@	���bH�E�H� H��H�dH�%    H������H��H�U�H�u�H�E�H���ӉE�}� tH��� �;  H�5b� H�=ӟ �c���H�E�H+E�H��H[]�UH��H���   H��X���H��P���H��H���H��`���H��P�K H��H���4���H��`���H�5�� H���T���H������H��`���H���1���H��X���H��uH�&� �@  H�5 H�=� �����H��P���H��uH��� �A  H�5�� H�=W� ����H��H���H��uH�д �B  H�5l� H�=0� �m���H��P���� ��uH��� �C  H�5?� H�=� �@���H��P����H��X����҉�   ��UH��H��H�}��u�H�_� �H  H�5�� H�=/� �����UH��H��pH�}�H�u�H�U�蒚 H�E�f�E�  f�E�  �E�    H�E�    H�E�    H�E�H�E�H�E�H�E�H�E�H��    H�E�H�H�E�H�}� uNH�E�H� H�� H� H�M�H�U�H�u�H�}��ЉE�}� tH��� �U  H�5>� H�=�� �?���H�E��H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� tH�d� �Z  H�5� H�=a� �����H�E�H+E�H��H�E�H�E�H;E�sH�E�H��    H�E�H��     H�E���UH��H�� H�}�H�u�H�U�H�� �e  H�5�� H�=�� ����UH��H��P  H������H�=8� �yf  H��������   H������H��P�K H��H���Y���H������H�5� H���y���H��H������H��H���  H������H������H���A���H��������H��tIH��`���H��P�K H��H�������H�EH��H��`���H��H���4  H���V���H��`���H�������贓 H��H������H��H���  ���UH��H��   H��X���腓 H��H��X���H��H���  H�E�H�=� �_e  H������tXH��`���H��P�K H��H���C���H��`���H�5� H���c���H��H�E�H��H���y  H������H��`���H���.���H�E���UH��H��   H��X���H��P����ڒ H��H��P���H��X���H��H���  H�E�H�=l� �d  H������t|H��`���H��P�K H��H������H��`���H�5�� H������H��H��X���H��H����  H�5� H������H��H�E�H��H���  H�������H��`���H���X���H�E���UH��SH��8H�}�H�u�H�U�H�E�H��w
�  �   H�E�H�P�H�E�H!�H��t�  �~�ّ H��H�U�H�E�H��H���O  H� H��H����  H�E�H�}� u�  �CH�E�H�P�H�E�H!�H��tH�� ��  H�5\� H�=�� �]���H�E�H�U�H��    H��8[]�UH��H�� H�}�H�u�H�U�H��� ��  H�5� H�=M� ����UH��H���}��u��}�u�}���  uH��`�K H���   ���UH����  �   ����]�UH��H��H�}�H�E��q  H���   ���UH��H�}��u�H�E��U�H�E�ǀ�	     H�E����	  =o  wH�E����	  �P�H�E�Hcҋ�H�E����	  �P�H�E�Hcҋ���1�i�e�lH�E����	  ��H�E����	  �H�E�Hc҉�H�E����	  �PH�E����	  �x����]ÐUH��H�}��E�    �E�߰�H�E؋��	  =o  �N  �E�    �}��   kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE�E����  H�E�Hcҋ��U���1E�����D����1�H�E؋U�Hc҉��E���E��   �}�n  kH�E؋U�Hcҋ�%   ����E��PH�E�Hcҋ�%���	ȉE��E������H�E�Hcҋ��U���1E������D����1�H�E؋U�Hc҉��E��H�E؋��	  %   ���H�E؋ %���	ЉE�H�E؋�0  �U���1E�����D��1�H�E؉��	  H�E�ǀ�	      H�E؋��	  �HH�U؉��	  H�U�H����E�E���1E�E���%�V,�1E�E���%  ��1E�E���1E�E�]ÐUH��H�� H�}�H�u��U�H�U�H�E�H��H��� ���H�E��U��H�E���UH��H�}�H�E�H�     H�E�H�@    H�E�H�@    H�E�H�@    H�E�H�@     H�E��@(    �]�UH��H�}�H�E�H��?]�UH��H��H�}�H�U��   �������tH�� �   H�5�� H�=(� �X������UH��H�}�H�E��    ��]�UH��H��PH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH��� �   H�5<� H�=e� ����f���E�H�E��.   H���~ H�E�H�E�H������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� �����J  �������  �M��ɪ �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   ��� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH�n� �&   H�5� H�=;� ����H�E�H;E�sbH�E�H�E�� �����-I  ������uBH�E�� ����0�*��^E��M��X��E��M��ԩ �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E��~�� fW��E��E���UH��H��@H�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH�S� �   H�5� H�=� �p���f���E�H�EȾ.   H���A| H�E�H�E�H�������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sZH�E�� �����G  �������  �M���� �Y��E�H�E�� ����0�*��M��X��E�H�E��H�}� ��   �R� �E�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH�)� �&   H�5Œ H�=� �F���H�E�H;E�sbH�E�H�E�� ������F  ������uBH�E�� ����0�*��^E��M��X��E��M���� �Y��E�뛐����H�}� tH�E�H�U�H��}� t�E��x� W��E��E���UH��H��pH�}�H�u�H�E�� <-���E�H�E�� <+tH�E�� <-uH�E�H�E�� <0u=H�E�H��� <xtH�E�H��� <XuH�� �   H�5�� H�=̑ �$������}�H�E��.   H����y H�E�H�E�H������H�P�H�E�H�H�E�H�}� u
H�E�H���H�E�H�E�H�E�H�E�H�E�H;E�sNH�E�� �����mE  ��������   �m��-p� ���}�H�E�� ����0�E��E��m����}�H�E��H�}� ��   �-8� �}�H�E�H�E�H�E�H��� <0u=H�E�H��� <xtH�E�H��� <XuH��� �&   H�5�� H�=�� ����H�E�H;E�sVH�E�H�E�� �����D  ������u6H�E�� ����0�E��E��m����m����}��m��-�� ���}�말����H�}� tH�E�H�U�H��}� t�m����}��m���UH��H��H�}�H�u�H�U�H�E�H��H���0  H�E���UH��}�H�E�   �E�H9E�vH��`-J �U�H���U�E�   �E�H+E�H��H�E�E�H+E�H�P�E��H�H!�H�E�H�E�H��H�E؋E�Hc�H�E�H�H�E؉�H��H��]�UH��H��@H�}�H�E�   H�E������_���H9E�����tG�E�    �E�H�U�H��H9�s#�E����3���H9E�����t�E��   �E���H�E�H���   H�E�H������H��?   H)�H��H�E�H�E�H�E�H�E�H��H�E�H�E�   ��H��H�E�H)�H��H�E�   ��H��H��H�H�P�H�E���H��H��H�E�H�U�H�E�H�H�E�H�H���ÐUH��H��H�}�H�u�H�E�H� H�U�H��H����   ��ÐUH��H��H�}�H�u�H�E�H� H�U�H��H���
  ��UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���  ��UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]�UH��H��0H�}�H�u�H�E�H�������H�E�H� H�U�H�M�H��H���J
  H�E�H���������UH��SH��xH�}�H�u�H�}� �D  H�E�H�E�H�E�H�PH�E�H��H���}
  H�U�H�E�H��H����
  H�E�H�}� uH��    H��uH�=V� �u��H�E�� ����   H�E�H�@H9E�tH��    H��uH�=�� ��t��H�E�H�PH�E�H��H���  H�E�H�P H�E�H�@H   H��H)�H�E�H�P H�E�H���  H�E�H� H�U�H�RH��   H�U�H�RH�� ���H��H��H���%� �    �   H�E�� ��tH��    H��uH�=E� �0t��H�E�H���6  H�E�H�E�H�E�H%  ��H��H�E�H9�tH��    H��uH�=i� ��s��H�E؋@HH�H��H��H��H�E�H�H��H�E�H�E؋@H�������H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=� �zs��H�U�H�E�H��H���  H�E�H�@PH�����E�H�E؋@L��uH��    H��uH�=�� �1s��H�E�H�ƿ   �3���H��H���w
  H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H���e
  ����t�   ��    ��tH��    H��uH�=�� �r��H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H���F
  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���X	  H�E�H���  �   H�E�H���  ����H��x[]�UH��SH��   H��x���H��p���H��p��� uHǅp���   H��p��� �  ��  H��p���H���Y����E�}�~H��    H��uH�=� �q���E�H�H��H��H��H��x���H�H��H�E�H�U�H�E�H��H���  H�E�H�@H���*  H�E�H�@H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=ƌ �)q��H�E�H�U�H��H���  ����tH��    H��uH�=� ��p��H�E�H� H��t$H�E�H�U�H�H��H���K  ����t�   ��    ��tH��    H��uH�=� �p��H�E�H�H�E�H�PPH�E؋@L�PH�E؉PLH�E�H�@PH���$  H�E�H�PH�E�H��H���	  H�E�H��H���	  H��H�E�H�P��  H�E�H���@  �U�H��x�����H����	  H�E�H�E�H�@PH�E�H�E�H��uH��    H��uH�=�� ��o��H�E�H�U�H��H���L  ����tH��    H��uH�=، �o��H�E�H� H��t$H�E�H�U�H�H��H���	  ����t�   ��    ��tH��    H��uH�=� �`o��H�E�H�H�E�H�PPH�EЋ@L�PH�EЉPLH��x���H�PH�E�H��H���Z  H��x���H�PH�E�H��H���
  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H����  H�E�H����
  H�E�H�@PH��uH��    H��uH�=�� �n��H�E�H�PH�E�H��H���M  H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���  H�E�H���S  H�]�H�E�H���  �   H��p���H�  H% ���H�E�H�U�H��x���H��H���M
  H�E�H��x���H�PH�E�H��H���  H��x���H�PH�E�H��H����  H��x���H�P H�E�H�@H   H��H�H��x���H�P H�E�H���  H�E�H�@H��H�E�H����  H��H�Ĉ   []�UH��SH��hH�}�H�u�H�U�H�}� uH�U�H�E�H��H���!���H����  H�}� uH�U�H�E�H��H�������    �  H�E�H�E�H�E�H�PH�E�H��H���&  H�U�H�E�H��H���m  H�E�H�E�H����  H�}� uH��    H��uH�=� �l��H�E�� ����   H�E�H�E�H�E؋@H������H�E�H�E�H;E�w	H�]��  H�U�H�E�H��H���C���H�E�H�}� u
�    ��   H�U�H�M�H�E�H��H������H�U�H�E�H��H������H�]��   H�E�� ��tH��    H��uH�=Ǌ ��k��H�E�H�@H9E�tH��    H��uH�=� ��k��H�E�H�@H9E�sH�]��WH�U�H�E�H��H������H�E�H�}� u�    �2H�E�H�PH�M�H�E�H��H���a���H�U�H�E�H��H�������H�]�H�E�H���   H��H��h[]�UH��H��`H�}�H�u�H�U�H�E�H�5�� H������H�E�H���<���H�E�H�M�   H��H���:���H�E�H�U�H�M�H��H����  H�E�H�������H�E�H����������UH��H��H�}�H�u�H�E�H�U�H�H�E��@ H�E�H���  ���UH��H��H�}�H�E��@��tH�E�H���  ��ÐUH��H�� H�}�H�u�H�E�H��H����  H�E�H�}� ��   H�E�H�@H9E�sH�E�H����  H�E���H�E�H�PH�E�H�@H�H9E�rH�E�H���  H�E��H�E�H�@H9E�rH�E�H�PH�E�H�@H�H9E�rH��    H��uH�=T� �i��H�E���    ��UH��H��0H�}�H�u�H�E�H���)  H�E�H�E�H���7  H�E�H�}� uH�U�H�M�H�E�H��H���4  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���g	  H�E�H�E�H���  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���I	  ���UH��H��H�}�H�E��@����tH��    H��uH�=� �h��H�E�H� H�������H�E��@ ��ÐUH��H�}�H�E�H�     �]�UH��H�}�H�u�H�E�H�E�H�E�H�@H9E�r H�E�H�PH�E�H�@H�H9E�s�   ��    ]ÐUH��H�� H�}�H�u�H�E�H���  H������tH�E�H�U�H��H����
  �   H�E�H����
  H�E�H�E�H�HH�U�H�E�H��H���5  ��tAH�E�H���M  H������tH�E�H�U�H�M�H��H���J  �VH�E�H���  H�E��H�E�H���a  H������tH�E�H�U�H�M�H��H���_  �H�E�H���2  H�E��\�����UH��H��0H�}�H�u�H�E�H���
  H�E�H�E�H����  H�E�H�}� uH�U�H�M�H�E�H��H���0  �iH�}� uH�U�H�M�H�E�H��H���  �IH�E�H���c  H�E�H�E�H���F
  H��H�M�H�E�H��H����  H�U�H�M�H�E�H��H���E  ���UH��H�� H�}�H�E�H���Z	  H�E�H�}� u�    �,H�E�H����	  H������tH�E�H����	  H�E���H�E���UH��SH��XH�}��u�H�E�H� �   H���u H�E�H�E�H�� H%  ��H�EЋE��������H�E�H�E�    H�}�   w
H�E�HE���H�}��� vH��    H��uH�=)� �e��H�E�H�ƿ�   设��H�ø   H+E�H�M�H�U�H�4�U���H��H���  H�]�H�E�    H�E�    H�E�H�@H9E�sHH�E�H�PH�E�H�H�ƿ   �H���H��H������H�]�H�E�H�U�H�H�E�H�E�H�E�HE��H�E�H�U�H�PPH�E�H��X[]�UH��H�� H�}�H�u�H�E�H���`  H������tH�E�H�U�H��H���]  �   H�E�H���2  H�E�H�E�H�HH�U�H�E�H��H����  ��tAH�E�H���  H������tH�E�H�U�H�M�H��H���f  �VH�E�H����  H�E��H�E�H����  H������tH�E�H�U�H�M�H��H���]  �H�E�H����  H�E��\�����UH��H��H�}�H�E��@��tH��    H��uH�=�� ��c��H�E�H� H������H�E��@���UH��SH��(H�}�H�u�H�E�%�  H��tH��    H��uH�=�� �yc��H�E�H� H�U�H��   H��H����r H�E�H�E�H�ƿH   �Z���H��H�E�H��   H�E�H���   H���  H�]�H�E�H��([]�UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���  �UH�E�� ��t%H�E�� ��tH��    H��uH�=�� �b��H�u�H�E�A�    A�   �    �
   H���C  ��ÐUH��H�}�H�E�H� ]�UH��H��H�}�H�E�H���m  H�@��UH��H��H�}�H�E�H���O  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���-  H�E�H�}� tH�]�H�E�H����  H�X H�}� tH�]�H�E�H����  H�XH�E�H����  �@(������t8H�E�H����  ��tH�E�H���  �@(   �H�U�H�E�H��H����  H�E�H�������H��uH�E�H������H9E�t*H�E�H�������H9E�uH�E�H�������H��t�   ��    ��tH��    H��uH�=�� ��`��H�E�H���9  H�E�H�}� uH�E�H�U�H��rH�E�H���g���H9E�����tH�]�H�E�H����  H�X�EH�E�H���X���H9E�����tH��    H��uH�=�� �z`��H�]�H�E�H���  H�XH�}� tH�]�H�E�H���o  H�H�E�H���`  H�@    H�E�H���L  H�@    H�E�H���8  H�     H�E�H���%  H�@    H�E�H���  H�@     H�}� tH�U�H�E�H��H���5  �H��H[]�UH��H��H�}�H�E�H����  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H��� ���H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���H  H�X�EH�E�H�������H9E�����tH��    H��uH�=�� ��^��H�]�H�E�H���  H�XH�]�H�E�H����  H�H�E�H����  �X(H�E�H����  �X(H�]�H�E�H���  H�XH�}� tH�]�H�E�H���  H�H�]�H�E�H���  H�XH�}� tH�]�H�E�H���s  H�H�E�H���}���H������tH�]�H�E�H���c���H���B  H�X H�E�H���K���H��H�E�H���#  H�XH�E�H���)  H��H�E�H���  H�X H�E�H���
  H������tH�]�H�E�H����  H����  H�XH�E�H����  H�@    H�E�H���  H�@    H�E�H���  H�     H�E�H���  H�@    H�E�H���s  H�@     H�U�H�E�H��H����  H�U�H�E�H��H���  �H��H[]ÐUH��H�}�H�E�H� ]ÐUH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=ɀ ��\��H�E�H�U�H�H�U�H�E�H��H���  H�U�H�E�H��H���  ���UH��H�}�H�u�H�U�H�E�H�PH�E�H�@H9���]�UH��H��H�}�H�E�H���  H�@��UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=g� �"\��H�E�H������H������tH��    H��uH�=�� ��[��H�]�H�E�H���&  H�XH�]�H�E�H���  H�H�E�H���T  H�E�H�}� tH�]�H�E�H����  H�X H�]�H�E�H����  H�XH�]�H�E�H����  H�X H�]�H�E�H���  H�XH�U�H�E�H��H���  H�U�H�E�H��H���  H�U�H�E�H��H���  �H��8[]�UH��H��H�}�H�E�H���O  H�@�ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=� ��Z��H�E�H������H������tH��    H��uH�=� �Z��H�]�H�E�H����  H�XH�]�H�E�H���  H�H�E�H���  H�E�H�]�H�E�H���  H�X H�]�H�E�H���  H�XH�]�H�E�H���q  H�X H�}� tH�]�H�E�H���V  H�XH�U�H�E�H��H����  H�U�H�E�H��H���B  H�U�H�E�H��H����  �H��8[]ÐUH��SH��HH�}�H�u�H�U�H�E�H���@  H�E�H�E�H���=  H�E�H�}� tH�]�H�E�H����  H�X H�}� tH�]�H�E�H���  H�XH�E�H���  �@(������t8H�E�H����  ��tH�E�H���p  �@(   �H�U�H�E�H��H���  H�E�H������H��uH�E�H�������H9E�t*H�E�H���i���H9E�uH�E�H������H��t�   ��    ��tH��    H��uH�=-{ �X��H�E�H���I  H�E�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���  H�X�EH�E�H��� ���H9E�����tH��    H��uH�=S{ �X��H�]�H�E�H���R  H�XH�}� tH�]�H�E�H���7  H�H�E�H���(  H�@    H�E�H���  H�@    H�E�H���   H�     H�E�H����  H�@    H�E�H����  H�@     H�}� tH�U�H�E�H��H����  �H��H[]�UH��H��H�}�H�E�H���  H�@�ÐUH��SH��HH�}�H�u�H�U�H�E�H����  H�E�H�E�H������H�E�H�E�H�������H�E�H�}� uH�E�H�U�H��rH�E�H���o���H9E�����tH�]�H�E�H���  H�X�EH�E�H������H9E�����tH��    H��uH�=*z �V��H�]�H�E�H����  H�XH�]�H�E�H���  H�H�E�H���  �X(H�E�H���  �X(H�]�H�E�H���  H�XH�}� tH�]�H�E�H���i  H�H�]�H�E�H���V  H�XH�}� tH�]�H�E�H���;  H�H�E�H���}���H������tH�]�H�E�H���c���H���
  H�X H�E�H���K���H��H�E�H����  H�XH�E�H���9  H��H�E�H����  H�X H�E�H���  H������tH�]�H�E�H���   H���  H�XH�E�H���  H�@    H�E�H���v  H�@    H�E�H���b  H�     H�E�H���O  H�@    H�E�H���;  H�@     H�U�H�E�H��H���
  H�U�H�E�H��H���#  �H��H[]ÐUH��H�� H�}�H�u�H�U�M�H�E�H�M�H�U�   H���  H�E��U�PHH�E��@L    H�E�H�@P    H�E�H��XH����������UH��H��H�}�H�u�H�E�H� H��tH��    H��uH�=x �&T��H�E�H�U�H�H�U�H�E�H��H���	  H�U�H�E�H��H����  ���UH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=�w �S��H�E�H���I���H������tH��    H��uH�=x �S��H�]�H�E�H���  H�XH�]�H�E�H���  H�H�E�H������H�E�H�}� tH�]�H�E�H���\  H�X H�]�H�E�H���H  H�XH�]�H�E�H���4  H�X H�]�H�E�H���   H�XH�U�H�E�H��H���  H�U�H�E�H��H���<  H�U�H�E�H��H���  �H��8[]ÐUH��SH��8H�}�H�u�H�U�H�E�H��uH��    H��uH�=ow �R��H�E�H���/���H������tH��    H��uH�=�w �RR��H�]�H�E�H���b  H�XH�]�H�E�H���N  H�H�E�H���U  H�E�H�]�H�E�H���+  H�X H�]�H�E�H���  H�XH�]�H�E�H���  H�X H�}� tH�]�H�E�H����   H�XH�U�H�E�H��H���_  H�U�H�E�H��H���  H�U�H�E�H��H���]  �H��8[]ÐUH��H�� H�}��u�H�U�H�M�H�E��U�H�E�H�U�H�PH�E�H�U�H�PH�E�H��H���������UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�}��   H�E�H�]�UH��H��H�}�H�E�H�������H�@ ��UH��H��H�}�H�}� u�    �H�E�H�������@(�����ÐUH��SH��XH�}�H�u�H�E�H���}����@(������tH��    H��uH�=�u �6P��H�E�H���s  H�E�H�}� �\  H�E�H������H9E�������   H�E�H������H������tH��    H��uH�=�u ��O��H�E�H���}���H��������@(��������   H�E�H���X���H�E�H�E�H���H���H��H�E�H��H���  H�E�H������H9E�����tH��    H��uH�=�u �LO��H�E�H���`����@(   H�E�H���M����@(   H�E�H�������H�E��  H�E�H������H9E�����tH��    H��uH�=�u ��N��H�E�H���o���H������tH��    H��uH�=�u �N��H�E�H���?���H�������@(������tzH�E�H������H�E�H�U�H�E�H��H���  H�E�H������H9E�����tH��    H��uH�=�u �;N��H�E�H���O����@(   H�E�H���<����@(   H�E�H������H�E�H�E�H������H����  ��tH�E�H������H���  ��t�   ��    ��toH�E�H��������@(������t+H�E�H��������@(   H�U�H�E�H��H��������  H�E�H�������@(   H�E�H�������@(   �  H�E�H���j����@(�E�H�E�H�������H9E������  H�E�H������H���i�����tH�E�H������H����  ��t�   ��    ��tQH�E�H���x���H�E�H�U�H�E�H��H���h  H�E�H��������@(   H�E�H��������@(   H�E�H�E�H�E�H���E���H�����������tH��    H��uH�=0t �cL��H�U�H�E�H��H���R  H�E�H���d����@(   �]�H�E�H���N����X(H�E�H�������H���7����@(   �M  H�E�H������H9E�����tH��    H��uH�=t ��K��H�E�H������H��������tH�E�H���Q���H���~  ��t�   ��    ��tQH�E�H���G���H�E�H�U�H�E�H��H���y  H�E�H�������@(   H�E�H���x����@(   H�E�H�E�H�E�H�������H����������tH��    H��uH�=�s �K��H�U�H�E�H��H���  H�E�H�������@(   �]�H�E�H��������X(H�E�H���k���H��������@(   ��H��X[]�UH��H��H�}�H�E�H������H� ��UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H���  ����uH�E�H������H�E��Ԑ���UH��H��H�}�H�u�H�E�H���x  ��ÐUH��H��H�}�H�u�H�E�H���g  ��ÐUH��H�� H�}�H�u�H�E�H���	  H�E�H�}� uH�E�H���#  �@(   �  H�E�H���  �@(   H�E�H����  �@(��������  H�E�H���L	  H�E�H�}� tH�E�H����  �@(��t�   ��    ��tH��    H��uH�=3r �NI��H�E�H�������H9E�uH�E�H������H����  ��t�   ��    ��tYH�E�H���L  �@(   H�E�H���9  �@(   H�E�H������H���  �@(   H�U�H�E�H��H��������  H�E�H������H9E�uH�E�H���%���H���U  ��t�   ��    ��tYH�E�H���  �@(   H�E�H���  �@(   H�E�H�������H���  �@(   H�U�H�E�H��H�������j  H�E�H������H9E�������   H�E�H�������H9E�����t;H�U�H�E�H��H���C  H�U�H�E�H��H����  H�E�H���  �@(   �&H�U�H�E�H��H���  H�E�H����   �@(   H�E�H����   �@(   �   H�E�H���N���H9E�����tH��    H��uH�=�p �LG��H�E�H�������H9E�����t;H�U�H�E�H��H���"  H�U�H�E�H��H���o  H�E�H���G   �@(   �&H�U�H�E�H��H���G  H�E�H���   �@(   H�E�H���   �@(   ����UH��H�}��X   H�E�H�]�UH��H�� H�}�H�u�H�E�H�E�H�}� t&H�E�H����  ����uH�E�H���  H�E��Ԑ���UH��H��H�}�H�E�H������H�@ ��UH��H��H�}�H�}� u�    �H�E�H���^����@(�����ÐUH��SH��XH�}�H�u�H�E�H���5����@(������tH��    H��uH�=_k ��E��H�E�H���s  H�E�H�}� �\  H�E�H���+���H9E�������   H�E�H���e���H������tH��    H��uH�=ak �dE��H�E�H���5���H�������@(��������   H�E�H������H�E�H�E�H��� ���H��H�E�H��H���q  H�E�H������H9E�����tH��    H��uH�=5k ��D��H�E�H�������@(   H�E�H�������@(   H�E�H������H�E��  H�E�H���v���H9E�����tH��    H��uH�=)k �tD��H�E�H�������H������tH��    H��uH�=Yk �DD��H�E�H�������H���t����@(������tzH�E�H������H�E�H�U�H�E�H��H���   H�E�H�������H9E�����tH��    H��uH�=<k ��C��H�E�H�������@(   H�E�H��������@(   H�E�H���%���H�E�H�E�H������H���%  ��tH�E�H���R���H���  ��t�   ��    ��toH�E�H�������@(������t+H�E�H���x����@(   H�U�H�E�H��H��������  H�E�H���M����@(   H�E�H���:����@(   �  H�E�H���"����@(�E�H�E�H���T���H9E������  H�E�H���9���H���i�����tH�E�H���v���H���1  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���Z  H�E�H�������@(   H�E�H�������@(   H�E�H�E�H�E�H�������H�����������tH��    H��uH�=�i ��A��H�U�H�E�H��H���D
  H�E�H�������@(   �]�H�E�H�������X(H�E�H������H��������@(   �M  H�E�H���p���H9E�����tH��    H��uH�=�i �nA��H�E�H���?���H��������tH�E�H�������H����  ��t�   ��    ��tQH�E�H�������H�E�H�U�H�E�H��H���k	  H�E�H���C����@(   H�E�H���0����@(   H�E�H�E�H�E�H���Y���H����������tH��    H��uH�=5i �@��H�U�H�E�H��H���
  H�E�H��������@(   �]�H�E�H�������X(H�E�H�������H�������@(   ��H��X[]�UH��H��H�}�H�E�H���w���H� ��UH��H�� H�}�H�u�H�E�H���[���H�E�H�}� uH�E�H�������@(   �  H�E�H�������@(   H�E�H��������@(��������  H�E�H�������H�E�H�}� tH�E�H�������@(��t�   ��    ��tH��    H��uH�=Oh �j?��H�E�H�������H9E�uH�E�H������H��������t�   ��    ��tYH�E�H���D����@(   H�E�H���1����@(   H�E�H������H�������@(   H�U�H�E�H��H��������  H�E�H������H9E�uH�E�H���T���H��������t�   ��    ��tYH�E�H�������@(   H�E�H�������@(   H�E�H������H�������@(   H�U�H�E�H��H�������j  H�E�H�������H9E�������   H�E�H�������H9E�����t;H�U�H�E�H��H���  H�U�H�E�H��H���  H�E�H��� ����@(   �&H�U�H�E�H��H���f  H�E�H��������@(   H�E�H��������@(   �   H�E�H���F���H9E�����tH��    H��uH�=�f �h=��H�E�H�������H9E�����t;H�U�H�E�H��H����  H�U�H�E�H��H���-  H�E�H���?����@(   �&H�U�H�E�H��H���  H�E�H�������@(   H�E�H�������@(   ����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��R H�E��E�    �E���~H��    H��uH�==f �<���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=f �<���E��P�U�H��D�-H�U�H�E�H��H���:���� 9E�����tE�E�    H�U�H�E�H��H������� �U�)�9E�����t�U�H�E���H��蒤���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���[����E��ڋE����E�}� x!�E�H��D���H�E���H���+����m��ِ��UH��H��H�}�H�}� u�   �H�E�H���*����@(�����ÐUH��SH��8H�}�H�u�H�E�H���*���H�E�H�}� tH�E�H������H9E�t�   ��    ��tH��    H��uH�=�d �:��H�E�H���)���H�E�H�E�H�������H�E�H�}� tH�]�H�E�H������H�H�]�H�E�H���p���H�XH�]�H�E�H���\���H�H�]�H�E�H���I���H�XH�]�H�E�H���5���H�H�}� uH�E�H�U�H��rH�E�H������H9E�����tH�]�H�E�H�������H�X�EH�E�H���~���H9E�����tH��    H��uH�=ed �9��H�]�H�E�H������H�XH�U�H�E�H��H���'���H�U�H�E�H��H�������H��8[]�UH��SH��8H�}�H�u�H�E�H������H�E�H�}� tH�E�H�������H9E�t�   ��    ��tH��    H��uH�=d ��8��H�E�H������H�E�H�E�H���'���H�E�H�}� tH�]�H�E�H�������H�H�]�H�E�H�������H�XH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H������H�H�}� uH�E�H�U�H��rH�E�H�������H9E�����tH�]�H�E�H���W���H�X�EH�E�H�������H9E�����tH��    H��uH�=�c � 8��H�]�H�E�H������H�XH�U�H�E�H��H������H�U�H�E�H��H���t����H��8[]�UH��H�}��    ]�UH��H�}��    ]�UH��SH��8H�}�H�u�H�E�H���8���H�E�H�}� tH�E�H���I���H9E�t�   ��    ��tH��    H��uH�=�a �<7��H�E�H������H�E�H�E�H�������H�E�H�}� tH�]�H�E�H���I���H�H�]�H�E�H���6���H�XH�]�H�E�H���"���H�H�]�H�E�H������H�XH�]�H�E�H�������H�H�}� uH�E�H�U�H��rH�E�H������H9E�����tH�]�H�E�H������H�X�EH�E�H���D���H9E�����tH��    H��uH�=a �B6��H�]�H�E�H���v���H�XH�U�H�E�H��H�������H�U�H�E�H��H��������H��8[]�UH��SH��8H�}�H�u�H�E�H������H�E�H�}� tH�E�H���T���H9E�t�   ��    ��tH��    H��uH�=�` �5��H�E�H���m���H�E�H�E�H���5���H�E�H�}� tH�]�H�E�H������H�H�]�H�E�H������H�XH�]�H�E�H������H�H�]�H�E�H���o���H�XH�]�H�E�H���[���H�H�}� uH�E�H�U�H��rH�E�H���|���H9E�����tH�]�H�E�H������H�X�EH�E�H������H9E�����tH��    H��uH�='` �4��H�]�H�E�H�������H�XH�U�H�E�H��H���I���H�U�H�E�H��H���6����H��8[]�UH��H��H�}�H�}� u�   �H�E�H���~����@(������UH��H�� �}��BG H�E��E���H�U�H�E���H����  �E�}� t�    ���[ H�E���H���\P ����UH��H�� �}���F H�E��E���H�U�H�E���H���  �E�}� t�    ��l[ H�E���H����P ����UH��H�� �}��F H�E��E���H�U�H�E���H���5  �E�}� t�    ��[ H�E���H���6Q ����UH��H�� �}��@F H�E��E���H�U�H�E���H����  �E�}� t�    ���Z H�E���H���Q ����UH��H�� �}���E H�E��E���H�U�H�E���H���  �E�}� t�    ��jZ H�E���H���FR ����UH��H�� �}��E H�E��E���H�U�H�E���H���3  �E�}� t�    ��Z H�E���H��� T ����UH��H�� �}��>E H�E��E���H�U�H�E���H����
  �E�}� t�    ��Y H�E���H���dT ����UH��H�� �}���D H�E��E���H�U�H�E���H���
  �E�}� t�    ��hY H�E���H����T ����UH��H�� �}��D H�E��E���H�U�H�E���H���1
  �E�}� t�    ��Y H�E���H���dU ����UH��H�� �}��<D H�E��E���H�U�H�E���H����	  �E�}� t�    ��X H�E���H����U ����UH��H�� �}���C H�E��E���H�U�H�E���H���	  �E�}� t�    ��fX H�E���H���,V ����UH��H�� �}��C H�E��E���H�U�H�E���H���/	  �E�}� t�    ��E����!
  ����UH��H�� �}��EC H�E��E���H�U�H�E���H����  �E�}� t�    ��E���������UH��H�� �}��C H�E��M�H�U�H�E���H���IC �E�}� t�    ��~W H�E���H���L ����UH��H�� �}��.C H�E��M�H�U�H�E���H����B �E�}� t�    ��+W H�E���H���L ����UH��H�� �}���B H�E��M�H�U�H�E���H���B �E�}� t�    ���V H�E���H����L ����UH��H�� �}��B H�E��M�H�U�H�E���H���PB �E�}� t�    ��V H�E���H���M ����UH��H�� �}��5B H�E��M�H�U�H�E���H����A �E�}� t�    ��2V H�E���H���N ����UH��H�� �}���A H�E��M�H�U�H�E���H���A �E�}� t�    ���U H�E���H����O ����UH��H�� �}��A H�E��M�H�U�H�E���H���WA �E�}� t�    ��U H�E���H���2P ����UH��H�� �}��<A H�E��M�H�U�H�E���H���A �E�}� t�    ��9U H�E���H���P ����UH��H�� �}���@ H�E��M�H�U�H�E���H���@ �E�}� t�    ���T H�E���H���8Q ����UH��H�� �}��@ H�E��M�H�U�H�E���H���^@ �E�}� t�    ��T H�E���H���Q ����UH��H�� �}��C@ H�E��M�H�U�H�E���H���@ �E�}� t�    ��@T H�E���H���R ����UH��H�� �}���? H�E��M�H�U�H�E���H���? �E�}� t�    ��E�����  ����UH��H��  H������H������H������H��H����  H������H�5�Y H����  H������H������H������H��H���  ��t
�   �X  H������H�5�Y H���  H������H������H������H��H����  ��t
�   �  H������H�5IY H���`  H������H������H������H��H���  ��t
�   ��  H������H�5Y H���  H������H������H������H��H���N  ��t
�   �  H������H�5�X H����  H������H������H������H��H���
  ��t
�   �H  H������H�5�X H���  H������H������H������H��H����  ��t
�   �  H�� ���H�5QX H���P  H�� ���H�����H������H��H���  ��t
�   ��  H�����H�5X H���  H�����H�����H������H��H���>  ��t
�   �|  H�� ���H�5�W H����  H�� ���H��(���H������H��H����  ��t
�	   �8  H��0���H�5�W H���  H��0���H��8���H������H��H���  ��t
�
   ��   H��@���H�5YW H���@  H��@���H��H���H������H��H���r  ��t
�   �   H��P���H�5W H����  H��P���H��X���H������H��H���.  ��t�   �oH��`���H��P�K H��H���$���H��`���H�5�V H���D���H��H������H��H���/���H�5�V H��� ���H���j���H��`���H��������    ��UH��H���}�H�u�H�0W �  H�5�V H�=�V 腉��UH��H�� �}��+; H�E��E���H�U�H�E���H����   �E�}� t�E���O H�E���H���-N ��UH��H�� �}���: H�E��E���H�U�H�E���H���y   �E�}� t�E���\O H�E���H���N ��UH��H���}�H�tV �  H�5�U H�=�U 蹈��UH��H���}�H�ZV �$  H�5�U H�=�U 菈��UH��H��`H�}���H�U��E��E��E��E���x H�E��@��t�U�H�E���    ��   H�E�H�E�H�E�H��H�E�H�E�H�E�H�E�H��H�E�f�E�  f�E�  �E�    H�E�H� H��H� H�M�H�U�H�u�H�}��ЉE��}� t�E��]H�U�H�E�H9�tH�YU �>   H�5�S H�=T 趇��H�U�H�E�H9�tH�-U �?   H�5�S H�=�S 芇���    ��UH��}��}�v�}�t�}�v�}��   w�   ��    ]�UH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�PH�E�H�� ��tH�E�H�@H�PH�E�H�P�Ԑ]�UH��H�}�H��H��H��H�E�H�U�H�E�H�PH�E�H9�t�    �LH�E�    H�E�H�@H9E�s1H�E�H�H�E�H��H�M�H�E�H�� 8�t�    �H�E����   ]�UH��ATSH���   H��H��H��H�� ���H�����H�E�    H�� �K H� H�U�H��H�H� H���F  H�� �K H� H�U�H��H�H�H�����H��H������H������    �=   H����  H�E�H�}����   H�� ���H��P�K H��H������H�� ���H�5�S H������H��H�����H����  I��H�����H����  H��H�E�L��H���8  H�U�H�E�H��H��H����  H�5�S H��觇��H������H�� ���H��脇���GH�U�H������    H���  H�E�H�U�H�� ���H�����H�E�H��H��������tH�E��H�E�����H������H���   [A\]�UH���� ������tRH�=� ��K ������t=��1 H�0H�=� �  H�=� �L H��� H�5w H����F H���	|��H�a ]�UH��H�� ����H�E�H�E�H����  H��H�� �K H� H9�������   H�E�H����  H�E�    H�� �K H� H�U�H��H�H� H��t+H�� �K H� H�U�H��H�H�E�H��H���  H�E��H�E�    H�U�H�E�H��H���	  H�E�H���J  H��H�� �K H�����UH��SH��HH��H��H��H��H��H�u�H�}�H�U��ȈE�����H�E�H�E�H����  H��H�� �K H� H9�����tH��f �>   H�5�Q H�=�Q �+���H�U�H�E�H��H������H�E�H�}��t&�}� ��   H�]�H�U�H�E�H��H����  H��fH�E�H����  H� H������tH�f �F   H�56Q H�=pQ 诂��H�]�H�E�H���  H�H�E�    H�U�H�E�H��H����  H�E�H���  H��H�� �K H��H��H[]�UH��SH��(H��H��H��H�E�H�U��f���H�E�H�E�H����  H��H�� �K H� H9�����tH�ve �Q   H�5�P H�=�P �����H�U�H�E�H��H���f���H�E�H�}��uH��    H��uH�=�P �V ��H�E�H����  H��vH�E�H���  H� H��t�   ��    ��tH��d �W   H�5�O H�=�P �n���H�E�H���  H�P�H�E�H��H���,  H��H�U�H�E�H��H���  H��H���v  H�E�H���  H�E�H���  H�     H�E�H���  H��H�� �K H��H��([]�UH��H��@H�}�H�U�H�E�H��H���|���H�U�H�E�H��H���:���H�E�H�}��u
�    �   H�� �K H� H�U�H��H�H�H�E�H��H���-���H�Eк    �=   H���O  H�E�H�}��uH��c �i   H�5�N H�=�O �@���H�E�H���m  H��H�E�H��H���UH��SH��8H�}�H�U�H�E�H��H������H�Eк    �=   H����  H�E�H�}��uH�Xc �q   H�5KN H�=O �����S���H�U�H�Eо    H���=  H�u�H��H��H��H�й   H��H��������    H��8[]�UH��ATSH��  H������H������������H������H�����H��H�������H������    �=   H���  H�E�H�}����   H�� ���H��P�K H��H������H�� ���H�5}N H���;���H��H�����H���  I��H�����H���  H��H�E�L��H���q  H�U�H�E�H��H��H����  H�5@N H�������H���*���H�� ���H��轀��dH�%    H�������   �������   H������H������H�����H�5�M H�Ǹ    ��O  ������tH��a ��   H�5�L H�=�M �	~��H�����H��uH�ya ��   H�5eL H�=�M ��}���m��������� ��D��H�����H������H�E�H��H���[���H�u�H�E�D��H��H��H��������    H��  [A\]�UH��H�� H�}�����H�U�H�E�H��H������H�U�H�E�H��H��������    �ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H�}��H�U؈E�H�E�H�E�H�E�H�@H9E�s#H�E�H�H�E�H�� 8E�uH�E��H�E���H������]ÐUH��H�}�H�E�H� ]ÐUH��H�}�H�E�H�@]�UH��H�� H�}�H��H��H��H�E�H�U�H�U�H�E�H��H���S  H�E���UH��H��0H�}�H�u�H�U�H�U�H�E�H�H�E�H�@H9�vH��    H��uH�=/L ���H�E�H�H�E�H�H�U�H�E�H��H���.  H�E�H�U���UH��SH��H�}�H�u�H�]�H�E�H���-  H�H�E�H�@    H�E�H�@    H�E�H�@    �H��[]�UH��H�� H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H�U�H�RH��H��舣����ÐUH��H�}�H�E�H�@]�UH��H�}�H�E�    H�E�H�@H9E�sH�E���H�E�H�@    �]�UH��H�� H�}�H�u�H�E�H�@H�PH�E�H��H���[  H�E�H�PH�E�H�@H��H�H�ƿ   �xr��H�U�H�H�H�E�H�E�H�@H�PH�E�H�PH�E��ÐUH��SH��(H�}�H�u�H�E�H�@H�PH�E�H��H����  H�E�H���   H��H�E�H�PH�E�H�@H��H�H�ƿ   ��q��H�H�E�H�E�H�@H�PH�E�H�PH�E�H��([]ÐUH��H�}�H�u�H�E�H�@H�U�H��H�]ÐUH��H�}�H�E�H�PH�E�H�@H��H��H�]ÐUH��H�}�H�E�H�@]�UH��H�}�H�E�H� ]�UH��H�� H�}�H�u�H�E�H�������H�E�H�E�H�������H��H�E�H�H�E�H������H��H�E�H����UH��H�� H�}�H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��H�H���a���H�E�H�E���UH��H��0H�}�H�u�H�E�H���p��H�M�H�U�H�E�H�0H�@H��H���H  H�E�H���q�����UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H�}�H�E�H� ]ÐUH��SH��8H�}�H�u�H�E�H�@H9E���   H�E�H�H�E�H�E�H�U�H��H��H��蝠��H�E�H�E�    H�E�H�@H9E�sHH�E�H�@H�U�H��H�H���X���H��H�E�H��    H�E�H�H�ƿ   �o��H�H�E��H�E�    H�E�H�@H9E�sH�E���H�E�H�U�H�RH��H���ݟ��H�E�H�U�H�PH�E�H�U�H�P��H��8[]�UH��H��PI��H��L��L��H��H�u�H�}�H�U�H�M�H�E�H�E�H�E�    H�E�H9E���  H�U�H�E�H�� �E�}�`v�}�zv�}�@v �}�Zw�E���H�E���H���~���q  �}�/v �}�9w�E���H�E���H���z~���K  �}� uH�E��    H���^~���/  �E��H�=%G � H������t�E���H�E���H���(~����   �}�\uH�E�H�5	G H���z����   �}�"uH�E�H�5�F H���z���   �}�'uH�E�H�5�F H���lz���   �}�
uH�E�H�5�F H���Nz���   �}�	uH�E�H�5�F H���0z���fH�E�H�5�F H���z��H�E�H�M��   H��H��诔���E�E�H�U�H�M�H�E�H��H���*   H�E�H���_n��H�E��}   H���*}��H�E��4������UH��H��@H�}�H�u�H�U�H�U�H�E�H��H���m��H�E؋ H�U�H�M�H�Ή��2y��H�E�H����m����ÐUH��H��H�}�H�u�H����K H�PH�E�H�H�E��@H    H�E��@L    H�E�H�U�H�PPH�E�H��XH���   H�E�H�@    H�E�H�@�   H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�@0    H�E�H�@8    H�E��@@    H�E��@D    H�E�H��H�=�� �7   ���UH��H���   H��H���H����K H�PH��H���H�H��H���H�P0H��H���H�@8H9�tFH��`���H��P�K H��H���3v��H��`���H�5X H���Sv��H���v��H��`���H���0v��H��H���H�@H��t��  H��H��H���H�@H��H���ܛ��H��H���H��H�=�� �!  H��X���H��X���H��H�=�� �I!  ���UH��H��H�}�H�E�H�������H�E��p   H���d���ÐUH��H��H�}�H�E�H�@PH��tH�E�H�@PH�U�H�������ÐUH��H���   H��(���H�� ���H�����H�����H�����H��uH��s �W   H�5"W H�=?W ��r��H��(���H���u  ������t
������%  H��(����@L����   H��(���H� H��(H� H�����H��8���H�� ���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��  H��8���H��uH��(����@D����H��(����PDH��8���H�����H��    �y  H��(����@@��tVH��(���H�@(H��tFH��@���H��Q�K H��H���5k��H��@���H�53V H���Uk��H���k��H��@���H���2k��H��(����@@    H��(���H�PH��(���H�@(H9��  H��(���H���
  �E��}� t�E���  H��(���H���  �E�}� t�E��  H��(���H���4  H��(���H� H��(H� H��(���H�RH��(���H�qH��0���H��(����ЉE��}� t!H��(����@D����H��(����PD�E��8  H��0���H��u1H��(����@D����H��(����PDH�����H�     �    ��   H��0���H��(���H�P H��0���H��(���H�P(H��(���H�PH��(���H�@(H9�rH�q ��   H�5xT H�=�T �1p��H��(���H�P(H��(���H�@H)�H��H�E�H�����H�E�H��H���   H� H�E�H��(���H�PH��(���H�@H�H�U�H�� ���H��H���Bx��H��(���H�PH�E�H�H��(���H�PH�����H�U�H��    �ÐUH��H��   H�����H�����H�����H�� ���H�����H��uH�p ��   H�5�S H�=�S �?o��H�����H����  ������t
������Q  H������@L����   H�����H�P0H�����H�@8H9�tH��o ��   H�5S H�=�S ��n��H�����H� H��0H� H�����H�� ���H�����H������ЉE��}� t!H������@D����H������PD�E��  H�� ���H��uH�+o ��   H�5�R H�=$S �Ln��H�� ���H�� ���H��    �e  H�����H�PH�����H�@H9�u@H�����H���2  �E�}� t�E��*  H�����H���&
  �E��}� t�E��
  H������@@��uVH�����H�@(H��tFH��0���H��Q�K H��H����f��H��0���H�5�Q H���g��H���hg��H��0���H����f��H������@@   H�����H�PH�����H�@H9�rH�	n ��   H�5qQ H�=LR �*m��H�����H�PH�����H�@H)�H��H�E�H�����H�E�H��H���  H� H��(����E� H������@L��u@H��(���H������
   H���N H�E�H�}� tH�E�H��H+����H��(����E�H��(���H��uH�Km ��   H�5�P H�=�Q �ll��H�����H���d	  H��(���H�����H�HH�����H�@H�H�����H��H���t��H�����H�P0H�����H�@8H9�trH�����H�PH�����H��0H��H���  H�H�����H�P0H�����H�PH��(���H�H�E�H�����H�P8H�E�H��H���M���H�H�����H�P8�6H�����H�PH�����H�P0H�����H�PH��(���H�H�����H�P8H�����H�P(H�����H�HH��(���H�H�E�H�E�H��H���ԓ��H�H�����H�P(H�����H�PH��(���H�H�����H�P�}� tH�����H���  ������t������H��(���H�� ���H��    �ÐUH��H��H�}����E�H�E�H�@H��uH�qk ��   H�5�N H�=�O �j��H�E�H�@H�P�H�E�H�PH�E�H�PH�E�H�@H��E���ÐUH��H��H�}��u�H�E�H�P0H�E�H�@8H9�tH�k ��   H�5_N H�=hO �j��H�E��U�PL�    ��UH��H�}�H�E�H�@    H�E�H�@     H�E�H�@(    H�E�H�P0H�E�H�P8�]ÐUH��H�� H�}�H�E�H�P8H�E�H�@0H9�tH�E�H����  �E��}� t�E��+H�E�H���  �E��}� t�E��H�E�H���_����    ��UH��H�� H�}�H�u�H�E�H� H��8H� H�U�H�}�H�Ѻ   �    �ЉE��}� t�E��)H�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H��    ��UH��H��@H�}�H�uЉU�H�E�H����  �E��}� t�E���   �}�ueH�E�H�@H��H�E�H�@ H)�H�E�H�H�E�H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� ��   H�E؋@D����H�E؉PD�E��|�}� t%�}�tH�%i �  H�5rL H�=�M �+h��H�E�H� H��8H� H�M��U�H�u�H�}��ЉE�}� tH�E؋@D����H�E؉PD�E��H�E�H��������    �ÐUH��H�� H�}�H�E�@H��t�    �_H�E�H� H��H� H�U�H�JHH�U�H��H���ЉE��}� t�E��/H�E�@H��uH�bh �%  H�5�K H�=8M �_g���    �ÐUH��H��H�}�H�E��@L��t�    �aH�E�H� H�� H� H�U�H�JLH�U�H��H���Ѕ�����t������/H�E��@L��uH��g �/  H�5$K H�=�L ��f���    �ÐUH��H��0H�}�H�E�H��������E��}� t�E���  H�E�H�P0H�E�H�@8H9�u
�    �  H�E؋@H��u\H�E�H� H��8H� H�U�H�R0H��H�U�H�R H��H)�H�U�H�}�H�Ѻ   �ЉE��}� t�E��S  H�E�H�P0H�E�H�P �_H�E؋@H��tH�g �B  H�5AJ H�=L ��e��H�E�H�P H�E�H�@0H9�tH��f �C  H�5J H�=L ��e��H�E�H�P H�E�H�@8H9���   H�E�H� H��0H� H�U�H�J8H�U�H�R H)�I��H�U�H�JH�U�H�R H�4H�U�H�}�H��L���ЉE�}� tH�E؋@D����H�E؉PD�E��`H�E�H��uH�?f �M  H�5cI H�=�I �e��H�E�H�P H�E�H�H�E�H�P H�E�H�P0H�E�H�H�E�H�P0�#����    �ÐUH��H���   H��8���H��8���H��������E��}� t�E���   H��8����@H����   H��8���H�@H��H��8���H�@ H)�H��H�E�H��8���H� H��8H� H��H���H�u�H��8���H�Ѻ   �ЉE�}� ttH��8����@D����H��8����PDH��P���H��P�K H��H���*f��H��P���H�5[J H���Jf��H�E��H���  H���f��H��P���H���f���E���    ��    ��UH��H�� H�}�H�E�H��������E��}� t�E��   H�E�@H��u4H�E�H�PH�E�H�@(H9�tH��d �m  H�5�G H�=�I �Xc��H�E�H�P0H�E�H�@8H9�tH�Sd �o  H�5kG H�=�G �$c��H�E�H�@    H�E�H�@     H�E�H�@(    �    ��UH��H�� H�}�H�E�H�@H��uH��c �x  H�5G H�=MI ��b��H�E�H�@H��u-�� H��H�E�H�@H��H�������H�E�H�E�H�U�H�P���ÐUH��H�� H�}��u�H�U�H�E�H�U�H��H������H����K H�PH�E�H�H�E��U�Pp��ÐUH��H�}�H�E��@p]ÐUH��H��   H��X���H��X���H�P0H��X���H�@8H9�tFH��`���H��P�K H��H����c��H��`���H�5rH H���d��H���hd��H��`���H����c��H��X����@p���= �E��}� t�E���    �ÐUH��H�� H�}�H�u�H�E�@pH�U�H�Ѻ   �    ���: �E��}� uH�E��    �    ��}�-  uH�E��    �    ��E���UH��H��   H��X���H��P���H��    H��u6H�@b ��  H�5,E H�=�G ��a��H��P����    �    �   H��X����@p���P����E��}� uH��P����    �    �h�}�"  uH��P����    �    �KH��`���H��P�K H��H���b��H��`���H�5_G H���b��H����b��H��`���H���b��������ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u����z �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�M�H�E�@pH�M�H�U�H�u����
 �E��}� t�E��H�E�H��H�E�H��    �ÐUH��H��0H�}�H�u��U�H�M�H�E�@pH�MЋU�H�u����1 �E��}� t�E���    �ÐUH��H�}��]ÐUH��H���   H��8���H�Q� H�E�H�E�H����  H��H���H�E�H���  H��@���H��@���H��H���H��H���"  ����   H��H���H���e  H�E�H�E�H��������E�}� tFH��P���H��P�K H��H���`��H��P���H�5�E H����`��H���a��H��P���H���`��H��H���H����  �]������UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���������UH��H��H�}�H�E�H�������ÐUH��H��H�}�H�u���
 H��H�E�H��H���  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��p  H������H������H�������+   H���b�  H�����E�H������� <ru�}� t�E�   �   �E�   �   H������� <wu�}� t	�E�   ��E�   �M�  �oH������H��P�K H��H���_��H������H�5sD H���5_��H��H������� ����H���  H�5aD H���_��H���V_��H������H����^��H������H������� ����   H������� <+u
H��������H������� <bu
H�������H������� <eu�M� @  H�������H��P���H��P�K H��H���=^��H��P���H�5�C H���]^��H��H������H��H���H^��H�5�C H���9^��H���^��H��P���H���^��H�������(���H�������M�H��������H���� �E�}� tdH�%    H������H�E��    �.� H��H�U�H������H��H���  H��tH����    ��UH��H��H�}�H�u��Q H��H�E�H��H���	  ���UH��H��H�}�H�E�H�ƿ    �����ÐUH��H�}�H�����]�UH��H��   ��\���H��P���H��`���H��P�K H��H����\��H��`���H�5tB H��� ]��H�5�B H����\��H���;]��H��`���H����\��� H��H�U�H��\���H��H���S  H��tH����    ��UH��H�� H�}�H�}� t
H�E�H����    H�E��E�    H�E�H���[���������t�E�����H�E�H� H��H� H�U�H���Ѕ�����t�E�����H�E�H�������E���UH��H��0H�}�H�u��U�H�}� t
H�E�H����    H�E��U�H�M�H�E�H��H�������E�}� tdH�%    H������H�E��������    ��UH��H��0H�}�H�}� t
H�E�H����    H�E�H�U�H�E�H��H��������E�}� t!dH�%    H������H�E�H�������H�E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H������������t�������    ��UH��H��H�}�H�E�H��������UH��H��@H�}�H�uЉU�H�M�H�}� t
H�E�H����    H�E��}�u@H�E��   H��������E�}� ��   dH�%    H������H�E�������   �}�u9H�E��   H�������E��}� t{dH�%    H������H�E��������a�}�u9H�E��   H���t����E�}� t<dH�%    H������H�E�������"dH�%    H�������   �������    ��UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E��    �    H���V���H�E�@<�����H�E�P<���UH��H�� �}�H�u�H�}� t
H�E�H����    H�E��E���H�E���H���+����E���UH��H�� H�}�H�}� t
H�E�H����    H�E�H�E�H���������UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H����~��H�E�H�E�H���  D� H�E�H������H������I��H�E�H�ƿx   ��M��H��L��D��H������H��H��8[A\A]]�UH��H�}�H�E�]�UH��AUATSH��8H�}�H�u�H�U�H�EȾx   H���7~��H�E�H�E�H���  D� H�E�H������H�������I��H�E�H�ƿx   �[M��H��L��D��H���!���H��H��8[A\A]]�UH��H���}��u��}���   �}���  ��   H�=�� ��   �    �    H�=�� �����H��� H�5�� H���G H����L���    �   H�=�� ����H�h� H�5�� H���G H���L���    �   H�=A� �f���H�5� H�5.� H���G H���`L��H�=�� �}���H�� H�5}� H�=t����:L�����UH����  �   �����]ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@ �]�UH��SH��(H�}�H�u�H�E�H��uH��    H��uH�=< ���H�E�H���3  H�E�H�U�H�E�H��H���+  �@��tH��    H��uH�=< �[��H�U�H�E�H��H����  H� H������tH��    H��uH�=.< �!��H�U�H�E�H��H���  H�@H������tH��    H��uH�=K< ����H�E�H�@H��uH�E�H���  H��H�E�H��HH�E�H�XH�U�H�E�H��H���T  H�XH�E�H���t  H��H�E�H�PH�E�H��H���*  H�H�E�H�U�H�PH�U�H�E�H��H���  �@H�U�H�E�H��H���3  H�E�H��([]�UH��H�� H�}�H�u�H�U�H�E�H��H����  �@����tH��    H��uH�=�; ����H�U�H�E�H��H����  H�E��ÐUH��SH��8H�}�H�u�H�E�H��uH��    H��uH�=�; ���H�U�H�E�H��H���=  �@����tH��    H��uH�=�; �j��H�U�H�E�H��H���  H���-  H�E�H�U�H�E�H��H����  H�@H�E�H�E�H��u9H�E�H�PH�E�H9�tH��    H��uH�=�; ����H�E�H�U�H�P�pH�E�H���  H��H�E�H��H���~  H�PH�E�H9�����tH��    H��uH�=�; ���H�]�H�E�H���3  H��H�E�H��H���0  H�XH�}� ueH�E�H� H���  H��H�E�H9�����tH��    H��uH�=�; �=��H�E�H���  H�E�H�E�H����  H��H�E�H��   H�U�H�E�H��H���  H� H���  H��H�E�H9�����tH��    H��uH�=�; ����H�U�H�E�H��H���d  H���  H�E�H�E�H���|  H��H�U�H�E�H��H���6  H�H�E�H���  H��H�E�H9�����tH��    H��uH�=�; �N��H�U�H�E�H��H����  H�     H�U�H�E�H��H����  H�@    H�U�H�E�H��H���  �@ H�E�H��8[]�UH��H�}�H�u�H�E�H�H�E�H� H9�sH�E��H�E�]�UH��H��H�}��u�H�U�H�E�H��H���  H�E���UH��H�� H�}�H�E�H� H���(  H��H�E�H��H���g  H�E��ÐUH��H�� H�}�H�E��    H���C  H�E��ÐUH��H��H�}�H�u�H�U�H�E�H��H���w  ����UH��H��H�}�H�E�H�H�E�H��H���r  H�H�E�H�H�E���UH��H�}�H�E�H� ]ÐUH��H��H�}����E�H�U�H�E�H��H���\  H�E���UH��H��H�}�H�u�H�}� t-H�E�H� H� H�U�H����H�M�H�E��p   H��H���\  ����UH��H�}�H�E�]�UH��H�}�H�E�]ÐUH��H��H�}�H�u�H�E�H���O  H��H�E�H��H���X  ��UH��H�}�H�E�H� ]ÐUH��H�}�H�u�H�E�H�U�H��]�UH��H��0H�}�H�u�H�E�H��� E��H�E؋ H�U�H�M�H�Ή��  H�E�H����E����ÐUH��H�}�H�u�H�E�H�H�E�H� H9���]�UH��H��H�}�H�u�H�E�H���   H��H�E�H��H���   ��UH��H��0H�}�H�u�H�E�H���jD��H�E�� ��H�U�H�M�H�Ή��v   H�E�H���2E����ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���   ���UH��H��H�}�H�E�H���  �ÐUH��H�}�H�u�X   H�E�H�]�UH��H��@�}�H�u�H�U�H�U�H�E�H��H���D��H�U�H�M��E�H�Ή��Y  H�E�H���D�����UH��SH��hH�}�H�u�H�U�H�}� �  H�}� �  vH�U�H�E�H��H���t����  H�E�H�E�H�E�H%  ��H�E�H�E�H�U�H��H���u�������tH��    H��uH�=�? ����H�E��@HH�H��H��H��H�E�H�H��H�E�H�E��@H���q��H�E�H�E�H�@H�U�H)�H�к    H�u�H��H��tH��    H��uH�=�? �j��H�U�H�E�H��H���~��H�E�H�@PH�����E�H�E��@L��uH��    H��uH�=�? �!��H�E�H�ƿ   �#B��H��H���g���H�]�H�E�H�@PH��t%H�E�H�U�H�RPH��H���U�������t�   ��    ��tH��    H��uH�=�? ���H�E�H�PPH�E�H�H�E�H�U�H�PP�}� tIH�E�H�PH�E�H��H���6���H�E�H�@H��tH�E�H�PH�E�H�@H�@H9�sH�E�H�U�H�PH�E�H���}����H��h[]�UH��H�}�H�E�]�UH��H�� �}�H�u�H�U�H�E�� ��u'�u�H�E�A�    A�   �    �   H���Y   �TH�E�� ��t%H�E�� ��tH��    H��uH�=�B ����u�H�E�A�    A�   �    �
   H���   ���UH��H��0H�}�u�U��M�D�E�D�ȈEԃ}� y=�E��؉E��M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ   H���xN��H���3�M�D�E؋}܋U��u�H�E�H��QE��A���Ѻ    H���   H�����UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��+ H�E��E�    �E���~H��    H��uH�=�G ����E���}���Hc�H�E�H���E��H�M�H��T��E���}��E��}� t맀}� t2�E���~H��    H��uH�=�G �4���E��P�U�H��D�-H�U�H�E�H��H���`F��� 9E�����tE�E�    H�U�H�E�H��H���:F��� �U�)�9E�����t�U�H�E���H���N���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���N���E��ڋE����E�}� x!�E�H��D���H�E���H���QN���m��ِ��UH��H��H�}�H����K H�PH�E�H�H�E�H���$�����ÐUH��H��H�}�H�E�H������H�E��x   H���7���ÐUH��H��H�}�H�8o ��   H�5H H�=OH �>F��UH��H�� H�}�H�u�H��    H��u<H�o ��   H�5�G H�=+H �G��dH�%    H�������   ������@H�U�H�E�H��H���f���E��}� tdH�%    H������H�E���������    ��UH��H�� �}�H�u��U�H�M�H�zn ��   H�5FG H�=�G �oE��UH��H�gn ��   H�5#G H�=]G �LE��UH��H��H�}�H�Dn ��   H�5�F H�=2G �!E��UH��H�� H�}�H�u�H�U�H�n ��   H�5�F H�=�F ��D��UH��H��H�}�H�u�H��m ��   H�5�F H�=�F �D�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���#  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L�����UH��H���   H��(���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H���K H� H��0���H��(���H��H���  ��L�����L�����UH��H�}��u�H�U�}���   �E�H��    H��D �H�H��D H���H�E��H�E���]H�E��H�E�f��NH�U�H�E�H��AH�U�H�E�H��4H�U�H�E�H��'H�U�H�E�H��H�E�H�U�H��H�E��H�E����]�UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��j �p  H�5RC H�=�C �{A��UH��H���   H��(���H�� ���H�����H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�����H�� ���H��(���H����  ��L�����L�����UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���  ��L�����L�����UH��H�}�H�E�H� � ]�UH��H�}�H�E��@�PH�E��PH�E�H� H�HH�U�H�
� ]�UH��H��   H�����H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�Hǅ0���    Hǅ8���    H�����H��0���ǅ���   ǅ���0   H�EH�� ���H��P���H��(���H�����H�� ���H��0���H��H���I  ��L�����L�����UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���u3  H�U�H�M�H�E�H��H���9  H�M�H�U�H�u�H�E�H��H���#9  H�E��ÐUH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H������H�E�H��tH�E�H� �U��҉�H���`���H�E�H��t�E���    ��UH��H�� H�}�H�E�H� H�U�H�u�H�Ѻ   H������H�E�H��tH�E�@�PH�E�PH�E�H��t�E���    ��UH��H��@H�}�H�u�H�U�H�}� t
H�E�H����    H�E�H�E�    H�E�    H�E�H�E�H�U�H�M�H�E�H��H���b$  ���UH��H��H�}�H�u�H���K H� H�U�H�M�H��H���8�����UH��H��H�}�H�u�H�Hf ��  H�5�> H�=? ��<��UH��SH��   H�}�H�u�H��x���H��p���H�}� u
�    �   H�M�H��p���H�H�VH�H�QH�FH�AH�E�H�P�H�M�H�E�H��H���3  H�U�H�M�H�E�H��H����=  H�M�H��x���H�u�H�E�H��H����=  H�]�H�E�H��H�E�H�E�H�PH�E�H��H�������H� H��  H�E�H�Ĉ   []�UH��H��`H�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�U�H�E�H��H���1  H�U�H�M�H�E�H��H���%D  H�M�H�U�H�u�H�E�H��H���4D  H�U�H�E�H��  H�E���UH��H�� H�}�H�u�H�U�H��d ��  H�51= H�=k= �Z;��UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�ed ��  H�5�< H�=Z= ��:��UH��H���   H��H���H��@���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��c ��  H�5A< H�=�< �j:��UH��H�� H�}�H�u�H�U�H��c ��  H�5< H�=�< �7:��UH��H�� H�}�H�u�H�U�H��c ��  H�5�; H�=|< �:��UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�Gc ��  H�5c; H�=< �9��UH��H���   H��H���H��@���H��8���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��b ��  H�5�: H�=�; �9��UH��H�� H�}�H�u�H�U�H�M�H��b ��  H�5�: H�=U; ��8��UH��H�� H�}�H�u�H�U�H�M�H��b ��  H�5}: H�=; �8��UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H�!b ��  H�5: H�=�: �.8��UH��H���   H��H���H��X���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�H��a ��  H�5�9 H�=.: �7��UH��H��H�}�H�u�H��a ��  H�5^9 H�=�9 �7��UH��H��H�}�H�u�H�ka ��  H�5/9 H�=�9 �X7��UH��H�� H�}�H�U�H�E�H�Ѻ   �   H���u  H�E�H�}�t�������E�����UH��H��0H�}�H�u�H�U�H�}� uH��` ��  H�5�8 H�=s9 ��6��H�E�    H�E�H��H9E�uH�U�H�E�H��  H�E��oH�E�H���L����E�}��u"H�}� tH�U�H�E�H��  H�E��?�    �8H�U�H�E�HЋU��}�
uH�E�H�PH�E�H��  H�E��
H�E��o�����UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���  H������t�������   ��UH��H���}�H�u�H�U��E�H�։�������UH��H��H�}�H�u�H�E�H���7?��H��H�U�H�E�H�Ѻ   H���  H������t�������   ��UH��H��H�}�H�u�H�U�H�E�H��H��������UH��H��H�}�H�E�H���	  ��UH��H��H�}�H�E�H���������UH��H���K H� H���o	  ]�UH��H���K H� H������]�UH��H�� �}�H�u��E�E�H�U�H�E�H�Ѻ   �   H���?  H������t�������E���UH��H���}�H�u�H�U��E�H�։�������UH��H���}�H���K H��E�H�։��s�����UH��H���}��E����������UH��H��@H�}�H���K H� H��tH���K H� H����    H�E�H�E�    H�E�H���=��H�E�H�E�H;E�sQH�E�H+E�H��H�M�H�E�H�4H�M�H�E�H���E���������t������NH�E�H��u������>H�E�HE��H�U�H�E�H�Ѻ   H�566 H�������������t�������   ��UH��H��H�}�H�l] �f  H�5"5 H�=�5 �K3��UH��H�� H�}��u�H�U�H�A] �g  H�5�4 H�=�5 �3��UH��H���}�H�u�H�] �h  H�5�4 H�=c5 ��2��UH��H��H�}�H�u�H��\ �i  H�5�4 H�=45 �2��UH��H��H�}��u�H��\ �j  H�5e4 H�=5 �2��UH��H��H�}�H��\ �k  H�5:4 H�=�4 �c2��UH��H��\ �l  H�54 H�=�4 �@2��UH��H���}�H�u�H�f\ �m  H�5�3 H�=�4 �2��UH��H���}�H�C\ �n  H�5�3 H�=`4 ��1��UH��H���}�H�u�H�%\ �o  H�5�3 H�=24 �1��UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���*  ��UH��H�� H�}�H�u�H�U�H�M�H�M�H�U�H�u�H�E�H���3  ��UH��H��H�}�H�u�H��[ �z  H�5�2 H�=83 �'1��UH��H��H�}�H�u�H�s[ �  H�5�2 H�=	3 ��0��UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�dH�%    H������� �E�H�}� t-H�E�� ��t"H���K H� H�U�H�53 H�Ǹ    �����E����P�  H��H���K H� H�5�2 H�Ǹ    �~������UH��SH���   H�����H�����H�����H����� t
H����� u"dH�%    H�������   H�������^  H�E�    H�E�    H�����H� H��tH�����H� H�E�H�����H� H�E�H�}� u��  �   H����W��H�E�H�E�   H�����H�M�H�E�H��H���R���H������tH��������   H�E�H����8��H�E�H�U�H�E�H�� 
H�E�H�PH�E�H��  H�� ���H��P�K H��H��� 1��H�� ���H�5�1 H���@1��H��H�E�H�PH�M�H�E�H��H��莱��H�U�H�E�H��H��H������H���V1��H�� ���H����0��H�����H�U�H�H�����H�U�H�H�E�H��H���   []�UH��H�� H�}�H�u��U�H�M�H��X ��  H�50 H�=S0 �B.��UH��H���   H��(���H�� ���H��`���H��h���L��p���L��x�����t )E�)M�)U�)]�)e�)m�)u�)}�ǅ0���   ǅ4���0   H�EH��8���H��P���H��@���H��0���H�� ���H��(���H��H���   ��L�����L�����UH��H��pH�}�H�u�H�U�H�M�H�u�H�H�VH�H�QH�FH�AH�E�H���%  H�U�H�M�H�E�H��H���<  H�M�H�U�H�u�H�E�H��H���<  H�E�H���%  H�U�H�E�H��  H�U�H�E�H�H�E���UH��H��   H��X���H��`���H��P�K H��H����.��H��`���H�5u/ H���/��H���K/��H��`���H����.�����UH��H��   H��X���H��`���H��P�K H��H���.��H��`���H�5J/ H���.��H����.��H��`���H���.�����UH��H��   H��X���H��`���H��P�K H��H���+.��H��`���H�5/ H���K.��H���.��H��`���H���(.�����UH��H�}�H�E��@<    �]�UH��H�}�H�E��@<��]�UH��H�}�H�E��@<��]�UH��H�� H�}�H�U�H�E�H�Ѻ   �   H�������H������t�������E�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H���w���������tHH������H��P�K H��H���,��H������H�5�- H���,��H���-��H������H���,���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H��茶��������tHH��@���H��P�K H��H���+��H��@���H�5�, H����+��H���,��H��@���H���+���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H��  H������H������H��x���H��p���H��p��� tH��p���H����    H�E�H������ t
H��x��� u
�    ��  H��������   H�E�    H�E�H;�x�����   H��x���H+E�H��H������H�E�H�4H������H�E�H���ظ��������tHH������H��P�K H��H���`*��H������H�5�+ H���*��H����*��H������H���]*���H������H��tH������HE��R����H�E��  H�E�    H�E�H;�x�����   H�E�    H�E�H;�������   H������H+E�H��H�E�H������H��H�E�H�H������H�4H������H�E�H������������tHH��@���H��P�K H��H���u)��H��@���H�5�* H���)��H����)��H��@���H���r)���H������H��tH������HE��@����H�E�H;�����sH�E��H�E��	���H��x�����UH��H�� H�}��u�H�U�H�kQ �b  H�5�( H�=�( �&��UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� �����)���������tbH�� ���H��� ��������������t
H�� �����H�����H�����������ܒ����������  H�����H��������H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� �����3�����tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H��P�K H��H���&��H�� ���H�51( H����&��H���'��H�� ���H���&��H�� ����T  H�� ���� <muSH������H��P�K H��H���Q&��H������H�5�' H���q&��H���&��H������H���N&��H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H�<' �H�H�0' H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H�' �H�H�' H����E�
   H�E�    H�����H��������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���[����E�륀}�0uHH�����H���U���H�����H���2����E׀}�xu!H�����H���.���H�����H�������E׀}�/~2�}�9,H�����H������H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H�������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H������H�E�H��H���E׃�AH�H�H�E�H�����H���K����E��;����}�/~S�}�7MH�����H���<���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H��������E�뭐����H�}� ��  H�U؋M�H�E���H���;����  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���\����E��H�}� �/  H�UȋM�H�E���H�������  H�E�    H�����H�������E��}�0uHH�����H������H�����H��������E��}�xu!H�����H�������H�����H��������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H���S���H�E�H��H���E���AH�H�H�E�H�����H�������E��C���H�}� ��  H�U��M�H�E���H���_�����  H�E�H�E�H�����H��������E��E�    �}� t�E���胊����u�   ��    ��tPH�����H������H�}� t�E�Hc�H�E�H��E��H�����H���j����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H�������E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H�������H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H���$��ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H�������E��}� te�E�;E�}]H�����H�������E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H�������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H���s����E��}�0uHH�����H���o���H�����H���L����E��}�xu!H�����H���H���H�����H���%����E��}�/~2�}�9,H�����H������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H�������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H������H�E�H��H���E���AH�H�H�E�H�����H���m����E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E���UH��H��  H�����H�� ���H�������E�    H�� ���� ����  H�� ���� �����j���������tbH�� ���H��� �����I���������t
H�� �����H�����H�����������������������  H�����H���0�����H�� ���� <%uH�� ���H��� <%uKH�� ���� <%uH�� ���H�����H���������_���H�� ���� 8�_�����  ������  H�E�    H�� ���� �����t�����tH�� ���H��� <$u�   ��    ��t
H�� ����gH������� ��/w0H������H�PH������� ��H�H��������JH�������
�H������H�@H�HH������H�JH� H�E�H�� ����E�    H�� ���� <*uH�� ����  H�� ���� <'uSH�� ���H��P�K H��H������H�� ���H�5r H�����H���]��H�� ���H������H�� ����T  H�� ���� <muSH������H��P�K H��H�����H������H�5. H�����H������H������H�����H�� �����
  H�� ���� </~_H�� ���� <9Q�E�    H�� ���� </~<H�� ���� <9.�U��������H�� ���� ����0ЉE�H�� ������E�   �E�
   H�� ���� ����0��J�3  ��H��    H��  �H�H��  H���H�� ���H��� <hu�E�    H�� �����   �E�   H�� �����   �E�   H�� �����   H�� ���H��� <lu�E�   H�� ����   �E�   H�� ����   �E�   H�� ����x�E�   H�� ����g�E�   H�� ����V�E�   H�� ����EH�� ���H��� <xtH�� ���H��� <Xu�E�   H�� �����E�   H�� ����H�� ���� ����X�� ��  ��H��    H��  �H�H��  H����E�
   H�E�    H�����H�������E׃}�
t�}�tj�}��s  ��  �}�/��  �}�9��  H�����H�������H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H���6����E�륀}�0uHH�����H���~���H�����H�������E׀}�xu!H�����H���W���H�����H��������E׀}�/~2�}�9,H�����H���*���H�E�H��H���E׃�0H�H�H�E��v�}�`~2�}�f,H�����H�������H�E�H��H���E׃�aH�H�H�E��>�}�@��   �}�F��   H�����H������H�E�H��H���E׃�AH�H�H�E�H�����H���&����E��;����}�/~S�}�7MH�����H���e���H�U�H��H��H�H�H���E׃�0H�H�H�E�H�����H��������E�뭐����H�}� ��  H�U؋M�H�E���H���|����  H�E�    H�����H�������Eǀ}�/~M�}�7GH�����H�������H�U�H��H��H�H�H���Eǃ�0H�H�H�E�H�����H���7����E��H�}� �/  H�UȋM�H�E���H��������  H�E�    H�����H��������E��}�0uHH�����H���@���H�����H��������E��}�xu!H�����H������H�����H�������E��}�/~2�}�9,H�����H�������H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H���|���H�E�H��H���E���AH�H�H�E�H�����H��������E��C���H�}� ��  H�U��M�H�E���H��������  H�E�H�E�H�����H�������E��E�    �}� t�E�����|����u�   ��    ��tPH�����H�������H�}� t�E�Hc�H�E�H��E��H�����H���E����E��E��}� t��E�;E�}댐H�}� �0  �E�H�H�PH�E�H��  �  H�E�H��x���H�����H��������E��E�    �}� u�E�   �}� ��  �E�;E���  H�����H������H��x��� t�E�Hc�H��x���H��E��H�����H�������E��E��H�� ����E�    H�� ���� <^u�E�   H�� ����M�H������  ��H������ƅ��� H�� ���� <-uH�� ����E��   )Ј�>����(H�� ���� <]uH�� ����E��   )Ј�n���H�� ���� <]��   H�� ���� ��u
�������  H�� ���� <-u\H�� ���� <]tNH�� ���H�� ���H��� �E�H�� ���� 8E�}&�E��   )��E���H�������E����E��ˋE��   )�H�� ���� ����H������H�� ����<���H�E�H��p����E�    H�����H��������E��}� te�E�;E�}]H�����H���;����E���H��������t8H��p��� t�E�Hc�H��p���H��E��H�����H�������E��E�떐H��p��� ��  �E�Hc�H��p���H��  �z  H�E�    H�����H���N����E��}�0uHH�����H������H�����H���'����E��}�xu!H�����H���q���H�����H��� ����E��}�/~2�}�9,H�����H���D���H�E�H��H���E���0H�H�H�E��n�}�`~2�}�f,H�����H������H�E�H��H���E���aH�H�H�E��6�}�@~G�}�FAH�����H�������H�E�H��H���E���AH�H�H�E�H�����H���H����E��C���H�E�H��h���H�U�H��h���H��:H�E�H��`���H��`��� t8H������PH��`�����#����
�������H�}� t�E�������H�� ����m����E��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H��H�}����E�H�E�H�H�E�H�Ѻ   �   H���Z���H�E�H�@H�PH�E�H�P���UH��SH��H�}�H�u�H�E�H�H�E�H���(��H��H�E�H�ٺ   H������H�E�H�����H��H�E�H�@H�H�E�H�P�H��[]ÐUH��H�� H�}�H�u�H�U�H�E�H�H�u�H�E�H�Ѻ   H������H�E�H�PH�E�H�H�E�H�P��ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    �]�UH��H�}����E�H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]�UH��H�}�H�u�H�E�    H�U�H�E�H�� ��t>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�밐]ÐUH��H�}�H�u�H�U�H�E�    H�E�H;E�s>H�U�H�E�H�H�E�H�H�E�H�@H���H�E�H�@H�PH�E�H�PH�E�븐]ÐUH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�PH�E�H�@    �]�UH��H�}����E�H�E�H�PH�E�H�@H9�sH�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P�]ÐUH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���e���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E�H�     H�E�H�@    H�E�H�@    �]�UH��H��0H�}�H�E�H�PH�E�H�@H9���   H�E�   H�E�H�@H�H�E�H�U�H�E�H��H����/��H� H�E�H�E�H��� ��H�E�H�E�H��uH��1 ��   H�5� H�=� ���H�E�H�PH�E�H�H�E�H��H���a��H�E�H� H���O��H�U�H�E�H�H�E�H�U�H�PH�E�H�PH�E�H�@H9�rH�/1 ��   H�5` H�=� �����ÐUH��H��H�}����E�H�E�H�������H�E�H�H�E�H�@H��E�H�E�H�@H�PH�E�H�P���UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t&H�U�H�E�H�� ��H�E��H���k���H�E��Ȑ�ÐUH��H��0H�}�H�u�H�U�H�E�    H�E�H;E�s&H�U�H�E�H�� ��H�E��H������H�E��А�ÐUH��H�}�H�E��@]�UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=
 �	���H��x���� <%uH�E��%   H����  H��x����  H�E�H�������H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�	 菢���H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=�	 �K����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=�	 � ����*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=�	 赡�������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=�	 �j���������E���tH��    H��uH�='
 �B����E���tH��    H��uH�=e
 � ���H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=�
 �⠸�H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=4
 �7���돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=:
 �ퟸ�H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=H
 諟��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H��������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=�	 � ���H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�	 葞���H�U�H�E�H��H���"  H�E�H�U�H��H��H����  H�E�H�������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=�	 ����H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�	 �˝���N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�	 �{���H�U�H�E�H��H�������H��x���� ���M�H�U�H�E�H���<  H�E�H���R���H��x���H�E�H���>����g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�= ����H��x���� <%uH�E��%   H����  H��x����  H�E�H������H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=� 虛���H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=� �U����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=� �
����*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�= 迚�������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=	 �t���������E���tH��    H��uH�=1 �L����E���tH��    H��uH�=o �*���H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=� �외�H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=> �A���돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=D �����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=R 赘��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H��������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=� �
���H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=� 蛗���H�U�H�E�H��H���,  H�E�H�U�H��H��H����  H�E�H�������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=� ����H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=� �Ֆ���N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=� 腖��H�U�H�E�H��H�������H��x���� ���M�H�U�H�E�H���z  H�E�H���\���H��x���H�E�H���H����g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���]  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�="� ����H��x���� <%uH�E��%   H���0  H��x����  H�E�H������H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=�� 裔���H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=� �_����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=	� �����*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=� �ɓ�������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=� �~���������E���tH��    H��uH�=;� �V����E���tH��    H��uH�=y� �4���H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=�� �����H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=H� �K���돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=N� ����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=\� 近��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���	  H�E�H�U�H��H��H����	  H�E�H��������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=� ����H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�� 襐���H�U�H�E�H��H���6	  H�E�H�U�H��H��H����  H�E�H��������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=�� �$���H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�� �ߏ���N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�� 菏��H�U�H�E�H��H�������H��x���� ���M�H�U�H�E�H���  H�E�H���f���H��x���H�E�H���R����g������UH��H�}�H�u�H�U�H�E�H�U�H�H�E�H�U�H�P�]�UH��H��   I��H��L��L��H��H�u�H�}�H��x���H��p���H��x���� ����  H��x���� <%tcH�E�   H��x���H�E�H�� ��tH��x���H�E�H�� <%tH�E���H�U�H��x���H�E�H��H���  H�E�H�x����  H��x���H��x���� ��uH��    H��uH�=,� �'���H��x���� <%uH�E��%   H���n  H��x����  H�E�H������H��x���� <-u6�E�H��x���H��x���� ��u�H��    H��uH�=� 譍���H��x���� <+u9�E�H��x���H��x���� ��u�H��    H��uH�=� �i����u���H��x���� < u=�E�H��x���H��x���� ���I���H��    H��uH�=� �����*���H��x���� <#u=�E�H��x���H��x���� �������H��    H��uH�=� �ӌ�������H��x���� <0u=�E�H��x���H��x���� �������H��    H��uH�=� 舌��������E���tH��    H��uH�=E� �`����E���tH��    H��uH�=�� �>���H��x���� <*ueH��x���H��x���� ��uH��    H��uH�=�� � ���H��p������/wH�P���Hʋ����H�PH�JH�H��E��~�E�    H��x���� </~cH��x���� <9U�U��������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=R� �U���돋E�E�H��x���� <.��  H��x���H��x���� ��uH��    H��uH�=X� ����H��x���� <*��   H��x���H��x���� ��uH��    H��uH�=f� �Ɋ��H��p������/wH�P���Hʋ����H�PH�JH�H��E�H�U�H�E�H��H���  H�E�H�U�H��H��H����  H�E�H��������   �E�    H��x���� </~H��x���� <9~H��    H��uH�=� ����H��x���� </~cH��x���� <9U�U���������H��x���� ����0ЉE�H��x���H��x���� ��u�H��    H��uH�=�� 诉���H�U�H�E�H��H���@  H�E�H�U�H��H��H����  H�E�H��������E�    H��x���� <l��   H��x���H��x���� ��uH��    H��uH�=�� �.���H��x���� <lu9�E�   H��x���H��x���� ��ujH��    H��uH�=�� �鈸��N�E�   �EH��x���� <zu7�E�   H��x���H��x���� ��uH��    H��uH�=�� 虈��H�U�H�E�H��H������H��x���� ���M�H�U�H�E�H����  H�E�H���p���H��x���H�E�H���\����g������UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H��������ÐUH��H��H�}����E�H�E�H� �U��H���0�����ÐUH��SH��H�}�H�u�H�E�H���5���H�E��@H�E�H���c�����H�E�H�ƿ   ������H��[]�UH��H��H�}�H�u�H�U�H�E�H��H����  H�E��ÐUH��SH��H�}�H�u�H�E�H������H�E��@H�E�H��躚���H�E�H�ƿ   �)�����H��[]�UH��SH��(  H��������H��������������������������E��3�	  ��H��    H�� �H�H�� H���H������H�XH������H������H��H������������H������H� ������H������I��H���  H������H���i����  H������H�XH������H�����H��H������������H������H� ������H�����I��H���  H�����H�������  H������H�XH������H��0���H��H���K���������H������H� ������H��0���I��H����#  H��0���H�������L  H�������@��tH� �*   H�5�� H�=�� �����H�������@��tH�� �+   H�5t� H�=z� ����H�������@��tH�� �,   H�5F� H�=_� �o���H�������@��tH�� �-   H�5� H�=G� �B��������� tH�] �.   H�5�� H�=:� ����H������H��H���r�����tH�' �/   H�5�� H�=0� �����H������H�dH�%    H������� ��趎  H��H��������  ������ tH�� �3   H�5`� H�=�� ����H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H��P�K H��H���5���H��P���H�5i� H���U���H����������H��襖��H�5n� H���2���H���|���H��P���H������H�� �;   H�5�� H�=<� �����H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���f�����ÐUH��H��H�}����E�H�E�H� �U��H��������ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H�t �H�H�h H���H������H�XH������H������H��H�������������H������H� ������H������I��H����   H������H���5����  H������H�XH������H�����H��H���x���������H������H� ������H�����I��H���[,  H�����H��������  H������H�XH������H��0���H��H������������H������H� ������H��0���I��H���3  H��0���H���s����L  H�������@��tH�� �*   H�5n� H�=c� ����H�������@��tH�� �+   H�5@� H�=F� �i���H�������@��tH�� �,   H�5� H�=+� �;���H�������@��tH�i �-   H�5�� H�=� ���������� tH�A �.   H�5�� H�=� �����H������H��H���>�����tH� �/   H�5�� H�=�� ����H������H�dH�%    H������� ��肊  H��H���!����  ������ tH��
 �3   H�5,� H�=u� �U���H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H��P�K H��H������H��P���H�55� H���!���H����������H���q���H�5:� H�������H���H���H��P���H�������H��	 �;   H�5P� H�=� �y����H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���������ÐUH��H��H�}����E�H�E�H� �U��H���$�����ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H� �H�H� H���H������H�XH������H������H��H������������H������H� ������H������I��H���0  H������H�������  H������H�XH������H�����H��H���D���������H������H� ������H�����I��H���+<  H�����H�������  H������H�XH������H��0���H��H�������������H������H� ������H��0���I��H���C  H��0���H���?����L  H�������@��tH�� �*   H�5:� H�=/� �c���H�������@��tH�� �+   H�5� H�=� �5���H�������@��tH�r �,   H�5�� H�=�� ����H�������@��tH�E �-   H�5�� H�=�� ����������� tH� �.   H�5�� H�=�� ����H������H��H���
�����tH�� �/   H�5S� H�=�� �|���H������H�dH�%    H������� ���N�  H��H�������  ������ tH�� �3   H�5�� H�=A� �!���H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H��P�K H��H�������H��P���H�5� H�������H����������H���=���H�5� H�������H������H��P���H������H�� �;   H�5� H�=�� �E����H��(  []ÐUH��H�� H�}�H�u�H�U�H�E�H� H�U�H�M�H��H���&�����ÐUH��H��H�}����E�H�E�H� �U��H���\�����ÐUH��SH��(  H��������H��������������������������E��3�	  ��H��    H�� �H�H�� H���H������H�XH������H������H��H���q���������H������H� ������H������I��H���q@  H������H��������  H������H�XH������H�����H��H������������H������H� ������H�����I��H����K  H�����H���l����  H������H�XH������H��0���H��H������������H������H� ������H��0���I��H���OS  H��0���H�������L  H�������@��tH�� �*   H�5� H�=�� �/���H�������@��tH�� �+   H�5�� H�=�� ����H�������@��tH�n �,   H�5�� H�=�� �����H�������@��tH�A �-   H�5}� H�=�� ���������� tH� �.   H�5U� H�=�� �~���H������H��H���������tH�� �/   H�5� H�=�� �H���H������H�dH�%    H������� ����  H��H��������  ������ tH�� �3   H�5�� H�=� �����H������H�@���/wH�P���Hʋ����H�PH�JH�HH�H�E�H������H� H�@��H�E��   H��P���H��P�K H��H������H��P���H�5�� H������H����������H���	���H�5�� H������H�������H��P���H���s���H�� �;   H�5�� H�=�� �����H��(  []�UH��SH��(H�}�H�u�H�E��@��t$H�E��@��tH�U�H�E�H��H���Q  �   H�E��@��tAH�E��@����t2H�E�H��������E�H�E�H���������H�E�H�ƿ   �"�����KH�E��@����t<H�E��@��t0H�E�H�������E�H�E�H��������H�E�H�ƿ   ������H�E�H�PH�E�H��H��H���P  �H��([]ÐUH��H��H�}�H�E��@����tH��    H��uH�=�� �gu��H�E���UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=�� ��t��H��x����@��tH��    H��uH�=�� ��t��H��x����@��tH��    H��uH�=�� �t��H��x����@��tH��    H��uH�=&� �yt��H�E�H�5w� H������H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���dO  �  H��x����@��tH��    H��uH�=�� ��s��H��x����@��tH��    H��uH�=.� �s��H��x����@��tH��    H��uH�=e� �s���}� tH��    H��uH�=�� �ps��H��x���H��H���5�����tH��    H��uH�=�� �?s���E�    H��x����@��9E�}H�E��    H���o����E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H���(����?  H��x����@��tH��    H��uH�=�� �r��H��x����@��tH��    H��uH�=�� �wr���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��� H�E�H�U�H�E�H��H���-L��H�E�H���V���E�H��x���H��H���������t!H��x���H��H���>���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H�������E�뽋E�E�H��x����@9E���  H�E��    H�������E��֋E�E�H��x����@9E�}H�E��    H���V����E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H�������E�뵃}�tH��    H��uH�=Q� �p��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�y� H�E�H�U�H�E�H��H����K  H�E�H���$L  �E�H��x���H��H���������t!H��x���H��H���U���� 9E�~�   ��    ��tH��x���H��H���+���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H�������E�뱋ẺE�H��x����@9E���   H�E��    H�������E��֋ẺE�H��x����@9E�}H�E��    H���]����E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H�������E��H��    H��uH�=�� �n������ÐUH��SH��H�}�H�u�H�E�H� H��H���:�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���M������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���	I  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���a�����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��� �����tH�E�H� H��H���u������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���I  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��������t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���(�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���YG  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H���&���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���P�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����G  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���������t'H�E�H� H��H���O���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���x�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���E  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��������t&H�E�H� H��H���v���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���5F  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H��� �H�H��� H���H�E��@��tH��    H��uH�=�� �i��H�E��@��tH��    H��uH�= � ��h���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=�� �h��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��������t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���?�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���>C  �W  H�E��@��tH��    H��uH�=�� ��f��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���(����}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �ff��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=�� � f��H�E��@��tH��    H��uH�=�� ��e��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �be��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=�� ��d��H�E��@��tH��    H��uH�=+� ��d��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=�� �d��H�E��@��tH��    H��uH�=� ��c��H�E�H��H��躿����tH��    H��uH�=9� ��c���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���c@  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���9>  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����=  �   �}� tH��    H��uH�=#� �Nb��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���>  �H��    H��uH�=� ��a�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5+� H�������H��    H��uH�=� �`a�����UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=|� ��`��H��x����@��tH��    H��uH�=�� ��`��H��x����@��tH��    H��uH�=�� �`��H��x����@��tH��    H��uH�="� �u`��H�E�H�5s� H���n���H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���o=  �  H��x����@��tH��    H��uH�=�� ��_��H��x����@��tH��    H��uH�=*� �_��H��x����@��tH��    H��uH�=a� �_���}� tH��    H��uH�=�� �l_��H��x���H��H���1�����tH��    H��uH�=�� �;_���E�    H��x����@��9E�}H�E��    H���˷���E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H��脷���?  H��x����@��tH��    H��uH�=�� �^��H��x����@��tH��    H��uH�=�� �s^���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��� H�E�H�U�H�E�H��H���)8��H�E�H���B���E�H��x���H��H���Ź����t!H��x���H��H���:���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H�������E�뽋E�E�H��x����@9E���  H�E��    H���޵���E��֋E�E�H��x����@9E�}H�E��    H��貵���E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H���`����E�뵃}�tH��    H��uH�=M� �\��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�u� H�E�H�U�H�E�H��H����7  H�E�H��� 8  �E�H��x���H��H���ܷ����t!H��x���H��H���Q���� 9E�~�   ��    ��tH��x���H��H���'���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H�������E�뱋ẺE�H��x����@9E���   H�E��    H�������E��֋ẺE�H��x����@9E�}H�E��    H��蹳���E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���c����E��H��    H��uH�=�� �Z������ÐUH��SH��H�}�H�u�H�E�H� H��H���6�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���Ե����tH�E�H� H��H���I������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���7  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���]�����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���q������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���37  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��膴����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���$�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���d5  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��譳����t&H�E�H� H��H���"���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���L�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���5  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���ֲ����t'H�E�H� H��H���K���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���t�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���3  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���������t&H�E�H� H��H���r���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��蜱����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����3  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�� �H�H�� H���H�E��@��tH��    H��uH�=�� ��T��H�E��@��tH��    H��uH�=�� ��T���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=�� �T��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��蘯����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���;�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H����0  �W  H�E��@��tH��    H��uH�=�� ��R��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H��脫���}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �bR��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=�� ��Q��H�E��@��tH��    H��uH�=�� ��Q��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �^Q��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=�� ��P��H�E��@��tH��    H��uH�='� ��P��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=�� �P��H�E��@��tH��    H��uH�=� ��O��H�E�H��H��趫����tH��    H��uH�=5� ��O���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���.  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���D,  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����+  �   �}� tH��    H��uH�=� �JN��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���=,  �H��    H��uH�=� ��M�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5'� H��脦���H��    H��uH�=� �\M�����UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=x� ��L��H��x����@��tH��    H��uH�=�� ��L��H��x����@��tH��    H��uH�=� �L��H��x����@��tH��    H��uH�=� �qL��H�E�H�5o� H������H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���+  �  H��x����@��tH��    H��uH�=� ��K��H��x����@��tH��    H��uH�=&� �K��H��x����@��tH��    H��uH�=]� �K���}� tH��    H��uH�=�� �hK��H��x���H��H���-�����tH��    H��uH�=�� �7K���E�    H��x����@��9E�}H�E��    H��艢���E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H���B����?  H��x����@��tH��    H��uH�=�� �J��H��x����@��tH��    H��uH�=�� �oJ���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH��� H�E�H�U�H�E�H��H���%$��H�E�H���.���E�H��x���H��H���������t!H��x���H��H���6���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���̠���E�뽋E�E�H��x����@9E���  H�E��    H��蜠���E��֋E�E�H��x����@9E�}H�E��    H���p����E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H�������E�뵃}�tH��    H��uH�=I� �|H��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�q� H�E�H�U�H�E�H��H����#  H�E�H���$  �E�H��x���H��H���أ����t!H��x���H��H���M���� 9E�~�   ��    ��tH��x���H��H���#���� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���Ӟ���E�뱋ẺE�H��x����@9E���   H�E��    H��裞���E��֋ẺE�H��x����@9E�}H�E��    H���w����E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H���!����E��H��    H��uH�=� �F������ÐUH��SH��H�}�H�u�H�E�H� H��H���2�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���С����tH�E�H� H��H���E������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���$  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���Y�����t&H�E�H� H��H�������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���������tH�E�H� H��H���m������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H����$  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H��肠����t'H�E�H� H��H�������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��� �����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���#  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��詟����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���H�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���!#  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���Ҟ����t'H�E�H� H��H���G���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���p�����tH�E�H� H��H����������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���R!  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���������t&H�E�H� H��H���n���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��蘝����tH�E�H� H��H���������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���q!  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H��� �H�H��� H���H�E��@��tH��    H��uH�=�� ��@��H�E��@��tH��    H��uH�=�� ��@���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=�� ��?��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��蔛����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���7�����tH�E�H��H���������   H�E��PH�u�H�E�A��A�ȉѺ
   H���z  �W  H�E��@��tH��    H��uH�=� ��>��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H���B����}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �^>��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=�� ��=��H�E��@��tH��    H��uH�=�� ��=��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=߷ �Z=��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=� ��<��H�E��@��tH��    H��uH�=#� ��<��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=ŷ �<��H�E��@��tH��    H��uH�=�� ��;��H�E�H��H��貗����tH��    H��uH�=1� �;���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H����  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���p  �   �}� tH��    H��uH�=� �F:��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H����  �H��    H��uH�=	� ��9�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5#� H���,����H��    H��uH�=� �X9�����UH��H��   H�}���H��x����M�L��p����E��E���pt��s�a  ��c�  �u  H��x����@��tH��    H��uH�=t� ��8��H��x����@��tH��    H��uH�=�� �8��H��x����@��tH��    H��uH�=� �8��H��x����@��tH��    H��uH�=� �m8��H�E�H�5k� H��莓��H��p������/wH�P���Hʋ����H�PH�JH�HH�H��H�E�A�    A�   �    �   H���  �  H��x����@��tH��    H��uH�=� ��7��H��x����@��tH��    H��uH�="� �7��H��x����@��tH��    H��uH�=Y� �7���}� tH��    H��uH�=�� �d7��H��x���H��H���)�����tH��    H��uH�=ج �37���E�    H��x����@��9E�}H�E��    H�������E���H��p������/wH�P���Hʋ����H�PH�JH�H���H�E���H��誑���?  H��x����@��tH��    H��uH�=�� �6��H��x����@��tH��    H��uH�=Ь �k6���}� ��  H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�ܬ H�E�H�U�H�E�H��H���!��H�E�H������E�H��x���H��H��轑����t!H��x���H��H���2���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@��tz�E�    �E�;E�};�E�Hc�H�E�H�� ��t'�E�Hc�H�E�H�� ��H�E���H���4����E�뽋E�E�H��x����@9E���  H�E��    H�������E��֋E�E�H��x����@9E�}H�E��    H���؏���E����E�    �E�;E��X  �E�Hc�H�E�H�� ���@  �E�Hc�H�E�H�� ��H�E���H��膏���E�뵃}�tH��    H��uH�=E� �x4��H��p������/wH�P���Hʋ����H�PH�JH�HH�H�E�H�}� uH�m� H�E�H�U�H�E�H��H����  H�E�H���  �E�H��x���H��H���ԏ����t!H��x���H��H���I���� 9E�~�   ��    ��tH��x���H��H������� �E�H��x����@����   �E�    �E�;E�}G�E�H�H��    H�E�HЋ ��t-�E�H�H��    H�E�HЋ ��H�E���H���;����E�뱋ẺE�H��x����@9E���   H�E��    H�������E��֋ẺE�H��x����@9E�}H�E��    H���ߍ���E����E�    �E�;E�}c�E�H�H��    H�E�HЋ ��tI�E�H�H��    H�E�HЋ ��H�E���H��艍���E��H��    H��uH�=ީ �2������ÐUH��SH��H�}�H�u�H�E�H� H��H���.�����t'H�E�H� H��H��裼��� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���̍����tH�E�H� H��H���A������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���P  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���U�����t&H�E�H� H��H���ʻ��� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H���i������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���o  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���~�����t'H�E�H� H��H������� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H��������tH�E�H� H��H��葺�����   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H���  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H��襋����t&H�E�H� H��H������� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H���D�����tH�E�H� H��H��蹹�����   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��H�}�H�u�H�E�H� H��H���Ί����t'H�E�H� H��H���C���� ��uH�}� u�   ��    ��uyH�E�H� �@��t�0   ��    H�E�H� H��H���l�����tH�E�H� H��H���������   H�E�H� �PH�E�H�@H�u�A��A�ȉѺ   H����  �H��[]ÐUH��SH��H�}�u�H�E�H� H��H���������t&H�E�H� H��H���j���� ��u�}� u�   ��    ��uxH�E�H� �@��t�0   ��    H�E�H� H��H��蔉����tH�E�H� H��H���	������   H�E�H� �PH�E�H�@�u�A��A�ȉѺ   H���  �H��[]�UH��SH��hH�}���H�U��M�L�E��E��E���X�� �c  ��H��    H�� �H�H�� H���H�E��@��tH��    H��uH�=�� ��,��H�E��@��tH��    H��uH�=�� ��,���}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E���   �}�u7H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��   �}�u4H�E����/wH�P���Hʋ����H�PH�JH�HH�H�E��S�}� tH��    H��uH�=�� ��+��H�E����/wH�P���Hʋ����H�PH�JH�H�H�H�E�H�E�H��H��萇����t$H�E�H��H������� ��uH�}� u�   ��    ����  H�E��@��t�0   ��    H�E�H��H���3�����tH�E�H��H��諵�����   H�E��PH�u�H�E�A��A�ȉѺ
   H���  �W  H�E��@��tH��    H��uH�=� ��*��H�E�H�E�H�E�H�E�H�E��@��tH�E��0   H��誅���}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=�� �Z*��H�E����/wH�P���Hʋ����H�PH�JH�H�H�EЉ�H�������]  H�E��@��tH��    H��uH�=�� ��)��H�E��@��tH��    H��uH�=� ��)��H�E�H�E�H�E�H�Eȃ}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H�������  �}� tH��    H��uH�=ۣ �V)��H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H���+����Y  H�E��@��tH��    H��uH�=� ��(��H�E��@��tH��    H��uH�=� ��(��H�E�H�E�H�E�H�E��}�uBH�E����/wH�P���Hʋ����H�PH�JH�HH�H�E�H��H���]����  H�E����/wH�P���Hʋ����H�PH�JH�H�H�E���H��������u  H�E��@��tH��    H��uH�=�� �(��H�E��@��tH��    H��uH�=�� ��'��H�E�H��H��讃����tH��    H��uH�=-� �'���}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���=	  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �  �}�ulH�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�pH�2H�E�A��A�   �
   H���  �   �}� tH��    H��uH�=� �B&��H�E��@��t�0   ��    H�E��HH�E����/wH�P�0��H�0���0�H�PH�rH�p�2H�E�A��A�   �
   H���y  �H��    H��uH�=� ��%�����H��h[]�UH��H�� H�}���H�U�M�L�E��E��E��E|"��G~��e��wH�E�H�5� H��褀���H��    H��uH�=	� �T%�����UH��H�� H�}�H�u�H�E�H��������E�H�E�H��������H�E�H�E�H���Ԝ����H�E�����UH��H�}�H�E�� ]�UH��H�� H�}�H�u�H�E�H��������E�H�E�H���������H�E�H�E�H��������H�E�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H����ÐUH��H�}�H�u�H�E�H�U�H�H�E�H�@    H�E�H�@H��    H�E�HЋ ��tH�E�H�@H�PH�E�H�P�͐]ÐUH��H�}�H�E�H�@]�UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H����  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���A  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����	  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���-  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H����
  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���6  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���"  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���+  H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���~  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H����  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H��0H�}�H�u��U܉M�D�E�D�ȈE�H�}� yAH�E�H��H�E��M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ   H���  H���4�M�D�Eԋ}؋U�H�u�H�E�H��QE��A���Ѻ    H���   H�����UH��H�� H�}��u�U��M�D�E�D�ȈE��M�D�E�}�U��u�H�E�H��QE��A���Ѻ    H���s  H�����UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���  H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��� H�E��E�    �E���~H��    H��uH�=Ġ �_���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�� �����E��P�U�H��D�-H�U�H�E�H��H���}��� 9E�����tE�E�    H�U�H�E�H��H����|��� �U�)�9E�����t�U�H�E���H����r���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���r���E��ڋE����E�}� x!�E�H��D���H�E���H���rr���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�
 H�E��E�    �E���~H��    H��uH�=� ����E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�� �E���E��P�U�H��D�-H�U�H�E�H��H���q{��� 9E�����tE�E�    H�U�H�E�H��H���K{��� �U�)�9E�����t�U�H�E���H���1q���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����p���E��ڋE����E�}� x!�E�H��D���H�E���H����p���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�c} H�E��E�    �E���~H��    H��uH�=u� ����M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=[� ����E��P�U�H��D�-H�U�H�E�H��H����y��� 9E�����tE�E�    H�U�H�E�H��H���y��� �U�)�9E�����t�U�H�E���H���o���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���[o���E��ڋE����E�}� x!�E�H��D���H�E���H���+o���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��{ H�E��E�    �E���~H��    H��uH�=՛ �p���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�� �����E��P�U�H��D�-H�U�H�E�H��H���*x��� 9E�����tE�E�    H�U�H�E�H��H���x��� �U�)�9E�����t�U�H�E���H����m���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���m���E��ڋE����E�}� x!�E�H��D���H�E���H���m���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�z H�E��E�    �E���~H��    H��uH�=-� �����E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=� �V���E��P�U�H��D�-H�U�H�E�H��H���v��� 9E�����tE�E�    H�U�H�E�H��H���\v��� �U�)�9E�����t�U�H�E���H���n���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���kn���E��ڋE����E�}� x!�E�H��D���H�E���H���;n���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�sx H�E��E�    �E���~H��    H��uH�=�� � ���E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=c� ����E��P�U�H��D�-H�U�H�E�H��H����t��� 9E�����tE�E�    H�U�H�E�H��H���t��� �U�)�9E�����t�U�H�E���H����l���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����l���E��ڋE����E�}� x!�E�H��D���H�E���H���l���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��v H�E��E�    �E���~H��    H��uH�=ޖ �y���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=Ė ����E��P�U�H��D�-H�U�H�E�H��H���;s��� 9E�����tE�E�    H�U�H�E�H��H���s��� �U�)�9E�����t�U�H�E���H���[k���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���$k���E��ڋE����E�}� x!�E�H��D���H�E���H����j���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�,u H�E��E�    �E���~H��    H��uH�=>� �����E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=� �g���E��P�U�H��D�-H�U�H�E�H��H���q��� 9E�����tE�E�    H�U�H�E�H��H���mq��� �U�)�9E�����t�U�H�E���H���i���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���|i���E��ڋE����E�}� x!�E�H��D���H�E���H���Li���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��s H�E��E�    �E���~H��    H��uH�=�� �1���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=t� ����E��P�U�H��D�-H�U�H�E�H��H����o��� 9E�����tE�E�    H�U�H�E�H��H����o��� �U�)�9E�����t�U�H�E���H����f���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���f���E��ڋE����E�}� x!�E�H��D���H�E���H���ff���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��q H�E��E�    �E���~H��    H��uH�=� ����E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=̑ ����E��P�U�H��D�-H�U�H�E�H��H���Cn��� 9E�����tE�E�    H�U�H�E�H��H���n��� �U�)�9E�����t�U�H�E���H���%e���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����d���E��ڋE����E�}� x!�E�H��D���H�E���H���d���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H�5p H�E��E�    �E���~H��    H��uH�=G� �����M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=-� �x���E��P�U�H��D�-H�U�H�E�H��H���l��� 9E�����tE�E�    H�U�H�E�H��H���~l��� �U�)�9E�����t�U�H�E���H���c���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���Oc���E��ڋE����E�}� x!�E�H��D���H�E���H���c���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��n H�E��E�    �E���~H��    H��uH�=�� �B���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�� ��
���E��P�U�H��D�-H�U�H�E�H��H����j��� 9E�����tE�E�    H�U�H�E�H��H����j��� �U�)�9E�����t�U�H�E���H����a���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���a���E��ڋE����E�}� x!�E�H��D���H�E���H���wa���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��l H�E��E�    �E���~H��    H��uH�=�� �	���E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=݌ �(	���E��P�U�H��D�-H�U�H�E�H��H���Ti��� 9E�����tE�E�    H�U�H�E�H��H���.i��� �U�)�9E�����t�U�H�E���H���c���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���kc���E��ڋE����E�}� x!�E�H��D���H�E���H���;c���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H�Ek H�E��E�    �E���~H��    H��uH�=W� �����E�Hc�H�E�H�H��H��H��H�E�H���E��H�M�H��T��E�Hc�H�E�H�H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=5� ����E��P�U�H��D�-H�U�H�E�H��H���g��� 9E�����tE�E�    H�U�H�E�H��H���g��� �U�)�9E�����t�U�H�E���H����a���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H����a���E��ڋE����E�}� x!�E�H��D���H�E���H���a���m��ِ��UH��H��pH�}��u��M�D�E�D�M��E�U��E�H��i H�E��E�    �E���~H��    H��uH�=�� �K���M��E��    ��Љ�H�E�H���E��H�M�H��T��M��E��    ��E��}� t뜀}� t2�E���~H��    H��uH�=�� �����E��P�U�H��D�-H�U�H�E�H��H���f��� 9E�����tE�E�    H�U�H�E�H��H����e��� �U�)�9E�����t�U�H�E���H���[`���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���$`���E��ڋE����E�}� x!�E�H��D���H�E���H����_���m��ِ��UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��g H�E��E�    �E���~H��    H��uH�=� ����E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=� �9���E��P�U�H��D�-H�U�H�E�H��H���ed��� 9E�����tE�E�    H�U�H�E�H��H���?d��� �U�)�9E�����t�U�H�E���H���^���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���|^���E��ڋE����E�}� x!�E�H��D���H�E���H���L^���m��ِ��UH��H�}�H�u�H�E�H�E�H�E�H�E�H�E�� ��tH�E�H�PH�U��H�E�H�HH�M����H�E��  H�E�]�UH��H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E�H;E�sH�E�H�PH�U��  H�E���H�E�]�UH��H��H�}�H�u�H�E�H���Sm��H��H�E�H�H�E�H��H�������H�E���UH��H��@H�}�H�u�H�U�H�E�H�E�H�E�H�E�H�E�H���m��HE�H�E�    H�E�� ��t.H�E�H;E�s$H�E�H�PH�U��H�E�H�HH�M��H�E���H�E��  H�E���UH��H�}�H�u�H�U�H�E�    H�E�H;E�sIH�U�H�E�H�� �E�H�U�H�E�H�� �E��E�:E�s�������E�:E�v�   �H�E�뭸    ]�UH��H�}�H�u�H�E�    H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H��H�}�H�u�H�U�H�E�H��H���k�����UH��H�}�H�u�H�U�H�E�    H�E�H;E�r�    �\H�U�H�E�H�� �E�H�U�H�E�H�� �E��}� u�}� u�    �'�E�:E�s�������E�:E�v�   �H�E��]�UH��H�� H�}�H�u�H�U�H�� �g   H�5u� H�=�� �na��UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s)H�U�H�E�H�� �U�8�uH�U�H�E�H��H�E��͸    ]�UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E��ă}� uH�U�H�E�H���    ]�UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H���N���H��t�   ��    ��tH�E��H�E����UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t=H�U�H�E�H�� ��H�E���H�������H������tH�U�H�E�H��H�E�뱸    ��UH��H�� H�}�u�H�E�H���7i��H�E�H�E�    H�E�H;E�w8H�E�H+E�H��H�E�H�� ��9E�uH�E�H+E�H��H�E�H��H�E�뾸    ��UH��H�� H�}�H�u�H�E�    H�U�H�E�H�� ��t$H�U�H�E�H�� ��H�E���H������H��u�   ��    ��tH�E��H�E����UH��H�}�H�u�H�E�    H�U�H�E�H�� ����   �E�H�E�    H�U�H�E�H�� ��tGH�U�H�E�H�� ��t-H�U�H�E�H�H�E�H��H�M�H�E�H�� 8�t�E� ��H�E�맀}� tH�U�H�E�H��H�E��h����    ]�UH��H��0H�}�H�u�H�U�H�E�H��uH��� ��   H�5� H�=A� �^��H�}� t
H�E�H�E��#H�E�H� H��tH�E�H� H�E��
�    �   H�E�� ��t$H�E�� ��H�E���H������H��t�   ��    ��tH�E���H�E�H�E�H�E�� ��t$H�E�� ��H�E���H���R���H��u�   ��    ��tH�E���H�E�� ��tH�E��  H�E�H�U�H��H��H�E�H�     H�E���UH��H��H�}�H�u�H�M�H�E�H��� H��H��������UH��H�}�u�H�E�    H�U�H�E�H�� ��t*H�U�H�E�H�� ��9E�uH�U�H�E�H��H�E���H�U�H�E�H�]�UH��H��H�}�H�u�H�� ��   H�5g� H�=�� �`\��UH��H��H�}�H�u�H�� ��   H�58� H�=q� �1\��UH��H��H�}�H�u�H�͏ ��   H�5	� H�=B� �\��UH��H�� H�}�H�u��U�H��� ��   H�5׋ H�=� ��[��UH��H�� H�}�H�u��U�H�y� ��   H�5�� H�=ދ �[��UH��H�� H�}�H�u��U�H�O� ��   H�5s� H�=�� �l[��UH��H�� H�}�H�u��U�H�%� ��   H�5A� H�=z� �:[��UH��H��H�}�H�u�H��� ��   H�5� H�=K� �[��UH��H�� H�}�H�u�H�U�H�ӎ ��   H�5ߊ H�=� ��Z��UH��H�� H�}�H�u�H�U�H��� ��   H�5�� H�=� �Z��UH��H�� H�}�H�u�H�U�H�}� ��   H�5y� H�=�� �rZ��UH��H��H�}�H�u�H�W� ��   H�5J� H�=�� �CZ��UH��H�� H�}�H�u�H�U�H�+� ��   H�5� H�=P� �Z��UH��H��H�}�H�u�H�� ��   H�5� H�=!� ��Y��UH��H��H�}�H�u�H�ݍ ��   H�5�� H�=� �Y��UH��H�� H�}�H�u�H�U�H��� ��   H�5�� H�=�� �Y��UH��H�� H�}�H�u�H�U�H��� ��   H�5S� H�=�� �LY��UH��H�� H�}�H�u�H�U�H�\� ��   H�5 � H�=Y� �Y��UH��H��H�}��u�H�6� ��   H�5� H�=+� ��X��UH��H��H�}�H�u�H�� ��   H�5È H�=�� �X��UH��H��H�}�H�u�H�� ��   H�5�� H�=͈ �X��UH��H��H�}��u�H� ��   H�5f� H�=�� �_X��UH��H��H�}�H�u�H��� ��   H�57� H�=p� �0X��UH��H��H�}�H�u�H�s� ��   H�5� H�=A� �X��UH��H�� H�}�H�u�H�U�H�G� ��   H�5Շ H�=� ��W��UH��H�}�u�H�U�H�E�H�E�H�E�    H�E�H;E�s6H�E�H��    H�E�HЋ 9E�uH�E�H��    H�E�H��H�E����    ]�UH��H��H�}�H��� �  H�5D� H�=}� �=W��UH��H�� H�}��u�H�U�H��� �  H�5� H�=K� �W��UH��}�E�-�  ��C�  ��H��    H�a� �H�H�U� H���H�-� H�E���   H�<� H�E���   H�D� H�E���   H�P� H�E���   H�]� H�E��   H�g� H�E��   H�u� H�E��   H�� H�E��   H��� H�E��sH��� H�E��fH��� H�E��YH��� H�E��LH�� H�E��?H��� H�E��2H�� H�E��%H�� H�E��H�%� H�E��H�:� H�E�H�E�]�UH��H��0�}�H�u�H�U؋E������H�E�H�U�H�M�H�E�H��H������H�E�H���_��H9E�����t�   ��    ��UH��H�� H�}�H�u�H�U�H�U�H�M�H�E�H��H����]��H��H�E�H���UH��H�� H�}�H�u�H�E�H���^��H�E�H�E�H�PH�M�H�E�H��H���z]��H�U�H�E�H���UH��H��0�}�H�u�H�U�H�M�H�u�H�U��E�H�H�M�A�    I��H�ƿ   �AI���E�Hc�H�E�H�H�E�H� H���u�������    ��UH��H��0�}�H�u�H�U�H�M�H�u�H�U��E�H�H�M�A�    I��H�ƿ   ��H���E����u�������E�Hc�H�E�H��    ��UH��H��0�}�H�u��U�H�M�H�u��E�Hc�H�U��E�H�A�    I��H�ƿ   �yH��H�E�H�E�H�}��u������H�E�H�U�H��    ��UH��H��0H�}�u�H�U�H�U�H�E�A�    A�    �    H�ƿ   �H��H�}� u�������U�H�E؉�    ��UH��H���}��E�H�A�    A�    �    �    H�ƿ   ��G���    ��UH��H�� H�}�u�H�U��M�H�E��H���K����E���t�E��������    ��   ��UH��H����� ������t-H�=�� �  ������tH�=�� �u  H�=�� �1  �|� ������t<H�=l� ��  ������t'H�=o� �d  H��H�=�� �q  H�=<� ��  �@� ������tDH�=0� �  ������t/H�=C� �  H�E�H�E�H��H�=�� �  H�=�� �  H�=�� ��  �ÐUH��H�� H�}�H�u�H�U�H�E�H��H����F��������tH�І �   H�5=� H�=f� �Q��H�E��ÐUH��H�� H�}�H�u�H�U�H�E�H�U�H��H���G��������tH�~� �!   H�5� H�=8� �XQ�����UH��H�}�H�E��     �]ÐUH��H��H�}�H�E�H����   H�E�H�ƿ   �H�����UH��H�}�H�E�]�UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H���   H�E�H�������H��H�E�H�ƿ�  �`H��H��H���   �H��[]�UH��H�}�H�E�]�UH��H�}�H�E�]�UH��SH��H�}�H�u�H�E�H����   H�E�H�������H�H�E�H�ƿ   ��G��H��H����   �H��[]�UH��H�}�H�E�]�UH��H�}�H�E��  �]�UH��H�}�H�E�H�Ƹ    �9   H��H���H��]ÐUH��ATSH��H�}�H�u�H�E�H�U�H�H�E�H��H���r���H�E�H��H���n   H�E�H�@     H�E�H��(�   I��H��xL���i   I�� H����H��[A\]ÐUH��H�}�H�E�H�     �]�UH��H�}�H�u�H�E�H�U�H��]�UH��H��H�}�H�E�H���N   H�}�:   ���UH��H��H�}�H�E�H������H�E�H�@    H�E�H��H���$   ���UH��H�}�]ÐUH��H�}�H�E�H�     �]�UH��H��H�}�H�E�H���   H�}�������UH��H�}�H�E�H�     �]�UH��H�}�H��p�K H�PH�E�H��]ÐUH��H��H�}�H�E�H�������H�E��   H����>����UH���B� ������tJH�=2� �i  ������t5H�=� ��  H�=� �  H�U� H�5�� H��tH H���E��H��� ]�UH��H�}��u�H�U�U�H�E��    ]�UH��H��� ]�UH��H�}����E�ЈE�H��p�K H�PH�E�H�H�E��U�PH�E��U��P	�]ÐUH��H�}�H�E��     H�E��@    �]�UH��H�}�H�E�� ]�UH��H�}�H�E��@]ÐUH��H�� H�}�H�u�H�E�H� � �E�H�E� ����   �E���x�U�H�E�P�-  �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    ��   �E�%�   =�   u�E�����H�E�PH�E��    �   �E�%�   =�   t/�E�%�   =�   tH�ӂ �'   H�5o� H�=�� �(L���   �q�E�%�   =�   tH��� �,   H�59� H�=�� ��K��H�E�@�����E���?	�H�E�PH�E� �P�H�E�H�E�H� H�PH�E�H��    �ÐUH��H��0H�}�H�u�H�U�H�E�H� � �E��}�vH�ہ �>   H�5�� H�=H� �hK��H�E�H� �U��H�E�H� H�PH�E�H�H�E�H� H�PH�E�H��    ��UH��H��H�}�H�E��    �   H���X���H��0�K H�PH�E�H���ÐUH��H��H�}�H��0�K H�PH�E�H�H�E�H���<�����ÐUH��H��H�}�H�E�H������H�E��   H���E;���ÐUH��SH��XH�}�H�u�H�U�H�M�H�E�� f��tH�(� �W   H�5� H�={� �[J��H�E�H�PH� H�E�H�U�H�E�H�������H�E�H���  ��tH�E�H���  ��t�   ��    ����   H�U�H�E�H��H�������E�}� t�E��   H�E�H������������t�H�U�H�E�H�H�E�H���o���������t�    �MH�E�H�H�E�H���L����H�E�H� H�PH�E�H��@���H�E�H������������t�   ��    H��X[]ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH�� �s   H�5W~ H�=0 �I��H�E�H�PH� H�E�H�U�H�E�H���x���H�E�H���F  ��tH�E�H���v  ��t�   ��    ����   H�U�H�E�H��H���s����E��}� t�E��   H�E�H���4���������t�H�U�H�E�H�H�E�H���$���������t�    �OH�E�H��������H�E�H� �H�E�H� H�PH�E�H��>���H�E�H�������������t�   ��    �ÐUH��H��PH�}�H�u�H�U�H�M�H�E�� f��tH�S~ ��   H�5} H�=�} ��G��H�E�H�PH� H�E�H�U�H�E�H���0���H�E�H�     H�E�H����  ��ttH�U�H�E�H��H���D����E��}� t�E��tH�E�H������������t�H�U�H�E�H�H�E�H�������������t�    �8H�E�H� H�PH�E�H��|���H�E�H������������t�   ��    ��UH��H��`H�}�H�u�H�U�H�M�H�E�� f��tH�} ��   H�5�{ H�=�| �F��H�E�H�PH� H�E�H�U�H�E�H���V  ��tH�E�H���f  ��t�   ��    ����   H�E�H� � �E؋E؅�u
�    �   H�E�H�E�H�E�H��H�E�H�U�H�M�H�E�H��H���x����E��}�tY�}� t�E��pH�U�H�E�H9�tH�@| ��   H�5,{ H�=| ��E��H�E�H� H�PH�E�H�H�U�H�E�H��"��������H�U�H�E�H� H9�t�   ��    ��UH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}�H�E�H�H�E�H�@H9���]ÐUH��H�}��   ]ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t2��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H��P�K H��H���pF��H��`���H�5${ H���F��H����F��H��`���H���mF���    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t ��T���/v��T���9w�   �[�    �T��T���vFH��`���H��P�K H��H���E��H��`���H�5�z H����E��H��� F��H��`���H���E���    ��UH��H��   H��X�����T�����T���wH��X���H���:�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���fv��T���@v��T���Fw�   �[�    �T��T���vFH��`���H��P�K H��H����D��H��`���H�5,z H����D��H���BE��H��`���H����D���    ��UH��H��   H��X�����T�����T���wH��X���H���\�����t�   ��    ��tD��T���/v	��T���9v$��T���`v	��T���zv��T���@v��T���Zw�   �[�    �T��T���vFH��`���H��P�K H��H����C��H��`���H�5�y H���D��H���dD��H��`���H����C���    ��UH��H��   H��X�����T�����T���wH��X���H���~�����t�   ��    ���r  ��T���!�W  ��T���"�J  ��T���#�=  ��T���$�0  ��T���%�#  ��T���&�  ��T���'�	  ��T���(��   ��T���)��   ��T���*��   ��T���+��   ��T���,��   ��T���-��   ��T���.��   ��T���/��   ��T���:��   ��T���;��   ��T���<t~��T���=tu��T���>tl��T���?tc��T���@tZ��T���[tQ��T���\tH��T���]t?��T���^t6��T���_t-��T���`t$��T���{t��T���|t��T���}t	��T���~u�   �[�    �T��T���vFH��`���H��P�K H��H����A��H��`���H�5�w H���
B��H���TB��H��`���H����A���    ��UH��H��   H��X�����T�����T���wH��X���H���n�����t�   ��    ��t ��T��� v��T���~w�   �[�    �T��T���vFH��`���H��P�K H��H���0A��H��`���H�5tw H���PA��H���A��H��`���H���-A���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T��� t	��T���	u�   �n�    �g��T���vYH��`���H��P�K H��H���v@��H��`���H�5
w H���@��H��T�����H���@��H����@��H��`���H���`@���    �ÐUH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��tD��T��� t-��T���	t$��T���
t��T���t��T���t	��T���u�   �[�    �T��T���vFH��`���H��P�K H��H���?��H��`���H�5hv H���?��H����?��H��`���H���?���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���v��T���~w�   �[�    �T��T���vFH��`���H��P�K H��H����>��H��`���H�5�u H����>��H���4?��H��`���H����>���    ��UH��H��   H��X�����T�����T���wH��X���H���N�����t�   ��    ��t ��T���`v��T���zw�   �[�    �T��T���vFH��`���H��P�K H��H���>��H��`���H�5Du H���0>��H���z>��H��`���H���>���    ��UH��H��   H��X�����T�����T���wH��X���H��������t�   ��    ��t ��T���@v��T���Zw�   �[�    �T��T���vFH��`���H��P�K H��H���V=��H��`���H�5�t H���v=��H����=��H��`���H���S=���    ��UH��H��   H��X�����T�����T���wH��X���H���������t�   ��    ��t��T���@v��T���Zw��T����� �U��T���vFH��`���H��P�K H��H���<��H��`���H�5#t H���<��H���	=��H��`���H���<����T�����UH��H��   H��X�����T�����T���wH��X���H���"�����t�   ��    ��t��T���`v��T���zw��T����� �U��T���vFH��`���H��P�K H��H����;��H��`���H�5�s H���<��H���Q<��H��`���H����;����T�����UH��H��� ]ÐUH��H�� H�}��E�    H�E�H�pH�U���   ��������u�
��uH�=�u ��.�����UH��H�}�H�E�H���    ��]�UH��H��   H��`���H��Q�K H��H���b2��H��`���H�5pu H���2��H��H�EH��H���   H���2��H��`���H���M2�����UH��H�� H�}�H�E�H�E�H�E�H������H�E�� ������tH�E�H���D����    ��   ��UH��H��H�}�H�E�H�E�H�E��   �H�E�H���������UH��H��H�}�H�u�H�U�H�E�H��H���   H�E���UH��H��0H�}�H�u�H�E�H���/��H�E�H� H�U�H�M�H��H���   H�E�H���0�����UH��H��`H�}�H�u�H�U�H�E�H�5dt H���53��H�E�H���a/��H�E�H�M�   H��H���_V��H�E�H�U�H�M�H��H���   H�E�H���0��H�E�H���
0�����UH��H�� H�}�H�u�H�U�H�E�� ��u(H�u�H�E�A�    A�   �    �   H���Z   �UH�E�� ��t%H�E�� ��tH��    H��uH�=�s �{շ�H�u�H�E�A�    A�   �    �
   H���   ���UH��H�� H�}�H�u��U�M�D�E�D�ȈE��M�D�E�}�U�H�u�H�E�H��QE��A���Ѻ    H���   H�����UH��H�ĀH�}�H�u��M�D�E�D�M��E�U��E�H��r H�E��E�    �E���~H��    H��uH�=�s �Է��E�Hc�H�E��    H��H�E�H���E��H�M�H��T��E�Hc�H�E��    H��H�E�H�}� t딀}� t2�E���~H��    H��uH�=�s �1Է��E��P�U�H��D�-H�U�H�E�H��H���]4��� 9E�����tE�E�    H�U�H�E�H��H���74��� �U�)�9E�����t�U�H�E���H���;4���E��U��E�9�}-�E�    �U��E�)�9E�}H�E��0   H���4���E��ڋE����E�}� x!�E�H��D���H�E���H����3���m��ِ�� H�a� H���t3UH��S��K H��D  ��H��H�H���u�H��[]�f.�     ������         r close.bmp /shell.lef /dev/mouse0 Error initializing freetype /montserrat.ttf  Error loading font from memory /montserrat.ttf FREETYPE_PROPERTIES              �@H     `OH     `dH      iH     �uH     @{H     �|H     ��H     ��H     ��H      �H     ��H      �H      �H     ��H      �H     `I     @I             properties kerning glyph-dict postscript-font-name sfnt-table tt-cmaps type42 truetype truetype-engine darkening-parameters hinting-engine adobe no-stem-darkening random-seed .resource/ resource.frk/ .AppleDouble/ % ._ cff type1    �B@     �B@     �B@      A@     0B@     �@     [�@     [�@     [�@      �@      �@     [�@     [�@     ��@     ��@     ��@     ��@     ��@     ��@     ��@     ��@     p�@     p�@     �@     �@     ��@     ��@             ��     G	           ��     8�     *�      �r      L9      �      S      )      �      �      �       s       9                                                                 ��@             P�@            ��@            P�@            ��@            p�@             �@            �@            P�@            /..namedfork/rsrfont-format interpreter-version Weight OpticalSize Slant sfnt .notdef TrueType multi-masters metrics-variations tt-glyf          ~A     �zA     ~A      ~A     0~A     @~A     P~A     �}A     $�A     $�A     $�A     $�A     $�A     $�A     �A     �A     �A     �A     ��A     w�A     X�A     /�A     �A     �A     !�A     �A     ��A     t�A     �A     ��A     �A     ؋A     ��A     ��A     ��A     �A     �A     c|A     ��A     ��A     �A     �{A     ��A     ۂA     A     �{A     �A     ٘A     `~A     Z�A     ΍A     x�A     ��A     =�A     ĄA     ĄA     ��A     ��A     l�A     l�A     ��A     ��A     TA     TA     g�A     V�A     ��A     ��A     ��A     ��A     ��A     ��A     #�A     *�A     ~�A     I�A     ��A     ��A     m�A     m�A     D�A     ڛA     ڛA     ԒA     ��A     ��A     ��A     x�A     U�A     2�A     �A     ܑA     ��A     {�A     Q�A     ,�A     וA     �{A     ��A     ~�A     t�A     @A     @�A     %�A     �A     �A     ԔA     ��A     ��A     {�A     4�A     �A     �A     �A     �A     �A     њA     њA     њA     њA     t�A     @A     @A     ��A     ��A     ��A     řA     K�A     ;�A     �A      �A     `~A     ��A     u�A     �{A     �{A     >�A     ߗA     ��A     `~A     `~A     �A     ��A     ��A     ��A     ��A     J�A     Q�A     ƘA     h�A     ��A     `~A     `~A     ��A     ��A                  
                                               "             
                                    X�    �      �;#(    ć      �D�    �      X�    �      �;#(    ć      �D�    �      ���    P      d    ��      c���    X      ���    P      �VY�    ��      �r�    E       N�b    P      d]j�    @y      )�Px    �      
�-    P      �2=    ��      ;�?�    �      &�_    P      �ɬ�    �~      ����          ���    P      ;�0Z    c�      &�    ~       ���    P      ��    ��      &�    ~       F��          �|�@    *�      �t�`    z       8��          ����    og      ��    �      ����           �H��    ��      p           ����           �Z
    9|     p                           U%�@    �       �X��    |                      R�3    �       *��&    j                      e�m    �      Knl    �$                      U%�@    �       ��Q�    |                      dv�    �       1(Ʀ    �                      ��-    �      3F`�    �                      Lw�@    �      ��\�    �                      ��=    A      fw�    �"                      �&iJ    �      FC4    �                      �4�    f      F�l    �"                      S�]    �      _Zt@    �"                      H�U�    �      �� 9                `       n0��    �X      *HC�    5       cpop                DFGirl-W6-WIN-BF    DFGothic-EB         DFGyoSho-Lt         DFHSGothic-W5       DFHSMincho-W3       DFHSMincho-W7       DFKaiSho-SB         DFKaiShu            DFKai-SB            DLC                 DLCHayMedium        DLCHayBold          DLCKaiMedium        DLCLiShu            DLCRoundBold        HuaTianKaiTi?       HuaTianSongTi?      Ming(for ISO10646)  MingLiU             MingMedium          PMingLiU            MingLi43                                ��		             P    "                    !!  !!!!!! !!!!!!              3!!                                                                        @   @   @               @             D                       	                         �       �.H                           ��@     ��@     pwA     p             0      �lA      A     `�@     P�@     A             @�A     ��@             �A     @JA     ��@     `1H     �1H     �1H      BH     �1H     �AH     �.H     �AH     �1H     �AH     8.H     PBH                     ��@            `kA                     PkA                             pkA                     �fA     peA      MA     �`A     `dA     `cA     �A     P�@     �wA     @A     pshinter StandardEncoding ExpertEncoding ISOLatin1Encoding eexec closefile FontDirectory CharStrings dup put %!PS-AdobeFont %!FontType postscript-cmaps psaux Regular Black Notice FullName FamilyName ItalicAngle isFixedPitch UnderlinePosition UnderlineThickness UniqueID lenIV LanguageGroup password BlueScale BlueShift BlueFuzz BlueValues FamilyBlues FamilyOtherBlues StdHW StdVW MinFeature StemSnapH StemSnapV ExpansionFactor ForceBold PaintType StrokeWidth FontBBox NDV CDV DesignVector FontMatrix Subrs Private BlendDesignPositions BlendDesignMap BlendAxisTypes WeightVector postscript-info               q�A     q�A     ��A     ��A     �A     ��A     ��A     ��A     <�A     �A     `�A     ��A     ��A     ��A     `�A     8�A     �A     ��A     ��A     8�A     �A     ��A     `�A     0�A     �A     ��A     ��A     ��A     ��A     ��A     8�A     ��A     ��A     ��A     X�A     0�A     �A     ��A     H�A     �A     ��A     ��A     ��A     P�A      �A     �A      �A     ��A     ��A     ��A     p�A     @�A     �A     ��A     8�A             x1H                                         CH                                        CH                                        CH                                        �1H                                         'CH                   (                     3CH                   0                     @CH                   2                     RCH                   4                     qQH                                         eCH                                         nCH                                        tCH                   �                     �CH                   �                     �CH                   p                     �CH                   x                     �CH                   |                     �CH        	                              �CH        	           (      
   	          �CH        	           <         
          �CH        	           X      
             �CH        	           �                    �CH        	           �                    �CH        	           �                    �CH        	           �         �          �CH        	           �         �          �CH                   �                     DH                   �                     �gH                                        DH                   �                    �BH                   �                    DH                                       +DH                                         4DH                   X                    8DH                   \                    <DH        	           �        �         IDH           ��A                            �BH           ��A                            TDH           ��A                            �BH           ��A                            ZDH           0�A                            bDH           ��A                            wDH           @�A                            �DH           ��A                            �DH           p�A                            �hH           �A                                                                                                  h       /H                           ��A     p�A     ��A     x      X       P      �B     p�A     pB     �B     ��A     ��A     ��A      �A     �B     `�A      B             V.H     PQH     K.H     `QH     `1H     /hH     �DH     �PH     8.H     �PH     C.H     �PH     �1H      QH                     �s@     Pv@     ��A             ��A     ��A     ��A     ��A     ��A                             ��A     pB     �B     ��A     `B      B     � B     �B             ��A     p�A             ��A     ��A     /FSType cff-load CFF CID                        WB     -WB     �VB     �VB     -WB     -WB       ( ) *                                                                                                  � �   � � � � � � � �    c � � � � � � � � � �   � � � �   � � �                	  
m n    !"#$%&'()*+,-./                                                                    012    34567  8    8    :;    <=>      � � � ?@ABCDE    F� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                                                                        	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _                                                                     ` a b c d e f g h i j k l m n   o p q r   s t u v w x y z   {   | } ~  � � � �   � �   � � � �                                 �   �         � � � �           �       �     � � � �            � � � � � �    c � � � � � � � � � �   � � � � � �  	
m n ,-.1:;� � � @ABCDEF� � � GHIJKLMNOPQRSTUVWXYZ                     � � � � � � � � � �    c � � � � � � � � � �   � � � � � � �  	
m n  !"#$%&'()*+,-./0123456789:;<=>� � � ?@ABCDEF� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                              	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _ ` a b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                                                                                        (                           0                           8                           <                                   �`B                  �                                   TB                  �                           �                           �                           �                                   �\B                  �                           �                                   @\B                          �[B                  �                                                     !                          "                          #                          $                           %  (                        &  0                                                      x              
            �                       	   8             
         	!  �                        
!  �                        !  �                        
   �                           �                        !  �                �     !                   �     !  �                        !  �                        !  �                        !  �                        !  �                        !  �                           �                           �                           �                        1          �`B                0  �                         $1                           %1  (                        0  8                        0          �[B                @          �\B                A          �`B                P                          P  x              
         P  �                       	P  8             
         	Q  �                        
Q  �                        Q  �                        
P  �                        P  �                        Q  �                �     Q                   �     Q  �                        Q  �                        P          @[B                P          @]B                P  �                                                     ���������������G�z�G�S㥛�  e�c]�F ��#��S  �Z�{c  �Ք��   0�y   }�%                          
       d       �      '      ��     @B     ���      ��     ʚ;                          h       /H                           `#B     �#B      dB     p      `       H       iB     �PB     �<B     �:B     �$B     P#B     0NB     � B             �NB     @;B     �9B     `1H     �QH     �1H     `fH     �1H      fH     �DH      gH     V.H     �fH     K.H     0gH     v.H     �fH     �QH     �fH     8.H     �fH     xQH     �eH                                      "B     �XB     @"B      .B     `.B                              "B                                                     "B                     �!B     �!B     �!B     �!B     �!B     �!B      #B     0#B     �s@     Pv@     `6B      !B     P!B     0'B     �'B                             7B     @8B     !B                             `dB      ,B     (       @ B     �#B     � B     � B                                                                     �B     �B     �B       B                                             CIDFontName StartData /sfnts (Hex) %ADOBeginFontDict t1cid CID Type 1 CIDFontVersion CIDFontType Registry Ordering Supplement UIDBase CIDMapOffset FDBytes GDBytes CIDCount SubrMapOffset SDBytes SubrCount lenBuildCharArray ForceBoldThreshold FDArray        %!PS-Adobe-3.0 Resource-CIDFont                       h       %hH                           ЏB     P�B     �B     x      `       H      @�B     ��B     ��B      �B      �B     ��B     @�B                             `�B             `1H     +hH     V.H     �jH     �DH     �jH     �QH     PjH     8.H     @jH                     �s@     Pv@     АB      �B     �B                             ��B     ��B                             `�B                     �gH                                           6hH                                          EhH                                          QhH                                          ZhH                                           chH                    (                      nhH                    �                      vhH                                         �hH                                          �hH                    $                     �hH                    (                     x1H                                          CH                                         CH                                         CH                                         �1H                                          'CH                   (                      3CH                   0                      @CH                   2                      RCH                   4                      qQH                                          DH                                         �BH                                        �hH                   @                     �hH                   H                     �hH                   8                     �hH                   �                      �hH                   �                      DH                   �                      eCH                                          nCH                                         tCH                   �                      �CH                   �                      �CH                   p                      �CH                   x                      �CH                   |                      �CH        	                               �CH        	           (      
   	           �CH        	           <         
           �CH        	           X      
              �CH        	           �                     �CH        	           �                     �CH        	           �                     �CH        	           �         �           �CH        	           �         �           DH                   �                      +DH                                          �hH            �B                             IDH           ��B                             �CH           p�B                                                                                             8�B     �B     ��B     ]�B     �B     �B     ��B     N�B     ��B     ��B     ��B     ��B     �B     �B                             �B            P�B             �B            ��B                                      :            $ ( , 0 4 8 < @ D H L P T X \ ` d h                       8       0wH                                           ��B     �      X       h      0�B     ��B                     0�B     ��B     `�B      �B                                     4wH     �vH     `1H     @wH                     пB     �B     ��B                             (        �B     ��B     ��B      �B                                             pfr pfr-metrics PFR %!PS-TrueTypeFont known Type 42                             x1H                                          CH                                         CH                                         CH                                         �1H                                          'CH                   (                      3CH                   0                      @CH                   2                      RCH                   4                      qQH                                          �gH                                         DH                   �                     �BH                   �                     DH                                        +DH                                          IDH           ��B                             �BH           ��B                             �BH           P�B                             hH           ��B                                                                                   @       .H                           �B     ��B     ��B     �      `       8      �C     0�B     ��B     PC     ��B     ��B     0�B                              �B     ��B     K.H     �|H     V.H     �|H     �DH     `|H     `1H     \wH                                     ��B     ��B     ��B     ��B             ��B      �B     @�B     Bold Italic winfonts Windows FNT                                      8       �|H                                           �C           X       0      @C     �C                                     �C                             �C     �C     `1H     �|H     �|H     �}H                     �C                     �C             �C     �C                                                              �    < L N P R T V X Z [ \ ^ ` b d f h j l m n o p x � � � � � � � � � �                                                                       (               �    
       n    h                   (   "                 @   :       Oblique SLANT WEIGHT_NAME SETWIDTH_NAME ADD_STYLE_NAME FAMILY_NAME RESOLUTION_X RESOLUTION_Y CHARSET_REGISTRY CHARSET_ENCODING 10646 8859 646.1991 IRV pcf bdf PCF                                                                         	                      	                                             
             
                                                       @       k�H                           �!C     �!C     0'C     P      X       0      BC     �(C                                     @#C                             @"C     �!C     o�H     ��H     `1H     s�H     8.H     ��H                     �!C     �!C     �!C     p)C     (         C       C     @ C     � C                                             COMMENT DEFAULT_CHAR FONT_ASCENT FONT_DESCENT SPACING ENDPROPERTIES %hd _XFREE86_GLYPH_RANGES  + STARTFONT STARTPROPERTIES FONTBOUNDINGBOX - CHARS ENDFONT ENDCHAR STARTCHAR SWIDTH DWIDTH BBX BITMAP BDF CHARSET_COLLECTIONS COPYRIGHT DESTINATION DEVICE_FONT_NAME FACE_NAME FONTNAME_REGISTRY FOUNDRY FULL_NAME ITALIC_ANGLE NOTICE RAW_ASCENT RAW_AVERAGE_WIDTH RAW_AVG_CAPITAL_WIDTH RAW_AVG_LOWERCASE_WIDTH RAW_CAP_HEIGHT RAW_DESCENT RAW_END_SPACE RAW_FIGURE_WIDTH RAW_MAX_SPACE RAW_MIN_SPACE RAW_NORM_SPACE RAW_PIXEL_SIZE RAW_POINT_SIZE RAW_PIXELSIZE RAW_POINTSIZE RAW_QUAD_WIDTH RAW_SMALL_CAP_SIZE RAW_STRIKEOUT_ASCENT RAW_STRIKEOUT_DESCENT RAW_SUBSCRIPT_SIZE RAW_SUBSCRIPT_X RAW_SUBSCRIPT_Y RAW_SUPERSCRIPT_SIZE RAW_SUPERSCRIPT_X RAW_SUPERSCRIPT_Y RAW_UNDERLINE_POSITION RAW_UNDERLINE_THICKNESS RAW_X_HEIGHT RELATIVE_SETWIDTH RELATIVE_WEIGHT RESOLUTION _MULE_BASELINE_OFFSET _MULE_RELATIVE_COMPOSE                       8       o�H                                           KC     8      X       0      `ZC     `OC                                      HC                             LC     �GC     o�H     ЇH     `1H     �H                     �GC     �SC     (        FC     @FC     `FC     �FC                                             ��������              �~   ~                         �                                                                         	       
                          
                                                         �H                   ��H                   ��H                   ΄H                   �H                   �H                   B�H                   1�H                   P�H                   .�H                   X�H                   8�H                   D�H                   �H                   U�H                   �H                   �H                   �H                   _�H                   e�H                   q�H                   q�H                   y�H                   ��H                    �H                   .�H                   <�H                   ��H                   K�H                   Z�H                   ��H                   ��H                   ��H                   ��H                   ʄH                   �H                   �H                   ��H                   �H                   �H                   *�H                   8�H                   G�H                   V�H                   e�H                   s�H                   ��H                   ��H                   ��H                   ��H                   ΅H                   �H                   �H                   �H                   �H                   (�H                   :�H                   Q�H                   i�H                   v�H                   ��H                   ��H                   �H                   $�H                   �H                   �H                   ��H                   ~�H                   ��H                   ��H                   ҅H                   �H                   ��H                   �H                   �H                   ,�H                   >�H                   U�H                   ��H                   �H                   m�H                   ��H                   ��H                                           8�C     @�C     P�C     h�C     p�C     �C      �C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     ��C     i�C     ��C     ��C     i�C     i�C     ��C     ��C     ��C     I�C     `�C     i�C     i�C     i�C     i�C     i�C     i�C     i�C     *�C     *�C     *�C     F�C     1�C     ^�C     �C     ^�C     ^�C     ^�C     �C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ^�C     ��C     �0D     �1D     �1D     �1D     X0D     �1D     �1D     �1D     "0D     �1D     �1D     �1D     �/D     �/D     �1D      2D              ,         ( * 0 8 @ H P                                    ����cinu    ����cinu       nmra       bmys   
   cinu      cinu      sijs        bg      5gib      snaw      ahoj                             $    
             " $ &                           
             "                    � �      
 x z | ~ �           h p                      N       
             ! " # $ % & ' ( ) 0 8 @ H P Q R S T V X Z \ ^ ` b                                ( 0 8                                                          6           , 4 	: 	; < =                                  6        " ( 0 8 @ H J L N P R T V X                                       
                �H     ��H      �H     ��H      �H     ��H      �H     ��H      �H                             (       P�C     0�C     ��C     ��C                                             ����                                            H       СC     ��C      �C     �C     @�C     ФC     ��C     ��C     @�C              D      �C                             P       ПC             ��C     @D                                                    ��C     ��C                             P       0�C             ��C      D                                                    p�C     ��C                             (       ��C              �C     `�C                                             
       ��C     �C                             (       ��C             ��C      �C                                                     �C      �C                             (       ��C             @�C     ��C                                                    �C     `�C                             P       ��C             ИC     �D                                                     �C     �C                             (       ��C             ��C     P�C                                                    ��C     ��C                             (       ��C             ��C     ��C                                                     �$D      �C                                            �1H                    �H                     P�C                             �C     `D     ��C     @�C     P�C     ��C     PD     ��C     �D     ��C     `D     ��C      �C     0�C     `�C     @�C     ��C     @D     P%D     �D      �C     ��C      D     ��C     ��C     ��C     ��C     ��C     0�C     ��C     ��C             k.H     ��H     V.H     x�H     K.H     ��H     o�H     `�H     v.H     p�H                     0�C     @�C     ��C     �)D     0123456789ABCDEF    �|���������W�D     �D     ��C      �C     @D     glyph-to-script-map fallback-script default-script increase-x-height warping autofitter 田 囗 ꘓ ꖜ ꖴ า ๅ ๐ ⵔ ౦ ౧ ꪒ ꪫ ௦ ᮰ ට 𐑴 ꢝ ꣐ 𐒆 𐒠 𐓂 𐓪 𐰗 ᱛ ߋ ߀ ဝ င ဂ ഠ റ ꓳ ᵒ ᴼ ⁰ ₒ ₀ o O 0 ໐ ೦ ಬ ᧡ ᧪ ០ ꤍ ꤀ ם ਠ ਰ ੦ ટ ૦ ο Ο 𐌴 𐌾 𐍃 Ⱅ ⱅ Ⴖ Ⴑ ⴙ ი ე ა ዐ 𐐄 𐐬 ठ व ट о О 𐠅 𐠣 Ⲟ ⲟ Ꭴ Ꮕ ꮕ 𐊫 𐋉 ᑌ ᓚ 𑄤 𑄉 𑄛 ᝋ ᝏ ০ ৪ ꛁ ꛯ 𐬚 ս Ս ل ح ـ 𞤌 𞤮                              #                      
                                                         ��������������������������������������������������������������������������������                                                          
                      *0  /0  �1  �1                     �  �.  �.   /  �/  �/  �/   0  ?0  @0  �0  �0  �0   1  /1  01  �1  �1  �1  �1  �1  �1  �1  �1  �1   3  �3   4  �M  �M  �M   N  ��  `�  �   �  ��  ��  ��   �  ��  �  �  0�  O�   �  ��   � ��  � _�    ߦ  � ?� @� �  � �                     5  5  7  7  9  9  >  ?  q  ~  �  �  �  �  �  �             �          �  �  �  �  �  �  %�  &�                   �  /�              <  <  ?  ?  A  D  M  V  b  c                                                  "  '  4  7  ;             O                           �  ?�                          0-  -                          1  1  4  :  G  N                                             >  @  F  V  b  c                               ��  ��  ��  ��  ��  ��  ��  ��  ��  ��          ��  ߪ          �  �  �  �  �  �          �  �          �  �  �  �                  �  �  �  �                  �  �  �  �                  �  �                          P          ��  ��  ��  Ũ                  ��  ߨ                          � �                         � �                           O                         P                            �  �          �  �          -  0  2  7  :  :  =  >  X  Y  ^  `  q  t  �  �  �  �  �  �  �  �  |�  |�                                     �  �  ��  `�  �              M  N  b  c                                       Ф  ��                          �   �   �   �   �   �   �  �  �  �  ,  a  x  x  �  �  p      },  },  p�  p�  ��  ��  \�  _�                          b  j  �   �   |,  |,          ^   `   ~   ~   �   �   �   �   �   �   �   �   �   �   �  �  �  �     o  �  �  �  �        >   >   ��  ��  ��  ��                                         �   �   �   �   �   �   �   �        �  O  P  �  �  �  �  �     o  �  �     +  k  w  y    �  �  �  �     �      o   �   �   �   �   P!  �!  `,  {,  ~,  ,   .  .   �  o�  q�  ��  ��  ��  0�  [�  `�  o�   �  �   � ��                                 �  �  �  �  �  �          �  �                          �  �                          �  �  �  �  �  �  �  �                  �  �          �  �  �  �  �  �  �  �  �  �  �  �                  �  �          &�  -�           �  /�                          �  �  �  �  �  �  �  �  �  �          �  �  �  O�                                  
  
  <
  <
  A
  Q
  p
  q
  u
  u
           
  
          �
  �
  �
  �
  �
  �
  �
  �
  �
  �
          �
  �
          z  z  �  �  �  �  �  �  �  �  �  �  �  �          p  �     �                  0 O          � /�          ,  _,   � /�                 �  �   -  --                  �  �          ]  _               �  �  �-  �-   �  /�                    O          	  	  :	  :	  A	  H	  M	  M	  S	  W	  b	  c	  �  �           	  ;	  =	  P	  S	  c	  f	  	  �   �   �  ��                  �  �  �-  �-  o�  �  ��  ��                                     �     /  �-  �-  @�  ��  �  �                            ?         �,  �,          �,  �,                          �  �  p�  ��                  � �                              �  �                     ' 4                   O         R  S          @  _                          �	  �	  �	  �	  �	  �	  �	  �	  �	  �	          �	  �	          �  �          ��  ��          9 ?           ?         Y  _          0  �  �  �                                           K  _  p  p  �  �  �  �  �  �  �  �  �  �  �  �  ��  ��  p�  p�  r�  r�  t�  t�  v�  v�  x�  x�  z�  z�  |�  |�  ~�  ~�             �  P  �  �  �  P�  ��  p�  ��   � ��                 D� J�          � _�                H       �H                   ��H     @;D     �;D     pbD                                                     �|D     8.H     ��H                     ��D     �D                            ��      @�D     �`D             �8D     p:D     ��D            �p      ��D     �VD             �8D     �8D     ��D     ��H     p�H     P�H     0�H     �H     ��H     ��H     ��H     ��H     p�H     P�H     0�H     �H     ��H     ��H     ��H     ��H     p�H     P�H     0�H     �H     �H     пH     ��H     ��H     p�H     P�H     0�H     �H     �H     оH     ��H     ��H     p�H     P�H     0�H     �H     �H     нH     ��H     ��H     p�H     P�H     0�H     �H     �H     мH     ��H     ��H     p�H     P�H     0�H     �H     �H     лH     ��H     ��H     p�H     P�H     0�H     �H     �H     кH     ��H     ��H     p�H     P�H     0�H     �H     �H     йH     ��H     ��H     p�H     P�H     0�H     �H     �H     иH     ��H     ��H     p�H     P�H     0�H                                     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H     ��H     @�H      �H     ��H                              �H     �H     @�H      �H                     S      8   �   
               R      7       
               Q      6       
               P      5       
               O      4       
               N      3   �   
               M      2   �   
               L      1   �   
               K      0   �   
               J      /   �   
               I      .   �   
               H      -   �   
               G      ,   �   
               F      +   �   
               E      *   �   
               D      )   �   
               C      (   �   
               B      '   �   
               A      &   �   
               @       %   �   
               ?      $   �   
               >      #   �   
               =      "   �   
               <      !   �   
               ;          �   
               :         �   
               9         �   
               8         �   	               7         �                  6         �                  5         �                  4         �                  3         �                  2         �                  1         �                  0         �                   /         �   
               .         �   
               -         �   
               ,         �   
               +         ~   
               *         z   
               )         t   
               (         n   
               '         g   
               &         g   	               %         g                  $         g                  #         g                  "         g                  !         g                            g                           g                           g                            d   
                        _   
                        X   
                        S   
                        P   
                        K   
                        E   
                        ?   
                        ?   	                        ?                           ?                           ?                           ?                           ?                           ?                           ?                           ?                            :   
                        5   
               
      
   .   
               	      	   +   
                        $   
                            
                           
                           
                           
                           
                        	   
                           
                              
                               8        �H     �H              �H                             7       P�H      �H             �DH                             6       ��H     `�H             �DH                             5       �H     ��H             �DH                             4        �H      �H             �DH                             3       @�H     0�H             (�H                             2       ��H     ��H             4�H                             1       `�H     P�H             @�H                             0       �H     ��H             D�H                             /       0�H      �H             L�H                             .       `�H     @�H             T�H                             -       ��H     p�H             X�H                             ,       ЦH     ��H             \�H                             +       �H     �H             `�H                             *        �H      �H             e�H                             )       @�H     0�H             m�H                             (       `�H     P�H             w�H                             '       ��H     p�H             ��H                             &       ��H     ��H             ��H                             %       ��H     ��H             /H                             $       ЧH     ��H             ��H                             #       `�H     �H             ��H                             "       ��H     ��H             ��H                             !       ��H     ��H             ��H                                     �H     ШH             ��H                                    `�H     P�H             ��H                                     �H     ��H             ��H                                    `�H     @�H              H                                     �H     �H             ƠH                                    ��H     p�H             ΠH                                    ЫH     ��H             ֠H                                    @�H     0�H             ڠH                                    ��H     `�H             �H                                    �H     ��H            �H                                    0�H      �H             �H                                    ��H     @�H             ��H                                    ��H     ��H            ��H                                    ��H     ��H             �H                                    �H     حH             �H                                     �H     ��H             "�H                                     �H     �H             .�H                                    P�H     H�H             2�H                                    ��H     `�H            <�H                                     �H     �H             H�H                                    `�H     P�H             N�H                                    ��H     p�H             X�H                             
       ��H     ��H             `�H                             	       ��H     ��H             l�H                                    �H     ЯH             v�H                                     �H      �H             ~�H                                    @�H     0�H             ��H                                    ��H     `�H            ��H                                    ��H     ��H             ��H                                    аH     ��H             ��H                                    �H     �H             ��H                                    ��H      �H             ��H                                     �H      �H             ��H                                     H                                       @8D     `jD            �p      0�D     �VD             P5D     7D     �D                   (   	   A       )      i      {       �      )      �      �       �      �   	   �             )           .      )      8     X      )      �     �     x     x      )      �     �     �  	   �      )           4      M      )           4      T  	   t      �     �      )      �     �      )      �     �      �     �  	   �      �      )      �           >  	   ^      )      ~     �      �     �      )      �     �        	                )      �     �     �     �      �      )      )     B      [  	   t      )      �           )      5  	   U      u     �      )      �     �      �  	         5     U      )      u     �      �  	   �      )      �           )      1     F      X     j  	   j      �      )      �  	   �      �     	      -	     )      �	     a	     A	     �	      �	     )      �	     �	      �	      )      Z
  	   r
      �
     �
      �
      )      �
  	   �
     �
            1      )      �  	   �      )      
     :
      )      �  	   �      �     �     �      )                 ,     :  	   J      Z      )      d     x      �     �  	   �      �      )      �     �           .  	   .      G      )      R     r      )      �     �      )      �  	   �           :      )      Z     r      �  	   �      )      )      �     �      )      �     �      )      �     �            &  	   N      v     �      )      �     �      )      �           )      "     ,      E      O  	   r      )      �     �      �      )      �           %      )      M     m      )      -     A      )      �     �      )      5     5      )      �  	   �      �                !      )      )      U     u      )      �     _      )      𞤌 𞤅 𞤈 𞤏 𞤔 𞤚 𞤂 𞤖 𞤬 𞤮 𞤻 𞤼 𞤾 𞤤 𞤨 𞤩 𞤭 𞤴 𞤸 𞤺 𞥀 ا إ ل ك ط ظ ت ث ط ظ ك ـ Ա Մ Ւ Ս Բ Գ Դ Օ Ւ Ո Դ Ճ Շ Ս Տ Օ ե է ի մ վ ֆ ճ ա յ ւ ս գ շ ր օ հ ո ճ ա ե ծ ս օ բ ը ի լ ղ պ փ ց 𐬀 𐬁 𐬐 𐬛 𐬀 𐬁 ꚧ ꚨ ꛛ ꛉ ꛁ ꛈ ꛫ ꛯ ꚭ ꚳ ꚶ ꛬ ꚢ ꚽ ꛯ ꛲ অ ড ত ন ব ভ ল ক ই ট ঠ ি ী ৈ ৗ ও এ ড ত ন ব ল ক ᝐ ᝈ ᝅ ᝊ ᝎ ᝂ ᝃ ᝉ ᝌ ᝀ ᝃ ᝆ ᝉ ᝋ ᝏ ᝑ ᗜ ᖴ ᐁ ᒣ ᑫ ᑎ ᔑ ᗰ ᗶ ᖵ ᒧ ᐃ ᑌ ᒍ ᔑ ᗢ ᓓ ᓕ ᓀ ᓂ ᓄ ᕄ ᕆ ᘣ ᕃ ᓂ ᓀ ᕂ ᓗ ᓚ ᕆ ᘣ ᐪ ᙆ ᣘ ᐢ ᒾ ᣗ ᔆ ᙆ ᗮ ᒻ ᐞ ᔆ ᒡ ᒢ ᓑ 𐊧 𐊫 𐊬 𐊭 𐊱 𐊺 𐊼 𐊿 𐊣 𐊧 𐊷 𐋀 𐊫 𐊸 𐋉 𑄃 𑄅 𑄉 𑄙 𑄗 𑄅 𑄛 𑄝 𑄗 𑄓 𑄖𑄳𑄢 𑄘𑄳𑄢 𑄙𑄳𑄢 𑄤𑄳𑄢 𑄥𑄳𑄢 Ꮖ Ꮋ Ꭼ Ꮓ Ꭴ Ꮳ Ꭶ Ꮥ ꮒ ꮤ ꮶ ꭴ ꭾ ꮗ ꮝ ꮿ ꮖ ꭼ ꮓ ꮠ ꮳ ꭶ ꮥ ꮻ ᏸ ꮐ ꭹ ꭻ Ⲍ Ⲏ Ⲡ Ⳟ Ⲟ Ⲑ Ⲥ Ⳋ Ⳑ Ⳙ Ⳟ Ⲏ Ⲟ Ⲑ Ⳝ Ⲱ ⲍ ⲏ ⲡ ⳟ ⲟ ⲑ ⲥ ⳋ ⳑ ⳙ ⳟ ⲏ ⲟ ⲑ ⳝ Ⳓ 𐠍 𐠙 𐠳 𐠱 𐠅 𐠓 𐠣 𐠦 𐠃 𐠊 𐠛 𐠣 𐠳 𐠵 𐠐 𐠈 𐠏 𐠖 Б В Е П З О С Э Б В Е Ш З О С Э х п н ш е з о с р у ф 𐐂 𐐄 𐐋 𐐗 𐐑 𐐀 𐐂 𐐄 𐐗 𐐛 𐐪 𐐬 𐐳 𐐿 𐐹 𐐨 𐐪 𐐬 𐐿 𐑃 क म अ आ थ ध भ श ई ऐ ओ औ ि ी ो ौ क म अ आ थ ध भ श ु ृ ሀ ሃ ዘ ፐ ማ በ ዋ ዐ ለ ሐ በ ዘ ሀ ሪ ዐ ጨ გ დ ე ვ თ ი ო ღ ა ზ მ ს შ ძ ხ პ ს ხ ქ ზ მ შ ჩ წ ე ვ ჟ ტ უ ფ ქ ყ Ⴑ Ⴇ Ⴙ Ⴜ Ⴄ Ⴅ Ⴓ Ⴚ Ⴄ Ⴅ Ⴇ Ⴈ Ⴆ Ⴑ Ⴊ Ⴋ ⴁ ⴗ ⴂ ⴄ ⴅ ⴇ ⴔ ⴖ ⴈ ⴌ ⴖ ⴎ ⴃ ⴆ ⴋ ⴢ ⴐ ⴑ ⴓ ⴕ ⴙ ⴛ ⴡ ⴣ ⴄ ⴅ ⴔ ⴕ ⴁ ⴂ ⴘ ⴝ Ⰵ Ⱄ Ⱚ Ⰴ Ⰲ Ⰺ Ⱛ Ⰻ Ⰵ Ⰴ Ⰲ Ⱚ Ⱎ Ⱑ Ⰺ Ⱄ ⰵ ⱄ ⱚ ⰴ ⰲ ⰺ ⱛ ⰻ ⰵ ⰴ ⰲ ⱚ ⱎ ⱑ ⰺ ⱄ 𐌲 𐌶 𐍀 𐍄 𐌴 𐍃 𐍈 𐌾 𐌶 𐌴 𐍃 𐍈 Γ Β Ε Ζ Θ Ο Ω Β Δ Ζ Ξ Θ Ο β θ δ ζ λ ξ α ε ι ο π σ τ ω β γ η μ ρ φ χ ψ ત ન ઋ ઌ છ ટ ર ૦ ખ ગ ઘ ઞ ઇ ઈ ઠ જ ઈ ઊ િ ી લી શ્ચિ જિ સી ુ ૃ ૄ ખુ છૃ છૄ ૦ ૧ ૨ ૩ ૭ ਕ ਗ ਙ ਚ ਜ ਤ ਧ ਸ ਕ ਗ ਙ ਚ ਜ ਤ ਧ ਸ ਇ ਈ ਉ ਏ ਓ ੳ ਿ ੀ ਅ ਏ ਓ ਗ ਜ ਠ ਰ ਸ ੦ ੧ ੨ ੩ ੭ ב ד ה ח ך כ ם ס ב ט כ ם ס צ ק ך ן ף ץ ಇ ಊ ಐ ಣ ಸಾ ನಾ ದಾ ರಾ ಅ ಉ ಎ ಲ ೦ ೨ ೬ ೭ ꤅ ꤏ ꤁ ꤋ ꤀ ꤍ ꤈ ꤘ ꤀ ꤍ ꤢ ꤖ ꤡ ꤑ ꤜ ꤞ ꤑ꤬ ꤜ꤭ ꤔ꤬ ខ ទ ន ឧ ឩ ា ក្ក ក្ខ ក្គ ក្ថ ខ ឃ ច ឋ ប ម យ ឲ ត្រ រៀ ឲ្យ អឿ ន្ត្រៃ ង្ខ្យ ក្បៀ ច្រៀ ន្តឿ ល្បឿ ᧠ ᧡ ᧶ ᧹ າ ດ ອ ມ ລ ວ ຣ ງ າ ອ ບ ຍ ຣ ຮ ວ ຢ ປ ຢ ຟ ຝ ໂ ໄ ໃ ງ ຊ ຖ ຽ ໆ ຯ T H E Z O C Q S H E Z L O C U S f i j k d b h u v x z o e s c n r x z o e s c p q g j y ₀ ₃ ₅ ₇ ₈ ₀ ₁ ₂ ₃ ₈ ᵢ ⱼ ₕ ₖ ₗ ₐ ₑ ₒ ₓ ₙ ₛ ᵥ ᵤ ᵣ ᵦ ᵧ ᵨ ᵩ ₚ ⁰ ³ ⁵ ⁷ ᵀ ᴴ ᴱ ᴼ ⁰ ¹ ² ³ ᴱ ᴸ ᴼ ᵁ ᵇ ᵈ ᵏ ʰ ʲ ᶠ ⁱ ᵉ ᵒ ʳ ˢ ˣ ᶜ ᶻ ᵖ ʸ ᵍ ꓡ ꓧ ꓱ ꓶ ꓩ ꓚ ꓵ ꓳ ꓕ ꓜ ꓞ ꓡ ꓛ ꓢ ꓳ ꓴ ഒ ട ഠ റ ച പ ച്ച പ്പ ട ഠ ധ ശ ഘ ച ഥ ല ခ ဂ င ဒ ဝ ၥ ၊ ။ င ဎ ဒ ပ ဗ ဝ ၊ ။ ဩ ြ ၍ ၏ ၆ ါ ိ ဉ ည ဥ ဩ ဨ ၂ ၅ ၉ ߐ ߉ ߒ ߟ ߖ ߜ ߠ ߥ ߀ ߘ ߡ ߠ ߥ ߏ ߛ ߋ ߎ ߏ ߛ ߋ ᱛ ᱜ ᱝ ᱡ ᱢ ᱥ 𐰗 𐰘 𐰧 𐰉 𐰗 𐰦 𐰧 𐒾 𐓍 𐓒 𐓓 𐒻 𐓂 𐒵 𐓆 𐒰 𐓍 𐓂 𐒿 𐓎 𐒹 𐒼 𐒽 𐒾 𐓵 𐓶 𐓺 𐓻 𐓝 𐓣 𐓪 𐓮 𐓘 𐓚 𐓣 𐓵 𐓡 𐓧 𐓪 𐓶 𐓤 𐓦 𐓸 𐓹 𐓛 𐓤 𐓥 𐓦 𐒆 𐒉 𐒐 𐒒 𐒘 𐒛 𐒠 𐒣 𐒀 𐒂 𐒆 𐒈 𐒊 𐒒 𐒠 𐒩 ꢜ ꢞ ꢳ ꢂ ꢖ ꢒ ꢝ ꢛ ꢂ ꢨ ꢺ ꢤ ꢎ 𐑕 𐑙 𐑔 𐑖 𐑗 𐑹 𐑻 𐑟 𐑣 𐑱 𐑲 𐑳 𐑴 𐑸 𐑺 𐑼 𐑴 𐑻 𐑹 ඉ ක ඝ ඳ ප ය ල ෆ එ ඔ ඝ ජ ට ථ ධ ර ද ඳ උ ල තූ තු බු දු ᮋ ᮞ ᮮ ᮽ ᮰ ᮈ ᮄ ᮔ ᮕ ᮗ ᮰ ᮆ ᮈ ᮉ ᮼ ᳄ ꪆ ꪔ ꪒ ꪖ ꪫ ꪉ ꪫ ꪮ உ ஒ ஓ ற ஈ க ங ச க ச ல ஶ உ ங ட ப ఇ ఌ ఙ ఞ ణ ఱ ౯ అ క చ ర ఽ ౨ ౬ บ เ แ อ ก า บ ป ษ ฯ อ ย ฮ ป ฝ ฟ โ ใ ไ ฎ ฏ ฤ ฦ ญ ฐ ๐ ๑ ๓ ⵔ ⵙ ⵛ ⵞ ⴵ ⴼ ⴹ ⵎ ꗍ ꘖ ꘙ ꘜ ꖜ ꖝ ꔅ ꕢ ꗍ ꘖ ꘙ ꗞ ꔅ ꕢ ꖜ ꔆ 他 们 你 來 們 到 和 地 对 對 就 席 我 时 時 會 来 為 能 舰 說 说 这 這 齊 | 军 同 已 愿 既 星 是 景 民 照 现 現 理 用 置 要 軍 那 配 里 開 雷 露 面 顾 个 为 人 他 以 们 你 來 個 們 到 和 大 对 對 就 我 时 時 有 来 為 要 說 说 | 主 些 因 它 想 意 理 生 當 看 着 置 者 自 著 裡 过 还 进 進 過 道 還 里 面        0 1 2 3 4 5 6 7               `BH                   ��H     ��D     � E                     �D      �D     0�D     raster1                        �       ��H                           @E                     ltuo    �+E     �-E     p+E     pE     ��H             ltuo    0+E      E     0E     �'E     �E                     /E     �/E     �/E     �/E     �/E     �/E     v/E     p/E            �       ��H                           P.E                     ltuo    0BE     0HE     �/E     �.E     ��H                    �       ��H                           P.E                     ltuo     BE     0HE     �/E     �.E     ��H                    �       �H                           P.E                     ltuo     BE     0HE     �/E     �.E     ��H             ltuo    �;E     0.E     @.E     �3E     �.E                     p;E     @;E      HE     �EE                     smooth-lcdv smooth-lcd smooth unknown compression method invalid window size incorrect header check need dictionary invalid block type invalid stored block lengths invalid bit length repeat oversubscribed distance tree incomplete distance tree invalid literal/length code invalid distance code incorrect data check      too many length or distance symbols     oversubscribed dynamic bit lengths tree incomplete dynamic bit lengths tree     oversubscribed literal/length tree      incomplete literal/length tree  empty distance tree with lengths                YE     `YE     �WE     �ZE     �ZE     �YE     �YE     !`E     �ZE     ZE     �ZE     �XE     �ZE      YE     �[E     s\E     �bE     �aE     ^E     Y]E     VaE     XcE     �_E     ]E     LdE     xfE     4gE     �dE     /eE     �eE     �gE     �fE     �fE     i[E                                        	      
                                                                        ?      �   �  �  �  �  �  �?  �  ��                              P     W    S     [    Q     Y    U  A   ]  @  P     X    T  !   \     R  	   Z    V  �   �  `  P     W  �  S     [    Q     Y    U  a   ]  `  P     X    T  1   \  0  R     Z    V  �   �  `  `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �                                                                   	   	   
   
                                               	            !   1   A   a   �   �     �                     0  @  `                                                                                                          p   p                         	   
                           #   +   3   ;   C   S   c   s   �   �   �   �                 0�E     0�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     0�E     P�E     P�E     P�E     P�E     P�E     0�E     P�E     P�E     P�E     0�E     P�E     P�E     P�E     P�E     P�E     P�E     P�E     0�E     P�E     P�E     P�E     0�E     P�E     0�E     ��E     ��E     ��E     ȬE     �E      �E      �E     ��E     ЩE     ��E     ��E     ��E     `�E     0�E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     �E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     x�E     ��E     ��E     ��E     ��E     P�E     ��E     ��E     ��E     �E     ��E     ��E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     ��E     ��E     @�E     �E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     @�E     �E     ��E     `F     ��E     F     �F      F     �F     �F     hF     @F     @F     �E     `F     ��E     h F       F     x�E     ��E     `F     �E     �E     ��E     �E     F     hF     ��E     �E     �E     ��E     @F     �F     �F     u�E     �F     �F     �F     �F     u�E     �F     �F     �F     �F     �F     u�E     �F     �F     �F     �F     �F     u�E     �F     �F     �F     �F     �F     u�E     u�E     �F     <F     �F     xF     jF     FF     FF     FF     6 F      F     �F     FF     FF     FF     �F     wF     .F     FF     FF     F     �F     mF     mF     �F     FF     �F     �F     mF     5F     wF     FF     �F     �F     �F     CF     h F     FF     �F     �F     6 F      F     �F     iF     �F     FF     �F     wF     .F     FF     FF     F     �F     QF     F     �F     FF     �F     �F     mF     5F     wF     FF     �F     �F     �F     CF     h F     FF     FF     �F     �F     F     F     ^F     �F     �F     �F     �F     �F     �F     �F     �F     	F     	F     �F     �F     �F     �F     �F     �F     uF     VF     &F     �F     wF     *F     �F     �F     �F                                               (        �E     @�E     P�E     `�E                                                             (       0�E     `�E     ��E     ��E                                                             8       �E     ��E     ��E     ��E                                                             8       ��E     ��E     ��E     ��E                                                             ������������������������������������������������ 	�������
 !"#������
 !"#�����               �BH                   �I                                                     �I     @I     �I     �I      �E     p�E     жE     @�E     �I     �I      I             ��E     P�E     `!F             кE     ��E     `�E     �E     ��E      �E     ��E     @�E     �I      I     �I     `I      �E      �E     p�E             ��E     ��E     p�E     `!F     ��E     ��E     ��E     ��E     ��E     ��E     @�E     ��E      �E     �E                     �E     ��E     ��E     `�E     p�E     �E     ��E     ��E     ��E     ��E     p�E     ШE     @�E                             ��E     p�E     ��E     0�E     0I     OI     YI     bI     �DH     wDH     bDH     sI     rI     dI     gI     qI     {I     �I     �I     �I     �I     �I     �I     �I     �I     �I     �I     I     I     CH     +DH     �gH     CH     I     &I     0I     =I     'CH     FI     II     MI     QI     UI     WI     eI     B�H     CH     qI     uI     I     �I     �I     >I     �I     �I     �I     �I     �I     �CH     �CH     	I     @CH     RCH     �I     �I     =hH     �CH     I     	I     I     I     I     I     I     I     �1H     �DH     "I     Ascender true StartFontMetrics AxisLabel AxisType B CH CapHeight CharWidth CharacterSet Characters Descender EncodingScheme EndAxis EndCharMetrics EndComposites EndDirection EndFontMetrics EndKernData EndKernPairs EndTrackKern EscChar IsBaseFont IsCIDFont IsFixedPitch IsFixedV KP KPH KPX KPY L MappingScheme MetricsSets PCC StartAxis StartCharMetrics StartComposites StartDirection StartKernData StartKernPairs StartKernPairs0 StartKernPairs1 StartTrackKern VV VVector W0 W0X W0Y W1 W1X W1Y WX WY XHeight psnames                              *I                   �I                     P1F                             �BH     �I                     �2F     4F     �/F     P0F      1F      1F     ��I     ��I                     #   &   5   ;   H                           Delta Omega fraction hyphen macron mu periodcentered space Tcommaaccent tcommaaccent            �  �  "  �   �  �  "  �                                4 j�?�}	�
���W��hXn GM�I� k �!7"�#�:
@zH�PmXh]=b�j[ros�z�������՞l�s�������̦���Q�A� A � � ����(9R[���E� � � � �����e�������n������l�������e� � �����l�������e� � � � � �����e���������c���������w������e����������e������e��c y����n����c(-�e�$������x� �BJU]iq����e���������w������e����������e������l�������e����e��������l���������c�d���������e� ������s� �����������c�������n������l����t������w�������n������e� ������l�����������e��i��������c�������������e����a��1����s��m?G����n� �������e��!�����k����g� �hpx����e������w� ����l�������l��a����e� ������l������������n�1B� B���
".6�����e�$���t�������t�����w�e����������c���������n�2�a�����k����������w���������e��"��������l�������l��b�����r��C� CU�������a]ho�������n�>���e���n���w����l���c������n������a� �������e�����l�����c���e�$������x���t�
������t�
����������l���h������������n�Ie#gs�����������������c���������c�'d)U�������r6J����������������c���������c����������������c����������n�C�����������������c�����������������������c��i����k���������������l�����������e��#��������n�Q����l��cD� D�
$`y���� 09Z������n��a�������n�4�����n��c.5>Y���n������a���cFK�e�$�����������w����t���thq�����t�
����w�e����������c�������c����a�"�����k�����k��i�������s����������e�������e�������l������������k�����������c���������w���������e��$������������l���s")���h����l��d�����r��z��CKp����n��eQe����������������c���������c����������c�E� E���Y����$^����	,	m	s����e� ������l�������e�c����O���n�����������e���������n�5��c���e�$������x� � +3?G����e������w��������w������e����������e������l�������e��������c�dak������e�������s� �w����l����t��������t�����w����������c�$����e� ������l���h���������n�7�������e��i����������n�!g�����������e���������������c�dl�������c���������n�!jm,HS����n�8@����e�����e��������c��������e��%nhs���������c�����������������c��g�J����������c�������������c��o������k���n�������n�������s��r���������c� ������d����������c�-s			!	%�������c�!����������������c��h�����l��et	4	N	\a��	<	F������n�8����s��h� �	T����l������e��	e����w���o� ��h��	|	�����n���������d��F� F	�	�	�	�	�	�

�����e�$���������t�e	�	���������n�V������c�����k��i	�	����������c�r������n�!d��������e��&�������n�!c����l��fG� G
3
=
k
s
�
�
�'4AZk������e�3�a
E
L
^���e����a��
T������n�����������c������e�c
}
�
�
����n�������a�"��c
�
��e�$������x����������t�"��t� 
������t� ��������c�h
�
�!���������n�Be
�
������������������c���������������c���������������c����k�����������n�3���������c�mGO����n� �������e��'���e���c����l��`sq����l��gz���k������e��H� H����(Mu������5����3�%ϴ3�%��1�%�����3�%�������e�3�a�� ����������������c������������������c���������������c�*b�r�&��������w�*c.7�����a�(��c?D�e�$������x�$dS]������s�&�tdm�����t�"����w�$��������e��(o���������n�@�������c������l��h����������t��������l���������e�3�I� I���%^�����0Vc�����������c�/J�2��������c�.����e� �����l�������e�,c-4T���n����c<A�e�$������x� �L����l���������c�dfp�������e�������s� ��������e�.�������c������l����t�0�������t�0����w��e��������������c���������c�������r�!����e� ������l�����������e��i �������c������������e�
������������c�m6K����n�*@�������c���������e��)���������n�;okv~�������c�����k�.�a�����������n���������s������s��s�����l��i����e������e�(�����w�,�����a���������c�t���������������c�vJ� J)5CO��������n�A���c �e�$������x�4��������c�����������n�K��������e��*����l��jK� Ks}�ALj�����������e�3�������e�3�a���������������������c��c����e�0������c�����������������c�������������c����a���������������c�����������������������c��c#,4���n�������a�6����e�$����������t�6�������w�2eR^��������n�T��������n�?hr~���������c�%�������c����k�����������c���������w�4��������e��+���a���������c������k��s����������c�n���l��kL� L	_�����J��L���a���e�9���a��c'.7R���n�=�����a�;��c?D�e�$�����������w�<���������t�;��t�?ir�����t�?����w�6|�����n�8����������n�<j�����������c�	��������w�:��������e��,s�����h�A�����l������l��lM� M��!:GS[d������e�3��c��n���
����l�����e�>�����e�$���t)2�����t�@����w�B���������n�D��������e��-����l��m�����d��u��N� N������!-:BTJ������e�Cc�������n�G�����a�E��c���e�$�����������w�J���������t�E��t�������t�D����w�F�������t���������n�!hj��	��������c�
��������w�H��������e��.���������n�F����l��n����e� �L����l���u��O� Ov���N��0E���5E�R|����l�������e� ������l���b������d���������c�����������������c�����e�Nc���D���n�������������e����c���e�$������x� � (4<����e���������w������e����������e������l�������e��������c�dVm��l]e����e�P����e�������s� �{��������c������l���������w��g����������l������e� ������l���h���"�������n�Um�!&o��������e���n��������e���������w������e����������e������e������������t�Pi��6�����������e�mOk������n�L[c����e�R����e�P��a�!&y����������c�`����k��������������c�zt�������������c�|���s������n�������s���������e��/������n�!`o������k��������n����n��s!(���h� �����e������l������l��o���������e��t;F�������c�~���e� �S[f����e�L�������s�N����l���P� P�����������e�T�����e�$���������t�Ve����������c���������n�J�����������������c��h��i����k��i������������n�S��������e��0si���������c�p���l��pQ� Q*3?�����e�$���������e��1����l��qR� R_w�����+aep�������n�L���e�Tc�������n�X�����a�V����e�$����������t�Vd��������e��t�������t�X����w�Z������n�\���������n�P������r�!�o���n������l�������������e���������w�^��������e��2����l��r5�������d��B�������r��S� Sg7���Tiu��Fu��Mw�0	��������ɱ���0�%����0�%����0�%����0�%����0�%<����0�%,����0�%4����0�%����0�%$1��鰰��0�% ����0�%����0�%a2	%-5=E����0�%b����0�%V����0�%U����0�%c����0�%Q����0�%W����0�%]����0�%\����0�%[3W_go����0�%^����0�%_����0�%Z����0�%T4
���������հ���0�%i����0�%f����0�%`����0�%P����0�%l����0�%g����0�%h����0�%d����0�%e����0�%Y5���	����0�%X����0�%R����0�%S����0�%k����0�%ja,���e�Z ��������t�d�������k��cCbk�����n�`NZ��������t�f����l��������a�^��a��u��������c�����������������c����c���e�$������x�\���������t���t�������t�`����w�b���������t�he����������n�M�������n�!fh"0;Ha�������n�G�������c�(����������c�)�������c�����������c����������c��iZ`��a�������n�!e��������e��3��������������c�,����l��s���������k��T� T��� `�����.�u����r�fc�������n�d�����a�b��c���e�$�����������w�p���������t�b��t�����t�j����w�le*5IR�������c�"����������������c�������n�!i����������c��hhn���a��oty�k���n� ������l����������n�!bi���������l������������n�O��������w�n��������e��4o���������n�9�e������e����x����o��������������k��s'��������c�&���������c����l��tw4@��������n�!k�����n�!aU� Ui{��EW����������e� �s����l�������e�lc������n����c���e�$������x� �������w�v����l���������c�#d��;�l������e�p����e�������s� ��"*3����e������w�rc���n��������c������e�������n������l���������w������e� �O����l���h]�ocm������e���n��|��������e���������w������e����������e������e������������t�p��������c��������������e���������c�xm�
����n�j���������c���������s�z�������e��5�����k�r�����n��15Zy�1��a;Q������������������k�������n���������s��g��������������k�����������l������s�����g�ns��������������c����l��u������t���������c���������������c������e�h������e�x����w�tV� V    < C O [ c�����e�$��������w�~e % 0�������c���������n�N���k����������e��6��������n�H����l��v����e�|W� W { � � � � �����e�����c � ��e�$������x�td � �������s���t � ������t������w������e����������e��7����l��wX� X � �!!!#!/�����e�$�d �!������s���������t�����������n�=i����������e��8����l��xY� Y!Q!t!�!�!�!�!�"("4"<"Da!W!h���e� �!`����l�����������c�b���c!}!��e�$������x�vd!�!�������s�x!�����l����t!�!������t������w���r!�!���������c�+����������������c������e�����k��!�����e��i"""�������n�E�������c����������n�R��������e��9����l��y����e���s"K"q��g"S"^�������c�j���������������c�l�����e"|"��������c�f���������������c�hZ� Z"�"�"�##Q#�#�#�a"�"��������n�6���e�yc"�"����n�}"�����l�����c"�"��e�$������x����t�{"�#�����t�{����w��e##!#L�������c�d#'#:���������������c����������������c���a���e#\#g#w#��������n�:������������c���������c�d#�#����������������c����������������c����������w����������e��:s#�#����l��z����e��a� a$&�''D'�'�((D(~(�)F)�*�*�+1�1�2 2�34`4�5{5�689929�9�1�'$2$r$�$�%%Z%�%�&&Z0�'!$J$N$R$V$Z$^$b$f$j$n0�'^1�'a2�'b3�'c4�'d5�'6�'e7�'f8�'g9�&`1�&$�$�$�$�$�$�0�&e1�&f2�&c7�'	8�'9�'2�&$�$�$�$�$�$�$�$�$�$�0�$`1�$a2�$b3�$c4�$d5�$e6�$f7�$g8�$h9�$i3�'$�$�$�$�%%%
%%%0�'v1�'w2�'x3�'y4�'z5�'{6�'|7�'}8�'~9�'4�'%2%6%:%>%B%F%J%N%R%V0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�5�'%r%v%z%~%�%�%�%�%�%�0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�6�'%�%�%�%�%�%�%�%�%�%�0�'�1�!�2�'�3�!�4�!�5�'�6�'�7�'�8�'�9�'�7�'%�%�%�%�&&&
&&&0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�8�'&2&6&:&>&B&F&J&N&R&V0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�9�'&r&v&z&~&�&�&�&�&�&�0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�2�'&�&�&�&�&�&�&�&�&�' 0�'&�&�&�&�&�&�&�0�'�1�'�2�'3�'P4�'R5�'n6�'p1�'2�'3�'4�'5�'6�'7�'8�'9�'"3�''' '$'(','0'4'8'<'@0�'#1�'$2�'%3�'&4�''5�&6�')7�'*8�'+9�',4�&'\'`'d'h'l'p't'x'|'�0�'-1�'.2�'/3�'04�'15�'26�'37�'48�'59�'65�''�'�'�'�'�'�'�'�'�'�0�'71�'82�'93�':4�';5�'<6�'=7�'>8�'?9�'@6�''�'�'�'�'�'�'�'�'�( 0�'A1�'B2�'C3�'D4�'E5�'F6�'G7�'H8�'I9�'J7�'(( ($(((,(0(4(8(<(@0�'K1�%�2�'M3�%�4�'O5�'Q6�%�7�%�8�%�9�'V8�'(Z(^(b(f(j(n(r(v(z1�%�2�'X3�'Y4�'Z5�'o6�'q7�'r8�'s9�'h9�' (�(�(�(�(�(�(�(�(�(�0�'i1�'l2�'m3�'j4�'k5�'t6�'u7�'[8�'\9�']a(�(�(�(�(�))������i�	����e� ����a�	�u(�(������i�
������i�
������������i�
>�������e�3��������n)*)4);������i�	����a�	>�������i�
�b)P)y)�)����������n)_)n�����������n�_�������a�	p�����i�	�������o�1���e�)�)�)�)�)�)�����e���������c���������w������e����������e������e��c)�)�*9*���n����c)�)��e�$������x� �*
***%*1����e���������w������e����������e������e����e� �*I*T*e*l*u�������b�c*Z*_�b���b����a�	T�����d��������b�A������c�0d*�*�*�*�*�������e�����������i�
q��a�	������s� �*�*��������c�������n���t*�*�����w�������n��e� �*�*�+����e�������n�1P�����n����i+!+5-�-�.1o0+'+.���8� ���1� ��0+>-V-�0	+R+f+�+�, ,^,�,�-1+Z+^+b7�8�9�2
+|+�+�+�+�+�+�+�+�+�0�1�2�3�4�5�6�7�8�9�3
+�+�+�+�+�+�+�+�+�+�0�1�2�3�4� 5�!6�"7�#8�$9�%4
+�+�, ,,,,,,,0�&1�'2�(3�)4�*5�+6�,7�-8�.9�/5
,6,:,>,B,F,J,N,R,V,Z0��1�2�3�4�5�6�7�8�	9�
6
,t,x,|,�,�,�,�,�,�,�0�1�2�3���4���5�06�17�28�39�47
,�,�,�,�,�,�,�,�,�,�0�51�Q2�63�74�85�96�:7�;8�<9�=8
,�,�,�,�- -----0�>1�?2�@3�A4�B5�C6�D7�E8�F9�G9
-.-2-6-:->-B-F-J-N-R0�H1�I2�J3�K4�L5�M6�N7�O8��9�R1-`-�-�-�0
-v-z-~-�-�-�-�-�-�-�0�S1�T2�U3�V4�W5�X6�Y7�Z8�[9�\�0�^4-�-�-�-�5�6�b7�r8�t9-�-�-�-�-�2���3�_4�c5�s6�u8-�-�3-�-�1���2��ȴ6�ٲ�9� �0..0� 1� �7..b/�/�0�1"1i3.".08.(.,1�j8�9.B.F.J.N.R.V.Z.^2�`3�a4�b5�c6�d7�e8�f9�g4.r.�.�//./f/�0.~.�.�.�.�0�h1�i3�7�9�!1
.�.�.�.�.�.�.�.�.�.�0�"1�#2�$3�%4�&5�'6�(7�)8�*9�+2
.�.�.�.�.�.�.�///
0�,1�-2�.3�/4�05�16�27�38�49�53///"/&/*0�61�72�83�94�:4	/B/F/J/N/R/V/Z/^/b0�@1�A2�B3�C4�D5�E6�F8�H9�I5	/z/~/�/�/�/�/�/�/�0�J1�K2�L3�M4�N5�O6�P7�Q8�R�0�G5/�/�/�0/�/�/�/�/�5��6�~7��8��9��1/�/�/�/�/�1�y2��3��4��9�ҳ4��60 00
0050s0��6� ��5���8��600!0%0)0-014��5��6��7��8��9��7
0K0O0S0W0[0_0c0g0k0o0��1��2��3��4��5��6��7��8��9��8
0�0�0�0�0�0�0�0�0�0�0��1��2��3��4��5��6��7��8��9��90�0�0�0��4��*5��+70�0�0�0�00�0�0��K5��10�0�0�6��7��8��3��5911
111113��4��5��6��7��8��9��81*1V1[01:1>1B1F1J1N1R0��1��2��3��4��6��7���9��41a1e1��2����9��61w1�1�11�1�1�1�21�1��8�!�9�!��2�!�71�1�1�3� ,4� -5� .��4� ���7�m���7��g1�1����e� �u1�1������i�
������i�
h1�1�������a�0B�������e��i22)202<2U2e2�b22�����i�	�������o�1���a�	��������c���u2C2L�����i�
������i�
������������i�
Hn2q2z2�2�2������c�9����������c���������������c��������������c�������������e���������n2�2�2�������i�	����a�	H�������i�
�k2�2�������a�0�2���������h��q����n�1Ol34G4Pe34Bf��3)323A3O3�3�4%43�����c�'�����������w��0����������c���h3U3����a3^3����e3h3q�����c�#����������c�������w3�3������c�%����������c�������w������������w��O�a3�3��������e3�3������c�"����������c�������a3�3�44�����c�I����������c���������������c��������������c�������������w��.�����������w��/�h�!5�����l�"L��a��4X����s��m4j4r4}4�����n��������e��A������d� &4�4���������e������l��&�����e�3�n4�4�575A�������o�1"g4�4�4�5/�������o�1$����������i�Z�e�" 4�5 5'������t4�5���t�05 �������l��?����t�0	5�������l��@���t�#)����t�#*����m�!+������a��u5G5S��������a�	R����a5_5i5p������i�	����a�	�������i�
������k�p5�5�5�a5�5���������e�3 ��n�$��������e5�5��������n�Z��d��p5�5��e����o5�5�����s�"Px5�5�����l�"H5�������e�"R�����������l�"Er66*6.6[��a66!������n�1������n�1�c�#i646B����������g���g� �6K6S����e������w���w6o6v6�797k7�7�8���h�!�d6~6�6���h6�6�6�6����n�!����t�!�����t�!��p�!��l6�6�6�6�6����h�!����n�!����t�!�����t�!��p�!���n�!�6�6�6����t�!�����t�!�����e�!�h6�70��d7	777(������d��������d���������d������d�������x������t�!�7F7W7c��l�!�7N�����e�!���������t�!�����e�!�����t�!�7{7�7�7���������e�!�����y�'��������t�!�����e�!���b7�7����t�!�����t�!��p�!�7�7�7�7�d7�7�n�!�7���e�!�������e�!����t�!�7������n�!�����t�!�����e�!������x���s88e8�8�8�c88S�i8&8=�����m� ^81��������e��>����e� ~8G��������e��^���t�Q8\�����d�R���l8n8y�������a�0A�������a�0�8���������h��g����s8�8�k� *8�8�8�a8�8�����������c�m����c�mm8�8���h�"�������e��
����l��am� B������r�������������������l�"Ct� @999"9*���e� ���������e�� ����l��k����d�Pu9@9Y9`9y9�9�b9F9O�����i�	�������o�1 ���a�	�u9g9p�����i�
������i�
����������������i�	�������������i�
L��������n9�9�9�������i�	����a�	L�������i�
�����������a�	=y9�9���������n�a�n��9�:�����������w�� �����w��b� b:.:�:�:�:�<<I<�>H>T>>�>�@@'@0a:>:H:`:g:�:�:�������i�	�������h� \:T��������e��<���a�	,�u:n:w�����i�
������i�
,h:�:�������a�0p����i�?�������a�0�r� |:���������e��\�������o�1�����e�$���t:�:������t�����w�e:�;;;�;�;������������������s�&lc;;���e�"5������c�1h;(;1;?;];������c�(����������c���i;E;T�����������c��������a�0y�e;d;q���������c�����i;y;������������c���������������c����������������c��m�������a�0���������n�bt��;�;�;�;�a��;�����������k�������h��1;������w��1�����w�����������w��Lh<<Ca<<#<*������i�	����a�	-�u<1<:�����i�
������i�
-��k�Si<U<`<k<y<��������a�0s�������a�0�����������k������������i�
�������e�31l<�>7>Ba<�>2�k<�<�<�=r=�=������e�%�d<�<������d�%�������������������e�%�l<�=Je<�=���������g<�=������r�%��������e�%���������������t=!=5���t�0=*�������l��;����t�0=?�������l��<���r=S=b�����������e�%�������������e�%�r=x=��������e�%������������g=�=�������r�%��������e�%�s=�=�=�m=�=���������e�%���������e�&;����e�%���r�&��p=�>�r=�=������������e�%�������������e�%�������g>>'������������e�%��������e�%��k�$#�������w���k�%���������e��Bo>\>i>t���������i��������a�0|�������a�0�����n�$�������e�3�r>�?�?�@�c>�?8e>�>�>��x������t� {>�>�>�>�>��t���m>�>��d����������e��[����l��[�p����������l��7����t� }??
? ?(?-�t���m??�d����������e��]����l��\�p����������l��8��t?@?j���t� [?O?T?Y?e�t����x�����������e��;�p�������t� ]?z??�?��t����x�����������e��=�p�����e��?�?�?��������b�.��b��������d?�?�?��������b�/��b���������b�a���e?�?��������b�*���������������b�:������r� �s@@����e��������r��������r��u@8@C@N�������a�0v�������a�0��l@U@s�t� "@^@h������e�%��������r�"���e�%�c� c@�AiAtA�A�B0C�D�E+E\HTH\HfHrH�a	@�@�@�@�@�@�@�A*A3�������n�n������i�	����e����a�	�u@�@������i�
������i�
������e�3���������uAAAA������i�	���b����a�	�������i�
������k�!�rA;AAA[��f�!�n��AJAU�������b�,��b�����������n�!��������o�1cA~A�A�A����n������a� �A�����e�	��cA�A��e�$������x�	��l�UdA�A��t�A������t������e�3�eA�A�����a� �A���b�'�t� �A�BBB%iA�B����e�!������r�����������e����������e����������r���hB<B{B�C>C�aBFBQB[Bb�������n�y������i�	����a�	�uBiBr�����i�
������i�
�������o�1eB�B�B�CCC%����������������c��cB�B�����k�'������c�GdB�B��������rB�B�����������������c���������c����������������c����������n�s�����������������c�����������������������c��i��CD���hCQCtC�C�aCWCf�����������n�2w����������n�2�����������n�2i�����n�1J����������n�2	oC�C��hC�C�C��nC�C�����i�
���i�������i�	�����i��k��iC�DC��cC�DDD&D4aC�D �����������n�2v����������n�2�����������n�2h�����n�1H����������n�2�����������n�2�cDJD��e�%�DWDbDgD�������y�"��t�"�pDmDs��s�"���������k�06���hD�D�������������k�%��������������k�%������x��D�D��������b�-��b�lD�D�E��r�#'��kD�D�D�D��������r�������l��������l����������x���b�&cE���tEE#����k�&c����e�&gmE3EAEL����������e�3��������e��C������������e�3�oEnEyE�F�G�G�H=HF�������n����n� :E�E�E���nE�E�����y� ������e��sE�E���n� ����l��U���������rE�E�������d����d��mE�F��a� ,E�F'F2F>F\FsaE�F	F���eE�E���b��������b�����t���rFF���c������n�]�������r�����������e���������dFKFV�������b���d��sFbFi���l��P������r��������dF~F��������b���d�����s�&<nF�F������t�"EtF�F�����������l�".��l�#F�F�F�F�G+GXGfGkGpGuG{G�G�G���K� BF�F��L� S� CF�F��N� R� DGG!G&CGGGG1� 2� 3� 4� �L� �E� EG7G;G@GEGJM� �Q� �T� �C� TGPGTB� X� FG^GbF� S� �S� �T� 	�F� 
��K� �S� SG�G�G�G�G�I� O� G�T� �X� �B� �N� �S� �T� ������t� �G�sG�G���s������f���rG�H,���������tG�H	���t�0G�G���������h��b�������l��A����t�0HH!��������h��c�������l��B�������������e�3�����e�3�����������e�3�����n�$�������o� ���������d���rHyH��yH�H���d�"��r�"�����y� ��rH�H�H�H�����e������x�������e������x���d� dH�JnK�K�LrMDM�N;NHNQNkN�N�O�O�O�O�PaH�IIIYI�I�I�I�J1J7JU�������n�d������i�	�dII&I,I:IJ�����c�6��a�	&����������c���������������c��������������c���gIaIrI���h��Ii�����w����r�  Iz��l� !uI�I������i�
������i�
&�������a�0`�������a�0�lI�I�I������c�/�t��I�I������h��3I������w��3�����w������������c�����aI�JJ�����c�O��������c�O���aJJ)����������c�L����c�L��a�	d��aJ?JH�����w�����������w�����������������������b��bJvKsK}l	J�J�KKKK&K8KFKQ����e���aJ�J�����������tJ�J����t�0
J��������l��=����t�0J��������l��>rJ�J������������������b�+��wJ�J����t�!�����t�!�����a�	e����e���K��b��������l�",������e� K2��b�3����������b�?�������d���������lK^Kd��r� �����������b�������o�1	�����e�3�cK�K�K�K����n������a���cK�K��e�$�����������w����t�dK�LL'LZaK�K�K�L ������i�	����a�	!�uK�K������i�
������i�
!lLL�����c������������c���������a�	\�aL0L:LA������i�	����a�	"�uLHLQ�����i�
������i�
"�tLaLj�����t�����w�eL�L�L�L�L�L�MM?cL�L�������������rL�L������c�k������n�k������c�4���e� ��iL�L������w�������a�0g������c���������a�0�lL�M��eL�M���t�#+����t�#&�a��M�����d����������������������������������i�	��h��hMJM|aMRM\Mc������i�	����a�	'�uMjMs�����i�
������i�
'��k�WiM�M�M�NNNaM�M�����������s��M���b�D���d�&fM���������e�&b�����s� �M�M�M�M�M�����e����������b�$��b�����e�������s���������a�0b�������a�0�������k�0�iN$N/�e� �N+s�"#��������h�"���������c�R�����e�%�lNWNb�������w������e�3�mNqNy����n��������e��D�����k�%�o
N�N�N�N�N�OOO'O�O���������i�������i��������a�0i�������a�0����r� $N�N�N�O �������r�����������e���������e��$sOO���l��i������r����g� ��������e�3&tO5OFO\OgO�O������t��O@��b������cOQOV�b�#��b�#�������a�0����sOpOti�1j���Oz���������k�����h�"���������e�%������������h��O������w�������kO�O��������b���d������n�$��������r���tO�O���l�V����r��uO�P�������a�0e�������a�0�z��PP(P;P`�����e��cP.P5���n����l��ePAPU����������������c���������c�U���������c�_e� eP�P�P�Q�Q�RR%R<RqS�TT�T�U|U�U�V$VYWW�W�W�X8aP�P����e� ���h�&AbP�P�P������i�	�������o�1���e�cP�Q)Q7QWQ�aP�Q#���aP�P�Q���a�	�������i�
���������nQQ���a�	E�������i�
���n�����������e�hQ=QH�������n�e�����������n����cQ_Qd�e�$������x� �QyQ�Q�Q�Q�Q�����e������w��������w������e����������e������e��������c�TdQ�Q�Q�Q�������e���a�	������s� ��t�Q�Q������t�����w��eQ�R	�������i�
������������i�
G��������c�DgR+R2���e� �������i�
�hRFRQR\Rf�������n�g�������o�1������a�0H�������e��iR{R�S�S��������o�1��t� 8R�R�R�R�R�SSSLSnSzS�S�S�S������c�h������i�	������e�$gR����������������f�'����a�	n��nR�R������e�$qpR�R����n�$�����d�$��uSS�����i�
������i�
nhS%S?aS+S6�������c�h�����u�0(���������d�&kiSRSd��������������n�2'������r� ���������e���������e��8pS�S����n�${�rS�S���d�$����n������n�!w�������r� x���i�X�����������e���������������c�ekS�S�������a�0�S���������h��toTT�����������i�
t���n�1TlT#T.Tk�������c�;eT4T;���t�"��nTETNTc�����e�$jpTTT[���n�$~����d�$�����n�!z�����s� &Tv�������l�"�mT�T�T�T�T�����n�T�T�����e�����e��������c�<���h� T��������l��1�������e��EpT�T�����������������n�[����t�"nUUUUEUeUt�������o�1#�������c�=dUU2��h� U'�������l��2���������������c��g�KUMUX�������o�1%���������c�������������c������e� oU�U�U�����k������n�1S��n�[U�U������d���������d�\U�U������d�^���k�]pU�U����n�$�����n��U�����s���uU�V�l� =U�V��������e��sVV���l��f������r� |�������e�"arV,V7VB�������o�1&�������c�@������d�XVN�������c�MsVgVrV�V�WW�������c�A����������������c��h��V�V�V�V����l����tV�V����a�	������������a�	F�����������p��������������d�����lV�V��������a�0G�������a�0�V���������h��j������d�!.������r���tW$W>WBWSW�a��W,W6������n�h����s��h� ����e��WK����w�����aW_WW�����hWiWr�����w�����������w�������w�����������w������d��uW�W������n�1a�o� ���������nW�W�W�������i�	����a�	G�������i�
�xW�X,���m� !W�W�XX$�������n�\dXX�l� <��n� �X����l�����������e������l��!��������l�"�h��XCXVXacXIXP���n����l���������d�����l��f� fX�X�X�X�X�Y]Ym[u[�[�]!])aX�X�X�X����a�	^�������i�
^�������t�!	��aX�X�X������c�N��������c�N��������c�K�������o�1�����e�$���������t�eX�YLYVhYYY-Y=�rYY���c�A�����n������������c���������������c��������������c���������c�����e�&@f�� YeYii��l��i��Y�Y�Y�Y�ZDZUZ]Zj����nY�Y������e�$npY�Y����n�$�����d�$��������h� ���dY�Y���x�%����t�%���lY�Y�ZZ!Z1��f��Y�Y������h��:Y������w��:�����w����m��Z�����w����n��Z�����w���e��Z(�����w������i��Z;�����w���������������e������e�%����������c�s�e� 5Z�Z�Z�Z�Z�Z�Z�[[#[/[:[[[c[n�����c�e������i�	������e�$dZ����������������f�'����a�	k������s�!]�uZ�Z������i�
������i�
k�aZ�Z��������c�e�����u�0%i[[��������������n�2$������r� ���������e���������e��5p[@[G���n�$x�r[N[T��d�$����n������n�!t�������r� u���i�Ul��[{���n��m[�[��������e��F�����e�3�o[�[�[�[��a[�[�����i����i���������i�O���l�" �r� 4[�[�\\!\(\A\\\~\�\�\�\�\�\������c�d������i�	������e�$c\���������������f�'����a�	j�u\/\8�����i�
������i�
j�a\H\S�������c�d�����u�0$i\b\t��������������n�2#������r� ���������e�����������������i�	��������e��4p\�\����n�$w�r\�\���d�$����n������n�!s�������r� tt\�]��n\�\������e�$mp\�] ���n�$�����d�$�h]]�i�T����������e������n�$��a]0]8����n� D�c� �g� g]a^+^B^^�_A`:`�`�aa'aCaYb"b8b�a	]u]]�]�]�]�]�]�^������i�	����e�����a�	f]�]�]�]������c������������c���������������c��������������c����u]�]������i�
������i�
�������a�0L�������a�0���a��^^���������l�c�������r�����������c��b^1^;������o�1���e�c^L^S^\^r���n�������a�#��c^d^i�e�$������x����������t�#��t�!^������t�!e^�^�^�^�^�_8�������c�3�������a�0R�������a�0����������������l�"Qr^�__��h^�^�^������������w�������w�������������w��������s� ������m_ _/�����������w�������w�������k�0h_M_�``*`0a_W_a_x_�������i�	�d_g_r�������n�r��a�	�u__������i�
������i�
�n_�_�_�_������c�:����������c���������������c��������������c���e_�_�` �����������������c���������������c���������������c���a``���a�	Z�������i�
Z��k�`������e�3�i`B`M`X�������a�0N�������a�0�m`^`i�������n�c�l��`r`������h��2`}�����w��2�����w�����������c�S�����l`�`��������������e�����p��`�`�`�`��������d����d���������d��`�`���d���������r�������e��a�������d��maa����n�!�������e��Goa-a8�������a�0T�������a�0��aaJaP��n�$������e�3�ra_a�aaeam����t�"�e� `a~a�a�a�a�a��������b�ca�a��b� ��b� ���a�	S�����d����������e��@������b�@����r� >a�a�a�b����l�"ea������s�"���������e��oa�bra�b���������t�"s���s�"w�������l�"g����l��esb(b0����t�a����e��ubBbMb�b��������a�0P�lbTbm����tb^be���t� �����t� �����lbwb~���t� 9����t� :�������a�0����������e�3������e�3�h� hb�eZe}e�e�gZgnhKhWhci�i�i�i�jjab�ccc7cPc�c�c�c�c�c�d6d?ab�c���������������c������������c��������i�	��ec c2��������������c���a�	9�uc>cG�����i�
������i�
9hcZcccqc������c�-����������c���icwc������������c��������a�0o�����������c�����������e�3*�������a�0�c���������h��������������i�
M��ac�c������c�!��������c�!���������r�1drdd������������c�J���ndd(���������p�!�����������p�!������e�3���fdId�e ����h��d]dbdpdyd�d��6��2dhdl3��f�������w�������������w��������������w�����������w�������s��d�d�d�d�d�d�d�b���8���4�������w�������������w��������������w�����������w������l��eee e%e.e=eM�7���4���0�������w�������������w��������������w�����������w��bebegeq�r�'������o�1��������w�+ce�e������a�)��ce�e��e�$������x�%de�e�������s�'�te�e������t�#����w�%e��e�e�ff�gg5g>gK��t�&ee����te�e�����k�&e����e�&a�����h��4f
�����w��4hf!f=fEfwf�f�af'f5����������c������c�G����w�������afPfo�tfWfc��������c�����������c�������c������������ef�f�����������c����������������c���if�f�������af�f�����������c�������c��������a�0x������af�f�����������c�������c���������������e�3{kgg&������a�0�g��������h��������������e�36�����k�g���������e�39t��gQ�����w�����k�fgc�������r��igxg�g�g���hg�g�g�g�ag�g������������n�2{����������n�2�����������n�2m�����n�1N����������n�2�������a�0r�������a�0�g���������h�����q��hhhhh.h>�4��2hh1��d�������w�������������w��������������w�����������w����������w����������e��Ho	hwh�h�h�iiini�i��������n�p�ih�h�����i�+�����a�0{�������a�0�h���������h�����m��h�h�h�h�h�h�h��9���6���2�������w�������������w��������������w�����������w�����������i�.oiidki(i4i:iP��������b�	��b�	������������������b�!����������������b�"������e�3Briti�iizi������c����������r� ���b��������s�&h��e�#����n�$��������r�������d�eui�i�i�i��������a�0u���������e�33�������a�0�i���������h������������t��j��b�v������n� -j'j2j>jU�������r�����������e��sjDjK���l��c������r�����o� i� ij�j�j�j�n{n�oo3o�o�o�ppiqqYqaqnq�q�rrF�cj�j���e� �������c�Obj�j�j������i�	�������o�1'���e�-cj�j�j����n����cj�j��e�$������x� �������c�Vdj�knPnq������e�	eknK�����hk k.k;m�nn n,����������e�2����������e�2��ckZkjk�llElblrl�l�l�mmFm�m�������������n�2?cktkk�k��������n�2:����������e�2����e�0ok�k�k���a�0k����t��d����������������n�27����������e�2�ek�k�k���������n�2/�������������n�2=�������������e�2�fl	l�����������n�2@ill;������ll*l3�����e�2�����n�26������n�2+hlKlV�������n�22��������e�2�������������k�0llzl�l����rl�l������e�2�����n�28��������e�2��������e�2�ml�l�el�l������������e�2��������n�2.�������n�2*��������n�24pl�l�����d�0���������e�2�rm	m9emmm+�������n�2C�����������n�29����������n�2>���������e�2�smRmom}m�m�emXme���������e�2�������n�2B����������n�23pm�m���e�0 ���������n�25tm�m��������n�21�������n�2;um�m������n�20�����������n�2<wm�m���������n�2,�������n�2-���o�0mm�n���������e�2���������e�2����������e�2���������e�2�wn2n?���������e�2���������e�2��a�	������s� �n^nf����e�/�������c��������w��en�n�n�������������c���������c�5��gn�n�n�n�an�n������������n�2u����������n�2�����������n�2g�����n�1G����������n�2gn�o ���e� �uoo�����i�
������i�
hoo(������a�0D�������e��ioEoOoZoaozo�o�o�������i�	��������c�8���a�	�uohoq�����i�
������i�
������������i�
@�����������e�������������c�9��������no�o�o�������i�	����a�	@�������i�
�j�3ko�o�������a�0�o���������h��r����n�1clpp
�e���������w��mpp^ap#p7pP���n�+p,�������c�����������������������l�"S����������i�
?�������e��Inpupp�p�p�������t�"�����y�"��������n�ktp�p�ep�p����l�"+p�p�p�bp�p�����m�#!t�#!�x���tp�p��p�# p�# �������n�")������e�3vp�p�q�����t�%������e�%���������e�&;oqq!q)�������c�Q����k�/�a��q4qIqQ�������s��qA����s������n�i����s������n�$����������i�
rsqxq�q�q����lq�q��������a�0C�������a�0�q���������h��h����������i�	�����e�h������r���tq�q�������nq�q��������a�0��������a�0����e�)q�����w�-urr�������o�1)�������c�N��������nr*r4r;������i�	����a�	?�������i�
������arQr\�������c�u���������������c�wj� jr�r�r�sss�s�s�s�s�ar�r�r�r��������n�q������i�	����a�	�ur�r������i�
������i�
�������o�1cr�r�r����n����cr�r��e�$������x�5���������l��������������e�_ess&sg�������c�X�ms1s:sHsX�����c�,����������c���������������c��������������c���hsmsv�����c������������c���hs�s�as�s�s�������i�	����a�	�us�s������i�
������i�
���������n�{�s�0��������e��J����n�$��������r��k� ktvnvyv�v�ww*x�yZygy�y�z<zRz_zvz�z�at/tOtet�t�uu,uEu�u�v8vUbt5tF�������������c�������i�	�ctUt[��e�1������c�:�etlt~��������������c���a�	f��t�t�t�t�t�t�t������c�C�����h��;t������w��;����������c��������w��������������c��������������c������������w��M�ut�u�����i�
������i�
huu������a�0K����������c���������a�0�u9��������h��vpuKu`�a��uR����������k������nuluzu�����������n�1qpu�u������������n�1����������n�1x���������������n�1y����������e�3su�u�vvv(�������ou�u������c�@������������������c�@�����������a�0�����e�3��avv�����c�P��������c�M������������c���������������������������h��p���������������������c���������o�1cv�v�v�v�av�v�������e�3���n�������a�7����e�$����������t�7�������w�3ev�v�w whv�v��������n��������a�0Q�������a�0�v���������h��y��������n�o������������a�0�����������c�8hw8w�w�w�x4x�awDwNwYw`wy������i�	��������c�E���a�	�uwgwp�����i�
������i�
hw�w�w�w������c�.����������c���������������c��������������c����������c���aw�w����a�	Y�������i�
Y����hw�xxx&aw�x �����������n�2x����������n�2�����������n�2j�����n�1K����������n�2
ox>xoxyx~�hxIxRx[xe�����i������i�������i�������i�������i�[�k������������i�������e�3�ix�x�x�x��������a�0M�������a�0�x���������h��w�ox�x�x������������e�3������������e�3�����e�3���kyy'y6y?yMay
y�����������n�2n����������n�2�����������n�2`�����n�11����������n�2 ���������n�13���������c�\lymyx�������w�5�����e�3�my�y�y�����������e�3��������e��K������������e�3�oy�y�y�z
zhy�y�������a�0S������e�3��ay�y�����i������a�0�y���������h��z��������e�3����������c��rzz2����������������l�2������b�C�azCzI��n�$������e�3����������c�otzezn�����e�3�����d��uz|z��������a�0O�������a�0�z���������h��x������e�3�������e�3�l� lz�|�}}V}|~~~-~E~W~�~�}�����az�z�z�{{{-|�������i�	����e�:���a�	2�u{{�����i�
������i�
2������������i�Em
{C|||=|K|^|n|�|�|�a{I{���f{U{c{�{�����������c�������a{m{�����e{w{�����������c����������������c�������w{�{�����������c����������������c����������������c������������e{�{�����������c����������������c�������c�D��a��|�����e���d��| |4�����h��<|+�����w��<�����w������������c������������������c���������������c�������������������c�������������������c����������������������c����e|�|����������c����m|�|����������������c���������������c�����������e�%�b|�}}
�r����t�l������o�1c}}%}.}I���n�>�����a�<��c}6};�e�$�����������w�=���������t�<��t�@}`}i�����t�@����w�7}s�����n�9e}�}�~�t}�}�������������b������������b��s� <}�}�}�~����l�"d}���������r�"���������e��o}�}�r}�}����������t�"r������r�"v�������l�"f����l��d�h�n�����k�%�������������x�mi~3~8�a� ����������n�lj��~K��������c�Yl���~c~{~�~�a~i~p���a�	3�������i�
��������w�;�����a�	4������c~�~�~�������i�	����a�	a��������n~�~�������i�	����a�	cm~�~�~����������e�k�������e��L�����e�3�o:EKu��������i�,����l"5��d�"'��t� �*�������d�#�r�"(�������i�%��s�����eUlc[g��������e��N�b�2�����d��M����e�%�����n�$�s������h�B����e�!������r��������e�%�����i�&������c���������i�	����a�	��������n��������i�	����a�	b������e�3�m� m�#�����Ă݄�(�_�}����/�H�Q�l��a�=�G�������ׂ3�L�Q�_�k�p������i�	�c�M����n� ��[�f�l�u�������b�1��b������d����������e�����e�?���a�	.�u���������i�
������i�
.h��������h���������w�����������w��������a�0~i��(�g���'�������a�����w����������i�����������i������i�K������������i����k�1�P�W��w�9�D�������i�����������i������i�H������������i���������t�s�~�������i������i�1t����������u�����������i������i�G�o���с���w�����������i�����������i������i�I������������i����i�����w����������i�����������i������i�J������������i�����������i�F�������a�0ނ@��������h����e�&B����������e�3G��������w���s�&Bs�v����������������w������e�3�b����������o�1�����e�3�c��������e�$����������e�3���t�̂������t�A����w�Ce��l�w�����ă�e��_m�����$�����c�E����������c���������������c����e�+�8���������c�����i�@�O�����������c���������������c��H���������e�3M�������a�0������������e�3~�������a�0დ��������h���m�ރ��������h��>�������w��>�����w����������n�t���a�ۃ������w�������a��������w�����������w�����������w��h����k�q������e�3�i�6�[����A�d�=�V���������������������h��e�t� ���m�i��������a�o�~�����������n�2r����������n�2�����������n�2d�����n�1Ap����a��������������n�1p��������n�2���������n�1n���������n�1o�������a�0�������a�0߄���������h����u��<s�"��&�/�5�������b� �����e�"���d�����s�"�e� 2�i�H�V����������e�3J�����e�3Il�e�t�����������d�p�����e�3�m����������������e�3��������e��M������������e�3�o���ԅ��� h����������a�0�������e�3��������a�0����������h���������e�3������i�!���������e�3��������e�3��a� �&��n�$������e�3�s�5�>�����e�3�������r��������d�ou� ��o�s�}���������ن�����X�b1� �������e�3��h����������r�"k���s�"j������e�3�g�������k�������e�3��������a�0��������a�0�����������h���l�߆������e�3�����y� �������e�3���h�������w�����������w��s��O�c�'�8�C�����e�&j�2��l�&k�������n�&m��������n�&o�����e�3�������e�3�������e�3�v�r����������e�3������e�3�w�������������e�3������e�3�n� n�ԈZ�r���͉��T������̋��F�4�<�U�]�=�G�Qa������!�,�E�Qb��������i�	��a�"���e�D���a�	(�u�������i�
������i�
(�������a�0j�������a�0ʈ9��������h�����������e�I�����e�3�b�`�j������o�1����e� �c�|���������n�H�����a�F��c�����e�$�����������w�K���������t�F��t���������t�E����w�Ge�Ո����������a�0m�������a�0͈���������h�������������n� �������e�3�g��Ia��)�0������i�	����a�	�u�7�@�����i�
������i�
�������i�h�Z�d������a�0���k�l�s���t�r��������x�si���2�=�w��n�����މ����#a���������������n�2o����������n�2�i�ŉ���������n�15���������n�2a����������n�16�����n�14�a���
����������n�1h��������n�2���������n�1g�����������n�1f�������a�0kk�C�[������a�0ˊO��������h�������t�e�p�������i������i�M�e� 9�������ǊΊ��$�0�;�\�d�o�����c�i������i�	������e�$h�����������������f�'����a�	o�u�Պ������i�
������i�
o�a����������c�i�����u�0)i����������������n�2(������r� ���������e���������e��9p�A�H���n�$|�r�O�U��d�$����n������n�!x�������r� yt�u����n�}�������e�$rp�������n�$�����d�$���i�Yj�̋���������c�Z�������a�0����������h���l�ҋ�����������g���������w�Im����������e��N�����e�3�n��=a���$������i�	����a�	#�u�+�4�����i�
������i�
#�����a�	)o�T�_�x���q�(�������a�0n�������a�0Όl��������h���n������������������e� ������i�����i��n�����Ɍ���$�_�����c�F����������c��������a�Ԍ������c������������c���������������c�������i�������������c���������������c��K�e�+�8���������c�����i�@�O�����������c���������������c��N��������������c���t�������̍؍��������s�"e���������t�"	���f�"	���l�"`������r�"o����r��������l�"q���s�"y��������l�"b���s�"n���������l�"pp���������l�"&������s�"��u������t�"������s�"������t�"���������n�v����n�$�s�B�K�����e�3�������r� ����e� �u���i�t�ŏ�������a�0lk�z��������a�0̎���������h����a������������i�	����a�	<�u���������i�
������i�
<m�ˎ�������n� #�َ���������e������l��_�r�������n�������k�t���������k�uo�!n��� �4�����h��@�+�����w��@�����w��������e�3�������e�3��a�Z�d�k������i�	����a�	�u�r�{�����i�
������i�
o� o���Đ�����;���ˑ������H�i����G�Sa�������e� ������i�-b�Ώ�������d�u�ڏ��������c�����������������c�������i�	�������o�1���e�Oc��c��a� �]���a�+�2�=���a�	�������i�
���������n�K�R���a�	I�������i�
���n����c�k�p�e�$������x� ���������������e���������w������e����������e������e��������c�>d�Ɛݐ���l�͐�����e�Q����e���a�	������s� ����������c��������w��e�S�
�����n�1Zg��*�1���k�ۑ$��b�(���e� �������i�
�h�E�P�Z���������n��������a�0Jo�`�j������e���n���y������������e���������w������e����������e������e������������t�Qi���������������e�k�ё�������a�0�����������h��u����n�1W�������w��m�
�&�-����������n�M������e�S����e�Q���a�	P��a�ɒ=�A�L�Z�j1���������c�a����������d�w������������c�{t�p������������c�}���s���������i�
�����n��������s���������e��O�e� 1�Ւޒ���(�1�J�l���������ٓ��������c�a������i�	������e�$`�����������������f�'�d����a�	g���������r� $�����h�![�����d����u�8�A�����i�
������i�
g�a�S�^�c�������c�a�f� ������u�0!i�r����������������n�2 ������r� ���������e�����������������i�	��������e��1p�������n�$t�r�̓���d�$����n��������r� �����n�!p�������r� ��h����i�Q��d�!So��2�Bg��(���k�������n��������i�
������������i�
K��n�Tp�P�W�b���n�$��������t�%����n�#%r�o��d�u���������e� ���������e� ��������l�"s���Ôԕ����t�������a�	������������a�	J���h� �������e�����l�ݔ��������a�0I�������a�0�����������h��k���������e��������r���t��)�������c����e� ��4�<����e�M�������s�O��������o�1!v�Y���r�`�����e� >�m����c�s���������e��J�b�d��������d��I�����y��L���y��K����e� ��������n���Õ�������i�	����a�	K�������i�
�p� p���{�������P�Z�R�e���ٝ\�d��<�X�ba��9�C�J�Q���������Ԗ���oa��+��������e�3�����������e�3+������i�	����e�U���a�	*g�W�ie�]�d���n�!��p�!�u�o�x�����i�
������i�
*�������a�0q����������i�/�������a�0�l�������������������������b��������������c������������n�1r�����a�������h� ����l�"%�n��t���t� (��,�1�6�A�M�d�i�����������c��>�t����x����������r� ���������e��s�S�Z���l��Y������r� }�p����������l��5����t� )�������������ӗ������������c��?�t����x����������r� ���������e��	s�����l��Z������r� ~�p����������l��6�������f�"s�����������w����������w������e�3���h���'�5�:�C�R�b1�-�11��d���a�������w�������������w��������������w�����������w����������w���������o�1�����e�$���������t�We�䘱���Иܘ�V�a�v�I�������c�?�����h��D�������w��D��������e�3;����������������w��Ch�����)�G�r��
���c�~�����n�z����w������������c��Wi�/�>�����������c��X�����a�0z�����������c��Y�������a�0������������������c��r�������1�>��������w��N���t� %�����������c�j��������e������l��ji����d� .�ϙڙ�����������n���������d� ���������h��a�������r�����������e��s�����l��R������r�����������������b�B���������r�"��������d� 0���a� �������e�3�h�b���a�j�t�{������i�	����a�	+�u���������i�
������i�
+i�ƚ�������1�����h���֚��a���������������n�2z����������n�2�����������n�2l�����n�1M����������n�2����n�x�������i�:����������k��o�%�*�D�k���h�1�:�����i�������i�����������i� i���`�4�?�J�X��p�p�����ϛݜa�v�������������n�2s����������n�2�i������������n�1v���������n�2ek��������������n�1r����n�1B����������n�2���s��k�������������n�1t����n�1D�����������n�1ut��&�����������n�1w����������n�1s�������a�0t�������a�0�����������k�����������n����s� +�s�~�����������b������e�"�m�������s� �o����d��������e��s�������l��b������r� zm�Ŝ��������e��P�����e�3�o���3�>�H�������a�0}����������x����)��������e�&��������e�&���������e�&������e�&�������a�0�������i��������k�0�U���e�0 ����n�$�r�l����e�r�z����s�"z��������n�!��e������d���������d� 5o�����������t�"������e�#���������a�0�p�͝�e�ӝ����r�#��u������t�"������t�"������n�"7���l�"s��3i�Ȟ��������c�q��������������������b�������e�3�u�B�M�������a�0w�������a�0�������e�3�������e�3�q� q�������ş̟؟��a�����០d������a�	X�������w��f�����������c�B����������c���������������c��������������c������s��������$�-�<��1� ��0��a��c��2��7��9���3���e�������w�������������w��q�B�����n�O�X�g�w�����w�������������w��������������w�����������w�������������w�����������w���������������w���������o�1�����e�$����k����������e��Q�f���������h��G�������w��G�����w������n�$�u���u����������e�&i���s���1�6�;�@�I�X�h�8���5���1�������w�������������w��������������w�����������w�������n� ?�����������r�������c������n�^���n� �������l�������k�~��������e������l��?��e�ء�3�P��l� "���������e� ���t� ��������e������e�0��������d�0����t� ���t� �(�������d� r�9�C������d� ���t� �Ln�I����l�Z�a���e� e� '�g��������e��r� r�������ף
��3�����٦��#�ŧЧ�Wa�����ơ͢��7�B�[�r���������n�|������i�	����e�Ud�סݡ���a�	0���l�"���x�������������e�3���������e�3������e�3��e��������w���u�%�.�����i�
������i�
0�������a�0��������a�0�O��������h����������������������i�	�m�x���������������������i�	�����n�d��o�"6�������o�1c�����¢����n�Y�����a�W����e�$����������t�Wd�ݢ�������e��t��������t�Y����w�[������n�]e��E�h������f��+���������k� ;����u�5�<���t�"������t�"������r�P�U�d� �s�[�a��s������f���h�p�����r�w�~���c�1�����n������������c���������a�0��������a�0죬��������h����h����������������w��H�����w��v������������e�"=�a���������w��������������w�����������t�#�������k�~�(�������d�h�9�Pa�?�I������i�	����a�	]o���Z�w���k�}�a�����d�{�l�������r������������k�����������d��i���̥�������l	���٤���$�2������a���������������n�2q����������n�2�����������n�2c����������n�1@k�������k�������n�1:���������n�1i����n�19����������n�1;p�:�Z�ia�@�N����������n�1l��������n�2�����������n�1?���p�r�{�����n�1<���������n�1k���������n�1=t���������������n�1>����������n�1j����������������n�1m��t�ԥ�����e�"t�������������b�������e�"��������a�0��������a�0���������h���n�$��g�ڦ.�9�?�������b�%��b�
���f�H�v���t���U�`�k�������n�Y�������b��������d������t�������������b�9�������d������������e�����������e�3Ql�����������w�_�����g�|�������d�z��������e��Ro�����������a�0��������a�0���������h���������i�#����n�$�r�+�O�ma�3�=�D������i�	����a�	1�������i�
\�h�V�_�����c������������c���������c�}������������i�	����a�	`�������i�
���������n������������i�	����a�	D�������i�
��������r���t�֧�����k�%�����d�y���������r��u����!�P�������a�0��������a�0���������h���p�'�J�e�.�<����������i�	�����������i�	���h������i�$������c�g�q�x��������i�	����a�	�������i�
���������n������������i�	����a�	C�������i�
�s� s�٪��ƫD�k�1�<�˳U�����]�����˶��ηx��a	�����T�m�x������������i�	����e�[� ��������t�ed��!�'�5�E�����c�5��a�	8����������c���������������c��������������c����u�[�d�����i�
������i�
8�������a�0U�������a�0�����������h��{����������������������������c������h�᩼�������h��A�������w��A�����w���a��0�8�j�ra�����!�)����i�2����i�A����m���������i�D������i�C����i�3���i�0����i�@i�@�X�ci�F�Q�������i������i�5�������i������i�4����i�Bu�z����e������e�����������i������i�7�������i������i�6���i�8����i�9�������o�1c�Ҫ��!�7���n�a����������t�g�����a�_��a�Y�����������c�����������������c�����k�Z��c�)�.�e�$������x�]���������t���t�L�U�����t�a����w�c�_��������t�ie	�������Z�u���߬�������������b�<c������d� 3������������e�����n� ��n���ƫԫ������c�3����������c���������������c��������������c�����l������#�2�B�M1��3��f���c�������w�������������w��������������w���������w�����������w��h�`�k�������n�}������a�0[�������a�0�����������h��~�i��������n� ;�����������c���������e������l��T�������������a�0�����������h����t���������e�3"������e�3#��n� 7��%�/�M�T�^�w�������˭���������c�g������i�	������e�$f�:���������������f�'����a�	m������s�!^�u�e�n�����i�
������i�
m�a�~���������c�g�����u�0'i������������������n�2&������r� ���������e���������e��7p�ѭ����n�$z�r�߭���d�$����n������n�!v�������r� wt��+��n�������e�$pp��#���n�$�����d�$���i�W�������n� �h�L�2�=�K��!��a�Z�e�o�z�	�"�������n�w������i�	��������c�Hd�����a�������������c�Q����a���������c��a��������c��^����������c��`����a�ˮ������c��b��������c��_e�%���������k�%�����t�%������m�%��a�	6�u�������i�
������i�
6������������w���������o�1����������c�Ie�U�������n�`�i�w�������c�4����������c���������������c��������������c���������c����l� ��������w� ��a���¯ѯ߯���1�ȯͱ5��5��2�ׯ�2��e�������w�������������w��������������w�����������w�����������c��i�'�2�������c��n��<����d�B������h��I�N�W�����w��Is�]�q�����t��,�h�����w��,����t��-�{�����w��-�������w�������w��s���������t��*�������w��*����t��+�������w��+��k��i�ݱ	��-�K�S�`���a�ð���1������l������������������k���������a�0W�������a�0��!��������h��|��q�5�>�����w�����������w������r�"<���������w���s�o�����αܱ�a�u�������������n�2t����������n�2�i������������n�1~���������n�2fk��������������n�1z����n�1E����������n�1{p������������n�2���������n�1}�����������n�1|x� 6�)�2�<�Z�a�z�����òβ��������c�f������i�	������e�$e�G���������������f�'����a�	l�u�h�q�����i�
������i�
l�a�����������c�f�����u�0&i������������������n�2%������r� ���������e���������e��6p�Բ����n�$y�r�����d�$����n������n�!u�������r� vt��O��n��:c������e�$o������������������������i�	�p�@�G���n�$�����d�$���i�Vl�[�o��h� /�c��������e����g��w��������t��m����������e�&:�������e��So���޳��/�:f��������������w��t�Ƴ������n� ������������c�L�������a�0]�������a�0�����������h������s���������������b�8��������������b�7�������i�)s�B�L�T������i�(����i������i�*�a�f�z���e�  �m���������c�  �e�&`�����t��������k�&`����e�&d��n�$�����e���Ǵմ����(�I�d�����������b�;c�ʹ�c�3�m�3����������������������l�%��������������l�%�k��	g�3�m�3��������l�3�l��#n�3��g�3�m�2�6�;�?g�3��l�3�m�3�������d�3������������������������l�%�����r�n���������������������l�%��������������������l�%������������l�%�������������������k�%�������e�3�s�Ѷ{a�۵���������i�	����a�	7�������i�
��g�
��&�4�C�Q�_�l����������n�1I����������n�1�����������n�1������������n�12����������n�1e����������n�1C���������n�1F�����������n�18������r���t���������g� �����������e������e�����������������b�6��������������b�5u�޶����H�R�V���t�"�����������l�"�������l�"�c������s�"{����t�"�������a�0Yk�%�=������a�0��1��������h��}�������c�R������n�"n�&<�����t�"��c�n�������l�"�������l�"�������e�3��������������e�3|t� t�����չd�����F�����������9��å��a
�ͷ׷���Z�k������������i�	��k�޷����n�"����t�"����a�	$�u��������i�
������i�
$h���-�K�����c�7����������c���i�3�B�����������c��������a�0_�����������c����������������e�3}�������a�0��x��������h�������������c�@u��v�긞������s��J��h��J�������w��J�����w��b�Ƹ��r�g������o�1
c������<�W���n�e���l�������a�c��h����-�����c������������c��{������������c��|�����������c��}��c�D�I�e�$�����������w�q���������t�cd�j�t������s���t�{�������t�k����w�me	�������ɺ�"�e�j���������c�B����������������c��h�Ϲع��,�U�������c�*����������c������i��������������c���������������c��i��#�����������c��������a�0f����i�6�E�����������c���������������c��m�[�}�����a�f�o�����c�)����������c���e�������������c�����i���������������c���������������c����������������c��s�������a�0ƺ���������h���l��������e�!!������k�&���a�������������w�������������w��n�,�5�H�]�����e�$i���������������n�2)p�N�U���n�$}����d�$�����n�!y�h��t�ػt���������h��8������w��8�����w�����������c����r���������w�����������w��h�ʼb�ܽ`��<a�ֻ�� �������i�	����a�	%�u��������i�
������i�
%l�������c�0����������c����������t�,�K�R��w�4�?�������i�����������i������i�L������������i���e�j����h�t�}���������c�+����������c���������������c��������������c����e���������s�"���e�"4�a���ʼ�1������������k��i��8���h���!�*a��������������n�2y����������n�2�����������n�2k�����n�1L����������n�2����n�B�K�����e�$lp�Q�X���n�$�����d�$�o�n����������������������i��k������������i��n� ��h������a����������i�����i�������i�������i�����d�ֽ��������c�����������r��������c�l������n�l��e� 3�)�2�<�Z�a�k�������;���"�*�5�����c�c������i�	������e�$b�G���������������f�'����a�	i������s�!\�u�r�{�����i�
������i�
i�a�����������c�c�����u�0#i������������������n�2"������r� ���������e�����������������i�	��������e��3p������n�$v�r�����d�$����n���������s� �������h�������n�!r�������r� ����i�S������e�3�i�V�a���6�B�s���������a�0ak�g�������a�0��s��������h�����t��������a���������������n�2p����������n�2�����������n�2b�����n�17����������n�2��e�ܿ��� ��(�������b�0c�����b���b���������b�`o��������r�"<��������b�4����������b�>��������e�"�p�H�f��a�P�Y�����w�����������w�����������i�
p�������������b�����������n���������w�o��������e��To���������`�l���������n�i�������a�0h�������a�0�����������h���n���R�We���?�F�L��r��#�-�6����a��������d�������d��������d�������d�������d�����e����x����o���s�������e�3'��������i������������������t�������t�0��������l��]�������l��9����t�0��������l��^�������l��:������i��a������������k����n�$�r���
�������k�!"��s�����s������f��������������k����g�%�*�/�4�n�%��f�%��t�%��p�%�s���E�l������i���O�c�����h��F�Z�����w��F�����w��e�r�}�������c�F�e��¡ª¹��12��e���b�������w�������������w��������������w�����������w�����������c�[������r���t���)�jÝa���	�������i�	����a�	�u�� �����i�
������i�
�h�4�=�K�[�����c�y����������c��g������������c��h�����������c��i�a�s�}Ä������i�	����a�	 �uËÔ�����i�
������i�
 ����d��uíø���������a�0d�������a�0�����������h�������l�����������a�0c�������a�0�����������h��ow��ne��;��e���3�����e�$kp�$�+���n�$����d�$�����n�!{��y�E�N�Y�����e�$s�������u�SDp�_�f���n�$�����d�$�o� 2ĎėġĿ����'�I�U�h�sŔŜŴ�����c�b������i�	������e�$aĬ���������������f�'�d������a�	h�t�����������r� %�����r� %���������l��0�u��������i�
������i�
h�a���������c�b�����u�0"i�-�?��������������n�2!������r� ���������e�����������������i�	��������e��2p�yŀ���n�$u�rŇō��d�$����n������n�!qsŢŪ����e��������r� ��hŻ���i�R���s�!Tu� u������W���ǁǑ���
�[�d�����_�{������e� �b������r�������i�	�������o�1(���e�mc�&�-�M���n����c�5�:�e�$������x� ��E����w�w������c�Cd�c�nƅƋ���������a�	Q�l�u�}����e�q����e���a�		������s� �ƟƧƯ��������e������w�scƵƼ���n��������c������e�������n��������w��g�������e� �u���������i�
������i�
	h���f������a�0Fo��(������e���n���7�?�J�R�^����e���������w������e����������e������e������������t�q�v�������c��������������e�kǙǱǼ������a�0�ǥ��������h��s�������c�y����n�1\m����a�������n�k�����������c���������s�{����������i�
A�������e��Un��G�������e� _�#�)�5�@��l� ��������e��?�������l��3���y��Oi�M�R�n�"*�����l�" �����k�sp�p�w�Ȏ�����n�$�����k�%������������w������n��Ȝȱȹ�������s��ȩ����s������n������s�����k�����������b���d��r������������i�
s��g�os���
�7�����������c�^���l���������a�0E�������a�0��+��������h��i������t�C�N�������c���������������c������e�i�k�s����e�y����w�uuɇɑɘɱ��������i�	����a�	
�uɟɨ�����i�
������i�

������������i�
B��������n������������i�	����a�	B�������i�
���������n����������i�	����a�	A�������i�
�v� v�3������˔˛���	�m�ůa�=�D�]�h���a�	5�u�K�T�����i�
������i�
5�������a�0�v���tʏʯʻ�����h��5ʁʆ�5��5�����w��5hʕʝ����w�����m��Kʦ�����w��K��������w����������w�������e�$��������w�e�����4�?�Eˈ�������c�2h�����%�����c������������c��k������������c��l�����������c��m�������a�0���s�&@�����l�P�V��r� |���e�c�n�y˂�������b��������b�)�����d����d����������n�~���k��iˣˮ���������a�0����a˹����������i�	����a�	M�������i�
�����a������������i�	����a�	�������i�
���������e��Vo���b�������n�x���d�%�I��������n�3�>�������a�0��������a�0��������a�0��V��������h����������a�0�����n�$�t�{̂���e�}����d��u̛̐�������a�0��������a�0�w� w��ͱͻ�����=�E�(�Q�]Шаз����a����������<�H�l���e��������n�1Y�������a�0�k���������a�0����������h�������n�1X����l�&�1�������a�0��������a�0���������e�3Wv�N�V����h�0������������������l��4w�t�}͋�����c�H����������c������������e͚ͣ�����c�$����������c���������e�3����c�����e�$������x�ud����������s���t���������t������w��e����3�������a�0���������s�!k�!�+������a�0�����n�1^������n�1]����e�����e�Z�cη��eϒ���������t�%�c�i�}����e�%��s������e�%������������tΎ΢���t�0Η�������l��C����t�0ά�������l��Ddν�������d�%�����������������������������d�%�����������g���������������e�%��������e�%��e��B���������g�'�7������������e�%��������e�%���������������t�V�]���t�0����t�0������������g�wχ������������e�%��������e�%�sϚϸ��mϠϬ��������e�%���������e�&:����e�%���r�&t�����������e�&������������������t�������t�0����t�0���������g��������������e�%��������e�%�i�.�9�������a�0�k�?�I������a�0�����n�1_��������e��Wo�g�rЋН�������a�0��������a�0����������h��fn� �Б��������e����������i�'����n�$����g���������r�������d����n��x� x��������!�.�2�>�F�������b�=�������o�1�����e�$�d��������s���������t�����������n�mi����������e��X����n�$��������r��y� y�s�J�a҉�g�oԀ�������������aыїѡѨѯѹ�������>��������e�3N������i�	����e� ����a�	/������n�1R�u���������i�
������i�
/�������a�0�k����������a�0�����������h�������n�1Q���������i�N����l��%�������a�0��������a�0��2��������h��l��������c�c���c�S�X�e�$������x�wd�g�q������s� ��t�xҁ�����t������w��eҙӡӪӼ���(�[hҫҴ�����-�=�xӊ�����c�J�����eҿ�������c������������c�������������c������������e��� �������c�&����������c���������������c��������������c���������������c����e�D�Q���������c�����i�Y�h�����������c���������������c��X��������������c����������������������c�������n�1Vn� �Ӱ��������e���o���������n�1U�������������n�1�r������������o���������w�����������w����������c�K����������������c�������g�5�>�N�����n�1�������������n�1����������n�1���������w������e�����k���x����e��iԌԗԢԫԳ�������n�u�������c�W�����n�1b����g�&/���������n����������e��Yo���"�-�7�]ՋՔd������������h��9�������w��9�����w����d�������w������������w���������a�0�������n�1�k�=�U������a�0��I��������h�������n�1[����l�g�r�������a�0��������a�0����������h��n�����k��y՚տaՠժ������n�1�kհո����n�1����i�"������i�p�������n�$�����������i�z���������b�Er������g���������r��t�����e������d��u�)�4�>�d���������a�0�������n�1�k�D�\������a�0��P��������h�������n�1`s�lֻ֒��g�t��������c�k���������������c�m�����e֝֨�������c�g���������������c�i���l�����������a�0��������a�0�����������h��m�e���������n�1�������n�1��a�	�������i�	����a�	_z� z�:�B�M�xؓٶ�"�L�X�dڀڈژڡa
�P�[�b�i�t���������������n�f���e�z���a�	[�������i�
[h�~ׇו׳�����c�8����������c���iכת�����������c��������a�0V�����������c����n���������c�2����������c����������a�0���f�������������w������������w����������w����n���%�9�����h��6�0�����w��6�����w���������o�1c�U�\�r���n�~��c�d�i�e�$������x����l����t�|؂؋�����t�|����w��eءج������ٱ�������c�7dز�����������������c����������������c���������a�0\�������a�0��o� 0�
���$�=�J�U�a�l�vفو�����c�`������i�	����a�	f�u�+�4�����i�
������i�
f���������c�`�������r� ���������e���������e��0������n���������r� p���i�P����hٔٝ٩�����r�����������r� ����e� �a��hټ���������o�1e���������������n�j������������c���������c�6d������������������c����������������c��i�*�5�@�������a�0X�������a�0���������w����������w����������e��Zo�j�u�������a�0^�������a�0�����n�$�������������k�������e��uڧڲ�������a�0Z�������a�0�                                                                    � �   � � � � � � � �    c � � � � � � � � � �   � � � �   � � �                	  
m n    !"#$%&'()*+,-./                                                                    012    34567  8    9    :;    <=>      � � � ?@ABCDE    F� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                                                                        	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _                                                                     ` a b c d e f g h i j k l m n   o p q r   s t u v w x y z   {   | } ~  � � � �   � �   � � � �                                 �   �         � � � �           �       �     � � � �         � &-5?JT_hmsz������������������������������ 
(2?KV`bdfhjlnprtvxz|~�����������������������+:=@GNXgqx�������������*17>AMT[^knw~����������������
!'+4BLS_ipv}�������������� $+2<CJV`gmt}���������������")3:FXgv��������� ,:HUcw������������				 	$	6	I	Y	h	s	z	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	



"
)
7
A
H
S
c
p
|
�
�
�
�
�
�
�
�
�
�
",9ER[er���������(6CP_n|����������
%1BQZfr~���������$,4<BGLRYag                  �    &-5�JT_hmsz������������������������������ 
(2?K�`bdfhjlnprtvxz|~��������������_p}���C`JVmgt}��������������G����qg�B�� >T  �) 3 ��@ L V ^ a A^j k~���p �x � ��� iv�[�@7�V?�� )2��+:=NXx��S�L��������� �$n�����*1Mw �<3��'+"��!+�
4���� � � � � � � � � � �                             .null nonmarkingreturn notequal infinity lessequal greaterequal partialdiff summation product pi integral Omega radical approxequal Delta nonbreakingspace lozenge apple franc Gbreve gbreve Idotaccent Scedilla scedilla Cacute cacute Ccaron ccaron dcroat .notdef space exclam quotedbl numbersign dollar percent ampersand quoteright parenleft parenright asterisk plus comma hyphen period slash zero one two three four five six seven eight nine colon semicolon less equal greater question at A B C D E F G H I J K L M N O P Q R S T U V W X Y Z bracketleft backslash bracketright asciicircum underscore quoteleft a b c d e f g h i j k l m n o p q r s t u v w x y z braceleft bar braceright asciitilde exclamdown cent sterling fraction yen florin section currency quotesingle quotedblleft guillemotleft guilsinglleft guilsinglright fi fl endash dagger daggerdbl periodcentered paragraph bullet quotesinglbase quotedblbase quotedblright guillemotright ellipsis perthousand questiondown grave acute circumflex tilde macron breve dotaccent dieresis ring cedilla hungarumlaut ogonek caron emdash AE ordfeminine Lslash Oslash OE ordmasculine ae dotlessi lslash oslash oe germandbls onesuperior logicalnot mu trademark Eth onehalf plusminus Thorn onequarter divide brokenbar degree thorn threequarters twosuperior registered minus eth multiply threesuperior copyright Aacute Acircumflex Adieresis Agrave Aring Atilde Ccedilla Eacute Ecircumflex Edieresis Egrave Iacute Icircumflex Idieresis Igrave Ntilde Oacute Ocircumflex Odieresis Ograve Otilde Scaron Uacute Ucircumflex Udieresis Ugrave Yacute Ydieresis Zcaron aacute acircumflex adieresis agrave aring atilde ccedilla eacute ecircumflex edieresis egrave iacute icircumflex idieresis igrave ntilde oacute ocircumflex odieresis ograve otilde scaron uacute ucircumflex udieresis ugrave yacute ydieresis zcaron exclamsmall Hungarumlautsmall dollaroldstyle dollarsuperior ampersandsmall Acutesmall parenleftsuperior parenrightsuperior twodotenleader onedotenleader zerooldstyle oneoldstyle twooldstyle threeoldstyle fouroldstyle fiveoldstyle sixoldstyle sevenoldstyle eightoldstyle nineoldstyle commasuperior threequartersemdash periodsuperior questionsmall asuperior bsuperior centsuperior dsuperior esuperior isuperior lsuperior msuperior nsuperior osuperior rsuperior ssuperior tsuperior ff ffi ffl parenleftinferior parenrightinferior Circumflexsmall hyphensuperior Gravesmall Asmall Bsmall Csmall Dsmall Esmall Fsmall Gsmall Hsmall Ismall Jsmall Ksmall Lsmall Msmall Nsmall Osmall Psmall Qsmall Rsmall Ssmall Tsmall Usmall Vsmall Wsmall Xsmall Ysmall Zsmall colonmonetary onefitted rupiah Tildesmall exclamdownsmall centoldstyle Lslashsmall Scaronsmall Zcaronsmall Dieresissmall Brevesmall Caronsmall Dotaccentsmall Macronsmall figuredash hypheninferior Ogoneksmall Ringsmall Cedillasmall questiondownsmall oneeighth threeeighths fiveeighths seveneighths onethird twothirds zerosuperior foursuperior fivesuperior sixsuperior sevensuperior eightsuperior ninesuperior zeroinferior oneinferior twoinferior threeinferior fourinferior fiveinferior sixinferior seveninferior eightinferior nineinferior centinferior dollarinferior periodinferior commainferior Agravesmall Aacutesmall Acircumflexsmall Atildesmall Adieresissmall Aringsmall AEsmall Ccedillasmall Egravesmall Eacutesmall Ecircumflexsmall Edieresissmall Igravesmall Iacutesmall Icircumflexsmall Idieresissmall Ethsmall Ntildesmall Ogravesmall Oacutesmall Ocircumflexsmall Otildesmall Odieresissmall OEsmall Oslashsmall Ugravesmall Uacutesmall Ucircumflexsmall Udieresissmall Yacutesmall Thornsmall Ydieresissmall 001.000 001.001 001.002 001.003 Black Bold Book Light Medium Regular Roman Semibold rb      P<F      >F     �=F     8=F     �;F     �=F     �=F     �<F     JBF     aCF     JBF     �AF     �AF     �CF     DF     DF     DF     �CF     �CF     FCF     �BF     �CF     �CF      0123456789abcdef       ../sysdeps/lemon/generic/lemon.cpp !(size & 0xFFF) libc panic! In function  , file  : 
 __ensure( ) failed      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       sys_anon_allocate  0123456789abcdef      0123456789abcdef  In function  , file  : 
 __ensure( ) failed  ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!        0123456789abcdef       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    ../options/ansi/generic/stdlib-stubs.cpp *string != '+' !negative !"Not implemented" mlibc: srandom() is a no-op i == j !"decode_wtranscode() errors are not handled" mlibc: Broken mbtowc() called wc mbs max_size *mbs MLIBC_DEBUG_MALLOC mlibc (PID ?): free() on    mlibc (PID ?): malloc() returns  mlibc (PID ?): realloc() on   returns  !(reinterpret_cast<uintptr_t>(p) & (align - 1)) ../options/internal/include/mlibc/strtofp.hpp   !"hex numbers in strtofp are unsupported"       ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:348: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:365: Assertion 'fra->type == frame_type::large' failed!       ../subprojects/frigg/include/frg/slab.hpp:366: Assertion 'address == fra->address' failed! 0x   ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       strtofp strtofp strtofp strtol rand_r abort     at_quick_exit   quick_exit system mktemp        bsearch abs labs llabs ldiv lldiv mblen mbtowc wctomb   mbstowcs        wcstombs lock   posix_memalign  strtod_l              $@       �           A               �                   �@                                            @        0123456789abcdef       ../options/internal/include/mlibc/charcode.hpp nseq.it == nseq.end wseq.it == wseq.end alnum alpha blank cntrl digit graph lower print punct space upper xdigit mlibc: wctype(" ") is not supported     ../options/ansi/generic/ctype-stubs.cpp !"Not implemented"      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       promote iswctype        towlower        towupper                ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"  0123456789abcdef  mlibc: environment string "     " does not contain an equals sign (=)   ../options/ansi/generic/environment.cpp environ == vector.data() !vector.back() ../options/ansi/generic/environment.cpp:84: Assertion 'k != size_t(-1)' failed! vector.size() >= 2 && !vector.back() s != size_t(-1)    !"Environment strings need to contain an equals sign" mlibc: environment variable " " contains an equals sign %s=%s     asprintf(&string, "%s=%s", name, value) > 0 string      ../subprojects/frigg/include/frg/string.hpp:72: Assertion 'from + size <= _length' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{     ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed! lock     assign_variable unassign_variable getenv putenv setenv           0123456789abcdef       ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"    mlibc warning: File is not flushed before destruction   ../options/ansi/generic/file-io.cpp max_size    mlibc: Cannot read-write to same pipe-like stream __offset < __valid_limit __dirty_begin == __dirty_end io_size > 0 && "io_write() is expected to always write at least one byte" __offset < __buffer_size chunk __offset       __dirty_begin == __dirty_end && "update_bufmode() must only be called before performing I/O"    whence == SEEK_SET || whence == SEEK_END _type != stream_type::unknown  _bufmode != buffer_mode::unknown        _type == stream_type::pipe_like __io_offset == __dirty_begin hit io_seek() error  __offset == __valid_limit __buffer_size       mlibc warning: File is not flushed before closing       Library function fails due to missing sysdep    mlibc: sys_isatty() failed while determining whether stream is interactive      mlibc warning: Failed to flush file before exit() Illegal fopen() mode ' ' Illegal fopen() flag '       [31mmlibc: fdopen() ignores the file mode [39m        ../subprojects/frigg/include/frg/list.hpp:104: Assertion 'element' failed!      ../subprojects/frigg/include/frg/list.hpp:106: Assertion '!h(borrow).in_list' failed!   ../subprojects/frigg/include/frg/list.hpp:107: Assertion '!h(borrow).next' failed!      ../subprojects/frigg/include/frg/list.hpp:108: Assertion '!h(borrow).previous' failed!  ../subprojects/frigg/include/frg/list.hpp:79: Assertion 'h(ptr).in_list' failed!        ../subprojects/frigg/include/frg/list.hpp:164: Assertion 'it._current' failed!  ../subprojects/frigg/include/frg/list.hpp:165: Assertion 'h(it._current).in_list' failed!       ../subprojects/frigg/include/frg/list.hpp:170: Assertion '_back == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:173: Assertion 'h(traits::decay(next)).previous == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:179: Assertion 'traits::decay(_front) == it._current' failed! ../subprojects/frigg/include/frg/list.hpp:183: Assertion 'traits::decay(h(previous).next) == it._current' failed!       ../subprojects/frigg/include/frg/list.hpp:188: Assertion 'traits::decay(erased) == it._current' failed! ../subprojects/frigg/include/frg/slab.hpp:397: Assertion '!"Pointer is not part of any virtual area"' failed!   ../subprojects/frigg/include/frg/slab.hpp:403: Assertion 'address == fra->address' failed!      ../subprojects/frigg/include/frg/slab.hpp:421: Assertion 'fra->type == frame_type::slab' failed!        ../subprojects/frigg/include/frg/slab.hpp:425: Assertion 'reinterpret_cast<uintptr_t>(slb) == (address & ~(slabsize - 1))' failed!      ../subprojects/frigg/include/frg/slab.hpp:429: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:436: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:439: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/slab.hpp:508: Assertion 'address >= current->address && address < current->address + current->length' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed!       ../subprojects/frigg/include/frg/slab.hpp:471: Assertion 'slb->contains(pointer)' failed!       ../subprojects/frigg/include/frg/slab.hpp:475: Assertion '((address - slb->address) % item_size) == 0' failed!  ../subprojects/frigg/include/frg/slab.hpp:482: Assertion 'slb->num_reserved' failed!    ../subprojects/frigg/include/frg/slab.hpp:485: Assertion '!slb->available || slb->contains(slb->available)' failed!     ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed! lock read write unget update_bufmode seek     _init_type      _init_bufmode   _write_back _reset      _ensure_allocation              determine_bufmode               ../options/internal/include/mlibc/allocator.hpp !"Implement AllocatorLock slow path"  0123456789abcdef  ../options/ansi/generic/stdio-stubs.cpp new_buffer count < limit !"Not implemented"     Library function fails due to missing sysdep    L���Z���i���v���������������    Functionality is not implemented max_size > 0 
 %s:  %s
 returns:       mlibc: File locking (flockfile) is a no-op      mlibc: File locking (funlockfile) is a no-op    mlibc: File locking (ftrylockfile) is a no-op   mlibc: fread() I/O errors are not handled       mlibc: fwrite() I/O errors are not handled do_scanf: ' not implemented! do_scanf: m not implemented!    ����������������������������������������������������������������������������������������������������������������]������������������������������������������������������������������������������������������������������������������������������#�������������������n��������������������������������������������������A����������������������������������������������������������������������������������X�����������������������������������../subprojects/frigg/include/frg/formatting.hpp:200: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:213: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:217: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:221: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:225: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:229: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:235: Assertion '!opts.always_sign' failed!      ../subprojects/frigg/include/frg/formatting.hpp:236: Assertion '!opts.plus_becomes_space' failed!       ../subprojects/frigg/include/frg/formatting.hpp:240: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:247: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:254: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:258: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:262: Assertion '*s >= '0' && *s <= '9'' failed! ../subprojects/frigg/include/frg/formatting.hpp:266: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:275: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:279: Assertion '*s' failed!     ../subprojects/frigg/include/frg/formatting.hpp:286: Assertion '*s' failed! ,���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q�������q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���q���`���q�������q�������q���q���q���q�������q���q���
���q���q���q���q���q������;���]���]�������]���]���]���]���]���]���]���>�������]���]���]���]�������]���]���]���]���#�����������]���]�������]�������]���]���;���!opts.fill_zeros !opts.left_justify !opts.alt_conversion opts.minimum_width == 0    szmod == frg::printf_size_mod::default_size !opts.precision     [31mmlibc: Unknown printf terminator ' '[39m !"Illegal printf terminator"     ../subprojects/frigg/include/frg/slab.hpp:256: Assertion 'index <= num_buckets' failed! ../subprojects/frigg/include/frg/slab.hpp:266: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:267: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:269: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:284: Assertion 'object' failed!       ../subprojects/frigg/include/frg/slab.hpp:285: Assertion 'slb->contains(object)' failed!        ../subprojects/frigg/include/frg/slab.hpp:287: Assertion '!"slab_pool corruption. Possible write to unallocated object"' failed!        ../subprojects/frigg/include/frg/slab.hpp:299: Assertion 'slb->available' failed!       ../subprojects/frigg/include/frg/optional.hpp:97: Assertion '_non_null' failed! ../subprojects/frigg/include/frg/formatting.hpp:299: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:300: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:301: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:302: Assertion 'opts.minimum_width == 0' failed! 0x     ../subprojects/frigg/include/frg/formatting.hpp:307: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:308: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:309: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:310: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:311: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:317: Assertion '!opts.fill_zeros' failed!       ../subprojects/frigg/include/frg/formatting.hpp:318: Assertion '!opts.alt_conversion' failed! (null)    ../subprojects/frigg/include/frg/formatting.hpp:341: Assertion 'szmod == printf_size_mod::long_size' failed!    (   n   u   l   l   )           ../subprojects/frigg/include/frg/formatting.hpp:364: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/formatting.hpp:374: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:375: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:384: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:396: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:413: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:419: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:420: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:432: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:437: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:438: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:454: Assertion '!opts.left_justify' failed!     ../subprojects/frigg/include/frg/formatting.hpp:455: Assertion '!opts.alt_conversion' failed!   ../subprojects/frigg/include/frg/formatting.hpp:456: Assertion '!opts.precision' failed!        ../subprojects/frigg/include/frg/formatting.hpp:470: Assertion 'szmod == printf_size_mod::default_size' failed! ../subprojects/frigg/include/frg/formatting.hpp:477: Assertion '!"Unexpected printf terminal"' failed! %f       ../subprojects/frigg/include/frg/formatting.hpp:494: Assertion '!"Unexpected printf terminal"' failed!  ../subprojects/frigg/include/frg/mutex.hpp:57: Assertion '_is_locked' failed!   ../subprojects/frigg/include/frg/slab.hpp:529: Assertion 'overhead < slabsize' failed!  ../subprojects/frigg/include/frg/mutex.hpp:51: Assertion '!_is_locked' failed!  ../subprojects/frigg/include/frg/slab.hpp:554: Assertion '!(area_size & (page_size - 1))' failed! !#$%&()*+,-./:;<=>?@[]^_`{|}~ \\ \" \' \n \t \x{      ../subprojects/frigg/include/frg/rbtree.hpp:344: Assertion '(!get_left(node) && get_right(node) == child) || (get_left(node) == child && !get_right(node))' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:352: Assertion 'get_right(parent) == node' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:292: Assertion 'node == get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:125: Assertion '!_root' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:135: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:136: Assertion '!get_left(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:160: Assertion 'parent' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:161: Assertion '!get_right(parent)' failed! ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:377: Assertion 'h(n)->color == color_type::black' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:386: Assertion 'get_right(parent)' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:390: Assertion 'n == get_left(parent)' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:398: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:399: Assertion 'get_left(parent)' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:403: Assertion 'n == get_right(parent)' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:437: Assertion 'isRed(get_right(s))' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:444: Assertion 'get_right(parent) == n' failed!     ../subprojects/frigg/include/frg/rbtree.hpp:456: Assertion 'isRed(get_left(s))' failed! ../subprojects/frigg/include/frg/rbtree.hpp:209: Assertion 'grand && h(grand)->color == color_type::black' failed!      ../subprojects/frigg/include/frg/rbtree.hpp:240: Assertion 'parent == get_right(grand)' failed! ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/rbtree.hpp:480: Assertion 'u != nullptr && get_right(u) == n' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:496: Assertion 'get_right(w) == u' failed!  ../subprojects/frigg/include/frg/rbtree.hpp:515: Assertion 'u != nullptr && get_left(u) == n' failed!   ../subprojects/frigg/include/frg/rbtree.hpp:531: Assertion 'get_right(w) == u' failed! remove rename    renameat        tmpfile tmpnam  freopen setbuf scanf    operator() vscanf       operator()      operator()      vsscanf fwprintf        fwscanf vfwprintf       vfwscanf        swprintf        swscanf vswprintf       vswscanf        wprintf wscanf  vwprintf        vwscanf fgets fgetwc fgetws fputwc fputws fwide getwc   getwchar putwc  putwchar        ungetwc fgetpos fsetpos lock    getdelim        operator() expand       fgets_unlocked  ������������ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������� ��� ��� ��� ��� ��� ��� ��� ��� ��� ���9������������������� ������� ��� ��� ���\�����������9��� ��� ���9��� ������� ��� �������_���_���_�����������������������������������������������������������������������������������������������������������������������_���_���_��������������������������������������������������������������������������������������������������������������������������������������������������b����������������������������������������������b�������������������b���������������$���l���b���������������������b�����������b���'���'���'���L���L���L���L���L���L���L���L���L���L���L���L���L���L���L���L�������L���L���L���L���L���L���L���L���L���L���e�������'���'���'���L�������L���L���L���������������e���L���L���e���L�������L���L�����������������������������������������������������������������������������	�����������������j���������
����B"��B"��B"��B"��B"��B"��B"��B"��B"��B"��B"����B"��B"��B"��B"����B"��B"��B"��B"��B"����B"��B"��B"��B"��B"�����B"��B"�����2���5���5���5���5���5���5���5���5���5���5���5���.���5���5���5���5���.���5���5���5���5���5���0���5���5���5���5���5��j3���5���5���1��F��BI��BI��BI��BI��BI��BI��BI��BI��BI��BI��BI��B��BI��BI��BI��BI��B��BI��BI��BI��BI��BI��D��BI��BI��BI��BI��BI���F��BI��BI��E��../options/ansi/generic/string-stubs.cpp !"Not implemented" m   Functionality is not implemented        Operation would block (EAGAIN) Access denied (EACCESS) Bad file descriptor (EBADF) File exists already (EEXIST) Access violation (EFAULT) Operation interrupted (EINTR) Invalid argument (EINVAL) I/O error (EIO)       Resource is directory (EISDIR)  No such file or directory (ENOENT) Out of memory (ENOMEM)       Expected directory instead of file (ENOTDIR)    Operation not implemented (ENOSYS)      Operation not permitted (EFAULT) Broken pipe (EPIPE) Seek not possible (ESPIPE) No such device or address (ENXIO) Unknown error code (?)    �v���w���w���w���v���w���v���w���w���w���w���w���w���w���w���w���w���v���v���w���w���w���w�� w��w�� w���w��0w���w���w���w���w���w���w���w���w���w���w���w���w���w��=w���w���w���w��Jw���w���w���w��dw���w��Ww���w���w���w���w���w���w���w���w���w��qw��~w���w���w���w���w���w��    strxfrm strtok_r wcstod wcstof  wcstold wcstol  wcstoll wcstoul wcstoull wcscpy wcsncpy wmemcpy wmemmove wcscat wcsncat wcscmp  wcscoll wcsncmp wcsxfrm wmemcmp wcschr  wcscspn wcspbrk wcsrchr wcsspn wcsstr wcstok wcslen     wmemset         ../options/internal/generic/allocator.cpp       !mlibc::sys_anon_allocate(length, &ptr) !mlibc::sys_anon_free((void *)address, length) map unmap                 0123456789abcdef       ../options/internal/generic/charcode.cpp        (uc & 0b1100'0000) == 0b1000'0000 || (uc & 0b1111'1000) == 0b1111'1000  (uc & 0b1100'0000) == 0b1000'0000       wc <= 0x7F && "utf8_charcode cannot encode multibyte chars yet" !st.__progress cps.it == cps.end        encode_wtranscode       operator()              decode_wtranscode_length        operator()      decode_wtranscode decode         0123456789abcdef       mlibc: charset::is_alpha() is not implemented for the full Unicode charset      mlibc: charset::is_digit() is not implemented for the full Unicode charset      mlibc: charset::is_xdigit() is not implemented for the full Unicode charset     mlibc: charset::is_alnum() is not implemented for the full Unicode charset      mlibc: charset::is_punct() is not implemented for the full Unicode charset      mlibc: charset::is_graph() is not implemented for the full Unicode charset      mlibc: charset::is_blank() is not implemented for the full Unicode charset      mlibc: charset::is_space() is not implemented for the full Unicode charset      mlibc: charset::is_print() is not implemented for the full Unicode charset      mlibc: charset::to_lower() is not implemented for the full Unicode charset      mlibc: charset::to_upper() is not implemented for the full Unicode charset      ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!        0123456789abcdef      __cxa_guard_acquire contention  mlibc: Pure virtual function called from IP  0x ../subprojects/frigg/include/frg/logging.hpp:51: Assertion '_off < Limit' failed!       ../subprojects/frigg/include/frg/formatting.hpp:136: Assertion 'fo.conversion == format_conversion::null || fo.conversion == format_conversion::decimal' failed!        ../subprojects/frigg/include/frg/formatting.hpp:86: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/formatting.hpp:92: Assertion 'k < 32' failed!  ../subprojects/frigg/include/frg/logging.hpp:40: Assertion '_off < Limit' failed!              zR x�        �t��I    A�CD     <   �t��2    A�Cm      \   �a��   A�C    |   �b���   A�C� $   �   �d���   A�CN�����   �   3i���
   A�C      �   xt��-    A�Ch         �t��    A�CL         xt��"    A�C]      @  zt��-   A�C(    `  �u��"    A�C]       �  �u���    A�CE��      �  4v���    A�C�     �  �r��>    A�Cy      �  |v��8    A�Cs        �r��    A�CP   $   $  xv��3    A�I�I ]AA ,   L  �v���   A�A�O�V
AAG   H   |   x���    B�B�D �A(�D0T
(D ABBFT(G DBB     �  Tx��&    F�SG�    �  hx��1          �  �x��H            �x��       ,      �x��k    B�A�D �D0X DAB(   P  y��X    B�D�D �IAB     |  @y��z          �  �y��/    A�m      �  �y���          �  \z��          �  hz��#    TN $   �  �z���    G�A��
DA   (     8{���    G�A��
AAYA   @  |��\       �   T  X|��7   j�E�F �E(�D0�A8�GPv
8D�0D�(B� B�B�B�DR8A0A(B BBBD������PP������G8G�0A�(B� B�B�B�YP������     �  �|���            |}��   A��
D[   0  l~���          D  �~���    H�y   (   `  \��>    B�A�A �vAB   `   �  p��u   B�E�B �B(�A0�A8�D`E
8A0A(B BBBAD8F0A(B BBB      �  ����<    A�\   D     �����    B�B�E �B(�D0�A8�D@�8A0A(B BBB   T  ���(          h  $���-       D   |  @���m    B�E�B �B(�A0�A8�D@Q8A0A(B BBB   �  h���          �  t���          �  p���             l���\            ����V          (  ���           <  ���P       H   P  L���Q   [�B�B �B(�E0�E8��0f(I BFBL������      �  `����      L   �  ���!   T�I�E �B(�A0�A8�G`�8A0A(B BBBH������ <      �����    L�I�E �A(�A0�Y(A BBBD�����L   @  L����   F�B�A �A(�# AGBI����h(����} ADB   �  ���          �  �����          �  ����D       $   �  �����    A�A�G �AA$   �  ����#    A�A�G SDA    	  ����          0	  ����w          D	  (���Y       <   X	  t���y    G�E�A �D(�D0W(A ABBF����      �	  ����!    D\    �	  ̋��#    D^ 4   �	  ���[    F�D�D r
AAFDCAH��      
  ���          
  ���          (
  ���    D8   <
   ���A    G�A�C �b
�A�B�HAABD���   x
  4���d    U�|G� ,   �
  ����}    B�A�A �X
ABA   @   �
  ،���   B�B�B �A(�A0�NP
0A(A BBBK$     $���    A�D�G PAA <   0  ����    J�A�D A
AAFbG�A�G ��   <   p  |���   B�B�E �A(�D0��
(A BBBF      �  L����          �  ���       D   �  �����    K�A�A �c
ABEI
CBJAFBG���  \      \����    K�B�A �A(�D0w
(A ABBHD
(F ABBIh����H0����    �  ����&          �  ����          �  ����^      L   �  Г���   B�B�A �A(�D0g
(A ABBI�
(A ABBK      P���p    dK$   $  �����    e�G pAC�` �     L  `����    D0R
J    h  Ԙ��i    D0`
A @   �  (����   ~�G�D �
CBDCADH���h ���P   �  Ԛ���    _�J�D �C(�J0N
(L� A�B�B�GD(F ABBA����        ���~          0  ����Q          D  ؛��3    R�UI� ,   `  ����i    B�D�A �D0V DAB$   �  <���u    A�D�D0iAA   �  �����       8   �  P����    b�D�G RG�A�Q ��_
CAE<     ԝ���    u�C�G0Q
F�A�ILFAE��h0�� (   H  �����    W�T
�E^
B`�H�4   t  ����c    _�H�J O
F�A�IDCAH��\   �  0����    `�E�E �D(�I0�`�(A� B�B�B�R0�����A(F BBBC�����L     `����    e�E�D �H(�J@^
(A ABBDD(F ABBI����  (   \  ����c    a�O [
ADDCI�  $   �  ���^    F�G |
AFI�  D   �  ����    G�A�A �F
FBIA
FBGKABB���  4   �  d���\    F�D�K r
AAGDCAA��  4   0  ����g    b�D�D �f
�G�B�GACB,   h  Ġ��E    F�D�G f
AAAG��     �  ���;    F�c
�GCE�  4   �   ���S    F�D�G g
C�A�DDCAH��4   �  (���S    F�D�G g
C�A�DDCAH��   ,  P���6          @  |���a          T  ء��6       L   h  ����    S�E�D �D(�D0�
(A ABBAD(C ABBA����    �  ����6       H   �  ���p    B�B�A �A(�D0J
(D ABBCD(C DBB       ���'    DU
GF   @   8  ����    K�B�D �D(�F0b
(A ABBEP����  d   |  p����   J�E�B �B(�A0�A8�D@p
8C0A(B BBBK�������F@������      �  ؤ��          �  Ԥ��            Ф��             ܤ��          4  ���:       d   H  ���L   d�B�B �B(�D0�A8�D`�8C0A(B BBBI������A`������U������    �  ����+          �  ���C    Ii
FF      �  H����       �   �  Ħ���   T�B�B �B(�A0�A8�G�h
8A0A(B BBBK�������F�������J������F�������      |   ���f       �   �  \���=   K�B�B �B(�D0�A8�D`�
8D�0A�(B� B�B�B�KV
8A0A(B BBBHD
8F0A(B BBBE������P`�������   ,   ����   K�B�B �B(�A0�D8�D@
8A0A(B BBBEJ
8C0A(B BBBB`������P@������T8J�0I�(B� B�B�B� h   �  (����    ]�E�D �C(�G0z
(A ABBHO(Q� A�B�B�S0����J(M� F�B�B� (   0  ����F    F�C�G dF�A�   0   \  ����    [�D�G hCAF��X ��   (   �  \����    S�D�G kAAE��    �  ���          �  ���          �  ����/          �  ����       4     �����    ]�D�D �uABA���R ���    D  H���F    Ipp    \  ����          p  ����       T   �  ����*   K�H�J �H(�G0�A8�D�E
8A0A(B BBBA�������    �  p���          �  l���       X     x����   B�L�E �I(�A0�D`8
0C(A BBBES
0C(A BBBK     `  ܼ���       D   t  �����    B�E�E �E(�D0�D8�FP�8A0A(B BBB   �  ���          �  ���(          �  8���       0   �  D���B    A�D�G \
CADJFA 4   ,  `���^    F�D�D f
CAHJFAG��     d  ����       H   x  ����}    B�B�A �A(�D0w
(A ABBID
(F ABBA   �  ����       (   �  ����h    A�C�D s
DAH       ����+    A�i   X      ���1   a�B�A �D(�G0f
(A ABBEt(A ABBF����@0���� $   |  ���4    A�D�G eAA    �  ���6    A�t      �  ,���          �  8���'          �  T���(          �  p���.            ����          $  ����       4   8  ����    A�D�G0u
CAKU
AAI  4   p  �����    A�D�D0U
AAHK
CAI l   �  D���$   B�E�E �D(�A0�G`�
0C(A BBBEN
0F(C BBBCS
0F(C BBBF  4     ����    A�D�D0U
AAHK
CAI 4   P  \����    A�D�D0\
AAIK
CAA 4   �  ����|    A�D�D0M
AAHK
CAA T   �  ����y   B�B�B �D(�C0�G@_
0C(A BBBC�
0F(C BBBF     $���&          ,  @���&       4   @  \���|    A�D�D0I
AADK
CAI L   x  �����   T�E�D �D(�H@�
(A ABBH�����V@����    �  4���    D S    �  <���    D T    �  D���h    D c     ����?    T j    (  ����       4   <  ����9   S�A�D0�
AAF_AAG��<   t  �����    J�D _
DGC
CJN
AQlFN�      �  ����    D U <   �  �����    [�A�A �D0l AABG���H0���          ���!              <���/       4   4   X���g    A�D�G i
DAFT
DAG  $   l   ����3    A�I�G0]CA T   �   �����    B�B�B �D(�D0�J@�
0D(A BBBJL0F(A BBB   0   �    ���D    A�L�G ^
AADDFA 0    !  <���D    A�L�G ^
AADDFA H   T!  X����    B�H�E �E(�D0�F8�DPm
8C0A(B BBBE  H   �!  �����    B�H�E �E(�D0�F8�DPm
8C0A(B BBBE  (   �!  ����f    K�I�G0AAD��  l   "  4���Z   B�B�B �A(�A0�D@�
0D(A BBBB|
0G(D BBBCD
0G(D BBBK  <   �"  $����    B�A�D �Dpf
 CABID HAB h   �"  t����    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   h   4#  �����    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   h   �#  �����    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   @   $  ����    K�A�A �D@�
 AABHD FABK���    P$  ����6    IPa 0   h$  ����x    B�D�A �G0U
 AABI t   �$   ����   [�B�B �B(�A0�D8�G`u
8A0A(B BBBD�8A0A(B BBBE������``������  H   %  X���   B�E�B �E(�D0�A8�Dp\
8A0A(B BBBCT   `%  ���6   d�B�B �B(�D0�A8�GPD
8A0A(B BBBD�������   \   �%  ����   g�B�B �B(�A0�D8�D`8A0A(B BBBJ������V`������    &  ����1    A�Y
FP (   8&  �����    A�Z U
DDv
AA@   d&  h���o    B�B�E �D(�D0�G@j
0D(A BBBC     �&  �����    A�Q |Ax   �&  ���9   B�B�B �B(�D0�A8�G`
8A0A(B BBBCL
8A0A(B BBBJD
8F0A(B BBBEH   D'  �����   B�B�B �B(�D0�A8�GP_
8C0A(B BBBA  0   �'  ���    A�A�D0c
AAELAA   �'  h���V    A�c pA X   �'  ����6   K�B�A �A(�D@C
(A ABBA�(A ABBB����H@���� `   @(  ����3   B�B�B �B(�A0�A8�D`�
8A0A(B BBBGD
8F0A(B BBBE P   �(  h���%   Z�M�B �F(�D0�J@S0A(A BBBH�����P@�����   �(  D���       H   )  P���>   B�B�E �H(�D0�A8�GPb
8C0A(B BBBE     X)  D���          l)  @���       H   �)  <���x   B�E�E �B(�A0�A8�Gp�
8C0A(B BBBD h   �)  p����   B�B�B �B(�D0�D8�J�i
8D0A(B BBBHS�M�Q�B�J�N�V�A� l   8*  ����C	   B�E�E �B(�A0�A8�G���L�\�A�V�L�U�B��
8A0A(B BBBJ    �*  ����>    IPg |   �*  ����F   K�B�E �E(�D0�I8�D��
8A0A(B BBBEh
8A0A(B BBBFT8A0A(B BBBJ������H   @+  ����   B�E�B �E(�A0�A8�G�w
8C0A(B BBBF   �+  p���F    IPu    �+  ����       H   �+  ����q   B�G�B �B(�A0�A8�DPy
8A0A(B BBBJ H   ,  ����c   B�G�B �B(�A0�A8�DPw
8A0A(B BBBA    P,  ����V    A�c pA    p,  <���       8   �,  H���x    B�B�D �D(�G0t
(D ABBH  (   �,  ����2    B�F�D �^AB      �,  ����O           -  ����,          -  ����          (-  ���.          <-   ���          P-  ,���F       d   d-  h���   K�B�A �D(�D0�
(A ABBDD
(C ABBDD
(F ABBI`����  8   �-  ���V    L�D�D �b
ABGACBJ���      .  4���          .  @���#          0.  \���          D.  X���	          X.  T���          l.  P���              �.  H���3    \�QC�     �.  l����    `�G0^AJ�     �.  �����          �.  t����          �.  @����          /  ���          /  ���          (/  ���          </  ���          P/  ���          d/  ���G          x/  ��M          �/  P��          �/  L��          �/  H��(          �/  d��\         �/  ���8          �/  ���8          0  ��          0  ��          ,0   ���         @0  ����       H   T0  8���   B�B�B �B(�A0�A8�GP6
8A0A(B BBBGL   �0  �
���   B�B�B �A(�D0��
(A BBBE
(A BBBB   �0  \��!          1  x��
          1  t��          ,1  p���       (   @1  L��)   A�A�D 
AAH   l1  P��S    A�u
JR    �1  ���    DT d   �1  ���   L�J�E �E(�D0�C8�KP�
8A0A(B BBBD\8C0A(B BBBA������ \   2  @���    B�B�B �E(�D0�D8�G@^
8A0A(B BBBFg8A0A(B BBBH   l2  ���+   B�B�B �B(�D0�D8�GP�
8A0A(B BBBH `   �2  ����   B�B�B �B(�A0�D8�D`
8C0A(B BBBC�8F0A(B BBB  `   3  ���   B�B�B �B(�A0�A8�G`�
8A0A(B BBBJ�
8A0A(B BBBD$   �3  ����    A�A�G �AA$   �3  ���    A�A�D �AA$   �3  |���    A�A�G �AA   �3  D��    A�P   4   4  H���    B�B�A �A(�G0�(A ABBL   L4  ���	   B�B�B �A(�A0��
(A BBBNA(A BBB   ,   �4  ���W    R�G�H �P0a AAB 4   �4  ���T   A�D�G0�
AAD�AA  8   5  ���   B�H�A �D(�D0�
(A ABBHP   @5  ���Y   B�B�E �A(�A0�z
(A BBBD�
(A BBBH  4   �5  �"��R    B�G�D �Q
ABG_HB      �5  �"��	       H   �5  �"���   B�B�B �B(�D0�D8�G`�
8A0A(B BBBD H   ,6  `$��X   B�D�B �B(�A0�A8�D`�
8D0A(B BBBB    x6  t%���    Q�n  (   �6  �%��-    B�D�D �_AB   (   �6  �%��0    B�D�D �bAB   $   �6  �%��9    A�D�G VAA    7  �%��&    A�P   H   07  &���   B�B�B �B(�A0�D8�D`6
8A0A(B BBBG   |7  �*��       <   �7  |*��   K�B�A �A(�G0�(A ABBE����   H   �7  \+���   B�B�B �B(�A0�A8�D��
8A0A(B BBBG8   8  �1���    B�E�D �A(�G@x
(A ABBG  `   X8  d2��   B�G�B �B(�A0�A8�D`z
8A0A(B BBBIE
8A0A(B BBBA H   �8   4��
   B�B�B �E(�D0�A8�Dpx
8A0A(B BBBJ  H   9  �8��4   B�B�E �B(�D0�A8�DPe
8C0A(B BBBK   T9  �;��/          h9  �;��|       <   |9  `<���    B�H�G �A(�A0�G@�0A(A BBBH   �9  �<��   B�B�B �B(�D0�A8�FPj
8A0A(B BBBI    :  �=��f          :   >��]          0:  l>���          D:  (?��7          X:  T?��<          l:  �?��:          �:  �?��7          �:  �?��7          �:  @��R          �:  P@��U          �:  �@���          �:  A���       H   �:  �A���   B�B�B �E(�A0�A8�G@g
8A0A(B BBBKH   D;  (D���   B�H�K �K(�F0�H8�Dp
8A0A(B BBBDH   �;  �E���   B�B�B �B(�A0�A8�G��
8A0A(B BBBKH   �;  �Q���   B�B�B �E(�D0�C8�I��
8A0A(B BBBB`   (<  4g���   B�D�F �B(�A0�A8�Dp

8G0D(B BBBG�8C0A(B BBB  H   �<  �h���   B�G�M �B(�D0�A8�Fp�
8A0A(B BBBE L   �<  4j��   B�B�B �B(�A0�A8�D�3
8A0A(B BBBA   L   (=  m���    B�D�A �G0I
 CABC\
 CABFQ CCB H   x=  �m���   B�B�E �B(�A0�A8�DPE
8A0A(B BBBHL   �=  (o��?   B�B�B �E(�A0�A8�G��
8A0A(B BBBG   d   >  z���   B�B�E �B(�D0�C8�F�I
8A0A(B BBBE�
8A0A(B BBBH  H   |>  `���c   B�E�B �E(�A0�A8�FPb
8A0A(B BBBFT   �>  �����    B�G�B �A(�C0�G@]
0A(A BBBEf
0A(A BBBB8    ?  ,���   B�E�D �A(�F0�
(A ABBD 8   \?   ���   B�E�D �A(�F0�
(A ABBD $   �?  Ԇ��7    A�H�G dAA H   �?  ���l   B�B�E �B(�D0�A8�DpA
8D0A(B BBBF D   @  ���   Q�B�A �A(�G0�(A ABBK����H0����   T@  ���
          h@  ���       \   |@  ����k   O�B�E �B(�A0�A8�D@�8H�0A�(B� B�B�B�N@������   H   �@  �����
   B�B�E �E(�D0�A8�J��
8C0A(B BBBE4   (A  4���b    B�I�D �Q
ABEkGF   @   `A  l���~    A�K�I X
CAG\
CAHG
CAE  $   �A  ����R    A�D�G0CAA   �A  �����    �RL   �A  x���:0   B�G�B �B(�A0�A8�G�D
8A0A(B BBBD   0   4B  h����    A�A�D0�
AAD^DAH   hB  ����   B�M�B �E(�A0�D8�G�]
8A0A(B BBBG\   �B  �����   B�J�E �E(�A0�D8�G�y�_�H�B��
8C0A(B BBBH      C  ����              ,C   ���)          @C  ���          TC  ���1          hC  D���          |C  @���          �C  <����          �C  ����n          �C  D���    D�V      �C  H���       \   �C  D����    B�B�E �E(�D0�A8�G@Y
8A0A(B BBBCR8A0A(B BBB   HD  ����          \D  ����x          pD  ����       $   �D  ����M    A�A�D BCAL   �D  ���   B�E�B �E(�A0�A8�J��
8A0A(B BBBG      �D  ����Q    A�G@GAP   E  ���   B�F�B �D(�D0�G�h�B�B�K��0D(A BBB   L   pE  ����T   B�B�D �A(�J�T�c�B�B�K��
(A ABBJ`   �E  �����   B�B�B �E(�D0�D8�DP{
8F0A(B BBBG�
8A0A(B BBBKH   $F  8���   B�G�B �B(�A0�D8�J�N
8A0A(B BBBDL   pF  ����   B�J�B �B(�A0�A8�J�g
8A0A(B BBBC   L   �F  l���   B�J�B �B(�A0�A8�J��
8A0A(B BBBF   $   G  ,���P    A�D�G }AA H   8G  T���   B�B�B �B(�A0�A8�D@�
8A0A(B BBBE�   �G  (����   B�E�B �B(�A0�D8�Dpd
8A0A(B BBBF�
8A0A(B BBBK|
8A0A(B BBBJ�
8A0A(B BBBJ  `   H  �����   B�E�E �E(�A0�A8�J�s�~�D�A�V��
8D0A(B BBBF  (   �H  ����Q   J�A�G 4AAH��L   �H  ���p    L�F�A �D(�F0s
(C ABBHD(C ABBA����  H   �H  0����   B�E�B �B(�A0�A8�Hp
8A0A(B BBBF8   HI  ����n    B�D�D �D(�G@t
(A ABBA  H   �I  ���&   B�G�B �E(�A0�A8�J��
8A0A(B BBBId   �I  �����   B�B�E �B(�D0�A8�D��
8A0A(B BBBHu
8A0A(B BBBI  |   8J  4��:   B�E�B �B(�A0�D8�D��
8A0A(B BBBDe
8A0A(B BBBAM
8A0A(B BBBA   4   �J  ���3   A�N�JP|
AAIK
AAC (   �J  ����    {�G�J POAA��    K  ���
       \   0K  ����    B�B�B �B(�A0�A8�D@w
8C0A(B BBBGd8F0A(B BBB`   �K  ���J	   B�B�A �A(�I@t
(D ABBD
(D ABBGd
(F DBBF     �K  ���%    D`    L   ���           L  ���      0   4L  ����    A�A�D@~
CAHDFAT   hL  ���    B�B�B �A(�A0�DP�
0C(A BBBBD0F(A BBB   X   �L  ����   B�B�B �A(�D0�G�g
0A(A BBBG�
0A(A BBBC   H   M  0��   K�G�B �B(�A0�A8��0A(B BBBA������   H   hM  ����   B�B�B �B(�A0�A8�G��
8A0A(B BBBA<   �M  X��c    B�B�E �A(�F0�DPF0A(A BBB    �M  ���1    A�C�kA      N  ���          ,N  ���<    A�r
EC (   LN  ���C    B�D�A �vCB      xN  ���H    A�G ~A    �N  ��9    K�fG� H   �N  8���    B�B�B �B(�D0�A8�DPx
8D0A(B BBBJ H    O  ���Y   B�E�B �B(�A0�A8�G�Y
8A0A(B BBBI<   LO  ����    B�F�D �G@M
 AABDi AAB L   �O  ��   B�K�G �B(�A0�A8�G��
8A0A(B BBBB   l   �O  �*���   B�B�B �A(�H0�G@%
0D(A BBBJ�
0G(D BBBKL
0G(D BBBC   LP  P/��          `P  \/��	          tP  X/��          �P  d/��;          �P  �/��F          �P  �/��          �P  �/��          �P  �/��3    \�QC�    �P  0��
          Q  0��!          Q   0��A          0Q  \0��
          DQ  X0��
          XQ  T0��
          lQ  P0��
          �Q  L0��
          �Q  H0��
          �Q  D0��	          �Q  @0��
          �Q  <0��          �Q  H0���          �Q  1��
          R  1��           R  1��          4R  1��x          HR  �1��          \R  �1��(    A�f   4   xR  �1���    B�E�A �A(�G0�(A ABB$   �R  2��T    A�A�D ICA   �R  T2���      (   �R  �3��Q    I�A�G zAAC��  4   S  4��~    U�I�G s
G�A�HDCAH��0   PS  L4��o    A�A�D b
AAFxDA H   �S  �4���   B�B�B �B(�A0�D8�DP�
8A0A(E BBBH H   �S  <8��
   B�B�A �D(�G0�
(D ABBHD(G ABB  0   T   9���    B�C�A �D0�
 AABE    PT  �9��;    _[ d   hT  �9���   B�B�B �B(�A0�A8�D�q
8A0A(B BBBG)
8A0A(B BBBE   H   �T  L<��   B�E�E �B(�A0�A8�G�v
8A0A(B BBBI    U  @���          0U  �@��K          DU  �@��       8   XU  �@���    B�B�A �A(�D0b
(A ABBF 0   �U  hA��&   B�C�A �D0J
 AABH 8   �U  dB��    B�D�A �A(�D@o
(A ABBG     V  HC��D    A�y
FC D   $V  xC���    B�B�B �B(�A0�D8�DP�8C0A(B BBBH   lV  0D���    B�B�A �A(�D0[
(G ABBOD(A ABB  `   �V  tD��D   B�B�B �B(�A0�D8�G` 
8C0A(B BBBHQ8A0A(B BBB   H   W  `E��>   B�B�B �B(�A0�D8�G�V
8D0A(B BBBI$   hW  TF��Q    A�D�G0DA `   �W  �F���   B�G�B �B(�A0�A8�D`�
8A0A(B BBBJj
8A0A(B BBBD @   �W  (H���    A�A�G@c
DAGF
DAER
DAA x   8X  �H���   B�F�E �B(�D0�D8�GP[
8A0A(B BBBEd
8A0A(B BBBJ�
8A0A(B BBBA0   �X  �I��Z    A�D�G0p
AABWAA    �X  �I��W    D l
H  l   Y  8J���
   B�B�B �E(�D0�C8�J�C
8D0A(B BBBD1�E�_�B���\�K�B�   tY  �T��V       `   �Y  �T���   B�B�B �B(�D0�A8�F`�
8A0A(B BBBHZ
8A0A(B BBBD$   �Y  @V���    A�K�G qAA@   Z  �V���   K�B�B �A(�D0�x(A BBBE�����      XZ  Y���    O~
ChP(   xZ  �Y���    B�F�A ��AB     �Z  Z��g    LVd   �Z  `Z���   B�E�B �B(�D0�A8�D`
8A0A(B BBBD4
8F0A(B BBBA  X   $[  �]���   B�B�B �A(�C0�D�j
0C(A BBBFn
0C(A BBBH     �[  �_��G    A�|
CF    �[  �_��7    A�f
IF (   �[  �_��b    B�F�A �UAB  $   �[  @`��q    Y�A�K IAA@   \  �`��r    B�F�A �O
ABE}
ABHAFB   l   X\  �`��^   O�B�B �B(�A0�A8�Dp&
8A0A(B BBBE\
8A0A(B BBBJ�������  d   �\  �c��U   B�G�B �B(�A0�A8�D��
8A0A(B BBBE�
8A0A(B BBBA  4   0]  �f��Y    B�I�D �Q
ABEbGB   X   h]  �f���    B�E�D �D(�F0@
(C ABBCm
(H ABBFL(L ABBL   �]  Hg���   B�F�E �B(�D0�I8�Q��
8D0A(B BBBC   t   ^  �j��E&   B�B�E �E(�A0�A8�J�{
8D0A(B BBBF��L�u�B���F�]�B�          �^  А��K    X�kE�    �^  ���          �^   ���x          �^  l���          �^  h���          �^  t���1          _  ����           _  ����.          4_  ����          H_  ����
       $   \_  ����M    A�A�D BCAL   �_  ؑ���   B�B�B �B(�A0�D8�G��
8A0A(B BBBI   `   �_  X���u   B�H�B �B(�A0�A8�G�t�g�A�A�R��
8D0A(B BBBF  <   8`  t����   K�B�A �A(�G0�(A ABBF����  8   x`  $���c   B�D�A �A(�D`�
(A ABBE 8   �`  X����    B�B�D �A(�D@_
(A ABBF    �`  ���
          a  ���<    A�r
EC    $a  (���4    A�r      @a  L���Y    A�G OA   `a  ����9    K�fG� L   |a  �����   B�B�B �E(�A0�A8�J�
8D0A(B BBBE        �a  @���V          �a  ����          �a  ����h          b  ����          b  ����5       @   0b  ����#   B�B�B �D(�A0�D@w
0A(A BBBB  8   tb  �����    B�D�A �A(�D@S
(A ABBK  `   �b  <����   B�B�F �B(�A0�A8�D`
8A0A(B BBBGI
8A0A(B BBBE$   c  �����    A�A�G tAA   <c  ���H    DCL   Tc  ����   B�B�I �D(�G@;
(A ABBGL
(F ABBI  <   �c  ����u    B�C�A �D0S
 AABGH AAB L   �c  غ���    B�E�D �D(�F@�
(A ABBIN
(A ABBD      4d  x���
       <   Hd  t����    B�B�E �D(�A0�i
(C BBBH       �d  Ի���    T�R
JhH�  4   �d  `���t    A�D�G k
CAEY
CAC  ,   �d  ����q    K�D�G {
AAEX�� H   e  ����2   B�E�I �H(�A0�A8�G�X
8D0A(B BBBJ L   `e  ����   B�B�B �B(�A0�A8�F��
8D0A(B BBBA   <   �e  �����   K�B�A �A(�G0}(A ABBG����  H   �e  ,���B   B�B�B �B(�D0�D8�I�M
8A0A(B BBBH    <f  0���          Pf  ,���1          df  X���          xf  T���          �f  P����          �f  ����       (   �f  ����_    B�D�A �TAB  (   �f  ,���_    B�D�A �TAB     g  `���            g  \���Q    V�J ZAE�   $   Dg  ����6    A�A�G0hCA (   lg  �����   J�A�G �AAH��   �g  d���/    A�`
GF d   �g  t����    P�E�M �E(�A0�A8�F@J
8A0A(B BBBED8C0A(B BBBA������ d    h  �����   B�B�B �B(�A0�G8�G��
8A0A(B BBBA,
8A0A(B BBBD 4   �h  4���   A�K�JP|
AADK
AAK    �h  ���
          �h  ���%    D`    �h  0���       H    i  <���"   B�E�B �B(�A0�A8�Dp!
8A0A(B BBBD�   Li   ����   B�B�E �B(�A0�D8�Dpd
8A0A(B BBBFt
8A0A(B BBBJ|
8A0A(B BBBJH
8A0A(B BBBF   H   �i  8���   B�D�B �E(�D0�D8�D@�8A0A(B BBB      0j  ���6    A�t   L   Lj  0����   B�B�B �B(�A0�A8�J�
8D0A(B BBBF      �j  ���           �j  ���          �j  ���/          �j  ���       $   �j  ���L    A�C�G |CA X   k  ���i   B�B�B �A(�A0�D@u
0A(A BBBGd
0F(A BBBG   (   pk  ���l    B�A�A �dAB     �k  ��
          �k  ���       <   �k  ����    A�D�G S
AAGn
KANMFAL   l  (��k   B�G�E �B(�A0�C8�M�C
8A0A(B BBBB   ,   Tl  H��A    F�A�G kAAE��         �l  h��          �l  t��          �l  ���y       (   �l  ����    C�l
aF
JE
G      �l  ���           m  ���          m  ���          (m  ���          <m  ���       $   Pm  ���N    A�A�G @CAL   xm  ����    A�A�D f
AABD
FAEB
CAJYFA   `   �m  d��=   B�B�B �A(�A0�
(A BBBFQ
(F BBBCq
(F BBBC  (   ,n  @���    J�M o
AIGAA�    Xn  ���
       H   ln  ����   B�B�A �A(�G0d
(A ABBIW(A ABB    �n  ��       P   �n   ��h    F�E�E �D(�D0�e
(C BBBJH(A GBBA�����       o  <��U    A�
HL (   @o  |���    A�G b
AEXA   0   lo  ����   B�D�D �G@i
 AABB  H   �o  |���   B�B�B �B(�D0�D8�J�k
8D0A(B BBBF l   �o  2��E   B�B�E �G(�D0�GP�
0A(A BBBJe
0A(A BBBCh
0F(A BBBK     \p  �3���          pp  �4���          �p  h5��          �p  t5��           �p  �5��          �p  �5��y       (   �p  �5���    C�l
aF
JE
J       q  �6��       $   q  �6��G    A�A�G yCA H   <q  �6���   B�G�B �B(�A0�A8�D@.
8A0A(B BBBE(   �q  $8���    A�C�D0g
AAG    �q  �8��)    J�ZD� 4   �q  �8���    B�J�A �D(�K@e(A ABB   r  �8��
          r  �8��y          0r  \9��g          Dr  �9���       8   Xr  D:���   B�B�A �D(�D0�(A ABB   (   �r  �<���    J�A�G �AAD�� d   �r  l=��'   B�B�E �B(�D0�D8�D`�
8A0A(B BBBB	
8C0A(B BBBA     (s  4@��4    A�f
IC 0   Hs  T@���    q�h
GQ
AF
HP
HPH� d   |s  �@���   B�B�B �B(�D0�D8�G`[
8A0A(B BBBD�
8A0A(B BBBJ   H   �s  hF��4   B�B�E �B(�A0�A8�J�r
8A0A(B BBBE    0t  \W���          Dt  �W��I       H   Xt  X��d   B�B�J �E(�I0�G8�G��
8C0A(B BBBDH   �t  8\���   B�H�B �E(�D0�C8�G�~
8C0A(B BBBGH   �t  �d��I   B�G�E �B(�A0�D8�O`�
8C0A(B BBBJ   <u  �q���          Pu  ,r��"          du  Hr��          xu  Tr���          �u  �r��          �u  �r��          �u  �r��          �u  s��3          �u  0s��$          �u  Ls��`          v  �s���          v  $t��R         ,v  pu��$          @v  �u��(       H   Tv  �u��'   X�I�D �A(��
 AHBJA
 FBBAM���� l   �v  �v��W   B�E�B �B(�A0�A8��
0E(B BBBHF
0A(F BBBEO
0E(B BBBDX   w  |w���   B�E�B �B(�A0�A8��
0A(B BBBEA
0C(B BBBD L   lw   z��P   B�B�B �B(�A0�A8�D�p
8C0A(B BBBF      �w   ���:    Dd
HI      �w   ���$          �w  <���I          x  x����          x  4���$          ,x  P���e       D   @x  �����    q�F�A �I(�{
 ADBEV ADBK����     �x  d���          �x  p���3          �x  �����          �x  8���          �x  D���       L   �x  P���	   T�J�A �A(�� AFBE����H(����G AFB  4   <y  ���!   B�D�A �A(��
 ABBK      ty  ���    DT    �y  ���          �y  ���          �y  (����       4   �y  ����	   B�D�A �A(��
 ABBK       z  |���    DT    z  ����          ,z  ����!          @z  ����          Tz  ����	          hz  ����          |z  �����          �z  L����          �z  ����       X   �z  t����    B�B�F �C(�D0j
(C ABBE`
(A ABBBD(J ABB 4   {  ����x    B�A�E �q
CBBQ
ADJ   L{  ����&          `{  ���          t{  ���          �{  ���       X   �{  ���   B�I�B �B(�A0�H8�1
0D(B BBBK�0A(E BBB      �{  ԋ���       p   |  p���-   [�B�B �B(�A0�A8��
0A(B BBBFA
0F(B BBBI�������H8������ X   �|  ,����   B�B�B �B(�A0�A8��
0A(B BBBDy
0F(B BBBA    �|  `���
       H   �|  \���E   B�E�B �B(�A0�I8�G`8D0A(B BBB      <}  `���/    A�m      X}  t���V       H   l}  �����   B�B�B �E(�D0�D8�Dp�
8D0A(B BBBA @   �}  d���t    B�I�D �G@R
 AABDe
 FABB   8   �}  ����u    B�E�A �D(�D@G
(C ABBA H   8~  ����   B�H�B �E(�D0�A8�Np�
8A0A(B BBBK 4   �~  H����    A�I�I0y
AABD
CAH @   �~  �����    B�I�F �D0�
 AABHD
 CABF  (      \���X    A�A�D0U
AAC  L   ,  �����    B�B�D �A(�D0�
(A ABBAD
(C ABBA   8   |   ����    B�D�D �a
ABBA
CBJ   �   �  t���P   B�J�B �B(�A0�A8�D@�
8J0A(B BBBFD
8C0A(B BBBHJ
8D0A(B BBBI�
8A0A(B BBBA   H   P�  ,���   B�E�H �B(�D0�A8�DP�
8D0A(B BBBF 8   ��  ����    B�G�A �h
ABKA
CBJ   T   ؀  T���B   B�G�B �A(�D0�G@[
0A(A BBBFR
0F(A BBBAH   0�  L����   B�B�B �B(�A0�D8�D`R
8A0A(B BBBC8   |�  ����   B�B�A �A(�G0v
(A ABBG  4   ��  d���
   B�B�D �A(�D0�(A ABB4   ��  <���q   K�A�A ��
ABC����      (�  ����)    A�g      D�  ����1    Z�TB�    `�  ����(    A�f   H   |�  Ц��-   B�E�E �B(�D0�D8�G`�
8D0A(B BBBF H   Ȃ  ����J   B�E�B �E(�D0�D8�G`�
8A0A(B BBBG    �  �����       H   (�  T���)   B�B�B �B(�A0�D8�G@�
8D0A(B BBBG    t�  8���
       H   ��  4����   B�E�B �B(�A0�I8�G`�
8A0A(B BBBB 0   ԃ  ���J    A�I�L N
AAJDPA H   �  ���Z   B�E�E �B(�A0�A8�G`g
8A0A(B BBBH  0   T�  ���J    A�I�L N
AAJDPA 8   ��  4����    B�G�I �A(�G0P
(C ABBF  (   Ą  ���t    A�F�G H
AAH x   ��  <���(   T�B�E �E(�D0�D8�F�d
8A0A(B BBBDD8F0A(B BBBE������F�������   H   l�  ���K   B�K�B �B(�A0�A8�DP%
8A0A(B BBBA    ��  ����   G��
GL
D L   ܅  ����   B�B�B �E(�A0�D8�G�
8A0A(B BBBH   H   ,�  @���v   B�F�E �E(�A0�A8�D`�
8C0A(B BBBAL   x�  t���	   B�I�E �B(�A0�A8�D��
8A0A(B BBBF   <   Ȇ  4����    B�B�B �D(�D0��
(C BBBD   H   �  �����   B�I�B �E(�A0�A8�GP�
8C0A(B BBBD<   T�  8����    B�B�E �D(�A0�^
(C BBBK   H   ��  ����j   B�B�E �B(�E0�D8�D`,
8C0A(B BBBHH   ��  ����2   B�E�B �F(�A0�D8�DP�
8C0A(B BBBF L   ,�  ����   B�F�B �B(�A0�A8�G�w
8C0A(B BBBH      |�  ����V           ��  ����U    y�D�VA       ��  8���?    a�D�XA       ؈  T���?    a�D�XA   0   ��  p���\    A�N�L N
AAEiAA H   0�  ����n   B�G�B �B(�A0�A8�G�`
8D0A(B BBBE p   |�  ����Q   B�B�A �A(�D0K
(C ABBCa
(C ABBGw
(C ABBA\
(F ABBI     ��  ����&       8   �  �����    B�B�A �A(�D@c
(C ABBK    @�  ���(    D c L   X�  4���r    B�A�A �D0p
 DABAS
 DABFD JAB   H   ��  d����   B�B�B �H(�A0�A8�G�l
8A0A(B BBBC 0   �  ����B    A�I�J N
AADDPA    (�  ���          <�   ���       L   P�  �����    B�G�I �A(�G0P
(C ABBF�
(L ABBI   L   ��  ����(   B�E�B �E(�A0�A8�G��
8A0A(B BBBJ   ,   ��  �����    B�H�D �w
CBF   L    �  ���+   B�B�B �B(�A0�A8�D��
8C0A(B BBBK   H   p�  ����
   B�B�B �B(�A0�A8�D�P
8D0A(B BBBE D   ��  ����   B�B�B �B(�A0�A8�j
0A(B BBBC     �  8��       @   �  D���   D�I�B �I(�E0�A8�v0A(B BBB    \�  �	���          p�  <
��w          ��  �
��3          ��  �
��          ��  �
��          ��  �
��       @   ԍ  �
���   D�I�B �E(�D0�A8��0A(B BBB    �  D���          ,�   ��H          @�  <��       L   T�  8���   B�B�B �B(�A0�A8�G��
8A0A(B BBBA   L   ��  ���m   B�B�E �B(�A0�A8�G�|
8A0A(B BBBA   L   �  ����	   B�K�B �B(�A0�A8�G��
8A0A(B BBBJ   H   D�  H ��8   B�B�E �E(�D0�C8�F`�
8A0A(B BBBI H   ��  <"���   D�I�B �B(�A0�D8�D`Y
8A0A(B BBBCH   ܏  �$���   B�B�B �B(�A0�A8�D@�
8A0A(B BBBE$   (�  D&��C    A�F�G cLA    P�  l&��       L   d�  h&��5   B�G�B �B(�A0�A8�D��
8A0A(B BBBG   H   ��  X+��U   B�B�B �E(�A0�A8�D@<
8A0A(B BBBA$    �  l/��<    A�F�G \LA (   (�  �/��"   A�A�D AA   ,   T�  �0��}    G�A�D �b�G�B�      ��  �0��
       $   ��  �0���   K�i
Lp�H� d   ��  l2��\   B�E�E �E(�A0�A8�I@}
8A0A(B BBBE[
8A0A(B BBBC      (�  d4��Q       (   <�  �4��   e�C��FN��H��$   h�  �7��I    A�L�[ WHA 0   ��  �7��K    A�D�M0M
AAG`AA L   Ē  �7���   B�G�B �B(�D0�D8�D�
8A0A(B BBBG   H   �  H?��   B�B�B �B(�D0�A8�GP�
8A0A(B BBBF H   `�  @��P   B�B�B �B(�A0�A8�Dp�
8A0A(B BBBA H   ��   C���   B�E�B �B(�D0�A8�D`Z
8A0A(B BBBHH   ��  �E��?   B�B�B �B(�D0�D8�Dpw
8A0A(B BBBK  L   D�  �H���   B�F�B �B(�A0�A8�G�h�
8D0A(B BBBF   ,   ��  �S��f    F�D�G0[
AABp�� 4   Ĕ  8T���   A�W �
AJe
AJJ
AE   X   ��  �U��4   B�E�B �K(�I0�D`x
0C(A BBBES
0C(A BBBK   \   X�  �X���   B�B�B �B(�A0�A8�L�j�D�F�A��
8A0A(B BBBK  L   ��  $\���   B�H�E �B(�A0�A8�G�{
8A0A(B BBBA      �  �d��       \   �  �d��=   B�H�B �B(�A0�A8�L��b�X�A�
8A0A(B BBBE    |�  pr��          ��  lr��    D Z    ��  tr��       8   ��  pr���   B�D�D ��
IBJ�
IBD  L   ��  �s��Z   B�I�E �B(�A0�D8�G���
8A0A(B BBBA  L   H�  �v���   B�B�E �B(�A0�A8�G�1
8A0A(B BBBA   H   ��  �{���    B�E�E �E(�A0�D8�D��
8A0A(B BBBA(   �  8|��g    B�A�D �q
CBC(   �  ||��l    B�A�D �|
CBHL   <�  �|��Z   B�I�E �B(�A0�D8�G���
8A0A(B BBBA  L   ��  ����   B�G�B �B(�A0�A8�G��
8A0A(B BBBA   H   ܘ  P���M   B�B�B �B(�A0�D8�G�x
8C0A(B BBBH (   (�  T���:    A�A�G kDA     (   T�  h����    f�A�QAG��H��   ��  ܍���       D   ��  �����   B�E�B �B(�A0�D8�
0A(B BBBF     ܙ   ���          �  ���          �  ���          �  ���9          ,�  @���9          @�  l����       $   T�  H���m    A�D�G ^AA4   |�  �����    B�E�A �D(�D0u(A ABB$   ��  ���C   @�F��AA��  \   ܚ  ����   P�I�G �E(�A0�A8��
0A(B BBBEP������H8������ `   <�  @���#   B�G�H �E(�G0�H8�J`Z
8A0A(B BBBE�
8A0A(B BBBJ8   ��  ����    B�E�A �A(�G@t
(A ABBF  @   ܛ  `����    O�A�C �G0R
 AABH] AABG��� <    �  ̙��t    B�D�D �D0]
 AABA AAB  (   `�  ���Q    B�A�D �`
ABF`   ��  @����   B�H�E �E(�D0�C8�Dpu
8A0A(B BBBBY
8A0A(B BBBEH   �  |����    B�G�D �D(�G0M
(A ABBEI(A ABB  ,   <�  ����V    B�D�D �G0@ AABH   l�  �����    B�B�B �B(�A0�A8�G��8A0A(B BBB      ��  t���Q       T   ̝  �����   Q�E�E �B(�E0�J8�Ip�
8A0A(B BBBE�������  8   $�  ����u    R�A�A �L
�A�B�MAAB   <   `�  <���O   B�B�B �A(�C0��
(A BBBE   <   ��  L����   B�E�E �A(�A0��
(A BBBK  T   ��  ����   B�B�B �E(�A0�I8�G`�h]pUhE`/8A0A(B BBB |   8�  $���"   M�B�B �E(�D0�A8�GpE
8A0A(B BBBG�������Hp������o
8A0A(B BBBG  H   ��  ԩ���   B�J�B �B(�A0�A8�G��
8A0A(B BBBC   �  h���       \   �  t���   M�B�B �B(�A0�A8�Gp�8A0A(B BBBJ������Hp������ $   x�  4����    A�A�K �AAt   ��  ����4   B�B�E �E(�D0�D8�FPs
8A0A(B BBBG�
8A0A(B BBBGa8A0A(B BBBX   �  �����    I�B�B �A(�A0�Q(A BBBI�����H0�����D(A BBB\   t�  �����    I�B�B �A(�A0�Q(A BBBI�����H0�����E(A BBB       ԡ  �����          �  �����          ��  `����          �  ,����          $�  �����       d   8�  d���    B�E�B �E(�E0�A8�G`<
8A0A(B BBBG�
8A0A(B BBBB   (   ��  ���a    B�D�D �SAB  H   ̢  `����   B�E�H �D(�G03
(A ABBE�(F ABBH   �  ���   B�B�D �H(�G0}
(A ABBFi(F ABB   d�  �����          x�  t���B          ��  ����!      4   ��  �����   B�B�A �A(�U
 ABBH      أ  T���          �  P���           �  L����       <   �  ����   B�B�B �A(�A0�y
(A BBBH      T�  ����          h�  ����          |�  ����          ��  ����!    GY    ��  ����          ��  ����       d   Ф  �����   B�E�E �B(�A0�A8�Dp�
8C0A(B BBBH�
8F0A(B BBBD   d   8�  ���+   B�B�D �D(�G0m8f@I8A0k
(A ABBGt
(F ABBIP8F@W8A0   �   ��  ����\   B�B�E �B(�A0�A8�D���G�G�B��
8C0A(B BBBDQ
8A0A(B BBBE�
8F0A(B BBBET�B�I�A�      D�  ����2   '���
A$   d�  ����9    A�D�G0hCA    ��  ����/       H   ��  ����$   B�B�I �B(�A0�A8�J�L
8A0A(B BBBG,   �  ����S    B�G�A �EAB         �   ���          0�  ����          D�  ����!    GY    \�  ���          p�  ���           ��  ���   J d
Bz
F     ��  ���/          ��  0����       $   ԧ  ����h    A�D0f
ADvAL   ��  ����{   B�B�B �B(�A0�A8�GЁ[
8A0A(B BBBA  T   L�   ����   k�A�G�-��P���L
AABS
CAI`��P���   (   ��  X���    A�G }
AJO
AH L   Ш  �����   B�B�B �E(�A0�A8�D��
8A0A(B BBBD       �  ���)    Dd (   8�  $���G    B�D�A �|AB   $   d�  H���9    A�D�G0hCA H   ��  `����   B�E�B �I(�A0�A8�J�L
8A0A(B BBBD   ة  ���          �   ���           �  ���       H   �  ���p   B�J�J �B(�I0�A8�G�<8A0A(B BBB     `�  <���*    DC b  H   |�  P���   B�V�D �E(�G��
(A ABBFt(A ABB   Ȫ  $���$    D_ (   �  <���S    B�G�A �EAB  L   �  p����   B�E�B �B(�A0�A8�G��
8A0A(B BBBB   $   \�  ����    A�D�G qAA   ��  H��R    Ry (   ��  ���~    X�A�G PCAD�� X   ȫ  ���2   B�J�E �B(�A0�A8��
0A(B FBEGK0F(B BBB   4   $�  ����    B�A�D �~
ABHMIB     \�  @��          p�  <��          ��  8��    H R    ��  @��    H R (   ��  H��.   A�C�G0Q
AAB  H   �  L��A   B�B�B �B(�A0�D8�GP}
8A0A(B BBBE P   ,�  P���   K�B�B �A(�C0�
(A BBBD������F0������   ��  �	��b   X�B�B �B(�A0�A8�D�

8A0A(B BBBHT
8F0A(B BBBE�
8A0A(B BBBHH�F�B�D�P���R�F�F�N�}������F���������Q�I�F�W�  L   \�  p#���   B�M�H �A(�G0�
(A ABBKP
(C ABBH  `   ��  �$���   B�B�E �D(�D0�e
(A BBBCo
(D BBBG[
(A EBBK      �  &��	       \   $�  &��   T�B�B �B(�A0�D8�JPN8A0A(B BBBG������HP������ T   ��  �(���    `�A�G�s
DAHI
AAED
FAEX��P���       0   ܯ  p)��c    A�I M
AHa
FIQA   (   �  �)���   A�A�G 
AAF0   <�  +���    R�D�S0]AAH��H0��     p�  �+��*          ��  �+���       P   ��  T,��$   T�B�B �A(�D0�JPt0A(A BBBE�����HP����� $   �  0-���    A�H�G �AA(   �  �-��L    B�A�A �DAB  H   @�  �-���   B�B�B �B(�A0�C8�G`C
8D0A(B BBBE L   ��  �1��,   B�B�B �E(�D0�D8�D@�
8D0A(B BBBC        ܱ  `3��)       D   �  |3��f   Z�B�A �A(�B����H(����\
 DBBD <   8�  �4��p    B�I�A �D0i
 AABCi CAB     x�  �4��c          ��  05���          ��  6��c    D^,   ��  d6��$   A�G �
ACn
AA   4   �  d7��/   A�D�D(
AADP
AAF    �  \9��	       8   4�  X9���   B�B�A �D(�G8�
(A ABBF `   p�  �:���    B�B�E �B(�D0�D8�F�[
8A0A(B BBBB�
8A0A(B BBBA   Գ  �;��       `   �  �;��q   B�E�B �A(�D0�J
(A BBBA�
(A BBBHx
(F BBBA     L�  �<���          `�  ,=��          t�  (=��0          ��  D=���          ��  >��0          ��  ,>��H          Ĵ  h>���          ش  ?��0          �   ?��P           �  \?��          �  h?��           (�  t?��1          <�  �?��1          P�  �?��%          d�  �?��          x�  �?��          ��   @��d          ��  \@��          ��  X@��)          ȵ  t@��          ܵ  p@��          �  l@���         �  XB��      @   �  TC���   B�D�A �D0�
 AABAv
 AABD4   \�  �E���   D��
Hi
GO
Ah
H{
E  $   ��  �G��f    Q�A�G JAA$   ��  �G��q    A�A�D hAA   �  (H��    A�X       �  ,H��(    A�f   <   �  @H���    B�A�A �D0o
 AABE^ AAB 4   \�  �H��g    B�E�D �I(�J@B(A ABBL   ��  �H���    B�E�I �G(�G@z
(A ABBBu
(A ABBE   <   �  �I���    L�C�A �G0o
 AABF` CAB (   $�  J��Y    A�D�G g
AAK  H   P�  <J���    B�B�B �A(�A0�Z
(A BBBGO(A BBBH   ��  �J��   B�B�B �B(�A0�A8�Dph
8D0A(B BBBEH   �  DN��]   B�B�B �B(�A0�A8�Dp�
8D0A(B BBBH    4�  XO��)    D` H   L�  pO��e   B�B�B �E(�A0�A8�J��
8A0A(B BBBJH   ��  �T��O   B�E�B �B(�D0�D8�J��
8A0A(B BBBDH   �  �U��E   B�E�E �B(�D0�A8�D`�
8D0A(B BBBD    0�  �V��     DW    H�  �V���       0   \�  �W���    B�E�D �G0G
 AABC     ��  X��x   E��
Ge
c    ��  xY���      (   Ⱥ  �[���   A�C��
AK�A(   ��  �]��    A�L
CG
IQ
GF    �  �]��x    A�G
Hg8   @�  L^��$   B�B�A �A(�G0(A ABB   8   |�  @_��8   B�G�A �A(�G0(A ABB   L   ��  D`���    U�E�A �A(�G0\
(C ABBID(F ABBA���� \   �  �`��   B�D�E �E(�D0�D8�NP�
8A0A(B BBBCD8F0A(B BBB8   h�  da���    B�I�E �D(�A0�e(D BBB     ��  �a��c          ��  b��x          ̼  �b��h       H   �  �b��{   B�B�E �E(�A0�C8�H`d
8C0A(B BBBF    ,�  d���          @�  �d��    A�R   ,   \�  �d��	   B�A�D ��
ABG       ��  �e���    D�T��E  l   ��  �f���	   B�B�B �B(�A0�D8�J���L�}�B�v
8A0A(B BBBEP�L�I�A�     �  ,p��          4�  8p��          H�  Dp��2          \�  pp��5          p�  �p��h          ��  �p��o          ��  Tq��>       (   ��  �q��Q    F�A�G uAAK��  x   ؾ  �q���   B�B�B �B(�D0�A8�Dpi
8A0A(B BBBD\
8F0A(B BBBEH8A0A(B BBB   H   T�  s���    B�H�B �E(�D0�A8�D`�
8A0A(B BBBF d   ��  �s��`   B�I�B �E(�H0�A8�G�q
8A0A(B BBBC�
8A0A(B BBBK      �  �x��j    A�G E
AB    ,�  �x��i    A�|
C,   H�  4y���    B�D�C ��
ABA   0   x�  �y���    B�D�D �Gpa
 AABJ P   ��  z���   B�B�E �E(�D0�D8�D`AhE`V
8A0A(B BBBH \    �  \{��6   B�E�E �E(�F0�G8�G�R�U���B��
8A0A(B BBBA   T   `�  <}���   B�E�B �E(�A0�D8�G���E�Y8A0A(B BBBE�     ��  �~��'          ��  �~��       <   ��  �~��T    B�D�I �G0M
 AABI_ AAB  4    �  ��J    R�D�D �W
ABDJ�A�B�   X�  $��'          l�  @��<       H   ��  l���    B�B�A �A(�D@�
(A ABBJt(F ABB  8   ��   ���F   B�D�D �[
ABH�
ABA     �  ���'          �  0���       (   0�  <���d    B�D�I �QAB  4   \�  ����J    R�D�D �T
ABGJ�A�B�H   ��  �����   B�E�B �B(�D0�A8�D`c
8A0A(B BBBG  H   ��  ���}    B�D�B �A(�A0�R
(C BBBKC(C BBB   ,�  @���       4   @�  L���U    B�D�A �w
ABGIAB      x�  t���b       L   ��  Є��h   B�B�B �B(�A0�A8�G�
8D0A(B BBBD   (   ��  �����    B�J�K ��AB     �  �����       H   �  ���x    B�B�D �D(�D0H
(A ABBBD(J ABB     h�  D���X       p  |�  ����;/   B�F�E �B(�A0�A8�Q��+
8A0A(B BBBI*��H��k��A�����R��_��B����Q��^��B��A��H��e��B���
��G��gb��G��f��B�����J��_��A��M��Q��a��A��V	��H��]��A��M��N��z��A��u
��A��Z���H��E��B�����B��J��B��y��Q��O��E��   �   ��  \���   B�E�E �B(�A0�D8�G�O�L�F�A�g�P�J�B���H�\�A�n
8A0A(B BBBF��L�I�A�    ��  ����7          ��  ����           ��  �����    A��
VP
A    ��  ���          ��  (���#          ��  D���
           �  @����   A��
AL
L   0�  ����      L   D�  �����   B�F�B �E(�D0�A8�J�l
8A0A(B BBBD      ��  ���&    A�d   4   ��  ���V    M�A�D �W
�F�B�OP���      ��  D���          ��  @���          �  <���       4   $�  8����    J�A�J �
AAALFAE��    \�  ����7    Dr    t�  ����              ��  ����          ��  ����       �   ��  �����   B�B�B �B(�A0�A8�DP
8A0A(B BBBHh
8A0A(B BBBFl
8F0A(B BBBED
8F0A(B BBBEl   H�  T����   B�B�B �A(�A0�D@�
0A(A BBBH�
0F(A BBBGD
0F(A BBBG   ��  �����    f�R@UA   ��  T���F    K�eH� |   ��  ����M   I�G�E �B(�A0�A8�K�}������G��������
8A0A(B BBBA�������L�������   t�  X���1    D l    ��  ����'    D b    ��  ����          ��  ����+    D f    ��  ����+    D f    ��  ����,    D g     �  ����%    D `        �   ���k       <   0�  \����    B�A�D �G0U
 AABI[ AAB8   p�  �����    R�E�E �G(�N0N
(A ABBK     ��  ����3    A�q      ��  ����           ��  �����    A�A��A  $    �  \���     D�LG FAA      (�  T���       H   <�  `���I   B�F�E �H(�G0�A8�GP8A0A(B BBB   T   ��  d���o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T   ��  |���o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB     8�  ����(    DK X  8   T�  �����    B�I�B �A(�A0�}(A BBB  0   ��  ����    H�F�E �A(�� ABB     ��  ����(    D c    ��  ����              ��  ����          �  ����          �  ����          0�  ����          D�  ����          X�  ����       �   l�  ����R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   �  h���m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        l�  }���>    A�CA�x   ��  s���    A�CM      ��  f���\    A�CW     ��  �����    A�C�     ��  ���    A�CZ      �  ���6    A�Cq      ,�  1����    A�C�     L�  ����    A�CN      l�  ����6    A�Cq      ��  ����    A�C      ��  ����;    A�Cv      ��  ����c    A�C^     ��  ����   A�C    �  ����    A�CF      (�  ����    A�CB      H�  ����#    A�C^      h�  ����    A�CV      ��  ����V    A�CQ     ��  ���)    A�Cd      ��  ���    A�CF      ��  ���)    A�Cd      �  ���(    A�Cc      (�  ���,    A�Cg      H�  $���    A�CF      h�  ���    A�CF      ��  ����4    A�Co      ��  ���E    A�C@     ��  5���C    A�C~      ��  X���&    A�Ca      �  ^���*    A�Ce      (�  h���J    A�CE     H�  �����    A�C�     h�  C����    A�C�     ��  ����U    A�CP     ��  �����   A�C�    ��  s���(    A�Cc       ��  |����    A�C�         �  ���    A�CZ      ,�  ���!    A�C          L�  ���   A�C    l�  ����   A�C    ��  ����)    A�Cd      ��  ����    A�CF      ��  ����)    A�Cd      ��  ����(    A�Cc      �  ����,    A�Cg      ,�  ����4    A�Co      L�  ���E    A�C@     l�  3���C    A�C~      ��  V���&    A�Ca      ��  \���*    A�Ce      ��  f���J    A�CE     ��  �����    A�C�     �  A����    A�C�     ,�  ����U    A�CP     L�  �����   A�C�    l�  r����    A�C�     ��  ���F    A�CA     ��  +���Z    A�CU     ��  e����    A�C�     ��  ����<    A�Cw      �  ~��     A�C[      ,�  ~���    A�C�     L�  ���   A�C�    l�  ���6    A�Cq      ��  ���Q    A�CL     ��  ��    A�CN      ��  ���B    A�C}      ��  ��    A�CQ      �  [���-    A�Ch      ,�  h���$    A�C_      L�  l���$    A�C_      l�  p���$    A�C_      ��  t���3    A�Cn      ��  ����%    A�C`      ��  ����9    A�Ct      ��  ����J   A�CE    �  ����+    A�Cf      ,�  ����G   A�CB    L�  ���+    A�Cf      l�  ���    A�CU      ��  ���+    A�C      ��  ���"    A�C]      ��  ���Z    A�CU     ��  Q���U    A�CP     �  ����V    A�CQ     (�  ����#    A�C      D�  ����)    A�Cd      d�  ����+    A�C      ��  ����    A�C      ��  ����    A�C      ��  ����*    A�C      ��  ����+    A�C      ��  ����+    A�C      �  �����    A�C�     ,�  ����   A�C    L�  ����*    A�C      h�  ����+    A�C      ��  ����+    A�C      ��  ����&    A�Ca      ��  ����/    A�C      ��  ����/    A�C       ��  	���   A�CE��      �  ����1   A�C,    <�  ����.    A�C      X�  ���=   A�C8    x�  )���3    A�C      ��  @����    A�C�     ��  ����    A�C�     ��  �����    A�C�      ��  V����    A�CE��      �  ����3    A�C      4�  ���M   A�CH    T�  ��L   A�CG    t�  ?��   A�C    ��  <	��)    A�Cd      ��  E	��    A�Cz     ��  �	���    A�C�     ��  �
��)    A�Cd      �  �
��(    A�Cc      4�  �
��0    A�Ck      T�  �
��+    A�Cf      t�  �
��E    A�C@      ��  �
��h   A�CE�^      ��  ���   A�CH��      ��  ���#   A�CE�      �  ���}    A�Cx      �   ��2    A�Cm      @�  ��'    A�Cb      `�  ���    A�C�     ��  ����    A�C�     ��  ^��O    A�CJ     ��  ���    A�CQ      ��  ���I    A�CD      �  ����    A�C�      �  ����    A�C�     @�  ��X    A�CS      `�  V��D   A�CE�:     ��  v���    A�C�     ��  J��L    A�CG      ��  v���    A�CE��      ��  ����    A�C�     �  n��    A�CL      (�  _��    A�CY      H�  ]��    A�CY       h�  \��a   A�CE�W     ��  ���    A�CY       ��  ����   A�CE��     ��    ��    A�CL      ��  ���j    A�Ce     �  < ��(    A�Cc      0�  D ��    A�CY       P�  B ��7   A�CE�-     t�  U!��    A�CY       ��  T!��7   A�CE�-      ��  h"��a   A�CE�W     ��  �$��    A�CY       ��  �$���   A�CE��      �  '��d    A�C_     @�  P'��j    A�Ce      `�  �'��7   A�CE�-      ��  �(��7   A�CE�-     ��  �)��K    A�CF     ��  �)��W    A�CR     ��  $*��    A�CQ      �  *��    A�CY      (�  *��1    A�Cl       H�  **���   A�CE��     l�  �/��    A�CX      ��  �/��H    A�CC     ��  �/��    A�CZ      ��  �/��    A�CZ      ��  �/��V   A�CQ    �  $3��    A�CQ      ,�  3��H    A�CC     L�  B3��    A�CY      l�  @3��1    A�Cl       ��  R3���   A�CE��     ��  �8��    A�CX      ��  �8��V   A�CQ    ��  $<���   A�C�    �  �=��1    A�Cl       0�  �=���   A�CE��      T�  :?���   A�CE��     x�  �@��    A�CJ      ��  �@��    A�CJ       ��  �@���   A�CE��      ��  B���   A�CE��      �  �C��1    A�Cl       �  &���/    A�Cj       @�  5���    A�CP          d�  fP��   A�C    ��  RQ��0    A�Ck      ��  C��V    A�CQ     ��  OC��V    A�CQ     ��  �C��V    A�CQ     �  �C��V    A�CQ     $�  �C��V    A�CQ     D�  'D��V    A�CQ     d�  ]D��V    A�CQ     ��  �D��V    A�CQ     ��  �D��V    A�CQ     ��  �D��V    A�CQ     ��  5E��V    A�CQ     �  kE��K    A�CF     $�  �E��J    A�CE     D�  �E��S    A�CN     d�  �E��S    A�CN     ��  &F��S    A�CN     ��  YF��S    A�CN     ��  �F��S    A�CN     ��  �F��S    A�CN     �  �F��S    A�CN     $�  %G��S    A�CN     D�  XG��S    A�CN     d�  �G��S    A�CN     ��  �G��S    A�CN     ��  �G��H    A�CC     ��  H���   A�C�    ��  �K��.    A�C       �  �K��Q    A�CL      �  L��Q    A�CL     @�  6L��*    A�C      \�  DL��*    A�C      x�  �M��R    A�CM      ��  �M��    A�Cz         ��  XW��*    A�Ce       ��  �M���   A�CJ���    �  ~O��o    A�Cj      �  �O���    A�C�      @�  zP��?   A�CE�5      d�  �Q��r   A�CE�h     ��  �R���    A�C�      ��  �S���    A�CE��       ��  T���   A�CJ���   ��  �U��>    A�Cy      �  .V��S    A�CN     0�  bV��    A�CL      P�  TV��    A�CM      p�  FV��6    A�Cq      ��  \V��r    A�Cm      ��  �V��P    A�CE�F      ��  �V��C    A�C~      ��  �V��    A�CM      �  �V��4    A�Co      4�  W��w    A�Cr      T�  \W���    A�CE�{      x�  �W��!    A�C\      ��  �W��%    A�C`      ��  �W��    A�CM      ��  �W��    A�CL      ��  �W��O    A�CJ     �  �W��I    A�CD     8�  X��I    A�CD     X�  *X��*    A�Ce      x�  4X��    A�CL       ��  &X���    A�CE��      ��  �X��   A�C    ��  �Z��N    A�CI     ��  [���    A�C�     �  �[���    A�C�     <�  �\��+    A�Cf      \�  �\��/    A�Cj      |�  �\���   A�C�    ��  ,`���   A�C�    ��  �d��m    A�Ch     ��  "e��T    A�CO     ��  Ve��?    A�Cz      �  ve��h    A�Cc     <�  �e��n    A�Ci     \�  f��   A�C    |�  g��    A�Cz     ��  fg���    A�C|     ��  �g���   A�C�    ��  �i��    A�C    ��  �j���    A�C�     �  Dk��u    A�Cp     <�  �k��E    A�C@     \�  �k��    A�CL      |�  �k���    A�C�     ��  ,l��h    A�Cc     ��  tl���    A�C�     ��  Hm��U    A�CP     ��  ~m��U    A�CP     �  �m��E    A�C@     <�  �m��    A�CF      \�  �m���    A�C�     |�  �n��4    A�Co      ��  �n��    A�CU      ��  �n��*    A�Ce      ��  �n��    A�CZ      ��  �n��    A�CL      �  �n��Q   A�CL    <�  �p��*    A�Ce      \�  �p��    A�CZ      |�  �p��    A�CL      ��  �p���    A�C�     ��  Bq���    A�C|     ��  �q��r    A�Cm     ��  �q��i    A�Cd     �  >r��I    A�CD     <�  gr��    A�CU      \�  ar��   A�C    |�  Zs��R    A�CM     ��  �s��B    A�C}      ��  �s��5    A�Cp      ��  �u��"    A�C]      ��  �u��*    A�Ce       �  �u���   A�CE��     @�  tw��a    A�C\      `�  �w���   A�CE��     ��  qz��+    A�Cf      ��  |z��(    A�Cc      ��  �z��3    A�Cn      ��  �z��#    A�C^      �  �z��(    A�Cc      $�  �z��2    A�Cm      D�  �z��    A�CL      d�  �z��*    A�Ce      ��  �z��G    A�CB     ��  �q��    A�CI      ��  �z��    A�CI   $   ��  �q���    A�CI���v      �  %r��    A�CI   $   ,�  r���    A�CI���v      T�  7z��    A�CI      t�  &z��0    A�Ck      ��  6z��    A�CL      ��  (z��    A�CU      ��  "z��C    A�C~      ��  Fz��"    A�C]      �  Hz��0    A�Ck      4�  Xz��G    A�CB     T�  �z��1    A�Cl      t�  �z��    A�CU      ��  �z��    A�CU      ��  �z��J    A�CE      ��  �z��<   A�CE�2     ��  �|��    A�CI      �  �|���    A�C�     8�  2}���    A�C�     X�  �}���   A�C�    x�  ��-    A�Ch      ��  ,��+    A�Cf      ��  p���    A�C�      ��  �p��    A�CP          ��  $���&    A�Ca      �  *���H    A�CC      <�  R���e    A�CE�[      `�  ����M    A�CH     ��  º��&    A�Ca      ��  Ⱥ��<    A�Cw      ��  ���g    A�Cb     ��  ,���c    A�C^      �  p���6    A�Cq       �  ����Q    A�CL     @�  ����S    A�CN     `�  ���O    A�CJ     ��  ���.    A�Ci      ��  *���	   A�C    ��  ���L    A�CG     ��  @���S    A�CN      �  t���O    A�CJ      �  �|��+    A�C      <�  �|���    A�C�     \�  Y}��5    A�C      x�  r}��#    A�C      ��  y}��+    A�C      ��  �}��3    A�C      ��  �}��2    A�Cm      ��  �}���    A�C�     �  E~���    A�C�     ,�  �~���    A�C�     L�  p���    A�C�     l�  ���x    A�C      ��  V����    A�C�     ��  ����    A�C�     ��  ����    A�CO      ��  v���0    A�Ck        �����    A�C�     (  >���}    A�Cx     H  ����b    A�C]     h  ނ��[    A�CV     �  ���`    A�C[     �  Y���/    A�Cj      �  h���/    A�C       �  {����    A�CH��       9����    A�C�     ( ����3    A�C      D ����x    A�C      ` ���x    A�C      | s���3    A�C      � ����3    A�C      � ����x    A�C      � ����x    A�C      � Y���7    A�C       t���7    A�C      $ ����x    A�C      @ ���x    A�C      \ G���/    A�C      x Z���/    A�C      � m���D    A�C      � �����    A�C�     � F���K    A�CF     � q���"    A�C]       s���P    A�CK     4 ����%    A�C`      T ����    A�CU      t ����    A�CU      � ����    A�CS      � ����    A�CS      � ����I    A�CD     � ����"    A�C]       ����$    A�C_      4 ����    A�CR      T �����    A�C�     t o���+    A�C      � ~���2    A�C      � ����.    A�C      � ����/    A�C      � ����.    A�C        ˉ��+    A�C       ډ��#    A�C      8 ���.    A�C      T ���*    A�C      p ���.    A�C      � ���2    A�Cm      � %���2    A�Cm      � 7���/    A�C      � J���/    A�C       ]���    A�CQ      $ S���    A�CO      D G���    A�CO      d ;����    A�C~      � �����   A�CH��     � 9���6    A�C      � S����    A�C�     � ����    A�C�      b���[    A�CV     $ ����[    A�CV     D ؍��[    A�CV     d ���    A�CQ      � 	���    A�CO      � ����    A�CO      � ���D    A�C      � ���;   A�C6     0���;   A�C6    $ K���2    A�C      @ ����    A�CM      ` A����   A�C�    � V���*    A�Ce      � `����   A�C�    � �����   A�C�    � ���*    A�Ce       	 �����   A�C�     	 ����*    A�Ce      @	 �����   A�C�    `	 X���*    A�Ce      �	 b����   A�C�    �	 ���    A�CK      �	 ����1    A�Cl      �	 ���)    A�Cd        
 ���N    A�CE�D      $
 D���)    A�Cd       D
 N���N    A�CE�D       h
 x����   A�CH��     �
 ,���1    A�Cl      �
 >���)    A�Cd       �
 H����   A�CH��     �
 ����1    A�Cl       ���)    A�Cd       0 ����   A�CH��     T ����1    A�Cl      t ����)    A�Cd       � �����   A�CH��      � �����    A�CE��      � t���;    A�Cv      � �����   A�C�      J����    A�CE��       @  ����    A�CE��       d �����    A�CE��       � h����    A�CE��       � ����    A�CE��       � �����    A�CE��       � �����   A�CE��      ���d    A�C_     8 W����   A�C�     X ����    A�CE��       | �����    A�CE��       � z����    A�CE��       � 0����    A�CE��       � �����    A�CE��        �����    A�CE��       0 J����   A�CE��     T ���d    A�C_     t ���   A�C�     � �
���    A�CE��       � ����    A�CE��       � B���    A�CE��         ����    A�CE��       $ ����    A�CE��       H `���    A�CE��       l ���   A�CE��     � ���d    A�C_     � ����   A�C�     � ����    A�CE��       � X���    A�CE��        
���    A�CE��       < ����    A�CE��       ` r ���    A�CE��       � (!���    A�CE��       � �!���   A�CE��     � k)��d    A�C_     � �)��J    A�CE      �)��    A�CL      , �)��J    A�CE     L �)��W    A�CR     l ,*��Y    A�CT     � f*��    A�CM      � X*���    A�C�     � �*��U    A�CP     � +��W    A�CR      C+��W    A�CR     , z+���    A�C�     L �+��U    A�CP     l .,��W    A�CR     � e,��W    A�CR     � �,���    A�C�     � -��U    A�CP     � P-��W    A�CR      �-��W    A�CR     , �-���    A�C�     L =.��U    A�CP     l r.��W    A�CR     � �.���   A�C�    � 10���   A�C�    � �1���   A�C�    � 83���   A�C�     �4���   A�C�    , H6���   A�C�    L �7���   A�C�    l O9���   A�C�    � �:���   A�C�    � _<���   A�C�    � �=���   A�C�    � f?���   A�C�     �@���   A�C�    , vB���   A�C�    L �C���   A�C�    l }E���   A�C�    � G��S    A�CN     � 8G���    A�C�     � �G��;    A�Cv      � �G���    A�C}      H��r    A�Cm     , nH��r    A�Cm     L �H��%    A�C`      l �H���    A�C�     � ,I��3    A�C      � CI��Y    A�CT     � |I��i    A�Cd     � �I��m    A�Ch      J��n    A�Ci     ( `J��p    A�Ck     H �J��m    A�Ch     h �J���    A�C�     � �K��*   A�C%    � �L��,    A�Cg      � �L��\    A�CW     � �L��/    A�C       �L��/    A�C        M��/    A�C      < M��2    A�C      X 1M��2    A�C      t GM��2    A�C      � ]M��2    A�C      � sM��/    A�C      � �M��3    A�C      � �M��3    A�C        �M��3    A�C       �M��/    A�C      8 �M��3    A�C      T �M��/    A�C      p N��/    A�C      � N��3    A�C      � 2N��3    A�C      � IN��3    A�C      � `N��.    A�C      � rN��/    A�C       �N��/    A�C      4 �N��.    A�C      P �N��/    A�C      l �N��/    A�C      � �N��3    A�C      � �N��f    A�Ca     � -O��+    A�C      � <O��2    A�C      � RO��@   A�C;     rP��]    A�CX     < �P��7    A�Cr      \ �P��H    A�CC     | �P��f    A�Ca     � 4Q��a    A�C\     � uQ��g    A�Cb     � �Q��W    A�CR     � �Q��:    A�Cu       R��C    A�C~      < �S��    A�CP      \ R���    A�C�     | �R��Q    A�CL     � S��R    A�CM     � ^S��,    A�Cg      � jS��    A�CI      � XS��    A�CI        FS��P    A�CE�F      @ rS��    A�CI      ` `S��    A�CI       � NS��P    A�CE�F      � zS��    A�CI      � hS��    A�CM      � ZS��%    A�C`        `S��{    A�CG��o    ( �S��    A�CQ      H �S��    A�CU      h �S��$    A�C_      � �S��7    A�Cr      � �S��
    A�CE      � �S��    A�CQ      � �S��$    A�C_        �S��    A�CQ          , vT��=    A�Cx      L �T��     A�C[      l �T��    A�CK      � �T��    A�CL      � vT���   A�C�    � �U��|    A�Cw     � �R��    A�CX        �R��+    A�Cf      ,  �R��g    A�Cb     L  *S��    A�CZ      l  )S��    A�CH      �  �U��7    A�Cr      �  �U��-    A�Ch      �  �U��+    A�Cf       �  �U��K   A�CE�A     ! �V��G   A�CB    0! X��   A�C    P! Y��X   A�CS    p! JZ��    A�CZ      �! JZ��    A�CZ      �! JZ��    A�CZ      �! JZ��    A�CZ       �! JZ��    A�CZ          " FZ��    A�CJ      4" 6Z���    A�C�     T" �Z���    A�C�     t" |[���    A�C�     �" :\���    A�C�     �" �\��   A�C    �" �^���    A�C�     �" �_���    A�C�     # 0`���    A�C�     4# �`���    A�C�     T# �a���    A�C�     t# "b���    A�C�     �# �b���    A�C�     �# Tc���    A�C�     �# �c��    A�CH      �# �c��J    A�CE     $ d��    A�CU      4$ �c��f    A�Ca     T$ Dd��J    A�CE     t$ nd��.    A�Ci      �$ |d��)    A�Cd      �$ �d��E    A�C@     �$ �d��}    A�Cx     �$ e���    A�C�     % �e��W    A�CR     4% �e���   A�C�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �@     �}F     �G     ��������        ��������        J     �J     �J     �J     �-J     �/J     EJ     &cJ     ��J     1�J     ��J                     �G     �G     B�F     ��F     D G     8G     �G     �G                                     F(H     F(H     F(H     F(H     F(H     F(H                     tH     �H     �H     H     bH     vH                                     F(H     F(H     F(H     F(H                                                            1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `  @�K     ��K     ��K     H�K     GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o      �             ]@     �      �@     I       :@     2       l@     -       �@            �@     "       �@     -      �@     "       @     �       �@     �       t@     8                       ,    �       �@     �                      ,    �C       `@     �                      ,    �      p�@     2                       ,    ��      ��@     &                       ,    `�      ��@     V�                      ,    Xm      @�A     p^                      ,    �E      �B     �o                      ,    �U      p�B     �$                      ,    i�       �B     R5                      ,    �o      ��B     %                      ,    �      �C     a                      ,    �R        C     U$                      ,    ��      `DC     �B                      ,    �        �C     ��                      ,    >	      �3D     *�                      ,    +N
      ��D     �<                      ,    ��
      �E     S*                      ,    P=      0.E     S                      ,    �      �HE     �0                      ,    �      `yE     �                      ,    |�      P�E     *�                      ,    �Z      �/F     &                      ,    �      �6F     �                      ,    �      �8F     ]                      ,    =�      @RF     �                       ,    ��      �UF     >                       �   ��      ;VF     �      YF            &YF     \       �YF     �       ZF            6ZF     #       ZZF            vZF     V       �ZF     )       �ZF            [F     )       ,[F     (       T[F     ,       �[F            �[F            �[F     4       �[F     E       \F     C       T\F     &       z\F     *       �\F     J       �\F     �       �]F     �       [^F     U       �^F     �      O`F     (       x`F     �                       ,    C�      ,aF     A                       �   l�      maF           YF            &YF     \       �YF     �       ZF            6ZF     #       ZZF            vZF     V       �ZF     )       �ZF            [F     )       ,[F     (       T[F     ,       �cF     )       �cF            �cF     )       �cF     (       dF     ,       �[F            �[F            �[F     4       �[F     E       \F     C       T\F     &       :dF     4       ndF     E       �dF     C       �dF     &       z\F     *       �\F     J       eF     *       FeF     J       �\F     �       �]F     �       �eF     �       afF     �       [^F     U       �fF     U       �^F     �      RgF     �      O`F     (       x`F     �       �hF     �                       ,    �      �iF     �                      ,    m      *kF     Q                       �   �      {kF     #      �}F             �}F     �       l~F     �      YF            &YF     \       �YF     �       ZF            <�F     6       r�F     Q       ÀF            րF     B       �F            6ZF     #       ZZF            vZF     V       .�F     M      {�F     L      ǅF           �cF     )       �cF            �cF     )       dF     ,       �F     )       �F            ��F     �       ��F     )       ��F     (       ܉F     0       �F     +       �[F            �[F            :dF     4       ndF     E       �dF     &       7�F     E       |�F     h      �F     �      ��F     #      eF     *       ��F     }       4�F     2       f�F     '       ��F     �       V�F     �       �F     O       b�F            x�F     I       F     �       ��F     �       r�F     X       ʙF     D      �F     �       �F     L       N�F     �       �eF     �       �F     �       ��F            ��F            ��F            ؝F     a      9�F            X�F     �      �F            ��F     j       `�F     (       ��F            ��F     7      ݤF            ��F     7      4�F     a      ��F            ��F     �      @�F     d       ��F     j       �F     7      F�F     7      ~�F     K       ɮF     W        �F            6�F            T�F     1       ��F     �      I�F            f�F     H       ��F            εF            �F     V      D�F            Z�F     H       ��F            ��F     1       �F     �      ��F            ҿF     V      (�F     �      ��F     1       �F     �      ��F     �      B�F            Q�F            `�F     �       �F     �      ��F     1       O`F     (       �hF     �                       \   Oi      ��F           &YF     \       ZF            ��F           ��F     0       6ZF     #       ZZF            �F     R       l�F            �cF     )       �cF            �cF     )       dF     ,       �[F            �[F            :dF     4       ndF     E       �dF     &       eF     *       �eF     �                       �   ?�      ��F     <	      r�F     Q       ÀF            րF     B       �F            YF            &YF     \       �YF     �       ZF            <�F     6       (�F     *       6ZF     #       ZZF            vZF     V       �F     R       R�F     S       �cF     )       �cF            �cF     )       ��F            ��F            ��F     6       dF     ,        �F     r       l�F            r�F     P       ��F     C       �F            �F     4       L�F     w       ��F     �       J�F     !       l�F     %       ��F            ��F            ��F     O       �F     I       �[F            �[F            :dF     4       ndF     E       M�F     I       �dF     &       ��F     *       ��F            �F            ��F     �       ��F     )       ��F     �       eF     *       ��F           |�F     h      ��F     (       �eF     �       �hF     �       ��F     N       4�F     2       f�F     '       ��F     �       V�F     �       �F     O       b�F            x�F     I       F     �       �F     �      FeF     J       ��F            �F     L       ��F            ��F            ؝F     a      9�F            X�F     �      �F            ��F     j       `�F     (       ��F            ��F     7      ݤF            ��F     7      ��F     �       r�F     X       ʙF     D      �F     �       N�F     �       afF     �        �F            6�F            T�F     1       ��F     �      I�F            f�F     H       ��F            εF            �F     V      D�F            ��F            Z�F     H       ��F            4�F     a      ��F     �      @�F     d       ��F     j       �F     7      F�F     7      ~�F     K       �fF     U       ��F     1       �F     �      ��F     �      B�F            Q�F            ��F            ��F     1       `�F     �       �F     �      �F     �      ҿF     V      RgF     �      ��F     1       O`F     (                           ��                      �   W�      $�F     �       YF            &YF     \       �YF     �       ZF            r�F     Q       ÀF            րF     B       �F            6ZF     #       ZZF            vZF     V       �G     "       G     *       ,G     �      �cF     )       �cF            �cF     )       dF     ,       �F            ��F     �       ��F     )       �G     a       *G     �      �ZF     )       �ZF            [F     )       T[F     ,       	G     +       �F     +       4G     (       ��F     (       \G     3       �G     #       �G     (       �G     2       G             G     *       JG     G       �G            �[F            �[F            �G            �G     0       �G            �G            :dF     4       ndF     E       �dF     &       |�F     h      �[F     4       �[F     E       T\F     &       
G     C       �F     �      NG     "       pG     0       �G     G       �G     1       G            4G            eF     *       4�F     2       f�F     '       ��F     �       V�F     �       �F     O       b�F            x�F     I       F     �       z\F     *       NG     J       ��F     �       r�F     X       ʙF     D      �F     �       �F     L       N�F     �       �G     <      �G            �eF     �       ��F            ��F            ��F            ؝F     a      9�F            X�F     �      �F            ��F     j       `�F     (       ��F            ��F     7      ݤF            ��F     7      �\F     �       �G     �       4�F     a      ��F            ��F     �      @�F     d       ��F     j       �F     7      F�F     7      ~�F     K        �F            6�F            T�F     1       ��F     �      I�F            f�F     H       ��F            εF            �F     V      D�F            Z�F     H       ��F            ~G     �       ��F     1       �F     �      ��F            ҿF     V      ��F     1       �F     �      ��F     �      B�F            Q�F            `�F     �       �F     �      RgF     �      G     �      ��F     1       O`F     (       �hF     �       �G     -       �G     +                       �   CT      G     /;      r�F     Q       ÀF            րF     B       �F            YF            &YF     \       �YF     �       ZF            <�F     6       (�F     *       4VG     &       ZVG     H       �VG     e       WG     M       VWG     &       |WG     <       �WG     g        XG     c       �XG     6       �XG     Q       YG     S       `YG     O       �YG     .       �YG     	      �ZG     L       4[G     S       �[G     O       6ZF     #       ZZF            �[G            vZF     V       �F     +       �[G     *       \G     �      �bG     *       
cG     �      	G     +       �iG     *        jG     �      �F            ��F     �       ��F     (       �cF     )       �cF            �cF     )       ��F     6       dF     ,       �pG     *       �pG     �      �[F            �[F            �wG            �wG     1       xG     )       .xG     N       |xG     )       �xG     N       �xG     �      �|G     1       �|G     )       (}G     �       �G     1       2�G     )       \�G     �      �F     �      :dF     4       ndF     E       M�F     I       �dF     &       4�G     1       f�G     )       ��G     �      g�G     �       �G            d�G     ;       ��G     �      z�G     �       T�G     �       *�G     �       �G     �       ڔG     �       ��G     �       ��G     �      ?�G     d        G     *       ��G     �      ~�G     �       X�G     �       .�G     �       �G     �       ިG     �       ��G     �       ��G     �      C�G     d       ��G     �      ��G     �       \�G     �       2�G     �       �G     �       �G     �       ��G     �       ��G     �      G�G     d       4�F     2       f�F     '       x�F     I       ��F     �       r�F     X       �F     O       ʙF     D      �F     �       �F     L       F     �       N�F     �       eF     *       ��F           ��G     �      ��G     �       `�G     �       6�G     �       �G     �       ��G     �       ��G     �       ��G     �      K�G     d       ��G     J       ��G            
�G     J       T�G     W       �F     R       ��F            ��G     Y       �G            �G     �       ��G     U       �G     W       �G     G       c�G     W       ��G     �       Y�G     U       ��G     W       �G     W       \�G     �       ��G     U       P�G     W       ��F            ��F            ݤF            4�F     a      ��F            ��F     �      �F            @�F     d       b�F            ��F     j       `�F     (       ��F            �F     7      ��F            F�F     7      ��F     j       ��F     7      ��F     7      ~�F     K       �eF     �       �hF     �       ��F     N       ��G     W       ��G     �       ��G     U       ��G     W       I�G     �      ��G     �      ��G     �      8�G     �      NG     J       ��G     �      ��G     �      0�G     �      ��G     �      w�G     �      �G     �      ��G     �      f�G     �      D�F            ��F            ��F     1       �F     �      ��F            Z�F     H       εF            ��F            ҿF     V       �F            9�F            f�F     H       6�F            �F     V      FeF     J       �G     �      ��G     �      ^�G     �      ��G     �      O`F     (       �G     �       ��F     1       `�F     �       �F     �      Q�F            B�F            I�F            T�F     1       �F     �      ��F     �      afF     �       ~G     �       �fF     U       RgF     �      G     �                      ,    O$      ��G     �                      ,    �6      ~H                           |   �:      �H     �      YF            H            .H     ,       ZH            hH            vH     P       �H            �H            �H     P       2H            @H            RH     %       xH     {       �H            
H            $H     $       HH     7       H     
       �H            �H     $       �H                            L   Z      �H     �       �H     =       �H             H            $H            6H     �      �H     |       <H     7       tH     -       �H     +       �H     K      H     G      bH           vH     X      �H            �H            H            .H            NH                            �   	p      nH     s      YF            &YF     \       �YF     �       ZF            6ZF     #       ZZF            vZF     V       �cF     )       �cF            �cF     )       dF     ,       �cF     (       �[F            �[F            :dF     4       ndF     E       �dF     &       �dF     C       eF     *       FeF     J       �eF     �       afF     �       �fF     U       RgF     �      O`F     (       �hF     �                       �   5�      �'H     B      YF            &YF     \       �YF     �       ZF            <�F     6       6ZF     #       ZZF            vZF     V       �ZF     )       �ZF            [F     )       $)H     )       T[F     ,       �[F            �[F            �[F     4       �[F     E       M)H     E       T\F     &       z\F     *       �)H     }       �\F     �       *H     �       �*H     W       +H     �      O`F     (       x`F     �                                       �       +	    W                   a  5   �  3  H   �  t  [   �i -  n   �i 4  	�   �  -  x  �   int �   X  �  �n     u   h  �     )   j  <   g  O   7  b   �  4�   �  P  ��  �    �  �   bpp 	�   �  �   
 �    ^� �n   	S  �
  &E E
  (	�  x 	�    y 		�   ��  	�   �  	�   �  	�   E? 	
�   B� 		�  �  	

�     
�   `  	  �  '  x 	�    y �    �  	  '  �  r  r �    g �   b �   a �    �  8  "�  �  �  #�   �  $�   ݖ %�   x  &�   
 �  �  n    �  �  '~  ()�   �  �  *�    ��  +
�   �  ,
�   E  -�   bpp .�   _  /�   �  0�   �  1
�   �  2
�   �  3�    �	  4�   $ �   5�  �
  �  $  
h  
�  |0  /  x �    y �   ��  �   �  �   ?1  �   �  /  �  �   l`  �  t2  	  (      �  ?  n   _ 2  �  {S @�  g
  �      	\  v  #	\  �  &	\  |
  )	\   h  ,	\  (�  -	\  0�	  2�   8�  5�   < 
�  �
  8"K    K�  
�  �  L�  �  M�  (�  Y  3  �    h  �   msg �   �U  �   �
  �     �  
  �  �q  
�  {  ��  �  ��   �  ��      ��   �	  [   �  A"�  
�     �  R   �h   �� �  �N �.  �6  �P   �  X  
  h  .  �  �      m:  
@  P  �  h   �  �\  
b  h  �  �  �   �   h   �  �"�  
�  �   PH-  2�  J�   �  Kn   pos Ln   �  NS  SF  OS   �1 P_  (=9 Q�  0R�  S�  8y�  T�  @�� U�  H �  �S  �\ ��   m  �h   o  �-  �  �k  
q  n   �  �  n   �  n    
5   2  �  
�  �  �     :�   �  L�  x N�   y O�   )  Q�  B   w1  M   y�   }  y�  V  z�  /  z�   t
  |�  k	  (�  �  [    ��  [   �  	�   B� 
�  L  H     5   s  5   v	  h    �  =  �  (Q,	  �  S�    Z�  T�   �  V,	  s  W�  [  X2	  ?1  Z�     
�  
�     \�  =  [   ��	  �   M
  pmoc5  stib	  ltuo|  tolp 	  �E	  �  ��  �
  ��   �  �H   �  ��   
  �[   �  ��   �  �     ��	  
�	  
  h   �  �.
  �U  �h     ��	   %  �
  �  $H
  
N
  �  +�
  �� -;
   �@ .;
  �U  /h   �  D�
  �; F;
   ��  G;
   L  I�
  �
  @<>  ��  >�   �  ?�  ~  A�  �  B�  �  C�   5  E�  (B  F�  0�  G�  8 �	  I�
  
   s�  �  u�	   ��  v�	  �  x�  �
  z�  (  {�   �  }K  �  �#�  
�  k  �  �"�  
�  %  K  � �  
�  �  ��  �   �	   �  �	  O  �	  C  �	  �  �	   d> �  (A  �  0T  �	  8  �  @�  !�	  H�  "�  PE-  $.
  X�!  )1  h:  +�	  �  ,�	  ��  -�	  ��  .�	  ��  0�	  �  1�	  �U  3�	  ��  4�	  �)�  6  ��  7�  ��� 8h  �K1 <�  �R�  =�  �Jy  >�  �%  @�
  ��	  B.
  �    Ch  ��8  E�  � L   �  
�    Xm  �  o�   E-  p.
  N qU  �8  r�  P �  $%  
  �  0\h  k  ^�   �  _�  �@ `  �^ a�	  E-  b.
   N d>  0�  e�	  pR  f�	  x�  g�  �ߣ  i�	  ��I k�  ��  l�	  �h  m�	  ��S  o8	  �4  q�	  �8  rb  �   th    �  u�    �  w�   o  x�   �L zh    �8  |z  ( �
  F#u  
{  W  A�  �  C�   = D�    E�	  d  F�	   �  [   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  #   `)�  
�  �   
�	  
�  
h  �
  �)�  
�  �   ~	  8HU  �
  J�	   (  K�	  �� M�	  �� N�	    P�  �  Q�   �  R�  (�  S�  0 y  U�    �$o  
u  �  �  �)�  
�     �   �  n    !�  �  	��K     �
  �B�  `  C�   ��  D?  pos E'  ��  F�  � t "fb I
�  	��K     !�   JP  	��K     !�  K�  	��K     �   R  n    !K  MB  	��K     !�  N'  	��K     !�  O�  	��K     !@  P�  	��K     !p  Q'  	��K     !d  S�  	��K     !  U�  	��K     !k  W�  	��K     !  X	�  	��K     !�  sr  	��K     !�  t�  	 �K     !�  v�   	(�K     #    $wT  �  |  �     $F  �  �  �    �    $��  !�  �  �     $,  *+  �  �    (   $�  ; 
  �  �    (   %d  L�  (    !    [    %�  P�  (  :  E    [    $B  Z  Z  j    [   (   %�  dN  �   �  �     %�  h�  (  �  �    [    %�
  }G  (  �  �     %[  ��  (  �  �     &�  ��   &0  ��  'num �[   (T (   
Z    
�  #   �  &�@ 	�   &�� 
�  'obj (  )�  �   w  }  �   (T (   
.  �  !�  wZ  	0�K     !�  x(  	H�K     *Z  h  +�  �@            �,�  �    -�  #  -0  �   ./D� �    0�  �  .  t@     8       �d  1�  �X2�  E  3�   4�  �@     )       5�  �h  6M  �@     >       ��  7<  ��   �l7  ��   �h 8!  �  �@     �       �	  9�  #  �X:pos P[   �T;�� S�  �h<2@     8       =i U[   �d  >�  (  @     �       �S  9�  #  �H:obj *(  �@;D� +�  �X ?e  d  n  -�  �   @S  �  �  �@     "       ��  1d  �h >�  �  �@     -      �7  9�  #  �H:pos h[   �D;�� n�  �h=obj r(  �XA�@     	         ;/� j(  �P <@     8       =i p[   �d  >�  V  �@     "       �r  9�  #  �h:pos L[   �d 8j  �  �@            ��  9�  #  �h ,g  �  �  -�  #   @�  �  �  l@     -       ��  1�  �h B�  ��   
@     �
      �;  ;C
  ��  �H;�  ��  �@;�  ��   ��;�   ��  ��;�  �;  ��;   ��   ��;�N  ��   ��A�@     O       �  =err �	�   �� <&@     s      Cmsg \Y  ��~A]@     7         Ci 
�   �l<o@            Cwin (  ��  A�@     
      �  Ci  �   �h<�@     �      Cwin !(  ��<�@     �       D�  *Y  ��~Dz  ,�   �dD�  -�   �`   A�@     �       �  D�  JY  ��~Dz  L�   �\D�  M�   �X A@     �       �  D�  aY  ��~ <@     &       Ci ��   �T<(@            Cj ��   �P    
�  E�  ��
  G@     �      ��  :win �(  ��;t  �'  �� Ef  ��  e@     �      �Y  ;�  ��   �L<�@     �      =j �
�   �l<�@     �      ;�  ��  �k;�  �?  ��~;  ��  �XA�@     D       5  =i ��   �d <O@     �       =win �(  �P    EQ  z'  ]@           �  ;�  {�   �T<�@     �       =i ~
�   �l<�@     �       ;�  	�  �k<�@     }       =j ��   �d<�@     e       ;�  �?  ��~;  ��  �X     
?    ?  7  A  -�  !   @&  �  d  :@     2       �m  17  �h F�  �  '  �@     I       ��  :l 0�  �h:r E�  �` G3   &   /  �  g&  $"  �@     �        X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �	  	N   �  B"]  c     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  Q  -      n�  �  �  Q  U    �  ��  �  U     Q  -   -   U    �  �")  /  �   PJ�  2�  L,   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S9  0R�  UQ  8y�  V,  @�� W,  H �  ��  �\ �-   m  �U    o  ��  �  �    @   ,    @   ,  @    2  �  2  F  L  W       :-   �  J�  x LW   y MW   )  Oc  	�  B   s�  M   uW   }  uW  V  vW  /  vW   t
  x�  k	  (e  �  N    ��  N   �  	G   B� 
,  L  0    2  s  2  v	  U     �  �  	e  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     �  )    Yw  �  =  N   �7  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "Q  W  �  %  <�  x >)   len ?0  *� @2   %  B\  	�    `�  �  �  G   G   �  U    �  �  q�  �  G     G   G   U    �      ,  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  �  0R   �U   8�  ��  @ r  �  �  �,  	�  �   �  �  G   �  U   �   D  �      #  D   �  ?0  6  K  D  ,  @    �  YX  ^  G   w  D  @   U    s  ��  �  G   �  D  �   �  W  0�  �  �7   e� ��  �� �#  �� �K  �� �w   �� �  ( �'  ��  �!  l2  �  �,  �  -  �2  	3  ?  �  ��   	J  �
  �)  �  �0  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   b   �	  xx ��   xy ��  yx ��  yy ��   a  ��  		  z'  �J	  m  �D   ss  �s   �  �	    �d	  j	  u	  U    �  ��	  �U  �U      �W	   %  �u	  �  $�	  �	  �   �	  �� "�	   �@ #�	  �U  $U    �  7$
  �; 9�	   ��  :�	   L  <�	  N   �t  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=�  ��  ?W   �  @W  ~  BW  �  CW  �  DW   5  FW  (B  GW  0�  HW  8 �	  Jt  
   sU  �  u[   ��  v[  �  xW  �
  zW  (  {W   �  }   �  �#o  u  k  `	�$  R�  	�Q   (  	�s  |  	�s  �  	�s  �  	�  �  	�H!  v  	�$
  �  	��  (�%  	�$  07&  	�X!  8G   	�s  X �  �"1  7  h  	p  �M 	/!   k  	b  R�  	Q   �  �"}  �  %  8	;�  �� 	=5!   �M 	>0    	?$
   r$  	@T  0 5  �$�  �  %  �	N  �� 	5!   �M 	B!  �  	7   �  	�  (�� 	
D  h�� 	w  p�� 	Q  x K  � [  a  �  �,"  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9s  8  :�  @�  <s  H�  =�  PE-  ?�	  X�!  D�  h:  Fg  �  G[  ��  H[  ��  I[  ��  K[  �  L[  �U  N[  ��  O[  �)�  Q|  ��  R"  ��� S�  �K1 Wp  �R�  XQ  �Jy  Y  �%  [$
  ��	  ]�	  �    ^U   ��8  `  � L   /  5    X�|  �  �N   E-  ��	  N �t  �8  ��  P �  *%�  �  �  0t�  k  vb   �  wN  �@ x|  ݖ y  E-  z�	   N |�  0�  }�  pR  ~�  x�  �  �ߣ  �7  ��I �e  ��  �s  �h  �s  ��S  ��  �4  �  �8  ��  �  �U    �  �-   �  �W  o  �W  �L �U    �8  ��  ( �
  L#�  �  W  H3  �  JN   = K�    Lg  d  Mg   �  N   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  3  #   g)    �   �	��  =  	�	   L  	��   $  	�s  0�  	��  8m  	�#)!  h�  	�   pآ  	�7  tG   	�s  x J  U  �  �
  �)�  �  �   H	��  �  	�U    "  	�|  �!  	�t   ~	  8ft  �
  hg   (  ig  �� k�  �� l�    nW  �  oW   �  pW  (�  qW  0 y  s�    �$�  �  �  0
'�  �N  
)s   ?1  
*g  }0  
+s  i/  
,s  � 
-	   �  �)�  �     H	�Y  ��  	�T   ?1  	�  (  	�  4  	�	  \  	��  0  	�U   @ +!  �  tag �   �U  �   �  Y  �  `  N   
�  w%   }#  �&  h  �  &     
�  E   9
1  � ;
�   ��  <
�  �  =
�  �  >
  �#  ?
   �  L
(>  �  �  N   �|  :   �   ^$  1  �!  �!   :  �D  �  ��  �#  ��  �  �  �  $   I$  ��  �  �  $   �&  ��  �  �  �  $  �   �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  ��  @ V  R  ��  	�  x  =d	  H  E#�  	�  �  @J-  �  L�   �  M7  �� O�  .� P�  �  Q   �  R�  (�!  S�  08'  TE  8   W!9  ?  -  (l�  k  nb   �M o�  ߣ  p7  �  q�   �  k  )�  �  �  �  -  |   w   .�  �  �  -   �  1�  �  �  -  �  �   	  K  6  	    -     �  �  :+  1  �  E  -  -   �  >�  "  Y]  c  �  �  �  |  |  �   �  _�  �  �  �  �  |  �  �   $  f�  �  �  �  |     �  l�  �  �    �  �  �   #  x�l  �� � �   �  � 7  H  � Q  P�  � �  X9!  � �  `l� � �  h  � l  p     �  	r  �  H
2�  �S  
4�   �  
5�  (  
6�  04  
7  88  
8�  @ �  
:�  �  �
=T  R�  
?Q   �  
@  n  
A  �  
B  1$  
C  2�  
E�  �� 
F�  `�L 
HU   � �  
J`  �  P   r  x  �  �    N  s  s  �   �  &�  �  �  N   �%  *�  �  �  �  "   �%  -�  �  �  "   {  1    �    |   �  4#  )  4  |   l  8@  F  �  Z  "  1   �  <f  l  �  �  "  �   �  @�  �  �  �  |  "    7   �  G�  �  �  �  N      �   �'  N�  �  �    N     �  S    �  ;  N      7  ;   �  &  ��  �� ��   i'  ��  H   ��  P  ��  X�A �f  `Y ��  h�#  ��  p�  ��  x�  ��  �  �  ���  ��  �U�  ��  ��!  ��  ���  �  ��  �4  �&  �Z  �   �A  	  �&  �<  A  �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }B  �  U'�  �  m  D   t   �  v�   A  w�  �  x�  &  y�   !  {�  �  �#   )   �  B   �    B    J	  �  �T   Z   j   �  B    �'  �v   |   �  �   �      �       �!  �   ��  )    ��  )H   �  )j    }  �   	�   O  ;!  _� =%!   ݰ  >%�   �   �  @�   !  �  �  	7  r  $  X!  @    �  h!  @    �  	�%  
�'  +  
;  +  
�  +  
V'  +  
6  +  
   +  
1  +  
�%  	+  
�  
+  
�'  �  
�  �  
!  �  
|  ~  
�  ~  
!   ~  
*  ~  
  �  
�  �  h"  ]"  @    	M"  �  	b"   /(  J!]"  	�-H     !�  d�  0@     &       ��"  "k  d!b         #R�  fQ  T   R   $>@     �%  �"  %U�U &F@     �%  %Us   !i  @�  �@     �       �$  "j  @"$  �   w   #� B�  �   �   #R�  CQ  b  Z  '#%  �@      �@     $       Y�#  (0%  �  �  )�@     $       *<%  +H%  �  �  &�@     �%  %Uv    ,�@     �%  $�@     �%  �#  %Us %T|  ,�@     $  &@     �%  %Us   b  -�  ��@     �      �%  .k  �*b  Z  R  /env ��  �  �  /p ��  �  �  /q ��  �  �      �%  ��| n  �%  ��} z  �%  ��~/i �
G   %    $@     �%  �$  %U	-H      &@@     �%  %Us %Tw %Q��}%R��~  �   #%  @   � 0�  �U%  1k  �'b  2� �$�  3cur �$U%   h"  4#%  �@     3       ��%  (0%      *<%  +H%  b  Z  &�@     �%  %Uv   5F'  F'  85'  '  	�5�  �   5�  �  	�5+  +   6�  �  M5K  K  	_ [l  U  x�  �4  $"  `@     �        Q�i :G  �@   QX  ^� �-   yint Q�i z${S @�   	g
  �    	   	G   	v  #	G   	�  &	G   	|
  )	G    	h  ,	G   (	�  -	G   0	�	  2S   8	�  5S   < �   Q�  .�   �
  8"c   c  K  �   c�  L  c�  M  QS  �9  A  1@   Q  2-    Q-  �[  �d  Q�  >   S   .k  �	  	Z   �R  l@   J)  m-   �  B"�  �  $   ��  	R   �a    	�� ��  	�N �  	�6  �@   �  Y  
  a     �  @      n*  0  5@  �  a    �  �L  R  a   p  �  @   @   a    �  �"|  �  �   PJ  2�  L   �  M-   Fpos N-   �  PC  SF  QC   �1 RO  (=9 S�  0R�  U�  8y�  V  @�� W  H i�  �C  j�\ �@   jm  �a    o  �  �  �[  a  -     p  -     -    �  Q�  2  �  �  5�  p     :@   $�  J�  ]x L�   ]y M�   )  O�  .�  $B   s-  	M   u�   	}  u�  	V  v�  	/  v�   t
  x�  ^�J  Z   ��  
�@   
�\  
0  
35  
G5  
8  
>  
�[  
F;   �X  �9  k	  (  �  Z    ��  Z   �  	S   B� 
  L  d    �  s  �  v	  a     �  �  .  �  (N�  �  PQ   Z�  QQ  �  S�  s  T�   [  U�  ?1  WS     �  Q    Y  .�  l<  ��  �  S   �  �  a    �  G  �  �:  '�  �  S     �  �  a    /\  G    S   7  �  �  �  a    oF  0t�  ��  v�   ��  w�  F� x�  �� y  �� {S    � |�  ( V  ~7  .�  R=  Z   ��  
�   3M
  pmoc35  stib3	  ltuo3|  tolp 	  ��  b   "  
  X�  %  <F  Fx >Q   Flen ?d  *� @�   %  B  .F    `e  k  5�  S   S   �  a    S  �  q�  �  S   �  S   S   a    �  �  �  5�  S   S   a    �  `�l  �  �l   �% �r  ?1  �S   �&  �X  !  �X   I  ��  ()  ��  0R   �a   8�  �-  @   x  {�  ��  .y  �   �  �  S   �  a   �   �  �  �  �  5�  �   �  ?�  �  5�  �    -    �  Y	  	  S   *	  �  -   a    s  �7	  =	  S   Q	  �  Q	   �  W  0��	  �  ��   e� ��  �� ��  �� ��  �� �*	   �� ��  ( �'  �W	  �!  l�  �  ��	  Q�  -  ��  .�	  �	  �L  �}  �  ��   .	
  �
  �Q  �  �d  �  �S   
  �Z   �  �@   \#  �-   )H  @   �   @   �  ,S   \&  7a   �0  DG   �H  Q4   b   ��
  Fxx �o
   Fxy �o
  Fyx �o
  Fyy �o
   a  ��
  .�
  z'  �0  m  ��	   ss  �2
   �  �    �J  P  5[  a    �  ��  �U  �a      �=   %  �[  �  $�  �  �   �  �� "�   �@ #�  �U  $a    tT   �  �  �  7  �; 9�   ��  :�   L  <�  |Z   5�m  
�   
  
�  
  
$  
K  
�%  
�%  
,#  
�  	
   

�$  
e#  
�  
�  
[%  
A#  
z"  
6  
�  
�  
�   
�"  !
Y  "
�  #
�#  $
_"  %
�  &
�"  '
H!  (
�  0
v  1
�  @
  A
l  Q
�   R
7  S
�$  T
�#  U
  V
   W
�  X
R  `
	  a
a  b
�"  c
�'  p
�  �
�  �
	  �
�  �
M  �
�  �
v  �
�  �
'  �
H%  �
  �
e!  �
�  �
'%  �
�   �
�  �
�  �
�$  �
�  �
g  �
  �
P  �
�  �
�  �
�  �
  �
�$  �
�&  �
N  �
�   �
  �
�  �
;$  �
�  �
#  �
�"  �
�  �
G  �
�  �
0  �
1  �
P  �
C&  �
:  �
_  �
A  �
^  � �
  @=�  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  Jm  
   sN  �  u
   ��  v
  �  x�  �
  z�  (  {�   �  }�  �  �#h  n  _k  `�  R�  ��   (  �2
  |  �2
  �  �2
  �  �>
  �  ��'  v  �  �  ��  (�%  �  07&  �(  8G   �2
  X �  �"*  0  h  i  �M �'   k  [  R�  �   �  �"v  |  %  8;�  �� =�'   �M >6"    ?   r$  @k  0 5  �$�  �  %  �G  �� �'   �M �'  �  �   �  �  (�� 
�  h�� *	  p�� [  x K  � T  Z  �  �,  �   .J
   �  /J
  O  1J
  C  2J
  �  4J
   d> 6�  (A  7�  0T  92
  8  :�  @�  <2
  H�  =�  PE-  ?�  X�!  D-  h:  F&
  �  G
  ��  H
  ��  I
  ��  K
  �  L
  �U  N
  ��  O
  �)�  Qu  ��  R  ��� S�  �K1 Wi  �R�  X�  �Jy  Yp  �%  [  ��	  ]�  �    ^a   ��8  `  � L   (  .    X�u  �  �G   E-  ��  N ��  �8  ��  P �  *%�  �  _�  0t�  k  v[   �  wG  �@ xu  ݖ y>
  E-  z�   N |�  0�  }o
  pR  ~o
  x�  �  �ߣ  ��  ��I �  ��  �2
  �h  �2
  ��S  ��  �4  �>
  �8  ��  �  �a    �  �@   �  ��  o  ��  �L �a    �8  ��  ( �
  L#�  �  W  H,  �  JG   = K�    L&
  d  M&
   R�  Z   ��  
�   3�  bmys3=  cinu3�  sijs3w    bg3O  5gib3p  snaw3M  ahoj3�    bg3�  sijs3�    bg3q  5gib3�  snaw3�	  ahoj3  BODA34   EBDA3�	  CBDA3  1tal3�  2tal3   nmra �	  ,  (0  O�  #   g)    �   ���  =  ��
   L  ��   $  �2
  0�  �$  8m  �#�%  h�  ��	  pآ  �k  tG   �2
  x 	
  N  �  �?  dZ  �
  �)�  �  �   H�  �  �a    "  �-  �!  ��   ~	  8f�  �
  h&
   (  i&
  �� ko
  �� lo
    n�  �  o�   �  p�  (�  q�  0 y  s    �$�  �  $�  0'�  	�N  )2
   	?1  *&
  	}0  +2
  	i/  ,2
  	� -�
   �  �)  	     H�l  ��  �k   ?1  �>
  (  ��	  4  ��
  \  ��  0  �a   @ +!  �  Ftag V
   �U  �
   �  l  �M  @W#  ?1  Y>
   �I  Z�	  N  [J
  SF  \�  Jy  ]p   K1 ^  (G  _2
  0G  `#  8 �  �O  b�  .)  R`  Z   
s  
w%   
}#  
�&  
h  
�  
&     
;  E   9
�  � ;
s   ��  <
J
  �  =
J
  �  >
>
  �#  ?
>
   �L  A
�  �  L
(�  �  R�  Z   �-  
:   
�   
^$  
1  
�!  
�!   :  ��  R�]  Z   ;`  
�>   
+V  
�H   �  ��
  �#  �x  ~  |
  �     I$  ��  �  5�     �&  ��  �  `  �    �   �   $�!  H�Y  	�  �V
   	S"  �J
  	   �Y  	�"  �o
  	�  �o
   	;  �r  (	%  �l  0	�   ��  8	��  ��  @ 
  R  ��  ._  x  =J  RT  Z   ��  
�L   
3A  
�<   �.  �}  H  E#�  .�  $�  @J7  	�  LJ
   	�  M�  	�� O�  	.� P�  	�  Q)   	�  R�  (	�!  S  0	8'  TO  8   W!C  I  $-  (l�  	k  n[   	�M o�  	ߣ  p�  	�  q�   �  k  )�  �  |
  �  7  u   w   .�  �  5�  7   �  1�  �  5�  7  �  �      K  6    5#  7  #   -  �  :5  ;  |
  O  7  7   �  >�  "  Yg  m  |
  �  �  u  -  �   �  _�  �  |
  �  �  u  �  �   $  f�  �  5�  �  u  #   �  l�  �  |
    �  V
  �
   $#  x�v  	�� � _   	�  � �  H	  � [  P	�  � �  X	9!  � �  `	l� � �  h	  � v  p �	    �  $�  H2�  	�S  4�   	�  5�  (	  6�  0	4  7>
  8	8  8�  @ �  :�  �(  :�  �  $�  �=k  	R�  ?�   	�  @>
  	n  A>
  	�  B>
  	1$  C�	  	2�  E�  	�� F�  `	�L Ha   � �  Jw  �  P   �  �  |
  �  p  G  2
  2
  #   �  &�  �  5�  G   �%  *�  �  |
  �     �%  -�     5      {  1      |
  .   u   �  4:   @   5K   u   l  8W   ]   |
  q     �   �  <}   �   |
  �     V
   �  @�   �   |
  �   u    >
  k   �  G�   �   |
  �   G  >
  >
  �   �'  N!  	!  |
  !  G  p   �  S)!  /!  |
  R!  G  >
  >
  k  R!   o
  $&  ��6"  	�� �_   	i'  �J
  H	   �J
  P	  �J
  X	�A �}  `	Y ��  h	�#  ��  p	�  ��  x	�  �   �	  �.   �	��  ��   �	U�  ��   �	�!  ��   �	��  �!  �	�  �K   �	&  �q   � �&  �B"  X!  }\  P&T"  Z"  XpR  qB  ik"  q"  5�"  H"  G  �"  �"   a   @   A  �"  �"  5�"  H"  a    4H  ��"  �"  5�"  H"  G   �U  ��"  �"  |
  #  H"  u    >
  k   $�*   �R#  	n*  �$�"   	�5  �$_"  	XO  �$�"  	��  �$�"   �4  �"^#  #  $�>  ��#  	'O  ��   	xC  �r   s/  �d#  .�#  3  �%�#  �#  �  0t$  �  v�
   a   w�
  �'  x�
  !  y�
  �#  z�
   �  {�
  ( �  }�#  �  U'+$  1$  Xm  $D   tx$  	�  vJ
   	A  wJ
  	�  xJ
  	&  yJ
   !  {6$  �  ��$  �$  |
  �$  $  >
  �$   0  �  ��$  �$  5�$  $  �$   �'  ��$  �$  |
  %  $  >
  �	  %   x$  �!  F%  ��  )�$   ��  )�$  �  )�$   }  %  .F%  O  ;�%  _� =%�%   ݰ  >%$   S%  �  @X%  �X  L*�%  �%  cA  �,�%  �%  $/  ��%  	�� ��   	�M ��%   ?<  �,�%  �&  $�5  P��&  	�  �V
   	�� ��&  	�Y ��&  	�H ��&  	U@ ��&   	�9 �#'  (	�A  �#O'  0	�^  �#z'  8	�^  �#�'  @	N7  �#�'  H .�%  (Z  ��&  �&  |
  �&  �%  �
   17  ��&  �&  5�&  �%   �G  ��&  �&  >
  �&  �%  }   %G  ��&  '  >
  '  �%  '   }  �@  �+'  1'  >
  O'  �%  �%  }  }   �;  �['  a'  �	  z'  �%  }  }   �W  ��'  �'  '  �'  �%  �   *;  ��'  �'  '  �'  �%  �  }   �T  ��'  _  �  0  |  -1  B|  1  (  2-    1p  (  2-    #(  �  2(  G   8(  |
  V(  G  >
  �
  >
   \(  >
  p(  G  �   }�  �%�	  Z  4o
  .}(  i�3   5�(  knum  72
  kstr  8�   +P   :�(  $�J   =�(  ]key  ?�(   	�U   @G    �7   D$�(  �(  O   H)  )  V
  )  )   �(  �Z   K-)  3)  �	  G)  )  )   $�S  ( O�)  	��  Q>
   	�   R>
  	�6  S>
  	�B   U�(  	3   V!)  	>)  X�)    �(  e-   \ �)  G)  ^�(  Z   !9:*  
x,   
�V  
�K  
*  	
�Z  
`Y  
�,  
/+  
�N  
�O  
 X  
�[  
�H  
�I  
�P  
�U  
�F  
r9   $�M  !Vo*  	�\ !X�	   	�  !Y�	  	x  !Z&
   �7  !\:*  .o*  �Y  "��*  �*  |
  �*  �  a    �J  "��*  �*  5�*  �  a   a    R�F  Z   #�*  
�D   
;?  
�O   
S  
�9   
W  #�*  �]  $*.+  m+  $J>  X$Xm+  	�P  $Z5   	2�  $\�	  @	�� $]�	  H	�D  $^�+  P	� $_|
  T ~+  ^\4  Z   $F�+  
�C   
 ]  
�]   RU  $Lr+  $bR  %,�+  	�[  %.
   	x  %/J
   �K  %1�+  OS  %6�+  �+  |
  ,  [  p  �   ,  ,   �   J
  ^+/  S   %<m,  l?V  ~lBN  
�G   
GR  
�.  
�S  
�2  
�B  
9,  
>@  
R   �>  %H,  $�V  %N�,  	�� %O�+   	� %Pm,   D  %Qy,  .�,  $�6  `&S�-  	�<  &Uo
   	�Q  &Vo
  	a(  &XJ
  	VA  &YJ
  	Q) &[&
   	nX  &\&
  "	�D  &^�-  (	�5  &_�-  8	M   &a
  H	}  &b
  J	V  &c
  L	/  &d
  N	7K  &f&
  P	>D  &g&
  R	�:  &i
  T	�3  &j
  V	=]  &k
  X 1J
  �-  2-    �5  &m�,  $�Q  8&��.  	�  &�o
   	�Z  &�
  	%?  &�
  
	L/  &�
  	�<  &�&
  	�Y  &�
  	�7  &�
  	�)  &�
  	�O  &�
  	�H  &�
  	vH  &�
  	^  &��.  	�>  &�
  $	�7  &�&
  &	0>  &�a   (	�+  &�a   0 1
  �.  2-    �H  &��-  �?  8&A�/  �  &Co
   �Z  &D
  %?  &E
  
L/  &F
  S.  &H&
  �W  &J
  �W  &K
  C  &L
  �O  &M
  �H  &N
  vH  &O
  ^  &Q�.  �>  &S
  $�B  &T&
  &0>  &Za   (�+  &[a   0 �]  &]�.  �B  �&|�1  ��  &~&
   �)  &
  �)  &�&
  �.  &�&
  U  &�&
  �V  &�
  
�0  &�
  �6  &�
  �C  &�
  U?  &�
  6P  &�
  �C  &�
  &L  &�
  *J  &�
  �L  &�
  HP  &�
  N*  &��1   [2  &�V
  0k2  &�V
  8.  &�V
  @{2  &�V
  HQ2  &��1  P�0  &�&
  Tp4  &�&
  VmU  &�&
  X�Z  &�
  Z ?  &�
  \:  &�
  ^�I  &�&
  `E8  &�&
  b�;  &�V
  h�;  &�V
  p�O  &�
  xDF  &�
  zfV  &�&
  |�9  &�&
  ~[9  &�&
  ��G  &�&
  �zQ  &�&
  � 1�	  �1  2-   	 1�	   2  2-    {D  &��/  �1  @&��2  �I  &�o
   6Y  &�o
  �^  &�
  S  &�
  )  &�V
  @3  &�V
   �0  &�V
  (4C  &�V
  0�C  &�V
  8 aM  &�2  �I  @&��3  �  &�o
   _7  &�V
  )  &�&
  �O  &�&
  �n &�&
  �T  &�&
  EF  &�&
  I  &�&
  �K  &��3  N:  &��3  ,L  &��3  4�E  &��	  :�Z  &��	  ;�Z  &��	  <^  &��	  = 1�	  �3  2-    1�	  �3  2-    1�	  �3  2-    eU  &��2  �9  (&7�4  ��  &9o
   a@  &:&
  b<  &;&
  
8  &<&
  .  &=&
  �H  &>&
  �Q  &?&
  X  &@&
  �.  &A&
  �;  &B&
  ))  &C&
  eH  &D&
  I_  &E&
  �B  &F&
   !3  &G&
  " �)  &I�3  R�(  Z   &e�4  
�-   
�D  
�1  
yA  
�>  
5  
�L  
}N   KK  &q�4  $�R   'FF5  ]tag 'HV
   	��  'Io
  	.� 'JJ
  	�P  'KF5   V
  DG  'M5  $f3   '��5  ]Tag '�V
   	Q  '�V
  	.*  '�V
  	�K  '�V
   gW  '��5  X5  �^   '6  k@  '&
   aE  '&
  p0  '&
  �>  '&
  H  '&
  �/  'V
  �� '6   �	  �F  '�5  9  '=6  �5  �<  '0|6  H  '2&
   �/  '3V
  �� '86   qS  ':C6  2R  ':�6  C6  A9  0'U7  ߣ  'W&
   �E  'X>
  �^  'Y>
  =Y 'Z7  <  '[>
  �=  '\7   Jy  ']p  ( #6  |6  rY  '_�6  �1  '~Q7  �.  '�&
   �L  '�&
   Z  '�^7  &7  �V  '��7  ��  '�&
   f>  '�&
  Y  '�Q7   �)  '�d7  �A  '/S8    '1�	   �  '2�	  �N  '3�	  o=  '4�	  D4  '5�	  �^  '6�	  `*  '7�	  �0  '8�	  �G  '9�	  �D  ':�	  	I:  ';S8  
 1�	  c8  2-    �@  '=�7  &
  �\  '��8  +  '�c8   Y�  '�c8  �
  '��	  (  '��	  �F  '��	  �C  '��	   <)  '��8  v8  �,  '39  �  '&
   AK  '&
  z8  'p8  V '39   99  �	  �R  '�8  	F  '.w9  �  '0&
   �P  '199   ">  '3L9  'I�9  m�K 'K?9  m`B 'Lw9   �[   'E�9  �z  'G�	   =Y 'N�9   �6  'P�9  O]  'a!�9  �9  X�(  7N  ('�\:  >) '�6   -N  '�6  V` '�6  TE  '�V
  �/  '�>
   �z  '��	  $ G  '��9  &8  '� v:  |:  _eS  p'o�>  �� 'q�   ^  'sL5  ��^  'uV
  [>  'v&
   �W  'w�5  (� 'y�-  0�=  'z�.  ��,  '|�4  ���  '~�	  ��(  '�/  �AK  '�&
  0XL  '�7  8Uos2 '� 2  hp�  '��2  �T  '�6  0#9  '�V
  8!H '��@  @�+  '��@  H@.  '�:A  P�E  '�A  X�P  '�A  `@  '�A  h$S  '�a   ps  '�a   xUmm '�a   �Uvar '�a   �Q  '�a   �<B '��7  �2Y '��3  �=  '�V
  �=  '��8  �UV  '��9  ��(  '�V
  =  '�6   /:  '�V
  (�?  '�6  0�]  '�V
  8Ucvt '��A  @�R  '��>  H5$  '��  P��  '��  `HT  '�V
  h�*  '�V
  p�J  '��	  x�+  '��	  y�  '��9  ��C  '�}  ��-  '��  �j7  '�>
  �kN  '�V
  ��F  '�V
  �#7  '�V
  ��(  '�6  �rE  '�6  �QZ  '�V
  �4  '�>
  ��@  '�V
  �:L  '�6  ��G  '�6  ��]  '�V
  ��W  '��A  ��/  '�>
  ��B  ' �A   �I  '6  s-  'V
  �*  '>
  ,  '}  ,  '}   Ubdf '	\:  (�T  'V
  P#F  'V
  X�U  'V
  `�K  'V
  h �=  '��>  �>  |
  �>  a    �Q  '�"�>  ?  _�\  x'c�@  �  'ei:   �  'fqB  )�  'gu  �V  'hk  :1  'jV
   �^ 'k>
  (Jy  'mp  0�  'n2
  8�  'p
  <�!  'q-  @R0  'r2
  `�  's2
  duN 't2
  h6  'u�	  lFpp1 'v�  pFpp2 'w�  �2�  'zLB  �Xc  '{LB  ��6  '}YB  )  '~6  �8  'V
   �L '�a   (C  '�2
  0��  '�2
  4Upp3 '��  8Upp4 '��  Hy�  '�6  X�� '�6  `U  '�  h �I  '��@  �@  |
  �@  i:  V
  p  F5    1  '�@  �@  |
  A  �>  >
  V
  >
   �M  '+%A  +A  |
  :A  �>   �<  ':GA  MA  5XA  �>   Ry*  Z   '=�A  
4   
�^  
J  
b8  
�T   lK  'HXA  
  >
  |T  @'?LB  R�  'A�   �  'B&
  n  'C
  
Z�  'D&
  �  'E
  Forg 'G�  Fcur 'H�  ��  'I�   s  'K6  ([  'Lp8  0c+  'N&
  8 R8  'P�A  RG  'T'fB  lB  X[  O  '_ ~B  �B  XLL    �  2
  �  6  $�C  h(*�B  	�� (,�'   	�Z  (.>
  8	�  (/�	  <	X;  (0�B  @	آ  (1k  ` 12
  C  2-    �D  (3C  �B  n)  )$C  *C  |
  HC    �  r  �	   �)  )$TC  ZC  |
  sC    �  a    $�;  ))�C  	�=  )+C   	z+ ),HC   .sC  �J  ))�C  �C  �Q  *(�C  �C  |
  �C  G  V
  J
  6  F5   �+  *2�C  �C  a   D  G  �4   �7  *:D  D  |
  BD  G  >
  F5  F5  F5   $�Y  *AwD  	$\  *C�C   	�5  *D�C  	�A *ED   .BD  ;=  *A�D  wD  FO  +)(  $Y  +,�D  	6 +.�D    .�D  �O  +,�D  �D  f.  ,&2(  <B  ,,V(  $�3  ,0E  	tW ,2!�D   	i�  ,3!�D   .�D  �?  ,0E  E  $&I  -:KE  	�8  -<V
   	ߣ  -=J
   `K  -?#E  'B  -CcE  iE  |
  }E  �  }E   KE  $b:  -G�E  	'�  -IWE    .�E  SQ  -G�E  �E  �N  . �E  �E  |
  �E  G  o
  2
  R!   $�I  .% F  	�2  .'�E    .�E  �8  .%F   F  $BY  /'2F  	/  /)�    .F  �*  /'CF  2F  ��S  	-�  (                                        1�,  �F  2-    .F  �V  ��F  	�0H     $(<  0jG  	  0l&
   	d  0m&
  	�Z  0n&
  	�9 0o&
  	�� 0q6  	��  0r>
   CS  0t�F  $&^  0�;G  	�� 0�6   	��  0�>
   KJ  0�G  1�(  WG  2-    .GG  EK  1WG  	 0H     H�9  ��G  �$ �)�  Յ �)�*  R�  �)�  R   �)a   %cur ��  ?�@ ��  �U  �a     7  }|
  ��@     V       ��H  �$ }&�  �  �  ��  ~&�*  '    R   &a   �  �  cur ��  K  C  � �|
  �  �  &�@            �@ ��  �  �  !�@     T|    H
0  \�H  �$ \�  D� ]�  AT  _�  ;  _�   H�Q  A(I  �$ A �  D� B �  AT  D�  ;  D�   6�@  '@�@     .       �{I  �$ ' �  UD� ( �  T;  *�  6  2   H�H  �I  �$ �  D� �  AT  �   I�]  ��  �I  !�$ ��  !�U  �a   (cur ��   )q]  �2
  ��@     O       �FJ  Bdst � �   r  l  Bsrc � �  �  �  �  � V
  �  �   )�?  ��
  `�@     2       ��J  R�  ��  <	  4	  Bstr ��  �	  �	  �4  ��J  

  
  "len �V
  k
  i
  |�@     �k �J  Us  ,��@     �J  U�UT�TR�Q  |
  )�3  ��
  ��@     x       �L  R�  ��  �
  �
   �r    �
  �  �V
  ~  t  �4  ��J  �  �  *� �|
  (p ��
  /�N  ��@      @T  ��K  �N  n  l  �N  �  �  �N      @T  J�N   �N  �  |  ��@     U�UTs    �@     �k Tv Qs   YF\  �3L  !R�  ��  AP �r   )�[  r�
  �@     �       ��M  R�  r�  �  �  Y  sJ
  �  �  �Y  tJ
  �    �2  uJ
  d  X  ��  va     �  �4  w�J  �  �  � y|
  �  �  :��@     5       FM  �)  ��
  V  T  *f;  �J
  *6^  �J
  ��@     U�UT�T�QRw   /L  x�@      @B  ��M  (L  }  y  L  �  �  ��@     U�UT�X  b�@     U�UT�R�T  )�6  \�
  ��@     o       ��N  R�  \�  �  �  Y  ]J
  :  0  �Y  ^J
  �  �  �2  _J
       ��  `a   �  �  �4  a�J  .  &  E� c|
  �L
�@     3L  �N  U�UTv Q} Rs X�XY�L I�@     �k U~ v "T0Qs �T  IkA  B�
  O  !R�  B�  !�  CJ
  !�4  D�J  *� F|
  *��  G�
   )�K  2�
  ��@     g       �P  R�  2�  �  �  �  3J
    �  �4  4�J  �  �  *� 6|
  *��  7�
  /�N  ��@      P>  7�O  �N      �N  :  .  �N  �  �  P>  J�N   �N  3  )  ��@     U�UTs    Ɍ@     �k T0Qs   s3  �}(  p�@     /       �_P  1  �}(  U 1  �}(  T� }(  �  �   6M<  �@�@     !       ��P  ;vec �%�  �  �  ss  �%o
  #    P�  �%}(  �  �  ,X�@     �R  U�UT�Q  6�3  �p�@     �       ��Q  ;vec �#�  �  �  ss  �#R!  I  ?  P�  �#�Q  �  �  �� �2
  =  7  Mv ��  �PUX  ɋ@        >  ��Q  fX  �  �   >  rX  i  c    ��@     �D �Q  Uu Tt 0(X  u  ŋ@     D Uu 0RW  u   }(  �K  �o
  `�@     �       ��R  ;vec �!�  �  �  �� �2
  =  5  Mv ��  �`UX  ��@       �=  �wR  fX  �  �  �=  rX    y    ��@     �D �R  Uu Tt 0(X  u  ��@     D Uu 0RW  u   6�8  � �@     9      �T  ;vec �!�  �  �  P�  �!}(  h   `   �� �2
  �   �   Mv ��  �P:��@     0       QS  �� �k  -!  +!   UX  u�@       p=  ��S  fX  d!  T!  p=  rX  7"  1"    UX  ��@      �=  ��S  fX  �"  �"  �=  rX  g#  a#    d�@     �D �S  Uu Tt 0(X  u  q�@     �C Uu Q�T0�W  u   H�0  i<T  `vec i�  P�  j}(   �5  T}(  ��@     ?       ��T  ;dx To
  �#  �#  ;dy Uo
  $  $  Mv W�  �`�@     �D �T  Uu Tt 0(X  u  ��@     D Uu 0RW  u   �L  Fo
  P�@     h       �V  P�  F}(  `$  Z$  Mv H�  �`T  W�@       W�@            K{U  .T  �$  �$  !T   %  �$  _�@     M Uw T�U  8> h�@       h�@     K       M0> )%  #%   %> &h�@     K       ;> }%  s%  F> �%  �%  Q> &  &  \> &  {&  g> �&  �&     �L  8o
  0�@            ��V  P�  8}(  �&  �&  Mv :�  �`8T  7�@       7�@            =.T  5'  /'  !T  �'  �'  ?�@     M Uw T�U   �6  *o
  �@            �EW  P�  *}(  �'  �'  Mv ,�  �`8T  �@       �@            /.T  �'  �'  !T  L(  J(  �@     M Uw T�U   a�Y  ��W  Avec �(�  *�5  �}(  (i �2
  (x �o
  (y �o
  *�?  �o
  (b �#o
  *�A  ��W   �(  az[  �X  Avec �&�  !�5  �&}(  (i �2
  (x �o
  (y �o
  *�?  �o
  (b �#o
  *�A  ��W   Z�M  �2
  UX  Avec � �  (x ��  (y ��  *�� �2
   ZR\  =o
  }X  Aval = o
  (s ?2
   d�N  �|
  0�@     �      �0Z  Jy  �0p  {(  o(  �S �00Z  )   )  �/  �0a   �)  �)  � �|
  3*  #*  y:  ��	  �*  �*  y�  �6  �+  �+  -�u  S��@     '�<  �Y  �\ �V
  �-  s-  o[  �2
  P.  @.  p �6  	/  �.  ' =  �Y  len �>
  �/  �/   $�@     �`  Uv   8~`  ��@      ��@     :       V�`  70  50  <�] ��@     #       �`  \0  Z0  7L  ��@       @=  O(L  �0  �0  L  �0  �0      {*  �P  �V
  ��@     |       ��Z  Jy  �%p  �0  �0  � �%�J  >1  21  �R  ��Z  �\p �6  �1  �1  E  �V
  d2  ^2  -�0  ��@     �@     Us Q�\R4  1�	  �Z  2-    �F  pV
  P�@     |       ��[  Jy  p#p  �2  �2  � q#�J  "3  3  �R  s�Z  �\p t6  �3  �3  E  uV
  H4  B4  -�0  ���@     ��@     Us Q�\R4  *  CV
  ��@     �       �\\  Jy  C%p  �4  �4  � D%�J  5  �4  �R  F\\  �]p G6  �5  �5  E  HV
  ,6  &6  -�0  e0�@     ��@     Us Q�]R3  1�	  l\  2-    -4  &
  0�@     �       �]  Jy  &p  6  w6  � &�J  �6  �6  �R  ]  �^p 6  ~7  r7  E  &
  8  
8  -�0  8��@     e�@     Us Q�^R2  1�	  .]  2-    >Q  �&
  p}@     �       ��]  Jy  �$p  c8  [8  � �$�J  �8  �8  �R  �]  �^p �6  b9  V9  E  �&
  �9  �9  -�0  �}@     �}@     Us Q�^R2  ?U  ��	  �|@            �o^  Jy  �"p  K:  ?:  � �"�J  �:  �:  E  ��	  i;  g;  -�0  �&}@      }@     Us Q�_R1  \  �V
  �|@            ��^  Jy  �$p  Up �6  �;  �;  E  �V
  �;  �;   RH  �V
  �|@            �%_  Jy  �"p  Up �6  <  <  E  �V
  m<  i<   �5  �V
  �|@     .       ��_  Jy  �$p  Up �6  �<  �<  E  �V
  �<  �<   �N  {&
  P|@     (       ��_  Jy  {%p  Up }6  6=  0=  E  ~&
  �=  �=   ?  h&
   |@     '       �6`  Jy  h#p  Up j6  �=  �=  E  k&
  >  >   iD  X�	   |@            �~`  Jy  X!p  UE  Z�	  J>  H>   HxL  :�`  Jy  :#p  ?R�  I�    )�3  �|
  @z@     1      �6b  Jy  �$p  |>  n>  .� �$V
  +?  ?  � �|
  @  @  �I  �V
  �@  �@  -�u  4.{@     9  R�  ��  �@  �@  �N  kz@      �9  �a  �N  %A  A  �N  �A  }A   �N  �9  �N  �A  �A  �N  TB  JB  �z@     U| Tv    L  �z@      �z@            	 b  (L  �B  �B   L  �z@     U|   9�z@     b  Us Rv  �z@     Us Q0R0   ��J  �z@     +       ��b  Jy  �&p  �B  �B  qI  �&�B  .C  (C  & z@            R�  ��  ~C  zC  #L  #z@       �8  �(L  �C  �C  L  �C  �C     )�*  �|
  �{@     4       �cc  Jy  �&p  D  D  .� �&V
  kD  gD  qI  �&�B  �D  �D  � �|
  �D  �D  �{@     �`  Us T�T  )�R  �V
  �y@     h       �#d  Jy  �!p  #E  E  B� �!6  �E  �E  .� �!V
  "F  F  �I  �V
  �F  �F  e�u  ��y@     9�y@     d  Us Q�TR�Q z@     �k U�TQv   )`I  w|
  y@     }       � e  Jy  w p  {G  qG  Bpos x V
  �G  �G  B� y 6  \H  TH  .� z V
  �H  �H  � ||
  @I  :I  �I  }V
  �I  �I  9;y@     �d  Uv Ts Q�QR}  �y@     �k U�QQ|   IE1  n|
  6e  !Jy  np  !B� o6  !.� pV
   IF  gV
  Te  !Jy  gp   I _  \|
  ~e  !Jy  \p  !3{  ]J
   I9  9|
  �e  !Jy  9p  Apos :V
  *� <|
   Y�U  1�e  !Jy  1p   Y�X  # f  !Jy  #)p  !2�  $)�	  !�  %)V
   )fQ  `|
  ��@     c      �h  �  `)G  �I  �I  �.  a)>
  5J  1J  �C  b)h  vJ  nJ  *� d|
  �R  e5  ii:  �J  �J   S  � r�6  CK  ?K  PS  R�  y�  {K  yK  Jy  zp  �K  �K  /~e  ��@       �S  ~1g  �e  �K  �K  �e  L  L  �S  �e  gL  aL  ��@     U} T Q0R0   / e  ��@       �S  �g  )e  �L  �L  e  �L  �L  e  	M  M  ��@     #d  U} T   NL  �@      �@            ��g  (L  AM  ?M  L  gM  eM  �@     U|   ��@     �M  U| T1Q0X0Y��     ;G  )I  -|
  p�@     q      �&j  �  -#G  �M  �M  Bidx .#>
  �M  �M  �D  /#&j  9N  1N  � 1|
  �N  �N  �Q  e5  6i:  �N  �N   R  � ;06  ,O  (O  0R  R�  A�  dO  bO  Jy  Bp  �O  �O  /~e  L�@       `R  FKi  �e  �O  �O  �e  P  �O  `R  �e  PP  JP  ^�@     U} T Q0R0   / e  ��@       �R  G�i  )e  �P  �P  e  �P  �P  e  �P  �P  ��@     #d  U} T   NL  ��@      ��@            I�i  (L  #Q  !Q  L  IQ  GQ  ��@     U|   8�@     �M  U| T1Q0X0Y��     G  )�/  $>
  �w@            �]j  S�  $$G  U C�Q  f�   P�@     �       ��k  R�  f(�  vQ  lQ  /  g(�  �Q  �Q  �O  h(�  �R  R  xI  j�   
S  �R  tmp k�  �S  �S  O  l�  �S  �S  �T  mG   T  T  � n|
  �Lu�@     �k ;k  Uv  ��@     �k Sk  U|  ��@     O  qk  Us Q�L ��@     �k �k  Uv T/ ˍ@     �k �k  Us T�TQ~ ܍@     �k �k  Us T|  �@     �k Us Tv   C�A  L|
  ��@     �       �On  k  L:[  DT  @T  R  M:�   �T  }T  �)  N:,  �T  �T  m-  P)  ���7  Qp  ���,  R�   RU  PU  � S|
  �U  vU  Jx  �@       �>  \:m  �x  �U  �U  �x  ]V  YV  vx  �V  �V  ix  �V  �V  \x  W  W  �>  �x  [W  WW  �@     $^ T Qv 0an  �U0{n  �T   � �@      �@     "       _+n  � �W  �W  � �W  �W  <DS �@            � �W  �W  /�e  �@       ?  ��m  �e  X  X  "�@     Uv   8L  "�@      "�@            	(L  2X  0X  L  WX  UX  -�@     U| Tv     �@     
 U�UT��Q��  =1-  
|
  o  k  
,[  Jy  ,p   L  ,�   �  ,k  �)  ,,  :  k  � |
  R(  k  �[  &
  %i S   =O  k  �F  k  �0  (k  /O  x   C}E  �|
  P�@     �       ��p  k  �-[  �X  zX  Jy  �-p  *Y  &Y   L  �-�   iY  cY  �+  �-,  �Y  �Y  �)  �-,  oZ  aZ  yM  ��   [  [  � �|
  �[  �[  R�  ��  
\  \  L  ��@      ��@            9p  (L  U\  S\  L  z\  x\  ��@     U| Ts   x�@     ]j  ep  U| T�QQ	 /H      ��@     �k  Uv Ts Q~   C�/  �|
  �@     �       ��q  k  �+[  �\  �\  Jy  �+p  M]  I]   L  �+�   �]  �]  �+  �+,  �]  �]  �)  �+,  �^  �^  yM  ��   >_  0_  � �|
  �_  �_  R�  ��  -`  '`  L  6�@      6�@            ��q  (L  x`  v`  L  �`  �`  A�@     U| Ts   �@     ]j  �q  U| T�QQ	/H      .�@     �k  Uv Ts Q~   C2  �|
   �@     D       ��r  k  �([  �`  �`  Jy  �(p  a  �`   L  �(�   @a  :a  �+  �(,  �a  �a  �)  �(,  b  b  yM  ��   �b  �b  R�  ��  �b  �b  <�@     ]j  T�QQ	�.H       C�F  �|
  p�@     D       ��s  k  �#[  c  c  Jy  �#p  Xc  Tc   L  �#�   �c  �c  �+  �#,  �c  �c  �)  �#,  ld  bd  yM  ��   �d  �d  R�  ��  Je  He  ��@     ]j  T�QQ	�.H       CaZ  r|
  P�@     �       ��t  k  r,[  ve  ne  Jy  s,p  �e  �e   L  t,�   f  f  �+  u,,  �f  yf  �)  v,,  �f  �f  � {|
  ��yM  |�   Mg  Gg  R�  }�  �g  �g  tO  ~J
  �g  �g  w�@     �k �t  U|  ��@     O  �t  TsQ�� ��@     �k T| Qs   C�E  N|
  ��@     �       �v  k  N-[  h  h  Jy  O-p  wh  sh   L  P-�   �h  �h  �+  Q-,  i  i  �)  R-,  �i  ~i  � W|
  ��yM  X�   �i  �i  R�  Y�  7j  5j  tO  ZJ
  aj  [j  �@     �k �u  U|  �@     O  �u  TsQ�� .�@     �k T| Qs   C)E  0|
  ��@     �       �tw  k  00[  �j  �j  Jy  10p  Zk  Vk   L  20�   �k  �k  �+  30,  �k  �k  �)  40,  �l  �l  yM  6�   Km  =m  � 7|
  �m  �m  R�  8�  :n  4n  L  ֓@      ֓@            G'w  (L  �n  �n  L  �n  �n  �@     U| Ts   ��@     ]j  Sw  U| T�QQ	/H      Γ@     �k  Uv Ts Q~   C=6  |
  P�@     &       �Jx  k  +[  �n  �n  Jy  +p  o  
o   L  +�   wo  qo  �+  +,  �o  �o  �)  +,  p  p  ��   k    ,l�@     $^ U�TT  Q�X0an  �U0{n  �Q  =�?  |
  �x  k  +[  Jy  +p   L  +�   �+  +,  �)  +,  �  
k   =�8  ��	  �x  k  �.[  1  �.>
   =d1  �m,  y  k  �6[  1  �6>
   6l5  �w@     �       �Mz  k  �![  mp  gp  Jy  �!p  �p  �p  �X  �!�   q  q  oM  �!,  Kq  Gq  �P  �!,  �q  �q  +  �!�J  �q  �q  i �2
  2r  (r  ~e  @w@      `8  �z  �e  �r  �r  �e  �r  �r  `8  �e   s  s  Tw@     U~ T0Q0R0   �w@     U T~ Q��RvxXs 3$} "  )ND  �|
  Щ@     x      ��  k  �+[  `s  Xs  Jy  �+p  �s  �s  ��  �+J
  7t  )t  y^  �+J
  �t  �t  Btag �+J
  Mu  =u  �[  �+�	  v  �u  S�P  �+�  � S.� �+,  �E� �|
  ��"i �S   pv  hv  "j �S   �v  �v  "cnt �S   �w  �w  YI  �S   x  x  7F  �J
  �x  xx  �;  �!J
  �x  �x  R�  ��  oy  ey  /� �J
  �y  �y  W  �,  Rz  Hz  "ref ��  �z  �z  -�u  Bx�@     /~e  ��@      �E  �R|  �e  �{  �{  �e  �{  �{  �E  �e  #|  |  �@     Us T Q0R0   ~e  '�@       F   �|  �e  _|  [|  �e  �|  �|   F  �e  �|  �|  @�@     Us T Q0R0   Te  Q�@      @F  U}  qe  }  }  ee  K}  G}  #~e  Y�@       pF  b�e  �}  �}  �e  �}  �}  pF  �e  '~  ~  ��@     Us T~ Q0R0    Te  ݫ@      �F  �}  qe  �~  �~  ee  �~  �~  #~e  �@       �F  b�e    �~  �e  R  L  �F  �e  �  �  ��@     Us T~ Q0R0    L  x�@      x�@            C	I~  (L  �  �  L  �  �  ��@     U��T}   4�@     .]  h~  Us T�� m�@     .]  �~  Us T�� ��@     .]  �~  Us T�� ��@     �Z  �~  Us T�� r�@     �M  �~  U��T@Q0X0Y�� Ϋ@     �Z    Us T�� E�@     .]  3  Us T�� ׬@     �M  c  U��T8Q0X0Y�� C�@     �k U} Q@R	0@       ,  �+  Vq(  �S   0@            ��  Oa �-�  UOb �-�  T )WB  3|
   ~@     $      �Ѓ  k  3*[  A�  9�  Jy  4*p  ��  ��  t6  5*J
  r�  d�  ��  6*,  "�  �  y^  7*,  ��  �  � 9|
  ��  ��  E�; :Ѓ  ��E�2  :Ѓ  �@�K  ;J
  �  �  )-  ;J
  _�  [�  )  ;&J
  ��  ��  R9  <S   ф  τ  [^  <S   ��  �  "i <(S   2�  .�  }Z  =J
  l�  j�  /~e   ~@      @:  B|�  �e  ��  ��  �e  �  �  @:  �e  9�  5�  1~@     Us T| Q0R0   / e  V~@      �:  F�  )e  s�  q�  e  ��  ��  e  ؆  Ԇ  [~@     #d  Us T| Q��R@  /~e  �@      �:  �L�  �e  �  �  �e  L�  H�  �:  �e  ��  ��  �@     Us T| Q0R0   / e  �@       ;  ���  )e  ��  ��  e  �  �  e  $�   �  �@     #d  Us T| Q�@R@  /Te  #�@      0;  �L�  qe  ^�  Z�  ee  ��  ��  #~e  +�@       `;  b�e  Ԉ  Ј  �e  �  
�  `;  �e  H�  D�  D�@     Us Tv Q0R0    /~e  x�@       �;  ���  �e  ��  ��  �e  ��  ��  �;  �e  ��  �  ��@     Us T| Q0R0   d�@     .]  Us T��  1�  ��  2-    )Q=  �|
  Pv@     �       ��  ~ �!  4�  0�  n  �!�  l�  j�  S�\ �!a   Qn� �|
   K1 �C  ��  ��  :�v@     @       ��  X;  ��B  ˊ  Ɋ  "val ��B  �  �   :�v@            ׄ  �Z  >
  �  �  val �A  =�  ;�   &�v@            �  �	  b�  `�  val �  ��  ��    �	  )v@  '|
  �s@     �      �&�  ~ '!  ��  ��  n  (!�  @�  >�  �\ )!r  q�  c�  �R  *!�	  �  �  n� ,|
   K1 -C  U�  I�  :�s@     !      ��  X;  6�B  �  ݍ  "x1 72
  0�  .�  "y1 72
  W�  S�  "x2 72
  ��  ��  "y2 72
  ��  ��  "x3 7 2
  �  �  "y3 7$2
  -�  )�  "x4 7(2
  h�  d�  "y4 7,2
  ��  ��  [dp :�B  ��&�s@     m       "s ?�  Ǐ  ŏ  [ep @�   ��(i AS   �s@     �k ݆  U~ T��Q: t@     �k U~ T��Q:   :u@     &       '�  "s ~�  �  �   '08  E�  �Z  ��A  +�  '�   :v@             ��  "s ��  c�  a�  "nsd �@   ��  ��  v@     �k U~ T0Q:  :�u@            ɇ  �  ��  ��  ��    8  آ  �k  ֐  А  &0v@            "s ��  3�  1�  ?v@     �k U~ T0Q:    WuJ  	�*  ӈ  �S  	,�B  C!  	-  �.  	2
  �-  	2
  �  	�  �0  	�  �I  	�  %c 	2
  %n 	2
  N� 	2
  OD 	�  ?k� 	82
    ;  	�|
  0o@     *      �;�  �S  	�'�B  b�  V�  �\  	�'�  �  �  h9  	�'�  [�  O�  �  	��  �  �  c 	�2
  !�  �  N� 	�2
  {�  o�  k� 	�2
  
�  �  V  	�2
  l�  f�  '02  ��  in 	��  ��  ��  Mout 	��  ��YK  	��  �  �  �� 	�#�  ڕ    �� 	�o
  �  �  �� 	�o
  ��  ��  WK  	�o
  �  �  l 	�-o
  )�  %�  q 	�0o
  g�  _�  d 	�3o
  "�  �  i 	�2
  ڙ  ҙ  j 	�2
  :�  8�  k 	�2
  c�  ]�  t> �p@      �2  	��  �> ��  ��   �> #FC �p@       3  �aC ۚ  ٚ   WC  3  kC �  ��  wC E�  C�     t> q@      �3  	�*��  �> o�  m�   �> #FC q@      4  �aC ��  ��   WC 4  kC ��  ��  wC  �  ��     t> �q@      p4  	��  �> =�  ;�  �> d�  b�  #FC �q@      �4  �aC ��  ��  WC ��  ��  p5  kC ٜ  ՜  wC �  �     t> �q@      �5  	�/��  �> Y�  W�  �> ~�  |�  #FC �q@      p6  �aC ��  ��  WC ȝ  Ɲ  �6  kC wC    t> -r@      p7  	��  �> �  �  �> �  �  #FC -r@      �7  �aC ;�  9�  WC b�  `�  �7  kC ��  ��  wC Ξ  ʞ     vp@     J2 0�  Uu  (r@     e? R�  T��Q�� tr@     e? |�  U��T��Q�� "s@     e? ��  U��T} Q��~ Js@     e? T} Q��~  7&�  }o@       2  	�8�  �  	�   2  E�  R�  _�  l�  y�  ��  ��  ��  ��  ��  \�  X�  �o@     �K Us     �L  	�|
  `s@            ���  �S  	�%�B  ��  ��  �\  	�%�  ՟  џ  ,hs@     ӈ  U�UT�TQ�T  H�-  	��  �S  	�,�  :  	�,�  %vec 	��  �� 	��   �  H�:  	�6�  ��  	�*�  :  	�*�  %xz 	��  %yz 	��   �Y  	�|
  �n@     F       ���  k  	�,[  �  �  �S  	�,�B  f�  `�  �O  	�,l  ��  ��  G  	�y  ���n@     ��  Qw   �]  	f|
  �m@     �       ��  k  	f)[  "�  �  �S  	g)�B  ��  ��  G  	h)�  �  �  � 	j|
  Z�  P�  9X  	k�  Ң  ̢  D� 	l�  $�  �  D�  /n@      /n@     8       	���  p�  ��  ��  c�  ��  ��  V�  ֣  ԣ  &/n@     8       }�  ��  ��  ��  5�  3�  \��  D�V �1  ��  _�  Y�     9'n@     
�  T|  un@     T|   y  6�?  	) m@     �       �1�  �S  	)$�B  Un 	+&
  ��  ��  N� 	,2
  ��  ��  k� 	,2
  K�  I�  '�1  ё  p 	:�  t�  n�  q 	;�  ť  ��  �8  	<�  �  �   &�m@     -       p 	K�   Y�  S�  q 	L�   ��  ��  &�m@            �8  	Q�   ��  ��     HcL  	�  �S  	,�  Y@  	,�  �K  	,�  %n 	&
  %vec 	�   H�,  	��  �S  	�+�  �9  	�+#  M   	��  }  	��  V  	��  /  	��  ?%vec 	��  �� 	��  ?%x 	��  %y 	��     _[  	�|
  �l@            �s�  k  	�![   �  �  �S  	�!�B  r�  l�  ,�l@     s�  T�T  M3  	�|
   l@     �       ���  R�  	�*�  Ƨ  ��  �S  	�*�B  -�  %�  L  (l@       (l@            	��  (L  ��  ��  L  ��  ��  0l@     Uv   L  <l@      <l@            	�d�  (L  �  �  L  �  �  Gl@     Uv   8L  Sl@      Sl@            	�(L  7�  5�  L  \�  Z�  ^l@     Uv    _  	�|
  Pk@     �       �=�  �% 	�'�  ��  �  �  	�'�B  	�  ��  }5  	�2
  ��  ��  K�k@     �k K�k@     �k K�k@     �k  �^  	e|
  �`@     f       ���  �S  	e"�B  �  �  �Bad 	��`@     �,  Z�  	i2
  "�  �  �  	j2
  j�  h�  �P  	k2
  ��  ��  end 	k2
  �  �  n 	l2
  7�  3�    E  	U|
  P�@            ���  k  	U [  u�  o�  �1  	V >
  Ǭ  ��  xW  	W 2
  �  �  �.  	X �B  k�  e�  ,]�@     ��  T�TQ�QR�R  W+  	+|
  �  R�  	+)�  �1  	,)>
  xW  	-)2
  �.  	.)�B  � 	0|
  >�0  	J )N  	3|
  �[@     �      ��  �S  	32�B  ˭  ��  �R  	42�  ��  ��  R   	52a   ��  ��  /_  	;�  ��  ��  E�C  	<�  ��~Ey>  	=�  ��oI 	?�  ��  ��  �� 	@�  a�  U�  s  	A�   �  �  � 	C|
  J�  8�  "n 	E2
  �  �  N� 	F>
  յ  ϵ  "tag 	G2
  /�  �  �� 	I2
  -�  %�  � 	J�  ��  ��  >��  	%>�u  	!e�S  	�	S^@     -�U  	�_@     p+  k� 	Y2
  w�  k�  :]@     ?       ��  [vec 	��  ��L]@     U��T��~  ' ,  )�  [vec 	��  ��Ep>  	��  ��9@^@     �  U T��Q��~ �^@     U��~T��Q��~  '@,  ��  E�(  	��  ��E�(  	��  ��'�,  ��  [vec 	��  ���_@     U��T��Q��R��~  �`@     U��T��Q��R��~  9�\@     ؙ  U��T��~ 9�^@     ��  U��T��~ �_@     U~ T��Q��~   �  �P  �|
  @[@     �       ��  )�  �'u  U�N  �'>
  T�)  �'�B  Q�W   '�A  R{0  '�B  Xg/  '�B  YWN  '�  � � |
  ;�  5�  &p[@     P       �.  �  ��  ��    �
  "D  ��  �Z@     C       �  k  �,[  ��  ��  E  ��  �  ��  @+  ~ �  Q�  O�  :[@            ��  YM  �$7F  v�  t�  [@     ��  T	�.H     Q0  [@     ��  U�UT	�.H        6�B  ��Z@     +       ��  k  �)[  U�8  �)>
  TU*  �)p  Q F'  d|
  pY@     L      ���  k  d [  ��  ��  R�  f�  .�  (�  >�u  �' +  �  m �>
  }�  {�  n �>
  ��  ��  �,  ���  ��&�Y@     G       ~ �  $�   �     ��  \�  Z�  �   ��  Z@     l �  T}  K)Z@     k�    L  yZ@      yZ@            �n�  (L  ��  ��  L  ��  ��  �Z@     U��T|   pZ@     ��  U|   1�  ��  2-    6�E  E0Y@     :       �.�  k  E$[  U�[  F$�B  T2  G$�B  Q�K  H$�B  R0  J2
  Ҽ  ̼  �  K2
  #�  �  �  L2
  t�  n�   +  |
  ��@     f       �  R�   �  ǽ  ��  j     .�  &�  k  [  ��  ��  � |
  �\�@     O  Us T
`Q�\  [  *W  |
  Y@            ���  k  %[  U K  �|
  �X@            ���  k  �-[  ��  �     �-Y  4�  0�  n  �-Y  q�  m�  �\ �-�  ��  ��  ,Y@     ��  U�UT�TQ�QR�RX1Y1  B(  �|
  �X@            �S�  k  �&[  �  �     �&Y  (�  $�  n  �&Y  e�  a�  �\ �&a   ��  ��  ,�X@     ��  U�UT�TQ�QR�RX0Y0  T1  �|
  �X@            ���  k  �&[  ��  ��     �&Y  �  �  n  �&Y  Y�  U�  �\ �&r  ��  ��  ,�X@     ��  U�UT�TQ�QR�RX1Y0  =�Q  g|
  ��  k  g%[     h%Y  n  i%Y  �\ j%a   `set k%�	  �R  l%�	  %cur n��  �� o��  P�  p`  YM  r�C  =>  z�	     d�:  ?|
   W@     �      ���  k  ?![  ��  ��  ~ @!  E�  9�  �(  cur I��  ��  ��  �� J��  >�  0�  7C�  �W@      @)  \Q�  ��  ��  @)  ^�  @�  :�  k�  ��  ��  x�  ��  ��  L  �W@      �W@     
       mˢ  (L  )�  '�  L  N�  L�  �W@     U} Ts   � �W@      �W@             f~�   s�  q�  7rG  �W@       �)  ��G  ��  ��  �G  ��  ��  �G  ��  ��  �G  �  �  �)  �G  �W@     `O Us T	 ;@     Rs     � �  �)  b��  �  e�  a�  �)  �  ��  ��  (�  ��  ��  5�  �  �  �I   X@       X@            )*�  �I  y�  w�  �I  ��  ��  & X@            �I  ��  ��    DB�  �)  C�  ��  ��  �H  0X@      @*  5��   I  %�  #�  �H  J�  H�  @*  I  I  @X@     O Uu Tv    L  @X@      @X@            6�   (L   L  GX@     U   7԰  GX@      p*  8�  t�  p�  p*  �  7D�  GX@      �*  �p�  ��  ��  c�  ��  ��  V�  .�  *�  �*  }�  h�  d�  ��  ��  ��  G��  vX@     D�V �*  ��  ��  ��          �W@     Us      WKM  �
  �  ~ '  �1  '�  t� '�	  E  �
  ?k  "[  %cur #��  �� $��    !,  r  0V@     '       ���  k  )[  �  �  T  )�  U�  Q�  ~   ��  ��  9V@     ��  U�UT�T  �R  �  �U@     p       �5�  k  �[  ��  ��     ��  �  �  PE  �   cur ���  Y�  W�  �� ���  ~�  |�  V@     l T|   d�  t|
  К@     �      �=�  k  t*[  ��  ��  �M u*=�  U�  G�  � w|
  ��R�  x�  ��  ��  ~ y  T�  >�  nn z>
  =�  9�  -�u  �x�@     -�0  �<�@     :ԛ@            �  K1 �i  w�  u�   :A�@     "       I�  9X  ��  ��  ��   R�  6�@      �@  ��  d�  ��  ��  �@  q�  �  �  ~�  c�  ]�  4��  ����  ��  ��  G��  �@     G��  �@     o��  �@  �  ��  i�  e�  Ű  ��  ��  {I  ��@      0A  B�  �I  ��  ��  �I  �  �  0A  �I  ɜ@     �N Uu T    ԰  ɜ@      `A  ��  �  X�  T�  `A  �  7D�  ɜ@      �A  �p�  ��  ��  c�  ��  ��  V�  �  �  �A  }�  L�  H�  ��  ��  ��  G��  ��@     D�V �A  ��  ��  ��       ��@     U| Ts�   L  �@       B  ]�  (L   �  ��  L  b�  \�  ��@     U| T   L�@     O  U| THQ��   L  c�@      c�@     
       �ת  (L  ��  ��  L  ��  ��  m�@     U} Ts   K�@     l �  T|  q�@     ��  �  Uv T  ��@     O  ,�  U} Q�� �@     Us   k  T�>  V��  ~ V  R�  X�  �M Y�'  k  Z[   �O  *|
  �U@     6       ��   *$u  ��  ��  Q,  +$-  y�  q�  k  -[  ��  ��  ,�U@     �  T�UQ�T  X]  �|
  �T@     �       �ޭ  k  �-[  �  �   �-u  ��  ��  Q,  �--  ��  ~�  � �|
  J�  <�  9X  ��  ��  ��  �'  D� ��  k�  _�  D�  �T@      0(  �*�  p�  ��  ��  c�  �  �  V�  @�  >�  0(  }�  e�  c�  ��  ��  ��  \��  D�V `(  ��  ��  ��     D�  U@       U@     5       ���  p�  ��  ��  c�  �  �  V�  9�  7�  &U@     5       }�  ^�  \�  ��  ��  ��  \��  D�V �(  ��  ��  ��     �T@     Tv Q| R0   �@  L|
  ��@           ��  k  L#[  �  ��  9X  M#�  ��  s�  G  N#>
  S�  I�  IE  O##  ��  ��  D� Q�  *�  &�  � R|
  n�  `�  l� T�  �  �  -�u  ��@     �I  $�@       �T  i�  �I  Y�  W�  �I  ~�  |�  �T  �I  ��  ��    D�@     �H  �  Tt  ��@     Uv   �A  @�  @T@     6       � �  k  @%[  Uߣ  A%�  T8D�  @T@      @T@     4       Ep�  ��  ��  c�  �  �  V�  @�  <�  &@T@     4       }�  z�  v�  ��  ��  ��  G��  tT@     <�V QT@            ��  ��  ��      T�S  R�  ~ "  k  [  R�  �  D�  �  ?�� ,�    =2X  �|
  ԰  ~ �  k  �[  R�  ��  � �|
  D� ��  >�u  >�0  ?�� ��  �M ��'    T9Z  ���  k  �([  9X  ��   =�M  ��  D�   �+u  �  �G  k  �[  E  ��   W6_  ��  ��  k  �([  ߣ  �(�  D� �(��  %cur ��  E  ��  -�u  �)T@     ?9X  ��    �  BX  �|
  �S@     6       ��  �  �  U�  �G  Y�  Q�   �9  nJ
  �P@     ^       ��  �� n#�  ��  ��  YM  p�E  5�  3�  �  qG  \�  X�  +�  rKE  �`:�P@            ϲ  ~ y  ��  ��  �O  y�
  ��  ��  �P@     T	v.H       �P@     Us Tw   !@  VV
  P@     c       ���  �� V(�  ��  ��  YM  X�E  ��  ��  �  YG  ��  ��  +�  ZKE  �`'P%  ��  ~ a  ��  ��  �O  a�
  �  �  BP@     T	v.H       OP@     Us Tw   �U  =|
  �O@     �       �ʴ  �  ="G  S�  G�  �P  >">
  ��  ��  ;tag ?"F5  {�  o�  ss  @"F5  �  �  YM  B|D  ��  ��  x  CV
  �H' %  ��  ~ K  ��  ��  �O  K�
  �  �  �O@     T	k.H       �O@     Us Tv Q| R�HX}   |;  &|
  �N@     �       ��  �  &"G  ��  q�  ;tag '"V
  ?�  /�  x  ("J
  ��  ��  B� )"6  ��  ��  ss  *"F5  y�  i�  YM  ,|D  +�  '�  '�$  ��  ~ 2  e�  a�  �O  2�
  ��  ��  /O@     T	k.H       @PO@     U�UT�TQ�QR�RX�X  �+  a   �N@     c       ���  �  #G  �  �  ;tag #�4  ��  ��  P>) a    YM  |D  W�  S�  'p$  ��  ~   ��  ��  �O  �
  ��  ��  �N@     T	k.H       @�N@     U�UT�T  �/  ��  �M@     �       ���  �  �$G  �  �  PE  ��   -�u  	cN@     �#  YM  ��D  ��  ��  '�#  ��  svc �
  /�  %�  @$  ~   ��  ��  �O  �
  ��  ��  GN@     T	V.H        @N@     U�U   �H  �|
  �L@     �       �ȸ  �  �"G  O�  ?�  �^ �">
  �  ��  B� �"�
  ��  ��  (5  �">
  q�  e�  � �|
  PYM  �E   �  ��  '#  ��  svc ��
  R�  J�  &�M@     "       ~ �  ��  ��  �O  ��
  ��  ��  �M@     T	K.H        @IM@     U�UT�T  �>  �>
  0L@     �       ���  �  �"G  J�  :�  la �"�  
�  ��  PE  �>
   �!  YM  �E  ��  ��  'p"  ��  svc ��
  #�  �  �"  ~ �  ��  ��  �O  ��
  ��  ��  �L@     T	K.H        @yL@     U�UT�T   �V  �'  0S@     S       ���  �  �(G  �  �  X6  �(V
  ��  ��  PE  �'   0'  �� ��  7�  3�  '�'  w�  �1  ��%  o�  m�  R�  ��  ��  ��  @nS@     Q�T  MS@     .V 0a s    �\  n'  �R@     S       �a�  �  n(G  ��  ��  �j o(V
  n�  b�  PE  q'   �&  �� v�  ��  ��  '�&  I�  �1  {�%  2�  0�  R�  |�  Y�  U�  @S@     Q�T  �R@     .V 0a s    p$.  S'  �R@     ;       ��  �  S)G  ��  ��  PE  U'   @&  �� Z�  )�  %�  'p&  ��  �1  _�%  a�  _�  R�  `�  ��  ��   �R@     .V 0a s    M  (2
  @R@     E       ���  �  (.G  ��  ��  �j ).V
  �  �  X6  *.V
  ��  ��  E  ,2
  �  
�  &  �� 1�  a�  ]�  :bR@            ߼  �1  6�%  ��  ��  pR@     Ts Qv   ]R@     .V 0a �U   p6  �>
  �Q@     g       �ν  �  �*G  ��  ��  �j �*V
  E�  ;�  X6  �*V
  ��  ��  PE  �>
   �%  �� �  =�  9�  �W  �%  {�  s�  '�%  ��  �1  �%  ��  ��   	R@     .V 0a s    \F  �|
  `K@     �       �Q�  �  �&G  U<M  �&>
  �  �  2�  �&#  .�  *�  � �|
  h�  d�  -�u  � L@      �W  �V
  pJ@     i       �+�  �  �G  ��  ��  �j �V
      �0  ��A  {  q  E  �V
  �  �  n�  �>
  0 ( &�J@     *       � �}  �\
H ��%  � � �J@     Us T�\   �2  qV
  �J@     u       �8�  �  q G  � � �0  r �A    E  tV
  _ W n�  u>
  �\8�  K@      �!  {�  W�  � � J�  � � �!  d�  ; 3 <�U K@            r�  � � K@     T0    1K@     Q�  Us T0Q�\  W)=  T>
  ��  �  T G  �j U V
  E  W>
  ?
H \�%    �3  |
  �@     3      �r�  �M �%  � � =R  �
  Z R ��  �  � � '1  !r�  @ 6 � #|
  ���  $G  � � R�  %�  � � 
H &�%  6 & -�0  J�@     -�u  D��@     �  �@      �D  K�  +�  � � �D  8�    E�  C A R�  i g L  ��@      �D  ��  (L  � � L  � � �@     Us   ��@     U~    9�@     O  5�  U Q�� 9d�@     Q�  U~ T�� ��@     �M  U T8Y��  �%  6�F  ���@     6      ��  
H ��%  � � D  �  �G  � � R�  ��  � � � �|
  �Li �2
  -	 !	 j �2
  �	 �	 `D  �2  ��  �	 �	 �  ��@      ��@     &       �  +�  +
 '
 &��@     &       8�  d
 b
 E�  �
 �
 R�  �
 �
 L  ��@      ��@     	       ���  (L  �
 �
 L  �
 �
 ��@     Us Tv   ��@     Uv    *�@     �M  T8Y�L    T�1  �`�  
H �#�%  �M ��%  �  �G  R�  ��   (6  �2
  �I@     Q       ���  �� �%�  Ui �2
  '   B2  �|
  �P@     �       �2�  �  �G  � � �� ��  S C cur ��    �� ��  o k Q@     �  Uv   �=  �|
  PI@     ~       ���  �  �#G  U= �#�  � � cur ��  � � �� ��  _ ] f�I@     �  �9  b|
  �H@     �       ���  �  b$G  � � � c$o
  9 + �9  d$2
  � � �I  e$R!  � } YM  gF  * & P� h|
   'p!  ��  ~ q  d ` �O  q�
  � � �H@     T	C.H       @I@     U�UT�TQ�QR�R  �-  |
  �F@     �      ���  �  G     �U  >
  � � B7  >
  u m �M  >
  � � �I  �  � � � |
  3 ) K1 i  � � '�   ��  3T  7�  � � :T  8�  e ] e? �G@      !  ?5�  �? � � �?  � v? k c !  �? � � �? �? "  �? � � �? � � �? | v   7e? �G@      @!  B�? � � �? ) # v? � � @!  �? � � �? �? F @ �? � � �? � � �? � �    t> )G@       �  2H�  �>  	 �> 1 / #FC )G@      0   �aC W U WC } { 0   kC � � wC  �    t> VG@      `   3��  �> �  �> � � #FC VG@      �   �aC � � WC � � �   kC   wC s o    G@     Us T�TQ�QRv   �6  �|
  PF@     i       �{�  �  � G  � � �<  � >
       �X  � >
  q  g  Mreq ��  �P�F@     ,�  Tw   �(  �|
  �E@     �       �,�  �  �!G  �  �  :  �!b
  >! 8! h6  �!b
  �! �! �2  �!>
  F" :" �2  �!>
  �" �" Mreq ��  �PF@     ,�  Tw   �Z  x|
  �D@     �       ���  �  x%G  Q# G# ;req y%�  �# �# � {|
  d$ Z$ �M |6"  �$ �$ -U }V
  �h��  pE@      pE@            �Q�  ��  :% 4% ��  �% �% ��  �% �% ��  & & &pE@            �  �  �  �E@     \G Us T�TRr    98E@     f�  T�T �E@     ��  ~�  Us  �E@     ��  Us   W�@  B|
  ��  �  BG  -U C2
  � E|
  �M F6"   6�=  ��@@     �      �_�  �  �(G  [& O& ;req �(�  �& �& N ��B  �' �' -�>  ) B@     0  w �J
  I( /( h �J
  x) X) �R  �J
  �* �* �R  �,J
  , �+ > �A@      p  �  0> - - %> P- L- p  ;> �- �- F> �- �- Q> /. +. \> k. e. g> �. �.   > �A@      �  ��  0> S/ M/ %> �/ �/ �  ;> �/ �/ F> \0 T0 Q> �0 �0 \> 1 
1 g> �1 ~1   t> WB@       �  -�  �> �1 �1 �> 2 2 #FC WB@      P  �aC ]2 [2 WC �2 �2 �  kC �2 �2 wC 
3 3    t> �B@      0  .��  �> G3 E3  �> #FC �B@      �  � aC WC m3 k3   kC �3 �3 wC �3 �3    > C@      �  %/�  0> �3 �3 %> 64 24 �  ;> r4 l4 F> �4 �4 Q> 5 5 \> O5 K5 g> �5 �5   g�B@     �  1�  Uu Tt  GC@     e? I�  Uz  bC@     e? U{    6P  �@?@     ^      ��  �  � G  U-U � V
  6 	6 N ��B  R6 F6 �� ��  �6 �6 > {?@      �  �I�  0> �7 �7 %> �7 �7 �  ;> H8 B8 F> �8 �8 Q> 9 
9 \> N9 D9 g> #: :   > �?@      �  ���  0> �: �: %> ?; 1; �  ;> �; �; F> y< i< Q> G= == \> �= �= g> �> �>   g�?@     �  ��  Tt  go@@     �  ��  Tt  ,�@@     �  Tt   h@C  ��@     �       �a�  �  �2G  UN �2�B  Tt> �@      0  ���  �> �? �? �> �? �? #FC �@      p  �aC (@ &@ WC N@ L@ �  kC �@ |@ wC �@ �@    t> �@      �  �V�  �>  A �@ �> &A $A #FC �@      0  �aC VA TA WC |A zA 0  kC �A �A wC �A �A    t> �@      `  ���  �> .B ,B �> XB RB #FC �@      p  �aC �B �B WC �B �B p  kC C C wC TC PC    7t> @      �  ��> �C �C �> �C �C #FC @      �  �aC D D WC BD @D 0  kC tD pD wC �D �D     6�D  u�>@     �       ���  N u6��  U�  v6�  �D �D �  x�  JE DE  �  WL  ;|
  7�  �  ;#G  `req <#�  �X  =#�	  5  >#F5  %i @2
  %w AJ
  %h AJ
  ?�� [�    �\  |
  �=@     �       ���  �    �E �E � |
  )F %F K1 i  kF aF R�  �  �F �F �  G  BG 8G D� �  �G �G �I  �=@      �=@             "9�  �I  H H �I  CH =H &�=@             �I  �H �H   �H  �=@      p  %��   I  �H �H �H  �H �H p  I  I  �=@     O Uu Tr    L  �=@      �=@            &��   (L   L  �=@     U}   >@     l U} Ts Q|   U/  �
|
  ��@     6      �e�  �  �
G  )I I �Y  �
e�  �I �I � �
|
  ��R�  �
�  J J K1 �
i  SJ QJ �M �
6"  zJ vJ �  �
  �J �J D� �
�  RK @K �8  �
�  L L >�u  �
L  ��@      ��@            9�  (L  �L �L L  �L �L �@     Uv T}   L  5�@      5�@             ��  (L  �L �L L  M M C�@     Uv T   {I  ��@      �@  �
��  �I  ;M 9M �I  `M ^M �@  �I  ��@     �N Uu Tt    �@     O  �  Uv Q�� *�@     O  /�  Uv THQ�� ^�@     O  T�  Uv THQ�� x�@     U}     A*  �
|
  �<@     �       ��  �  �
G  �M �M � �
|
  �M �M K1 �
i  @N >N R�  �
�  eN cN D� �
�  �N �N �I  =@      =@            �
X�  �I  �N �N �I  �N �N &=@            �I  O O   �H  ;=@      @  �
��   I  7O 5O �H  \O ZO @  I  I  J=@     O Uu Tr    L  J=@      J=@            �
��   (L   L  R=@     U|   `=@      U| Ts Qv   }K  �
|
  �<@            �N�  �  �
G  U �:  g
|
  0�@     �       ��  �  g
$G  �O �O IE  h
$�  �O �O Jy  j
p  �X� k
|
  WP OP K1 l
i  �P �P �M n
6"  
Q Q >�u  �
� ��@       ��@     6       �
��  � CQ AQ � jQ fQ <DS ��@     1       � �Q �Q /�e  ��@      P?  ���  �e  �Q �Q ��@     U|   8L  ˔@      ˔@     	       	 (L  L  �Q �Q Ԕ@     Us T|     f�@     
 ��  Ts Q�X ��@     Uv T|   )  ^  Q
|
  �@     6       ���  �  Q
 G  R R OF  R
 �  lR dR j�  T
)  ��6�@     N�  U�UTw   ��8  	|
   �@     C	      ���  k  	/[   S �R ��  	/��  UU -U �  	/J
  W �V �H  	/��  �W �W -  	/�	  DX "X � 	|
  ��|K1 	i  �Y �Y R�  	�  �[ �[ Jy   	p  ��|�  !	G  ��|D� "	�  6] $] �7  #	�	  ^ �] cur $	��  �^ �^ �� %	��  K_ C_ -�L  �	��@     -pW  �	$�@     -�0  4
i�@     -lE  �	��@     -�u  :
�@     '�J  ��  G  Q	2
  �_ �_ G  R	#  �_ �_ �@     �  U��|T��|Q} R��|  '�K  e�  G  s	2
  O` I` G  t	#  �` �` ~e  5�@       �K  �	 �  �e  �` �` �e  a a �K  �e  ~a za N�@     U��|T0Q0R0   � -�@       -�@     1       �	�  � �a �a � �a �a <DS 6�@     (       � b b /�e  >�@      L  ���  �e  =b ;b H�@     Us   8L  Q�@      Q�@     	       	(L  bb `b L  �b �b Z�@     Uv Ts     ��@     �  >�  U T��|Q} R��| ��@     �c U��|Q��|R��|  :��@     2       ��  �  �	  ��~��@     ��  T��~  :�@     �       ��  i �	2
  �b �b 0K  �� �	�  �b �b   ' N  �  �8  
  c 
c  {I  T�@       K  �	_�  �I  Hc Dc �I  �c ~c  K  �I  b�@     �N Uu Tt    � ��@      ��@     4       �	@�  � �c �c � �c �c <DS ��@     /       � d d /�e  ��@      `K  ���   �e  Ϸ@     Us   8L  ޷@      ޷@     	       	 (L  L  2d 0d �@     Uv Ts     ��  ��@      @L  �	 �  ��  id Ud ��  De :e ��  �e �e ��  Bf @f ��  qf gf @L  ��  �f �f ��  ��@      ��@     �       �G�  3�  g }g &�  �g �g �  �g �g �  �g �g &��@     �       4@�  ��~M�  h h Z�  \h Th g�  �h �h \t�  ~e  ��@      �L  U��  �e  �i �i �e  �i �i �L  �e  �i �i Ϲ@     Us T0Q0R0    e  ��@      �L  Y�  )e  j j e  Fj @j  e  	�@     #d  Us T0Q��|R�  ��@     ��  U��|Ts R��|X��|   ��  ��@      M  	��  <�  �j �j /�  -k %k "�  �k �k  �  �  	l �k M  I�  �l �l V�   m m c�   n �m 4n�  ��}4{�  ��~4��  ��}��  �n �n ��  o �n 4��  ��}4��  ��|� H�@       H�@     A       ���  � zo xo � �o �o <DS M�@     <       � �o �o /�e  U�@      �M  ���  �e  p p m�@     U��|  8L  �@      �@     
       	(L  Tp Rp L  yp wp    �x  ��@      �M  �!�  �x  �p �p �x  q q  L  ɽ@      ɽ@            �	s�  (L  <q :q L  aq _q н@     U~   ��@     y  ��  Us R��}X��|Y��} �@     
 ��  U~ T��}Q��| C�@     ��  U~ R��|X��|   �@     ��  U��|Ts Q0R��|X��|   � غ@      غ@     -       �		�  � �q �q � �q �q <DS �@     $       � �q �q /�e  �@      �M  ���  �e  �q �q �@     Us   8L  ��@      ��@     	       	 (L  L  r r �@     Uv Ts     � '�@       '�@            c	K�  � Cr Ar � hr fr  ��@     
 p�  Us Tv Q��| 8�@     O  ��  U��|THQ��| y�@     @ ��  T0 �@      ��  U��| K
�@     k�  K�@     k�   6  G  �?  	|
  `�@            ���  k  	&[  �r �r ��  	&��  �r �r �  	&J
  	s s �H  	&��  Fs Bs ,k�@     ��  U�UT�TQ�QR�RX1  =QT  �|
  ��  k  �'[  Jy  �'p  �  �'J
  �H  �'��  ��  �'��  � �|
   =?^  {|
  ��  k  {5[  Jy  |5p  �  }5J
  �H  ~5��  ��  5��  R�  ��  � �|
  %i �>
  �8  ���  �P  ���  +  ���  �K  ��	  A+  ��	  m-  �)  �7  �p   1�   ��  2-    1J
  ��  2-    1|
  ��  2-    =/?  H|
  ~�  k  H[  Jy  Ip  �  JJ
  �H  K��  � M~�  � N|
  FJ  OJ
  x  OJ
  >�u  u 1�  ��  2-    CRW  |
  P�@     �      �K�  k  [  �s s Jy  p  >u $u /U  J
  [v Wv �  J
  �v �v �H  ��  [w Ww R�  �  �w �w � |
  sx Ux ��  J
  ��y^  J
  ���P  ,  ��.� J
  ��' G  ��  �N  6J
  �y �y K�  %�@      pG  9��  ��  %z z ��  �z �z ��  s{ k{ w�  �{ �{ j�  D| 6| ]�  �| �| pG  ��  �} |} ��  S~ A~ 4��  ����  "  ��  � � ��  ��  l� `� G�  ��@     ~e  E�@       H  ���  �e  �� � �e  2� .�  H  �e  l� h� c�@     Us T} Q0R0   ~e  �@       @H  �B�  �e  �� �� �e  � ށ @H  �e  � � �@     Us T} Q0R0    e  \�@      �H  ���  )e  V� T� e  }� y� e  �� �� a�@     #d  Us Q| R   L  ��@      ��@     <       ���  (L  � � L  � � ״@     U��~T|   ��@     �Z  �  Us T�� Ү@     �c X�  Uv Ts Q| R��~0V�  00c�  0 4�@     O  �  U��~T Q�� ��@     ��  Uv T| Q R0Y��~   7L  ��@       �H  ;(L  A� 9� L  �� �� ϯ@     Uw    �  �@       0I  %v�  c�  � �  V�  I�  �� �� <�  � � /�  څ ȅ "�  �� �� 0I  4p�  ��}�  �� �� ��  ^� J� ��  L� 0� ��  �� r� ��  9� 7� ��  r� \� ��  f� T� ��  P� ,� ��  ׎ Î ��  �� �� ��  �� �� G
�  Ͱ@     G�  �@     ~e  ��@       �I   s�  �e  ِ Ր �e  � � �I  �e  M� I� L�@     Us Tv Q0R0   ~e  =�@       0J  :��  �e  �� �� �e  ڑ ֑ 0J  �e  � � �@     Us T��~Q0R0    e  
�@      `J  �`�  )e  P� L� e  �� �� e  � � �@     #d  Us R'��~20��~#������������������+(   L  \�@      \�@            ���  (L  � � L  8� 6� j�@     U��~T   j�@     �Z  ��  Us T�� u�@     O  �  U��~T��~Q�� �@     �Z  !�  Us T�� 2�@     .]  @�  Us T�� ��@     ��  Uv T R0X	/H     Y��~   L  Ͱ@      �J  '��  (L  a� ]� L  �� �� �@     Uw T~   ��@     �  ��  Uv Ts Q�QR��X�� ׭@     Mz  "�  Uv Ts XTSOPY1 �@     Mz  Uv Ts XtnfsY0  =�+  �|
  �  k  �'[  Jy  �'p  �P  �',  o;  �'J
  �  �'J
  �H  �'��  R�  ��  �5  �6  � �|
  �T  �V
  �O  �J
  �4  �S   �-  �J
  >�u   =.8  �|
  �  k  �'[  Jy  �'p  �P  �',  o;  �'J
  �  �'J
  �H  �'��  � �|
  R�  ��  }U  �6  %i �S   � �S   ?1  �S   %len �V
  J0  �V
  cN  �V
  �1  �"V
  �O  �V
  /� �V
  >�u  �>w\  � =�S  �|
  ��  k  �1[  Jy  �1p  �  �1J
  G  �12
  G  �1#  �H  �1��  � �|
  R�  ��  x  �V
  ss  �V
  %pos �V
  �/  ��	  QI  �6  >�u  �?�;  �|
    =\C  H|
  ��  Jy  H+p  �  I+J
  x  J+F5  ss  K+F5  �/  L+�  � N|
  eT  O&
  �P  PJ
  %tag QV
  %i RS    C(Q  |
  ��@     F      ���  k  '[  � Փ 2�  '6  �� �� �  'V
  g� W� �  'J
  (� � �,  '�  � ۖ �H  '��  <� ,� ��  	)  ��� 
|
  �� � Jy  p  �� �� R�  �  � � ��  ��@      PN  \�  ��  '� #� ��  s� o� ��  �� �� ��  � � ��  W� Q� PN  4��  ����  ��  �� �� \�  �e   �@      �N  �9�  �e  � � �e  ,� *� �e  Q� O�  �@     O  U TPQ��   �e  ��@      ��@            5��  �e  v� t� ��@     Us   L  ��@      ��@            6��  (L  �� ��  L  ��@     U Ts   L  ˿@      �N  =�  (L  ě �� L  � � տ@     U Tv   Q�@     ��  ]�  U} T��~ m�@     ��  U} T��Qw R| X0  =
H  �|
  �  k  �+[  2�  �+6  �  �+V
  =9 �+�  �/  �+�  � �|
  R�  ��  Jy  �p  >�u  � p  q-9  �P@     /       ���  Jy  �#p  =� 7� R�  ��  �� �� 7L  T@       �   �(L  �� ��  L    ?W  �|
  �@     F       �U�  k  �'[  ڜ Ԝ �S �'�	  .� &� �]  �'J
  �� �� �  �'J
  �� �� �H  �'��  f� ^� ��  �)  ��J�@     ��  U�UTw Q�RR�XX1  5*  ~|
  p�@     >       ��  k  ~[  ˞ Ş SF  �  � � �  �J
  �� � �H  ���  ן џ ��  �)  ����@     ��  U�UTw Q�QR�RX1  C�E  |
  ��@           �O K1 i  /� #� �/  �  �� �� �7  �	  "� � �  J
  _� [� G  2
  �� �� G  #  � �� �H   ��  � R�  "�  >� :� �M #6"  x� t� �  $G  ¢ �� �8  %  �� �� � '|
  ��	*  '|
  ;� 9� >�0  g: �@     I       i�  i @S   `� ^�  )  �@       @  j   D �� �� 7 ݤ Ӥ  @  Q ��@     [M ��  U~ Ts  �@     [M ��  U~ Ts  c�@     [M U~ Ts    L  Ø@      P@  mL  (L  P� L� L  �� �� ј@     Us T   L  ј@      ј@            n�  (L  å �� L  � � ߘ@     Us T~   ��@     O  �  Us Q�� 
�@     O  �  Us T�Q�� 9��@      T~ Q���R} X�� 9Ø@     ' U~  3�@     � ? Uu  ��@     U0  =3I  ��  � �  �+G  N� ��  %end ��  %cur ��   C�T  �|
  �@     z       �� �  �"G  UN� ��  � � cur ��  8� 0�  T�^  � K1 �i   q33  Q ;@           �) R�  Q�  �� �� �  RG  � � K1 Si  �� �� �M U6"  � ާ rG  A;@      0  b �G  � � �G  *� (� �G  O� M� �G  �� {� 0  �G  ];@     `O Us�T	p@     Qv R}    ) v;@      v;@            m~ D Ҩ Ш 7 �� �� &v;@            Q �;@     [M Us Tv    � �;@       `  tW �  � � � �� �� DDS �  � ߩ ۩ /�e  �;@      �  � �e  � � �;@     U|   8L   <@       <@     
       	(L  <� :� L  a� _� 
<@     U~ T|     L  �;@      �;@            }� (L  �� �� L  �� �� �;@     Uv   L  �;@        � (L  Ԫ Ϊ L  &�  � @�;@     U�UT�T  K5;@     B 9v;@      Us  �;@     Us   TZ  7l �  7 G  R�  8 �  %n :2
  ?
H B�%    h9J  !p@     X       �� R�  !�  z� r� �  "  � ٫ K1 #i  F� @� L  �@       �@            - (L  �� �� L  �� �� �@     Uv   L  �@      �   .j (L  � ܬ L  4� .� @�@     U�UT�T  9�@     ~ Us  �@     Us   �J  |
   k@     F       �� �  G  �� �� ��  V
  � �� :1  k  X� N� �^ >
  Ю ʮ 8�  k@      k@            � W�   � � J�  [� Y� &k@            d�  �� ~� <�U k@            r�  Я ί #k@     T�T    ,@k@     � U�UQ�Q  7  �|
   a@     =      �� �  �G  	� � �^ �>
  � � :1  �k  $� � � �|
  @� $� K1 �i  j� `�  �u  � ݴ k  �[  t� n� P�	   �	   �%    ȵ �� e5  i:  :� $� -�6  ��b@     >�u  '@0  '	 �� J-  *� $� �6  K�	  {� w� �g@     l 	 U|  �g@      l T	/hH       '�/  �	 Zy  i R#  �� �� '�/  �	 �8  }  ܷ ط $  ~2
  � � ve@     U Ts R~ Xv   e@     Us Q~   '`-  �
 N ��B  C� ;� e? �b@       �-  �!g
 �? �� �� �? � � v? /� '� �-  �? �� �� �? �� �� �? 8� 2� �? �� �� �? ʺ º �? 3� -�   7e? c@       �-  �!�? �� � �? �� �� v? �� �� �-  �? i� _� �? � ߼ �? !� � �? �� �� �? ɽ �� �? 2� ,�    '�-  j �8  �  �� ~� 0.  9X  ��  Ӿ ; ��  _c@       p.  �!) �  $� � �  $� � p.  �  s� m� )�  Ŀ �� 6�  %� � 8D�  {c@      {c@     +       �p�  �� �� c�  �� �� V�  ,� $� &{c@     +       }�  �� �� ��  �� �� \��  D�V �.  ��  0� ,�      ��  �c@      �.  �	� �  i� g� �  �� �� �.  �  )�  �c@     �H Uu T|    1�  �f@       /  �� Y�  �� �� L�  �� �� ?�  �� �� /  f�  )� #� q�  u� s�   ��  h@      @/  �L ǎ  �� �� ��  �� �� @/  Ԏ  �  h@     �J U} T|    �c@     Ts Q| R|    'p/  � �� �-  � �� f"d@     ��  6d@     E Us Q0  � =a@      �,  � � |� z� La@     A Us   � �e@      0  �O � �� �� � �� �� 0  � � � � W� Q� � �� ��   9�b@     o Us Q~ Rv  �e@     =�  U}   TK  ��  �0u  �(  �0�	  N ���  �� ��  u� ��   6�4  �<@     �       �B �  �!G  U:  �!�  !� � � �!�  q� m� �8  �  �� ��  6�M  d`:@     �       �@  d$u  �� �� �  K1 hi  e� ]� R�  i�  �� �� �� ju  Z� P� cur ku  �� �� L  �:@      �  � (L  b� \� L  �� �� @�:@     T�U  9�:@     * Us  �:@     � Us    �D  /|
  Е@     �      �� �  /$G  �� �� a/  0$� �� �� � 2|
  ��K1 3i  <� :� �M 46"  a� _� R�  5�  �� ��  6u  �� �� -�u  Z.�@     l E�@      �?  H$ ~ �� �� �?  � �� �� � L� D� � �� �� 4� ��� � �� G� ��@     �0 "�@      �?  /� �0 �� �� �0 �� �� �?  �0  � � 4�0 ��'�@     O  U~ T�Q��   z�@     O   U~ THQ�� ��@     U|    L  ;�@      ;�@     
       L	| (L  l� j� L  �� �� E�@     U} T|   �@     O  � U} Q�� ;�@     � U|   u  h:/  07@     }       ��  $u  �� �� K1 i  � � �M 6"  W� U� R�  �  � {� L  x7@      x7@            '{ (L  �� �� L  �� �� �7@     U|   (. �7@       �7@            #	� 5. � � K�7@     7R  9X7@     � Us  `7@     A Us   T�G  �  �%u   T)  �|
  P�@     x       ��  �,u  .� &� �  �,V
  �� �� R�  ��  �� �� � �|
  �\L  ~�@       ~�@            �� (L  0� .� L  U� S� ��@     Uv   ��@     O  Uv T| Q�\  6�U  �@:@            �E  �*u  ~� x� B� �*6  �� �� Q:@     A Us   6ZJ  N�7@     �      �A  N1u  &� � �� O1-  �� �� �\  P1�  7� +� �S  R�B  �� �� �I S�B  z� t�   U�  �� �� C!  W-  ���B  X�  |� v� M  Y�  �� �� �=  Z�  	� � �� Z�  X� R� ��  [�  �� �� �  [�  �� �� �  [�  E� ?� -�e  �X8@     �  �7@      `  i� ��  �� �� ��  �� �� `  ��  ��  ��  Β  �8@     �G Tw    09@     ,l  Uw T�@Qs  j9@     ,l U��T�HQs   H{X  :l  :+u  ?R�  >�    =�;  |
  �  $u  K1  i  �M !6"  R�  "�  � #|
  �8  $�  >�u  4 Y�:  �
 !Jy  �p  !�Z  �2
  ?*R�  ��    )2  �|
  `�@     Z      �� k  �'[  "� � ��  �'��  �� �� �/  �'�  !� � E� �|
  �LR�  ��  �� �� Jy  �p  � �� e�u  ��@     N�e  ��@       ��@     ,       �� �e  �� �� �e  �� �� �e  � �  NL  �@      �@            �T (L  7� 5� L  \� Z� #�@     U~ Tv   /L  /�@      �>  �� (L  �� � L  �� �� j�@     U~   ��@     O  � U~ TPQ�L L�@     9l Uv   b%[  �P6@            �G pw  �%+  � � � �%|
  K� E� �P  �G �� �� a6@     Fl U�UT1  A  )�7  �2
  @6@            �~ Spw  �#+  U bU  z 6@            �� Spw  z*+  US2�  {*�	  TS�� |*�	  QS�D  }*�+  R )�*  b�
  �5@     [       �\ K[  b+�#  �� �� �1  c+�  I� =� E  e�
  �� �� �5  f�#  (� "� �5@     l Tv   �X  G5 �5@     #       �5 ;num G 2
  u� q� x�  H �)  �� �� hk J�(  �� �� 8� �5@       �5@            O 4� 0�   &�5@            " o� m� �5@     B$ U	�U����T�T    G   d\  :5 `5@     !       �� ;key :$�  �� �� x�  ;$�)  �� �� hk =�(  � � 7� `5@      p  B Q� M�   p  " �� �� i5@     B$ U�UT�T    =�B  .5 / `key .�(  x�  /�)  %np 1�)   �4  |
  ��@            �� ;num "2
  �� �� �U   "G   �� �� x�  !"�)  -� )� R�  ""�  j� f� %hk $�(  ,ǩ@     � U	�U����T�TQ�QR�R  �,  |
  ��@            �� ;key $�  �� �� �U  $G   �� �� x�  $�)  !� � R�  $�  ^� Z� %hk �(  ,��@     � U�UT�TQ�QR�R  VW+  �|
  p�@     >      ��  Bkey ��(  �� �� �U  �G   �� �� x�  ��)  �� �� R�  ��  � � "nn ��(  � u� "bp ��)  �� �� � �|
  V� T� -�u  
��@     �# ��@      PE   |  �# }� y� �# �� �� PE  �# �� ��  $ -� '� $ x� v� $ �� �� !$ �� �� 4,$ ��G8$ ��@     /L  |�@      �E  �*  (L  � � L  O� K� ��@     U~ T   3�@     �M  f  U~ T8Q0R
| 1$����X0Y�� l�@     B$ Ts    ��@     B$ �  U| Ts  Ҩ@     O  U~ T@Q��  bUP  ��4@     y       ��! x�  � �)  �� �� R�  � �  �� �� @  "sz �>
  W� S� "bp ��)  �� �� "i �>
  �� �� NL  5@       5@            �	�! (L  �� �� L   � �� 5@     Uv   rL  25@      25@            �(L  %� #� L  K� I� @5@     Uv Ts     )�-  �|
  @�@     V       ��" x�  � �)  t� n� R�  � �  �� �� #~# J�@       �C  ��# � � �# f� d� �# �� �� �C  J�# �4�# �l��@     �M  U�TT8Q0R�X0Y�l    )�-  �|
  `�@     V       �~# x�  � �)  �� �� R�  � �  � � #~# j�@        T  ��# n� h� �# �� �� �# �� ��  T  J�# �4�# �l��@     �M  U�TT8Q0R�X0Y�l    Z�3  �|
  �# !x�  ��)  !�E  ��	  !R�  ��  (sz �>
  *� �|
   Z�P  �|
  B$ !x�  ��)  !R�  ��  (obp ��)  (bp ��)  (nbp ��)  (i �>
  (sz �>
  *� �|
  ��u  � V�0  j�)   @     k       ��$ Okey j�(  �Xx�  k�)   � � "res mV
  p� l� "bp n�)  �� �� "ndp o�)  �� �� 9@     �$ U�X @@     T�X  V3  _�	  �@            �"% Oa _")  UOb `")  T V�)  S�	  P@     #       �v% Ba S")  
� � Bb T")  G� C� Ki@     l  V�X  BV
  �@     H       ��% Okey B!)  U"num DV
  �� �� "res EV
  �� ��  Vg\  3V
  `@     1       �'& Okey 3!)  U"kp 5�  �� �� "res 6V
  �� ��  �=  
m|
   �@     �      ��' �  
m.k  <� 4� �% 
n.k  �� �� � 
p|
  
� � 2]  
q>
  p� h� [  
r>
  �� �� '�B  �' out 
x�B  � � in 
y�B  /� -� �- ڢ@       C  
�.' . Z� T�  C  . �� �� . �� ��   ��@     �k H' Q�� ��@     �k `' Q  ��@     �k �' Q
} ����1$ ^�@     �k �' Q  o�@     �k Q   I�@     �* Us T Q}   6o+  
H�4@     Y       �q( ��  
H'k  U2�  
J�  R� P� �� 
K�  y� w� �V  
M2
  �� �� a=  
N2
  �� �� n 
O2
  � � f�4@     q(  6�A  
8 4@     w       �[) ��  
8+k  U�� 
:�  A� ?� �- 4@        
A�( . i� g�   . �� �� . �� ��   8�, `4@      `4@            
B- �� �� &`4@            - �  � $- )� '�    aG  
|
  ��@            ��* ��  
2k  Y� O� `W  
2>
  �� �� R�  
�  � � � 
|
  �\�:  
>
  O� E� �<  
>
  �� �� 2�  
 �  � �� �� 
!�  �� �� -�u  
1��@     �, &�@      �C  
.{* - � � �C  - S� O� $- �� ��   �@     �M  T0Rs ����Y�\  )],  
�|
  ��@     9      ��, ��  
�/k  �� �� Z�  
�/>
  �� �� �  
�/>
  �� �� R�  
��  l� d� E� 
�|
  ��2�  
��B  �� �� �� 
��B  �� �� J}  
��	  {� o� �:  
�>
  � � �<  
�>
  �� �� -�u  
t�@     �- .�@      .�@     F       

�+ . b� `� &.�@     F       . �� �� . �� ��   y�@     �M  ,, U} T@Q��R~ Y�� ��@     �M  ^, U} T1Q��R~ Y�� �@     �M  �, U} T2R| ����Y�� ��@     P. �, Us  �@     �M  �, U} T@Q
 1$����R
v 1$����Y�� �@     Rl Q��4$  afP  
�1- !��  
�4k  *2�  
��  *�� 
��   )g?  
�|
  P�@     �       ��- ��  
�/k  �� �� E� 
�|
  �lR�  
��  (� &� /�- ��@      pB  
��- . N� L� pB  . s� q� . �� ��   u�@     �M  T@Q0X0Y�l  a�A  
�(. !��  
�1k  *2�  
��B  *�� 
��B   Y60  
�P. !��  
�(k  ?*R�  
��    bd^  
i�2@     �       �p0 ��  
i)k  �� �� R�  
k�      NL  �2@      �2@            
n�. (L  9  7  L  ^  \  �2@     Uv   NL  �2@      �2@            
o8/ (L  �  �  L  �  �  3@     Uv   NL  3@      3@            
p�/ (L  �  �  L  �  �  3@     Uv   NL  %3@      %3@            
q�/ (L    L  < : 03@     Uv   NL  <3@      <3@            
r+0 (L  a _ L  � � G3@     Uv   #p0 �3@      P  
z}0 � � P  �0 � � �0      YC  
X�0 !��  
X*k  *2�  
Z�  *�� 
[�   I�:  
F|
  �0 !R�  
F(�  !*R  
G(�0 *��  
Ik  *� 
J|
   k  -  �2
  �1@     �       ��1 oT  ��  ] Q n/  ��    bX  ��  � � hX  ��  � � ax ��  + # ay ��  � � 9@  ��  � � �@  ��  5 3 �5  ��  Z X  V  �2
  �1@            �J2 oT  �"�  Un/  �"�  � } bX  �"�  QhX  �"�  � � � ��  � �  02  }  �/@     �      �g3 ��  "�  Ux_ 
k  @ : y_ k  � � b k  � � z k   � x }  R L y }  � � u }  	 � v }  (	 $	 l }  p	 ^	 sx 2
  3
 +
 sy 2
  �
 �
 ��  2
  �
 �
  6]  �/@     �       �w4 ��  �1�  9 1 :  �1�  � � C�  �1J
  � � xz ��  ? 9 yz ��  � � val �J
  � � =/@     e?  4 Uv Qz  S/@     e? >4 U} Qz  h/@     e? \4 Uv Qz  z/@     e? U} Qz   6)S  ��-@     !      �W6 ;a �0�  [ S ;b �0�  � � C�  �0J
   	 xx �o
  ] [ xy �o
  � � yx �o
  � � yy �o
  � � val �J
  > 6 #.@     e? \5 Uv T��Qz  =.@     e? �5 U~ T| Qz  T.@     e? �5 Uv T Qz  i.@     e? �5 U~ T} Qz  �.@     e? �5 U~ T��Qz  �.@     e? 6 Us T| Qz  �.@     e? 66 U~ T Qz  �.@     e? Us T} Qz   �1  �|
  +@     �      ��9 :  �!�  U� ��  � � xx ��  � � yy ��  � o t>  +@       0  �M7 �> n l �> � � #FC  +@      �  �aC � � WC � � �  kC    wC G C    t> F+@         ��7 �> � � �> � � #FC F+@      �  �aC � � WC � � �  kC   wC ] Y    > v+@      �  �Q8 0> � � %>  � �  ;> � � F> K ; Q>    \> � � g> � �   > �+@      @  ��8 0>   %> � s @  ;> ? / F>  � Q>  � \> g> U Q   > �+@      �  �39 0> � � %>   �  ;> � � F> � � Q> \> g>   �   7> �+@      �  �0> @ 6 %> � � �  ;> 8  (  F> �  �  Q> \> 4g> P   68[  ��)@     Q      �> ;a �)�  �! �! �b �)�  Txx �o
  " �! %xy �o
  yx �o
  �" �" %yy �o
  t> �)@      P  �
�: �> F# D# �> l# j# #FC �)@      �  �aC �# �# WC �# �# p	  kC �# �# wC 8$ 4$    t> &*@       
  �
%; �> u$ s$ �> �$ �$ #FC &*@      �
  �aC �$ �$ WC �$ �$    kC % % wC R% N%    t> 1*@      �  �
�; �> �% �%  �> #FC 1*@      0  �aC �% �%  WC �  kC wC    t> 1*@      0  �
< �> �% �% �> & �% #FC 1*@      �  �aC '& %& WC M& K& p  kC u& q& wC �& �&    t> 1*@        �
�<  �> �> �& �& #FC 1*@      �  �aC ' �& WC '' %' P  kC O' K' wC �' �'    t> �*@      �  �
	= �> �' �' �> �' �' #FC �*@      p  �aC 
( ( WC 0( .( p  kC wC    t> 1*@      �  �
�= �> Y( W( �> �( }( #FC 1*@     ! `  �aC �( �( WC �( �( �  kC %) !) wC h) d)    7t> �*@      `  �
�> �) �) �> �) �) #FC �*@      �  �aC �) �) WC * * �  kC E* A* wC �* �*     I5<  �J
  t> Aa_ �J
  Ab_ �J
  %s  2
  %a �  %b �  %q �  %q_ J
   I
.  �J
  �> Aa_ �J
  Ab_ �J
   )�=  �J
  �(@     V       �e? Ba_ � J
  �* �* Bb_ � J
   + + Bc_ � J
  �+ �+ "s �2
  �+ �+ "a ��  �, �, "b ��  �, �, "c ��  - - "d ��  t- p- "d_ �J
  �- �-  IjO  �J
  �? Aa_ �J
  Ab_ �J
  Ac_ �J
  (s �2
  (a ��  (b ��  (c ��  (d ��  (d_ �J
   )@:  �o
  P�@            �=@ Bx �o
  �- �- By �o
  A. =. [v ��  �`e�@     �Q  Uw   )Q  jo
  p(@            �l@ Oa jo
  U )X  ao
  `(@            ��@ Oa ao
  U )\  Xo
  @(@            ��@ Oa Xo
  U I�M  q|
  _A !�  qG  !�S r>
  !.� s>
  !?1  tk  ![5  uR!  *� w|
  *�� y!  (num {>
  (end {>
  (nn {>
  *��  |2
   )tV  K|
   j@     �       ��B �  KG  �. z. n�  L>
  {/ e/ ?1  Mk  }0 e0 �,  NR!  �1 z1 �� P!  �2 �2 '01  �B � _|
  �2 �2 /�B �j@      @1  d�B �B 	3 3 "C ^3 X3 C �3 �3 
C �3 �3 @1  .C :C ,�j@     hF U�U#�T�RQ1R�Q0�B �U   ^j@     Us T} Q1Rv X|   ,�j@     �@ U�UT�TQ1R�QX�R  ZM-  |
  FC !�  'G  !\-  'R!  !.� '>
  !?1  'k  *��  o
  (nn !>
   Z�6  �k  �C Aa �k  Ab �k  (ret �.  (tmp �.   �W  �@     �       �D �W  ,4 "4  �W   �W  �W  �4 �4 �W  �4 �4 �W  @6 .6 �W  7 �6  X  �7 �7 
X  �7 �7  EW  `@     �       ��D  RW   RW  ^W  �8 �8 jW  �9 �9 tW  �9 �9 ~W  9; ); �W  �; �; �W  N< H< �W  �< �<  X  ` @     \       ��D  (X   (X  4X  �= y= >X  �= �= HX  O> E>  ��  � @     7      �hF �  �> �> �  s? _? +�  b@ J@ 8�  wA _A E�  �B tB R�  C C _�  l�  y�  ��  ��  D��  p  R�  �C �C E�  �C �C 8�  AD -D +�  ,E E �  F F �  �F �F p  _�  9G 1G l�  �G �G y�  �G �G ��  7H 3H ��  sH mH ;!@     l 
F Ts  9^!@     %F T	8.H      s�!@     MF T�QQ�RR���� @�!@     T�QQ�R    �B  "@     �       �\G 
C �H �H C  I I "C rI lI  �B .C �I �I :C �I �I #e? Q"@         3�? J 	J �? dJ ^J v? �J �J   �? KK ?K �? �K �K �? vL lL �? �L �L �? LM @M �? �M �M    ��  �"@           ��G ��  0N (N ��  �N �N ��  �N �N +��  R�  O 	O �  �O �O �  �O �O D'�  P  (�  IP AP   �  �#@     �       ��H ��  �P �P +��  T��  Q Q ��  UQ QQ ��  �Q �Q Β  �Q �Q <ے  �#@     Q       ܒ  +R )R �  PR NR <��  �#@     #       ��  yR sR �  �R �R    ��  @$@     �       ��J +�  U�  �R �R �  )�  0S &S t> @$@      �  	�
pI �> BT @T �> hT fT #FC @$@        �aC �T �T WC �T �T   kC �T �T wC 4U 0U    t> j$@      �  	�
�I �> qU oU �> �U �U #FC j$@         �aC �U �U WC �U �U    kC V V wC NV JV    t> }$@      �  	�
nJ �> �V �V  �> #FC }$@        �aC �V �V  WC   kC �V �V wC W W    7t> �$@      p  	�
�> [W WW �> �W �W #FC �$@      �  �aC �W �W WC �W �W �  kC %X !X wC hX dX     ��  �$@     >       ��K ��  �X �X ǎ  �X �X Ԏ  4Y 2Y �  YY WY 8��  �$@      �$@            	��  ~Y |Y �  �Y �Y &�$@            �  )�   %@     �H Us T|     &�  %@     u      �M 8�  �Y �Y 4E�  ��R�  1Z -Z _�  pZ lZ l�  �Z �Z y�  [  [ ��  �[ �[ ��  �[ �[ ��  \ \ ��  =\ 7\ ��  �\ �\ �  !%@       !%@            	&�L ��  �\ �\ ��   ] �\ &!%@            ��  ��  ��  Β  )%@     �G U{ Tw    <È  �%@     �       Ĉ  :] 6]   T  �&@     <       �[M +!T  U.T  x] r] �&@     �C Uu Tt Q�T0�W  u   ) �&@     �       ��N 7 �] �] D ^ ^ Q l^ h^ t\ �&@     D       �N ] �^ �^ 8�  �&@      �&@     3       E+�  �^ �^ &�&@     3       8�  �^ �^ E�  _ _ R�  ;_ 9_ L  !'@      !'@            ��N (L  `_ ^_ L  �_ �_ /'@     U Tv   !'@     Uv     8L  C'@      C'@            J(L  �_ �_ L  �_ �_ O'@     U~    {I  p'@     (       �O +�I  U+�I  T�I  �_ �_  �H  �'@     -       �`O +�H  U+ I  TI  ` ` I  @` >`  rG  �'@     m       �YP �G  i` c` �G  �` �` �G  a a �G  _a Ya �G  �a �a <�G  �'@     "       �G  b b �G  7b 5b L  (@      (@            �=P (L  _b [b L  �b �b (@     Uv   �(@     } Uv Q~    e? �(@     \       ��P v? �b �b �? c c �? �c yc �? �c �c �? �d �d �? �d �d �? e e �? �e |e �? �e �e  t> @)@             ��Q �> �e �e �> 7f 3f rFC @)@      @)@            �aC tf pf WC �f �f &@)@            kC �f �f wC g g    > `)@     P       ��Q %> Zg Tg +0> T;> �g �g F> *h (h Q> Qh Mh \> �h �h g> �h �h  p0 �2@     D       �7R +}0 U�0 i i �0 *i (i  (. �3@     #       ��R 5. Xi Pi DA. �  B. �i �i /L  �3@      �  
��R (L  �i �i L  Gj Cj @�3@     T�U  �3@     P. Us    (. �3@            �S 5. �j }j ,�3@     7R U�U  � p6@     A       ��S � �j �j � �k xk �  � l l /�e  �6@      �  ��S �e  _l [l �6@     Us   7L  �6@         	(L  �l �l L  �l �l @�6@     T�U    uA �6@     d       ��T O )m !m :�6@     *       PT ] �m �m 7L  �6@      0  A(L  �m �m L  �m �m   <A �6@            O 9n 5n <�S �6@            ]    ��  �>@     &       �U ��  xn rn ��  �n �n ��  o o +��  R�  �  �  ,�>@     \G U�UT�TQ�Q�Rr   ��  pD@     p       ��U ��  no ho ��  �o �o J��   ��  D��  �  ��  ,p $p ��  �p �p �  4��  P��  �p �p s�D@     �U T	�T $ & K�D@     _�     8�  0J@     3       �.V J�  Iq Aq W�  �q �q d�   r �q &BJ@            r�  Mr Kr OJ@     T�T   O pQ@     \       ��V  a  a n tr pr { �r �r � �r �r K�Q@     �   D�  �S@     a       ��V +V�  U+c�  T+p�  Q}�  7s 3s J��   �'  ��  us ms   ��  `V@     �       ��W ��  �s �s ˥  At 9t إ  �t �t �  %u u t��  �V@     @       �W إ  ru pu ˥  �u �u ��  �u �u &�V@     @       �  �u �u <�  �V@     @       �  7v 3v  �  pv nv �  �v �v �V@     T|     �V@     Uv T|   �@ @h@     �      ��Y �@ �v �v �@ �w �w �@ �x �x �@ �y �y A �z �z JA  #A /A �{ �{ ;A ~| n| GA RA D�@ p0  A P} @} �@ 
~ �} �@ �~ �~ �@ F 8 �@ � � p0  A �� �� #A � � /A ;A GA Z� T� RA �� �� /�B xi@      �0  ��Y �B Ӂ ˁ "C =� 5� C �� �� 
C � � �0  .C :C ,�i@     hF U�U#�T�XQ�QR�R0�B �U   9�h@     �Y U| Ts Q R} Xv  ;i@     � U| Ts Q}     �  �l@            �MZ ��  p� j� +��  T��  ��  ��  Β  ,�l@     �G U�UTt   1�  �l@     /       ��Z ?�  �� �� +L�  T+Y�  Qf�  �� �� q�  K� I�  ��  �n@            ��Z +�  U�  t� n� �  )�  ,�n@     �H Uu T�T  ��  o@            �O[ ��  Ƅ �� ǎ  � � Ԏ  �  ,o@     �J U�UT�T  &�  ps@            ��[ 8�  j� d� E�  R�  _�  l�  y�  ��  ��  ��  ��  J��   ,�s@     �K U�U  �e   x@     (       ��[ +�e  U+�e  T+�e  Q �e  0x@            �+\ �e  �� �� @@x@     U�U  ~e  Px@     B       ��\ �e  � � �e  �� �� J�e   kx@     Us Tv Q0R0  Te  �x@     ^       �!] ee  *� � qe  χ Ň #~e  �x@       �8  b�e  L� D� �e  �� �� �8  �e  C� A� �x@     Uv Ts Q0R0    6e   y@            �D] +Ge  U  e  �y@            ��] e  k� g� e  �� �� )e  �� �� ,�y@     #d  U�UQ�TR�Q  u~`  �{@     6       �$^ �`  N� H� &�{@            �`  �� �� 7L  �{@       :  O(L  ׊ Պ L  �� ��    On  Ђ@     y      ��` nn  A� 5� �n  Ӌ ɋ �n  T� H� {n  ތ ܌ an  � � �n  4� 0� 4�n  �L�n  n� j� �n  �� �� �n  �� �� �n  I� E� �n  �� � �n  �� �� Jo  Te  %�@      �;  )|_ qe  �� �� ee  6� 2� #~e  -�@        <  b�e  p� l� �e  �� ��  <  J�e   F�@     Us Tv Q0R0    Te  ȃ@      @<  A` qe  �� �� ee  8� 4� #~e  Ѓ@       p<  b�e  r� n� �e  �� �� p<  �e  � � ��@     Us Tv Q0R0    �@     �Z  4` Us T�L �@     �Z  R` Us T�L h�@     .]  p` Us T�L ��@     �Z  �` Us T�L �@     �Z  �` Us T�L 1�@     �Z  Us T�L  Jx  ��@     &       �ea \x  "� � ix  c� [� vx  ȑ  �x  � � �x  l� f� ��x   ,��@     $^ U�TT Q�X0an  �U0{n  �Q  T   �@            ��a +!T  U.T  �� �� ,
�@     M Uu T�T  �0 �@     3       �b �0 � 
� �0 b� \� �0 �� �� 4�0 �\+�@     O  Us T�Q�\  �N  ��@     1       ��b �N  � � �N  A� ;� �N  �� �� �N  �� �� �N  b� Z� ��@     U�UT�T  ��   �@     %      ��c ��  ʕ �� ��  F� <� ��   �� ɖ  >� 4� ֖  D��  �D  ɖ  �� �� ��  � �� ��  =� 9� ��  y� s� �D  4֖  �LG�  ٧@     ��@     �M  nc Uv T@Q0R~ X0Y�L ͧ@     �M  �c Uv T1Q0R~ X0Y�L �@     s�  �c Uv Ts  *�@     �M  Uv T2Q0R|  $ &X0Y�L    �   �@           �i /�  ֘  <�  �� �� I�  7� /� p�  �� �� c�  � � V�  � � 4}�  ����  =� 7� ��  �� �� ��  Ϝ �� ��  � � ��  {� m� ��  )� � G��  ��@     ��  >�@      O  �/g 7�  �� � *�  �� �� �  N� B� �  �� � �  �� |� O  4D�  ��Q�  -� � ^�  ֣ ʣ k�  j� Z� x�  � � Te  ��@      �O  c
�e qe  �� �� ee  ̥ ȥ #~e  ��@       �O  b�e  � � �e  V� R� �O  �e  �� �� ��@     U Tv Q0R0    Te  ~�@       @P  k(�f qe  ̦ Ȧ ee  � � #~e  ��@       pP  b�e  B� >� �e  �� x� pP  �e  � ܧ ��@     U T~ Q0R0    C�@     �Z  �f U T�� ��@     .]  �f U T�� o�@     �Z  �f U T�� ��@     �Z  g U T�� ��@     �Z  U T��   6e  1�@      �P  �Xg Ge  H� D�  o��  �P  �g ��  �� ~� 7~e  [�@       Q  ��e  �� �� �e  � �  Q  �e  � � u�@     U Tw Q0R0    ~e  ��@       PQ  �Bh �e  Z� V� �e  �� �� PQ  �e  Ω ʩ ��@     U T~ Q0R0    e  A�@      �Q  ��h  )e  e  � � e  -� +� S�@     #d  U Qv R��  L  ��@      ��@     '       ��h (L  R� P� L  w� u� ��@     U��Tv   *�@     O  "i U��T��Q�� ��@     ��  U} Tv Q��Rs 0s 0,( X'hH     /H     ���0.( Y��  L  ��@            ��i L  �� �� (L  �� � @��@     U�UT�T  �I  ��@     ,       �j +�I  U+�I  T�I  D� @�  {I   �@            �Mj +�I  U+�I  T�I  ,/�@     �N Uu Tt   �H  p�@            ��j +�H  U+ I  TI  I  ,�@     O Uu Tt   �H  ��@     F       �+k +�H  U+�H  T�H  ~� z� �H  �� �� <�H  ��@            �H  � � �H  +� )� &��@            �H  �H     rG  P�@            ��k �G  T� N� �G  �� �� �G  �� � �G  J� D� �G  ,_�@     `O U�UT�TQ�QR�R  L�O  �O  22v�D  �D  1 vi0  _0  1 L�\  �\  2&L�9  �9  2L�S  �S  2L_T  _T  3XL�\  �\  3.LBi  Bi  2L�,  �,  4OL�+  �+  2(wSX  SX  =w�<  �<  !EL+A  +A  #L�Z �Z 2 �   �  �  v_  $"  p�@     2       [�  X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �  B"P  V     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  D  -      n�  �  �  D  U    �  ��  �  U     D  -   -   U    �  �"  "  �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S,  0R�  UD  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��    @       @     @    %  �  2  9  ?  J       :-   �  Jz  x LJ   y MJ   )  OV  	z  B   s�  M   uJ   }  uJ  V  vJ  /  vJ   t
  x�  k	  (X  �  N    ��  N   �  	G   B� 
  L  0    %  s  %  v	  U     �  �  	X  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     z  )    Yj  �  =  N   �*  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "D  J  �  %  <�  x >)   len ?0  *� @%   %  BO  	�    `�  �  �  G   G   �  U    �  �  q�  �  G   �  G   G   U    �    
    G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  ��  0R   �U   8�  ��  @ e  �  �  �  	�  �   �  �  G   �  U   �   7  �        7   �  ?#  )  >  7    @    �  YK  Q  G   j  7  @   U    s  �w  }  G   �  7  �   �  W  0��  �  �*   e� ��  �� �  �� �>  �� �j   �� ��  ( �'  ��  �!  l%  �  �  �  -  �%  	&  2  �  ��   	=  �
  �)  �  �0  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   b   � 	  xx ��   xy ��  yx ��  yy ��   a  ��  	 	  z'  �=	  m  �7   ss  �f   �  �	    �W	  ]	  h	  U    �  ��	  �U  �U      �J	   %  �h	  �  $�	  �	  �   �	  �� "�	   �@ #�	  �U  $U    �  7
  �; 9�	   ��  :�	   L  <�	  �
  @=�
  ��  ?J   �  @J  ~  BJ  �  CJ  �  DJ   5  FJ  (B  GJ  0�  HJ  8 �	  J$
  
   s  �  uN   ��  vN  �  xJ  �
  zJ  (  {J   �  }�
  �  �#  %  k  `	��  R�  	�D   (  	�f  |  	�f  �  	�f  �  	�r  �  	��  v  	�
  �  	�z  (�%  	��  07&  	��  8G   	�f  X �  �"�  �  h  	   �M 	�   k  	  R�  	D   �  �"-  3  %  8	;z  �� 	=�   �M 	>�    	?
   r$  	@�  0 5  �$�  �  %  �	�  �� 	�   �M 	�  �  	*   �  	Q  (�� 	
7  h�� 	j  p�� 	�  x K  �     �  �,�  �   .~   �  /~  O  1~  C  2~  �  4~   d> 6G  (A  7G  0T  9f  8  :M  @�  <f  H�  =S  PE-  ?�	  X�!  D�  h:  FZ  �  GN  ��  HN  ��  IN  ��  KN  �  LN  �U  NN  ��  ON  �)�  Q,  ��  R�  ��� S�  �K1 W   �R�  XD  �Jy  Y  �%  [
  ��	  ]�	  �    ^U   ��8  `�  � L   �  �    X�,  �  ��   E-  ��	  N �$  �8  �Y  P �  *%9  ?  �  0t�  k  v   �  w�  �@ x,  ݖ yr  E-  z�	   N |�
  0�  }�  pR  ~�  x�  z  �ߣ  �*  ��I �X  ��  �f  �h  �f  ��S  ��  �4  �r  �8  �1  �  �U    �  �-   �  �J  o  �J  �L �U    �8  ��  ( �
  L#�  �  W  H�  �  J�   = K�    LZ  d  MZ   �  N   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  #   g)�  �  �   �	�G  =  	� 	   L  	�z   $  	�f  0�  	�:  8m  	�#�  h�  	�  pآ  	�7  tG   	�f  x =    �  �
  �)f  l  �   H	��  �  	�U    "  	�,  �!  	�$   ~	  8f$  �
  hZ   (  iZ  �� k�  �� l�    nJ  �  oJ   �  pJ  (�  qJ  0 y  s�    �$>  D  �  0
'�  �N  
)f   ?1  
*Z  }0  
+f  i/  
,f  � 
- 	   �  �)�  �     H	�	  ��  	��   ?1  	�r  (  	�  4  	� 	  \  	�z  0  	�U   @ +!  4  tag �   �U  �   �  	  4  `  N   
  w%   }#  �&  h  �  &     
G  E   9
�  � ;
   ��  <
~  �  =
~  �  >
r  �#  ?
r   �  L
(�  �  �  N   �,  :   �   ^$  1  �!  �!   :  ��  �  ��  �#  �Q  W  �  f  �   I$  �r  x  �  �   �&  ��  �  9  �  �  �   �   �!  H�2  �  ��   S"  �~     �2  �"  ��  �  ��   ;  ��  (%  �E  0�   �f  8��  ��  @ I  R  ��  x  =W	  H  E#b  	Q  �  @J�  �  L~   �  M*  �� O2  .� PX  �  Q�   �  Ru  (�!  S�  08'  T�  8   W!�  �  -  (l,  k  n   �M o,  ߣ  p*  �  qz   ]  k  )>  D  �  X  �  ,   w   .d  j  u  �   �  1�  �  �  �  �  �   	  K  6�  �  �  �  �   �  �  :�  �  �  �  �  �   �  >>  "  Y    �  ,  z  ,  ,  �   �  _8  >  �  \  z  ,  �  �   $  fh  n  �  z  ,  �   �  l�  �  �  �  z  �  �   #  x�  �� � 8   �  � *  H  � �  P�  � ,  X9!  � \  `l� � �  h  �   p �    ��  �  H
2x  �S  
4�   �  
5�  (  
6�  04  
7r  88  
81  @ �  
:)  �  �
=�  R�  
?D   �  
@r  n  
Ar  �  
Br  1$  
C  2�  
Ex  �� 
Fx  `�L 
HU   � �  
J  �  P       �  A    �  f  f  A   �  &M  S  ^  �   �%  *j  p  �    �   �%  -�  �  �  �   {  1�  �  �  �  ,   �  4�  �  �  ,   l  8�  �  �     �  �   �  <    �  &  �  �   �  @2  8  �  V  ,  �  r  7   �  Gb  h  �  �  �  r  r  �   �'  N�  �  �  �  �     �  S�  �  �  �  �  r  r  7  �   �  &  ���  �� �8   i'  �~  H   �~  P  �~  X�A �  `Y �A  h�#  �^  p�  �  x�  ��  �  ��  ���  �&  �U�  �V  ��!  ��  ���  ��  ��  ��  �&  �   � �&  ��  �  �  0t:  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�  �  U'S  Y  m  D   t�  �  v~   A  w~  �  x~  &  y~   !  {^  �  ��  �  �  �  G  r  �   =	  �  ��  �  �  G  �   �'  �    �  /  G  r    /   �  �!  n  ��  )�   ��  )�  �  )�   }  5  	n  O  ;�  _� =%�   ݰ  >%G   {  �  @�  �  8  �  	�    �  �  @    D  �  @    �  	�%�  __  +�  M   �  +$�  !E  -�  "!~ 1�  !�O  1�    #�,  �  p�@     #       �$�   �  �� �� %E  �   &u�@            '~ "�  խ ӭ '�O  "�  �� �� (��@     )T	`1H         d"   1  �  *`  $"  ��@     &       ��  X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �  B"P  V     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  D  -      n�  �  �  D  U    �  ��  �  U     D  -   -   U    �  �"  "  �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S,  0R�  UD  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��    @       @     @    %  �  2  9  ?  J       :-   �  Jz  x LJ   y MJ   )  OV  	z  B   s�  M   uJ   }  uJ  V  vJ  /  vJ   t
  x�  k	  (X  �  N    ��  N   �  	G   B� 
  L  0    %  s  %  v	  U     �  �  	X  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     z  )    Yj  �  =  N   �*  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "D  J  �  %  <�  x >)   len ?0  *� @%   %  BO  	�    `�  �  �  G   G   �  U    �  �  q�  �  G   �  G   G   U    �    
    G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  ��  0R   �U   8�  ��  @ e  �  �  �  	�  �   �  �  G   �  U   �   7  �        7   �  ?#  )  >  7    @    �  YK  Q  G   j  7  @   U    s  �w  }  G   �  7  �   �  W  0��  �  �*   e� ��  �� �  �� �>  �� �j   �� ��  ( �'  ��  �!  l%  �  �  �  -  �%  	&  2  �  ��   	=  �
  �)  �  �0  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   b   � 	  xx ��   xy ��  yx ��  yy ��   a  ��  	 	  z'  �=	  m  �7   ss  �f   �  �	    �W	  ]	  h	  U    �  ��	  �U  �U      �J	   %  �h	  �  $�	  �	  �   �	  �� "�	   �@ #�	  �U  $U    �  7
  �; 9�	   ��  :�	   L  <�	  N   �g  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=�  ��  ?J   �  @J  ~  BJ  �  CJ  �  DJ   5  FJ  (B  GJ  0�  HJ  8 �	  Jg  
   sH  �  uN   ��  vN  �  xJ  �
  zJ  (  {J   �  }�  �  �#b  h  k  `	�  R�  	�D   (  	�f  |  	�f  �  	�f  �  	�r  �  	�c!  v  	�
  �  	��  (�%  	�  07&  	�s!  8G   	�f  X �  �"$  *  h  	c  �M 	J!   k  	U  R�  	D   �  �"p  v  %  8	;�  �� 	=P!   �M 	>K    	?
   r$  	@�  0 5  �$�  �  %  �	A  �� 	P!   �M 	]!  �  	*   �  	�  (�� 	
7  h�� 	j  p�� 	�  x K  � N  T  �  �,  �   .~   �  /~  O  1~  C  2~  �  4~   d> 6�  (A  7�  0T  9f  8  :�  @�  <f  H�  =�  PE-  ?�	  X�!  D�  h:  FZ  �  GN  ��  HN  ��  IN  ��  KN  �  LN  �U  NN  ��  ON  �)�  Qo  ��  R  ��� S�  �K1 Wc  �R�  XD  �Jy  Y  �%  [
  ��	  ]�	  �    ^U   ��8  `�  � L   "  (    X�o  �  �A   E-  ��	  N �g  �8  ��  P �  *%|  �  �  0t�  k  vU   �  wA  �@ xo  ݖ yr  E-  z�	   N |�  0�  }�  pR  ~�  x�  z  �ߣ  �*  ��I �X  ��  �f  �h  �f  ��S  ��  �4  �r  �8  �t  �  �U    �  �-   �  �J  o  �J  �L �U    �8  ��  ( �
  L#�  �  W  H&  �  JA   = K�    LZ  d  MZ   �  N   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  &  #   g)    �   �	��  =  	� 	   L  	�z   $  	�f  0�  	��  8m  	�#D!  h�  	�  pآ  	�7  tG   	�f  x =  H  �  �
  �)�  �  �   H	��  �  	�U    "  	�o  �!  	�g   ~	  8fg  �
  hZ   (  iZ  �� k�  �� l�    nJ  �  oJ   �  pJ  (�  qJ  0 y  s�    �$�  �  �  0
'�  �N  
)f   ?1  
*Z  }0  
+f  i/  
,f  � 
- 	   �  �)�  �     H	�L  ��  	��   ?1  	�r  (  	�  4  	� 	  \  	�z  0  	�U   @ +!  w  tag �   �U  �   �  L  w  `  N   
�  w%   }#  �&  h  �  &     
�  E   9
$  � ;
�   ��  <
~  �  =
~  �  >
r  �#  ?
r   �  L
(1  �  �  N   �o  :   �   ^$  1  �!  �!   :  �7  �_  N   ��  �`   `  }`  �_  �_  �`   p`  �|  �  ��  �#  ��  �  �  �     I$  ��  �  	     �&  �    �  /    /   �   �!  H��  �  ��   S"  �~     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  �	  @ I  R  �5  x  =W	  H  E#�  	�  �  @J^  �  L~   �  M*  �� O�  .� P�  �  QP   �  R�  (�!  S(  08'  Tv  8   W!j  p  -  (l�  k  nU   �M o�  ߣ  p*  �  qz   �  k  )�  �  �  �  ^  o   w   .�  �  �  ^   �  1    "  ^  "  �   	  K  64  :  J  ^  J   �  �  :\  b  �  v  ^  ^   �  >�  "  Y�  �  �  �  �  o  o  �   �  _�  �  �  �  �  o  "  �   $  f�  �  	  �  o  J   �  l    �  4  �  �  �   #  x��  �� � �   �  � *  H  � �  P�  � �  X9!  � �  `l� � 	  h  � �  p �    �4  �  H
2�  �S  
4�   �  
5�  (  
6�  04  
7r  88  
8t  @ �  
:�  �  �
=�  R�  
?D   �  
@r  n  
Ar  �  
Br  1$  
C  2�  
E�  �� 
F�  `�L 
HU   � �  
J�  
  P   �  �  �  �    A  f  f  �   �  &�  �  �  A   �%  *�  �  �       �%  -    "     {  1.  4  �  C  o   �  4O  U  `  o   l  8l  r  �  �    $   �  <�  �  �  �    �   �  @�  �  �  �  o    r  7   �  G�  �  �    A  r  r  �   �'  N    �  2  A     �  S>  D  �  g  A  r  r  7  g   �  &  ��K  �� ��   i'  �~  H   �~  P  �~  X�A ��  `Y ��  h�#  ��  p�  �  x�  �"  �  �C  ���  ��  �U�  ��  ��!  �  ���  �2  ��  �`  �&  ��  � �&  �W  m  �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }]  �  U'�  �  m  D   t&   �  v~   A  w~  �  x~  &  y~   !  {�  �  �>   D   �  ]   �  r  ]    =	  �  �o   u   �   �  ]    �'  ��   �   �  �   �  r    �    &   �!  �   ��  )2    ��  )c   �  )�    }  �   	�   O  ;1!  _� =%1!   ݰ  >%�   !  �  @!  7!  �  �  	*  �    s!  @    �  �!  @     �  	�%�  !�`  s�  ��@            ��!  "k  s*U  U"�`  t*�  T !�_  h�  ��@            �"  "k  h3U  U"r� i3  T #SX  \��@     	       �a"  $Min \!a"  U$Max ]!a"  T" ^!o  Q J   �z  D  �  ��  $"  ��@     V�      ��  :G  �9   X  ^� �L   �i int �i {S @	�   g
  	�      	 	@   v  	#	@   �  	&	@   |
  	)	@    h  	,	@   (�  	-	@   0�	  	2S   8�  	5S   < �   �  	�   �
  	8"c   
  	K  �   
�  	L  
�  	M  S  .�  
�A  -  �[  
�T  �  >   
S   �	  
	Z   �  B"�  �     ��  R   �a    �� ��  �N ��  �6  �   �  Y�  �  a   �  u  9      n�      u  a    �  �  #  a   A  u  9   9   a    �  �"M  S  �   PJ�  2�  LP   �  ML   pos NL   �  P  SF  Q   �1 R   (=9 S]  0R�  Uu  8y�  VP  @�� WP  H �  �  �\ �9   m  �a    o  ��  �  �,  2  L   P  A  L   P  L    V  �  2  j  p  {  A   .|  YS    :9   �  J�  x L�   y M�   )  O�  	�  B   s  M   u�   }  u�  V  v�  /  v�   t
  x�  �J  Z   �`  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  Z    ��  Z   �  	S   B� 
P  L  T    V  s  V  v	  a     �  `  	�  �  (NT  �  PA   Z�  QA  �  ST  s  T�   [  UZ  ?1  WS     �  A    Y�  �  =  Z   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  �s  b   "�  �  �  %  <  x >A   len ?T  *� @V   %  B�  	    `,  2  L  S   S   L  a      �  q_  e  S   ~  S   S   a    �  �  �  �  S   S   a    �  `�3  �  �3   �% �9  ?1  �S   �&  �  !  �   I  �R  ()  �~  0R   �a   8�  �  @ �  ?  �  ��  	@  �   _  e  S   y  a   y   �  �  �  �  �  �   �  ?�  �  �  �  P  L    �  Y�  �  S   �  �  L   a    s  ��    S     �     M  W  0��  �  ��   e� �R  �� ��  �� ��  �� ��   �� �  ( �'  �  �!  lV  �  ��  	�  �  -  �V  	�  �  �L  �h  �  ��   	�  �
  �A  �  �T  �  �S   
  �Z   �  �9   \#  �L   Qd  A  )H  9   �   9   �  ,S   \&  7a   �0  D@   �H  Q-   Q}  b�	  x d.	   y e.	   r  g�	  b   � 
  xx �H	   xy �H	  yx �H	  yy �H	   a  ��	  	 
  z'  �=
  m  ��   ss  ��   �  �
    �W
  ]
  h
  a    �  ��
  �U  �a      �J
   %  �h
  �  $�
  �
  �   �
  �� "�
   �@ #�
  �U  $a    tT   �
  �
  �  7*  �; 9�
   ��  :�
   L  <�
  Z   %�z  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=�  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  Jz  
   s[  �  u�   ��  v�  �  x�  �
  z�  (  {�   �  }  �  �#u  {  k  `�*  R�  �u   (  ��  |  ��  �  ��  �  �
	  �  ��"  v  �*  �  ��  (�%  �*  07&  ��"  8G   ��  X �  �"7  =  h  v  �M �"   k  h  R�  u   �  �"�  �  %  8;�  �� =�"   �M >�     ?*   r$  @�  0 5  �$�  �  %  �T  �� �"   �M �"  �  �   �  �  (�� 
�  h�� �  p�� �  x K  � a  g  �  �,(  �   .	   �  /	  O  1	  C  2	  �  4	   d> 6�  (A  7�  0T  9�  8  :�  @�  <�  H�  =�  PE-  ?�
  X�!  D  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R(  ��� S�  �K1 Wv  �R�  Xu  �Jy  YA  �%  [*  ��	  ]�
  �    ^a   ��8  `  � L   5  ;    X��  �  �T   E-  ��
  N ��  �8  ��  P �  *%�  �  �  0t�  k  vh   �  wT  �@ x�  ݖ y
	  E-  z�
   N |�  0�  }H	  pR  ~H	  x�  �  �ߣ  ��  ��I ��  ��  ��  �h  ��  ��S  �`  �4  �
	  �8  ��  �  �a    �  �9   �  ��  o  ��  �L �a    �8  �  ( �
  L#�  �  W  H9  �  JT   = K�    L�  d  M�   �  Z   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  9  #   g)    �   ���  =  � 
   L  ��   $  ��  0�  �?!  8m  �#�"  h�  ��  pآ  �[  tG   ��  x �  [  �  �?  dg  �
  �)�  �  �   H�  �  �a    "  ��  �!  ��   ~	  8f�  �
  h�   (  i�  �� kH	  �� lH	    n�  �  o�   �  p�  (�  q�  0 y  s  �a  �;    �$�  �  �  0'  �N  )�   ?1  *�  }0  +�  i/  ,�  � - 
   �  �)       H�y  ��  ��   ?1  �
	  (  ��  4  � 
  \  ��  0  �a   @ +!  �  tag "	   �U  b	   �  y  �  `  Z   
�  w%   }#  �&  h  �  &     
�  E   9
Q  � ;
�   ��  <
	  �  =
	  �  >

	  �#  ?

	   �  L
(^  �  �  Z   ��  :   �   ^$  1  �!  �!   :  �d  �  �b	  �#  ��  �  U	  �  *   I$  ��  �  �  *   �&  ��    �    *     �   �!  H��  �  �"	   S"  �	     ��  �"  �H	  �  �H	   ;  �9  (%  ��  0�   ��  8��  ��  @ �  R  �  x  =W
  T  Z   ��  �L   3A  �<   �.  ��  H  E#  	�  �  @J{  �  L	   �  M�  �� O�  .� P�  �  Qm   �  R  (�!  SE  08'  T�  8   W!�  �  -  (l�  k  nh   �M o�  ߣ  p�  �  q�      k  )�  �  U	  �  {  �   w   .      {   �  1$  *  ?  {  ?  m   
  K  6Q  W  g  {  g     �  :y    U	  �  {  {   �  >�  "  Y�  �  U	  �  �  �  �  m   �  _�  �  U	  �  �  �  ?  m   $  f    &  �  �  g   �  l2  8  U	  Q  �  "	  b	   #  x��  �� � �   �  � �  H  � �  P�  � �  X9!  � �  `l� � &  h  � �  p �    �Q  �  H2  �S  4`   �  5T  (  6T  04  7
	  88  8�  @ �  :�  �(  :3  �  �  �=�  R�  ?u   �  @
	  n  A
	  �  B
	  1$  C�  2�  E  �� F  `�L Ha   � �  J�  9  P   �  �  U	  �  A  T  �  �  �   �  &      T   �%  *  %  U	  4  (   �%  -@  F  Q  (   {  1]  c  U	  r  �   �  4~  �  �  �   l  8�  �  U	  �  (  Q   �  <�  �  U	  �  (  "	   �  @�  �  U	    �  (  
	  [   �  G    U	  ;  T  
	  
	  T   �'  NG  M  U	  a  T  A   �  Sm  s  U	  �  T  
	  
	  [  �   H	  &  ��z   �� ��   i'  �	  H   �	  P  �	  X�A ��  `Y ��  h�#  �  p�  �4  x�  �Q  �  �r  ���  ��  �U�  �  ��!  �;  ���  �a  ��  ��  �&  ��  �   ��  	z   �&  ��   �  a   �>  ��   'O  �   xC  �9   s/  ��   	�   �  0t?!  �  vb	   a   wb	  �'  xb	  !  yb	  �#  zb	   �  {b	  ( �  }�   �  U'X!  ^!  m  D   t�!  �  v	   A  w	  �  x	  &  y	   !  {c!  �  ��!  �!  U	  �!  L!  
	  �!   =
  �  ��!  �!  "  L!  �!   �'  �"  "  U	  4"  L!  
	  �  4"   �!  �!  s"  ��  )�!   ��  )�!  �  )"   }  :"  	s"  O  ;�"  _� =%�"   ݰ  >%L!   �"  �  @�"  �"  �  �  =  �  -1  B�  *  �"  L    �  #  L     �  �%�  �(  Z   9�#  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  V�#  �\ X�   �  Y�  x  Z�   �7  \�#  	�#  �6  `S�$  �<  UH	   �Q  VH	  a(  X	  VA  Y	  Q) [�   nX  \�  "�D  ^�$  (�5  _�$  8M   a�  H}  b�  JV  c�  L/  d�  N7K  f�  P>D  g�  R�:  i�  T�3  j�  V=]  k�  X 	  �$  L    �5  m�#  �Q  8��%  �  �H	   �Z  ��  %?  ��  
L/  ��  �<  ��  �Y  ��  �7  ��  �)  ��  �O  ��  �H  ��  vH  ��  ^  ��%  �>  ��  $�7  ��  &0>  �a   (�+  �a   0 �  �%  L    �H  ��$  �?  8A�&  �  CH	   �Z  D�  %?  E�  
L/  F�  S.  H�  �W  J�  �W  K�  C  L�  �O  M�  �H  N�  vH  O�  ^  Q�%  �>  S�  $�B  T�  &0>  Za   (�+  [a   0 �]  ]�%  �B  �|)  ��  ~�   �)  �  �)  ��  �.  ��  U  ��  �V  ��  
�0  ��  �6  ��  �C  ��  U?  ��  6P  ��  �C  ��  &L  ��  *J  ��  �L  ��  HP  ��  N*  �)   [2  �"	  0k2  �"	  8.  �"	  @{2  �"	  HQ2  �)  P�0  ��  Tp4  ��  VmU  ��  X�Z  ��  Z ?  ��  \:  ��  ^�I  ��  `E8  ��  b�;  �"	  h�;  �"	  p�O  ��  xDF  ��  zfV  ��  |�9  ��  ~[9  ��  ��G  ��  �zQ  ��  � �  )  L   	 �  /)  L    {D  ��&  �1  @��)  �I  �H	   6Y  �H	  �^  ��  S  ��  )  �"	  @3  �"	   �0  �"	  (4C  �"	  0�C  �"	  8 aM  �<)  �I  @��*  �  �H	   _7  �"	  )  ��  �O  ��  �n ��  �T  ��  EF  ��  I  ��  �K  ��*  N:  ��*  ,L  ��*  4�E  ��  :�Z  ��  ;�Z  ��  <^  ��  = �  �*  L    �  �*  L    �  �*  L    eU  ��)  �9  (7�+  ��  9H	   a@  :�  b<  ;�  
8  <�  .  =�  �H  >�  �Q  ?�  X  @�  �.  A�  �;  B�  ))  C�  eH  D�  I_  E�  �B  F�   !3  G�  " �)  I�*  	  �  I,  F@ K�   I�  L	  K�  M	   ԃ  O�+  �b  hh^,  `h  j
	   m�  k
	  dh  l^,   ,  n,  L    ��  n),  �j  0��,  F@ ��   I�  �H	  def �H	  K�  �H	  tag �"	   c  �
	  ( )�  �z,  �  �-  �  ��   c  �
	  Cg  �
	   �~  ��,  z�   �r-  `h  �
	   m�  �
	  L�  �
	  dh  �r-  e  �x-   �,  -  J�  �#-  �R   F�-  tag H"	   ��  IH	  .� J	  �P  K�-   "	  DG  M�-  f3   � .  Tag �"	   Q  �"	  .*  �"	  �K  �"	   gW  �,.  �-  �^   �.  k@  �   aE  �  p0  �  �>  �  H  �  �/  "	  �� �.   �  �F  2.  �<  0�.  H  2�   �/  3"	  �� 8�.   qS  :�.  A9  0Um/  ߣ  W�   �E  X
	  �^  Y
	  =Y Zm/  <  [
	  �=  \s/   Jy  ]A  ( �.  �.  rY  _�.  �1  ~�/  �.  ��   �L  ��   Z  ��/  �/  �V  ��/  ��  ��   f>  ��  Y  ��/   �)  ��/  ��  ��0  �  ��   ��  ��  ~  ��  �  ��  �  ��  5  ��  
B  ��  �  ��   �w  �
0  �A  /?1    1�   �  2�  �N  3�  o=  4�  D4  5�  �^  6�  `*  7�  �0  8�  �G  9�  �D  :�  	I:  ;?1  
 �  O1  L    �@  =�0  �  �\  ��1  +  �O1   Y�  �O1  �
  ��  (  ��  �F  ��  �C  ��   <)  ��1  b1  �,  2  �  �   AK  �  z8  \1  V 2   %2  �  �R  �1  	F  .c2  �  0�   �P  1%2   ">  382  !I�2  "�K K+2  "`B Lc2   �[   E�2  �z  G�   =Y Np2   �6  P�2  O]  a!�2  �2  �(  �-#4  `h  /
	   �  0�  �  1�  6~  3G  ;�  4o	   �~  6�  (��  9�  0ux  :�O  8˄  <�  @��  =�  Al  >U	  D܀  ?�Q  H�  A�  Phx  B�  Q3p  CU	  Tk  D�Q  X�}  F!R  `��  H
	  h�t  I�  pte  K
	  xl  L�-  �(�  N"	  � 7N  (��4  >) ��.   -N  ��.  V` ��.  TE  �"	  �/  �
	   �z  ��  $ G  �#4  &8  � �4  �4  eS  po�8  �� q�   ^  s�-  ��^  u"	  [>  v�   �W  w .  (� y�$  0�=  z�%  ��,  |�+  ���  ~�  ��(  �&  �AK  ��  0XL  �y/  8#os2 �/)  hp�  ��)  �T  ��.  0#9  �"	  8!H ��:  @�+  �;  H@.  �d;  P�E  �B;  X�P  �B;  `@  �B;  h$S  �a   ps  �a   x#mm �a   �#var �a   �Q  �a   �<B ��/  �2Y ��*  �=  �"	  �=  ��1  �UV  ��2  ��(  �"	  =  ��.   /:  �"	  (�?  ��.  0�]  �"	  8#cvt ��;  @�R  ��8  H5$  ��
  P��  �  `HT  �"	  h�*  �"	  p�J  ��  x�+  ��  y�  ��2  ��C  �h  ��-  �  �j7  �
	  �kN  �"	  ��F  �"	  �#7  �"	  ��(  ��.  �rE  ��.  �QZ  �"	  �4  �
	  ��@  �"	  �:L  ��.  ��G  ��.  ��]  �"	  ��W  ��;  ��/  �
	  ��B   �;   �I  �.  s-  "	  �*  
	  ,  h  ,  h   #bdf 	�4  (�T  "	  P#F  "	  X�U  "	  `�K  "	  h �=  �9  9  U	  9  a    �Q  �")9  /9  �\  xc�:  �  e�4   �  f�@  )�  g�  �V  h�  :1  j"	   �^ k
	  (Jy  mA  0�  n�  8�  p�  <�!  q  @R0  r�  `�  s�  duN t�  h6  u�  lpp1 v�  ppp2 w�  �2�  zv<  �Xc  {v<  ��6  }�<  )  ~�.  �8  "	   �L �a   (C  ��  0��  ��  4#pp3 ��  8#pp4 ��  Hy�  ��.  X�� ��.  `U  �*  h �I  ��:  �:  U	  ;  �4  "	  A  �-    1  ;  $;  U	  B;  9  
	  "	  
	   �M  +O;  U;  U	  d;  9   �<  :q;  w;  �;  9   y*  Z   =�;  4   �^  J  b8  �T   lK  H�;  �  
	  |T  @?v<  R�  Au   �  B�  n  C�  
Z�  D�  �  E�  org GT  cur HT  ��  IT   s  K�.  ([  L\1  0c+  N�  8 R8  P�;  �  P�<  �;  RG  T'�<  �<  $[  P��@  �  ��4   �  ��@  R�  �u  � �U	  top �	   �m  �	  (4� ��+  0��  �	  8�l  �	  @zp0 �v<  Hzp1 �v<  �zp2 �v<  �%pts �v<  &�~  �v<  H&�  �	  �&N ��  �&�  ��M  �%GS �EL  &B�  ��  x&� ��.  �%IP �	  �&-d  �	  �&6f  ��  �&ss  ��  �&*o  ��  �&T�  �"	  �%cvt ��+  �&�k  �
	  �&�w  ��.  �&}w  �
	  �&1�  �
	  �&�w  �FM  �&vt  �
	  �&�  �
	  �&yt  �FM  �&�{  �
	  �&�  �
	  �&7�  ��  �&by  ��  �&qq  �CO  �&b<  ��   &8  ��  &�a  ��L  &��  ��  8&�^ ��+  @&/y  �;	  H& t  �;	  P&A�  �;	  X&�r  ��  `&Br  �EL  h&aa  ��  �&Qy  ��  �&f  �	  �&|o  ��M  �&Mr  �VN  �&�z  �VN  �&_�  �VN  �&�  �*N  �&  �*N   &�t  ��N  &t  ��N  &Yg  ��N  &y  ��N   &�g  ��  (�m  q�  )Ho  v�  *h�  {�  +�e  �  ,�f  ��  -y�  ��  .x�  �"	  0�l  �"	  8�x  �"	  @6v  �"	  H O  _ �@  �@  LL   BB  �� �   N �C  X��  �  `��  �M  �-U "	  �� "	  ��s  $
	  ��s  %
	  ��s  &FM   5�  (
	  �}  )
	  9�  *FM  ��  ,
	  �v  -
	  �a  /�L   #GS 1EL  P�]  3"	  �#cvt 4�+  ��c  6�  ��^ 7�+  ��~  9v<  �-�  ;�<  G�  ?U	  $|  @U	   }  �/9  Y�  E[B  aB  U	  �B  A  �4  �  �  �   ��  k[B  �y  ��B  �B  �B  �4   �m  ��B  �B  U	  �B  �4  "	  	  �.  �-   t�  "�B  �B  U	  "C  �4  "	  
	  
	  A  "C  (C   �  �0  ن  @;C  AC  U	  ZC  �4  Q  �-   �}  ZgC  mC  U	  �C  �4  "	  �C   �  kp  s�C  �C  U	  �C  �4  
	  �C   �  T�  ��C  �C  U	  �C  �4  A  �   �m  ��C  �C  D  �4  �  
	  �;  \1   1z  �)D  /D  U	  HD  �4  �  �C   �a  �UD  [D  �  yD  �4  �  yD  yD   �  sz  ��D  �D  U	  �D  �4  A   �w  �B  �m  !�D  �D  �  �D  �4  
	  
	   3b  �2�F  !H 4"�:   �A 6"OB  �M 7"�B  Y 8"�B  ��  9"�   K ;"�B  (�; ?"D  0|G @"�C  8H A"D  @"I B"D  H�Y C"D  P�Z D"D  X�S F"D  `�< G"�D  h�9 J"D  p7B L"D  x-Y M"D  �(K Q"D  �Z S"�B  ��i  V"�C  �s  W"�D  �U�  \"�D  ��@ b"D  �x> c"�C  ��j  e"D  ��w  f"�D  ��V h".C  ��= i"ZC  ��D k"�C  �tW m"D  ��9 n"HD  � ��  p�D  ~c  t�F  �F  ��  '�F  �F  U	  �F  T  �F   n,  jd  +�F  �F  U	  G  T  G   G  ~-  �g  /*G  0G  U	  IG  T  
	  �+   �{  6UG  [G  U	  tG  T  
	  �    l  =*G  �n  BUG  �x  G�G  �G  U	  �G  T  
	   1j  K*G  �}  P�G  �G  U	  �G  T  �;  �G  �G  G   �  ��  W  ��  ZH  	H  �b  PZ�H  h  \�F   �v  ]G  ��  ^tG  ��  _�G  .�  `�F   �  aIG  (V�  b�G  0��  c�G  88�  f�G  @��  g�G  H i   '�H  �H  U	  �H  T  
	  yD   4�   ,�H  \�   1�H  �l   8�H  ~�   =�H  ŋ   B�H  �w   G�H  H�   N  �r   Q6I  	%I  ȅ  @ Q�I  ��   S�H   ��   T�H  �n   U�H  Rs   W�H  ��   X�H   F}   YI  (�|   ZI  0��   \I  8 5l  !'�I  	�I  BY  !'�I  /  !)�    �  " �I  �I  "	  J  T  
	  �-   ��  "$J  	J  Y�  "$/J  �{  "&�I    n)  #;J  AJ  U	  _J  *    9  �   �)  #$kJ  qJ  U	  �J  *    a    nk  #)�J  	�J  �;  #)�J  �=  #+/J   z+ #,_J   
�'  $�   �z  '"�J  �J  ��  �KK  �� M�"   Xc  Ov<  8Nz  Q
	  x Zo  6�  xj  `AEL  rp0 C�   rp1 D�  rp2 E�  |a  G�	  hc  H�	  
Ό  I�	  D�  K	  +{  L;	   �l  M�  (ׄ  O�  ,g  P;	  0.�  Q;	  8zs  R;	  @,�  S�  Hō  T�  J1h  V�  L�i  [�  MT�  \�  P�{  ^�  T�{  _�  V{�  `�  X �|  b&K  	EL  �k  Z   ��L  �   �b  o  ��   fe  ��L  2�  ��.   �  �	   ��  ��L  �k  ��L  �L  �L  L    ]p  (�:M  �a  ��   �S �	  end �	  opc �
	  �  ��  $a  ��  �w  �"	    �s  ��L  �r  �RM  �L  bz  P��M  �  �	   �d  �	  :� �  B� 	  �� H	   �c  �M  (pw  �  H=f  	�  I4�  
�  J ;	  �M  L    �u  XM  y  5N  N  ;	  *N  �<  ;	  ;	   ^�  ;6N  <N  VN  �<  �<  �  ;	   �c  BbN  hN  ;	  �N  �<  �  �   �  H�N  �N  	  �N  �<   G  L�N  �N  ;	  �N  �<  "	   z�  R�N  �N  �N  �<  "	  ;	   }d   [1O  t  ]�   �d  ^	  ��  _	  Def a1O   :M  sc  c�N  !�  cOO  �N   x  �"QL  Le  )�O  A�  +H	   ��  ,H	   -�  .!�O  bO  �  :�O  �|  <�   �t  =�O   J�  ?�O  �O  �  BP  �  D
	   Kw  E
	  7�  F�;  ~  H�;   k�  K$P  �O  ��  O_P  ��  QH	   �  RH	  �w  SH	   r  UkP  *P  Bh  X�P  �{  Z_P    �t  \�P  qP  �e   `�P  ��  b
	   k  cP  �q  e�   q  f
	  y|  g�P   u�  i�P    iQ  �P  -m  l@Q  U{  n
	   �n  o�;  ]c  p�;   -r  rQ  �e  rXQ  Q  �a  8}�Q  �{  �P   �  �@Q    '�  ��Q  ^Q  ߐ  ��Q  tag �"	   �n  ��  ]c  ��  
�  ��   k�  ��Q  �Q  o{  0�!R  |  ��   �{  ��P  �D ��Q  ( {�  �-R  �Q  �  Z   [\R  'w   �'�b   p'em  � �z  Z   m�R  '�   �'h   @'Hk    'c   'ֈ  � Z   %��T  |m   �  ��  j  zn  �r  ��  �q  �`  �h  	�  
�p  э   �  ��  �j  �y  ˑ  ��  �y  !g  ˉ   ai  !k  "�f  #߃  $It  %�t  &��  '��  (�p  0��  1�j  @�  A,}  Qς  R�p  S�f  T�a  UN�  V�  W��  X-n  `\�  a_b  b[|  c�  p�v  �I�  ��v  ���  ��u  ���  �Ha  ��  ��u  ��  �p  �7q  ��b  ���  �o  �Cb  ��g  ��c  ��q  �Yf  ���  ��d  ��`  ��  ��z  ��y  �)�  �&t  ��m  �m  �a  �	q  �d  �G�  �
d  ��v  ��a  �2�  ��g  �W  �J�  ��o  �`u  �%u  �v  ��o  � y  � (�c  ��J  	PBH     )�k  �H  	 BH     )�|  �1I  	�AH     )d�  .�I  	�AH     )��  J  	�AH     �   XU  L    	HU  )�v  #XU  	@AH     *�J  q	�@H     ��  (n�U  ��  p	   �q  q�  k�  r�  
�{  s"	  :s  t�  ?1  u�  C�  v"	    'w  x�U   �  egV  ��  g	   C�  h�  �q  i�  
vb  j�  {q  k�  �f  l�   Fp  nV  ��  (q�V  p  s"	   ,�  tH	  Nx  uH	  �  vH	  ?1  w�   �>  x�  " ��  ztV  +UO  7	 @H     �  W  L   � 	�V  )��  {W  	 ?H     �  3W  L   � 	#W  )ls  �3W  	 >H     E�   s�W  {  uT   �j  vT  ��  wT  �  x
	   v�  zOW  �k  z�W  OW  >x  �W  Q  "	   �K  "	   �|  
�W  	�W  ,Ǝ  k�.  `X  -�  k(�4  -:� l(
	  -n�  m(
	  .nn o
	  /E  p�.  /�@  q"	  /�� r�.   0�j  Z�X  -�  Z�4  /Jy  \A  /R�  ]u   ,Oi  
U	  :Y  -�  
!�4  -Jy  !A  /� U	  /R�  u  .nn 
	  /ȃ  
	  /x-  "	  /�@  "	  .p �.  /�� �.  1�u  O1�0  R ,�e  �U	  �Y  -�  �!�4  -Jy  �!A  /� �U	  />k  �"	  1�u  � ,^n  �U	  �Y  -�  �!�4  -Jy  �!A  /� �U	  />k  �"	  1�u  � 2��  >U	  �	A     �       �g[  3�  > �4  &� � 3Jy  ? A  �� �� 4� CU	  � � 4R�  Du  @� <� )>k  E"	  �H5�u  o�
A     6x
A     -       �Z  7cur _�;  |� v� 4�� `�;  ɯ ǯ 8�
A     �x 9U|   :�	A     �Z  9Us 9T tvc9Q| 9R�H ;N
A     �x [  9Uv 9T29Q09X09Y�D ;p
A     �x 4[  9U|  ;�
A     �x L[  9U|  8�
A     H�  9Us 9T|   0i  !�[  -�  !�4  /Jy  #A   <�{  �"	  ��@     �       �1\  =�  �#�4  U>n�  �#
	  �� � =�Y  �#�;  Q?�} �"	  �� z� ?�} �"	  � � @p ��.   � � ?3o  ��.  �� ��  A1a  >U	  �\  B�  >!�4  BJy  ?!A  C� AU	  C>k  B"	  C�� C�  D�u  �EC5�  �"	  C� � .  C�� � .  Fpos �	  C��  �	  C;�  ��  EC-�  �	     2m�  �U	  A            �%]  3 ��  ?� ;� GA     �x  H'f  s��@            �T]  I�  s*  U 2r  NU	  ��@     
       ��]  I�  N*  U4K1 S�J  z� x�  2na  �U	  ��@     )      ��_  3�  ��@  �� �� 3D|  ��  � � 4�  ��4  �� �� 44  ��C  ۴ մ J�_ �@      �@     #        �^  K�_ 1� -� K�_ m� k� L�@     #       M�_ �� �� M�_ � ޵   J�_ D�@      D�@            !�^  K�_ � � K�_ F� D� LD�@            M�_ x� t� M�_ �� ��   N�_ r�@      U  E_  K�_ �� �� K�_ !� � OU  M�_ n� j� M�_ �� ��   N�_ ��@      @U  #�_  K�_ � � K�_ � � O@U  M�_ G� C� M�_ �� ��   P��@     �x PH�@     �x Pq�@     �x P��@     �x  Hy�  �P�@            �.`  3�k  �(  ˸ Ÿ 4�  ��@  � � 8Y�@     �a  9Us   2�d  �U	  `�@     !       ��`  I�k  �(  U4�  ��@  k� i� Q� �U	    ,n  cU	  �`  -�  c$�@  -�  d$�  /� fU	  1�u  �E.i t
	  /�  u�4    ,n�  �U	  �a  -'�  �#(  -�  �#�  /� �U	  /�  ��@  /�  ��4  /R�  �u  /�~  �  /'I �a  1�u  ZRwa  /�  "�a   E/k  Fh    �+  �M  H�  �`�@     �       ��b  3'�  �#(  �� �� 4�  ��@  � � 4�  ��4  4� 2� 4R�  �u  Z� X� P��@     @�  ;��@     �x +b  9Uv  ;��@     �x Cb  9Uv  ;��@     �r  \b  9Us� ;��@     �x tb  9Uv  8�@     �x 9Uv   2�o  �U	   �@     �      ��d  3�  ��@  �� }� 3�  ��  �� �� 4�  ��4  :� 6� 4�6  ��<  t� p� 4� �U	  �� �� J
�  ��@      ��@            �qc  K;�  � � K/�  � 	� K#�  0� .� K�  V� T�  J��  ��@      ��@            ��c  K��  {� y� K��  �� ��  N�  ��@      0X  ��c  K�  Ƽ ļ K�  � � O0X  M)�  � �   NH�  ��@      �X  �Rd  Km�  b� `� Ka�  �� �� KU�  �� �� O�X  Mx�  ӽ ѽ   ;H�@     5�  vd  9Us 9T| 9Qv  S��@     9Us   ,�c  )U	  �d  -�  )�@  -�  *�  /�  ,�4  /�6  -�<  /� .U	  E/4  D�C  /�  E�a    T�  � A           ��f  3e5  �T  � �� 4�  ��4  h� `� 4R�  �u  ɾ Ǿ 4Jy  �A  � � 4$S  ��F  � � Ng[  mA      �Z  ��e  Ku[  8� 6� O�Z  M�[  ]� [� 8�A     �x 9Ts�	   N`X  �A      �Z  �Af  KnX  �� �� O�Z  M{X  �� �� M�X  ο ̿ P�A     �x 8�A     �x 9U| 9Ts�	   :mA     Uf  9Us  ;�A     �x mf  9U}  ;�A     �x �f  9Uv 9Ts� ; A     �x �f  9Uv 9Ts� 8A     ��  9Us   2|  BU	  �lA     �
      �Vp  3Jy  B A  �� � 3e5  C T  �� o� 3�  D �  L� H� 3G  E �  �� �� 3G  F �  o� ]� 4� HU	  l� 6� 4k  Ih  �� �� 4$S  J�F  �� �� 4�  K�4  f� T� 1�u  �1�  �U�q  �g  4� �
	  5� -� ;�tA     ��  �g  9Us  8�tA     P 9Us   N�p  �mA      `o  �
j  K q  �� �� VFr  �mA     ,       �
yh  WWr  L�mA     ,       Xyr  8nA     y 9U| 9T~    Yq  0nA      �o  �
K q  @� 6� Op  MDq  �� �� ZQq  ��~M^q  W� I� Mkq  � �� Mxq  �� �� M�q  M� ?� M�q  �� �� M�q  � � Y�q  qA      `p  �K�q  ;� 7� K�q  {� u� N�q  >qA       �p   j  Kr  �� �� Kr  s� m� O�p  M#r  �� �� M/r  � �� M;r  h� `� ;SqA     �x �i  9U��~9T}  ;�qA     y �i  9U}  ;�qA     %y �i  9U��~ 8�qA     �x 9U��~   S#qA     9Us 9R0     N�X  �oA      �p  ��k  W�X  K�X  �� �� O�p  Z�X  ��~M�X  3� +� M�X  �� �� M�X  �� �� Z�X  ��~MY  �� {� MY  �� �� MY  �� �� ['Y  RsA     [0Y  �sA     :�oA     �j  9Us 9Txmdh9Q 9R��~ ;BrA     2y k  9U 9Q}  ;�rA     �x Kk  9U| 9T19Q09R	��~�
��9X09Y��~ ;�sA     �x kk  9U��~9T}  8uA     �x 9U| 9T19Q09R09X09Y��~   N�Y  1pA      @q  �=l  W�Y  K�Y  � � O@q  M�Y  Z� R� Z�Y  ��~[�Y  �tA     :IpA     l  9Us 9Tmgpf9Q��~9R��~ 8�tA     2y 9U��~9Qs�   N:Y  gpA     	 pq  ��l  WYY  KLY  �� �� Opq  MfY  �� �� ZsY  ��~[�Y  <uA     :pA     �l  9Us 9Tperp9Q��~9R��~ 8:uA     2y 9U��~9Qs�   \Vp  �q  ��m  Whp  O�q  Mup  X� V� X�p  Z�p  ��~M�p  �� |� M�p  �� �� M�p  =� 1� ]�p  wA     D       �m  M�p  �� �� Z�p  ��~;2wA     ?y �m  9Us 9T} 9Q��~9R8 8TwA     Ly 9U��~9T	�1H       8�uA     �[  9Uu 9T~ 9Qq    J&Q �pA      �pA     ?       �n  K4Q �� ��  N1\  �sA      r  ��o  WN\  KB\  � � Or  MZ\  ~� r� Zf\  ��~Mr\  �  � [~\  stA     ^�\  pr  o  M�\  �� �� M�\  �� �� M�\  � � M�\  Y� U� M�\  �� �� M�\  �� �� ]�\  �vA     "       �n  M�\  5� 3�  8�vA     Wy 9U��~  :�sA     7o  9Us 9Tfylg9Q��~9Rs� :tA     do  9Us 9Tacol9Q��~9R��~ ;itA     2y �o  9U��~9Qs�	 8�vA     Wy 9U��~   ;mA     dy �o  9T	�1H      ;,mA     qy �o  9U~ 9T0 :JmA     p  9U~ 9Ts 9Q��~�9R| 9X}  :�mA     9p  9U��~9Ts 9Q��~�9R| 9X}  8#pA     �Y  9Us 9T��~  ,N�  ��  �p  -e5  �$T  /E  ��  /�  ��4  /�Y  �
	  .i �"	  /�^  "	  /.� 
	  E/� U	  .buf �p    �   �p  L    ,�~  ��  q  -�  �!T   ,hg  �  �q  -�  *�4  )�a  !�q  	`7H     /�z  �"	  /�z  ��q  /�r  ��  /�n  ��  /ߊ  �#�  .i ��  .j �S   .k �S    �W  �q  L   L    	�q  S   �q  L    A��  �"	  �q  B�  �$�4  _i �$�   A�z  �h  Fr  BJy  �&A  Bss  �&"	  C� �U	  C�z  �h  Fi �
	   Arv  ��  �r  BF@ �+�  (+�  ��r  	@<H     Fnn �
S    �   �r  L   L    	�r  A�s  pU	  �r  BR�  p#u  Bb<  q#�  B8  r#�  BXc  s#�<  C� uU	   `2�  F��@     �       ��s  >Xc  F$�<  ^� X� ?R�  Hu  �� �� ;��@     �x Ls  9Uv  ;�@     �x ds  9Uv  ;�@     �x |s  9Uv  ;)�@     �x �s  9Uv  8=�@     �x 9Uv   a�j  �U	  pyA     :0      ��  bexc ��<  � �� 4�  �"	  � � 4��  �"	  �� �� 7i ��  �� �� 5�l  .!�A     5o�  1!�A     5��  !	|A     5s  (!~A     U�s  �  4��  ��+  e� !� 46f  ��  � L� Nu�  ��A      0u  L Pu  K��  Z� X� K��  �� }� O0u  M��  �� �� M��  M� E� M��  �� �� M��  � �� M˧  s� i� M֧  �� �� [�  ��A     :�A     >u  9U  SȚA     9U    N��  �{A      �u  B�u  K��  � � K��  X� T� O�u  M��  �� ��   N��  ڛA      �u  ��w  K��  �� �� K��  J� B� O�u  M��  �� �� M��  � � M̼  �� �� ^��  @v  kw  M��  �� �� M�  �� �� ]�  ��A     Z       �v  X�  N�_ ��A      pv  �v  K�_ Q� O� K�_ |� t� Opv  M�_ �� �� M�_ =� 9�   N�_ ߧA       w  �v  W�_ W�_ O w  M�_ |� x� M�_ �� ��   S�A     9U   J�_ ]�A      ]�A            
Zw  K�_ �� �� K�_ #� !� L]�A            M�_ J� F� M�_ �� ��   S]�A     9U   ]׼  k�A     <       �w  Mܼ  �� �� M�  �� �� S��A     9U   S8�A     9U    J��  g|A       g|A     	       "x  K��  � � K��  9� 7�  N�  E�A      pw  � fx  K�  b� \� K��  �� �� Opw  M�  �� �� M�  Z� T� M(�  �� ��   N�  TA      �w  {@y  K+�  *� $� K�  y� s� O�w  Z8�  ��ZD�  ��~ZQ�  ��~Z]�  ��~Mi�  �� �� Mv�  � �� ;�A     ̸  y  9U 9T��~9Q��~9R��9X��~ 8V�A     ~�  9Uu 9Ty 9Qq 9Rr 9Xx    J��  �A      �A            \ �y  K�  e� c� K�  �� �� 8�A     J�  9Uu 9Tt   J��  �A      �A     #       ��y  K��  �� ��  Nڱ  �A      �w  �|  K��  �� �� K�  �� �� O�w  M�  3� 1� M�  Y� W� M�  � }� M'�  �� �� M3�  �� �� M?�  � � ML�  ]� S� MY�  �� �� Me�  � � Mq�  �� ~� M~�  �� �� M��  �� �� M��  %� � M��  �� �� X��  ;��A     ~y �z  9U��~9T��~9Q@ ;�A     ~y {  9U��~9T��}9Q@ ;*�A     ~y >{  9U��~9T��}9Q@ ;I�A     ~y i{  9U��~9T��~| 9Q@ ;ըA     ~y �{  9U	��~��~9T��~9Q@ ;�A     ~y �{  9U| ��~9T��}9Q@ ;	�A     ~y �{  9U| 9T��~9Qv  8�A     ~y 9U| 9T��~9Qv    J4�  �A      �A            �T|  KB�  �� �� 8&�A     �  9Uu   JN�  7�A       7�A     !       ��|  K\�  �� �� K\�  �� �� Ki�  �� ��  Jw�  `�A       `�A     !       ��|  K��  � � K��  � � K��  <� :�  J/�  ��A      ��A     1       *�}  K=�  a� _� K=�  a� _� KJ�  �� �� c�_ ��A      ��A     "       �"K�_ �� �� K�_ �� �� L��A     "       M�_ �� �� M�_ =� 9�    JX�  ��A       ��A            &�}  Kf�  z� x� Ks�  �� ��  J��  ƂA       ƂA            >/~  K�  �� �� K�  �� ��  J�  ۂA      ۂA     !       :�~  K,�  � � LۂA     !       M9�  5� 1�   JE�  ��A      ��A            6�~  KS�  n� l�  Jk�  �A      �A            .�~  Ky�  �� ��  J��  $�A      $�A     S       �[  K��  �� �� L$�A     S       M��  �� �� M��  �  � M��  '� %�   J��  w�A      w�A     3       �R�  K��  N� L� K��  s� q� Lw�A     3       M��  �� �� M��  �� �� M��      Y��  �A       x  DK�  Z  T  K�  Z  T  K��  �  �  K��  �  �  O x  X�  8��A     �v 9Q�9R�d�  �     J��  ��A      ��A     =       �I�  K�  / - K��  T R L��A     =       M�  { w M�  � � M(�  � � Y��  ��A      Px  )K�  ; 5 K�  ; 5 K��  � � K��  � � OPx  X�  8ԃA     �v 9Q�9R�d�  �     JP�  �A      �A     $       ���  Kk�    K^�  5 3 8��A     ��  9U 9R�  Jy�  �A      �A     >       ��  K��  Z X K��   } ;"�A     ��  �  9U 9R� 8@�A     �  9U   J��  I�A      I�A     5       �|�  K��  � � K��  � � LI�A     5       M��  � �   JR�  ~�A      ~�A     5       �݂  Km�  ) ' K`�  N L L~�A     5       Mz�  s q   J�  ȄA       ȄA     u       g��  K4�  � � K'�  � � LȄA     u       MA�    MN�  - ) M[�  e c :��A     j�  9U  :�A     ��  9U 9Ts  S$�A     9U 9T� 9Qv 
��   N��  =�A      �x  be�  K��  � � O�x  M��  � � cD�  ~�A       ~�A     !       �Kp�  � � Kc�  � � KV�  � � L~�A     !       X}�  8��A     �c 9U 9Tt 9Qq      N��  ��A      �x  ^܄  K��    K��  _ W O�x  M��  � � M��   
 M��  _ Y 8F�A     ��  9Uu    N�  x�A       y  Zх  K6�  � � K)�  	 	 O y  MC�  x	 p	 MN�  �	 �	 M[�  P
 B
 [h�  x�A     ^q�  Py  e�  Mr�     YD�  1�A      �y  KKp�  O I Kc�  � � KV�  � � O�y  X}�  8I�A     �c 9U 9Tt 9Qq      J��  ^�A       ^�A     9       R?�  K�    K�  5 3 L^�A     9       M!�  Z X M.�  � }   JG�  ��A      ��A            ���  KU�  � � KU�  � �  N��  ��A      �y  ��  K̲  � � O�y  Mٲ    M�  A = e�  :i�A     �  9U  S�A     9U 9Ts 9Qv 
��   Ni�  ��A      �y  ���  K��  ~ z Kw�  � � O�y  M��  � � M��  @ > :�A     k�  9U  :�A     ��  9U 9T�9Q|  S٥A     9U 9T�9Q|    N��  g�A      z  ��  KǶ  g c K��  � � Oz  MԶ  � � M�    M�  Q K M��  � � e�  ;��A     =�  6�  9Uy  ;ˉA     =�  N�  9Uy  ;��A     ~�  x�  9Uu 9Qq 9Rr 9Xx  8/�A     ~�  9Uu 9Qq 9Rr 9Xx    N��  ��A       @z  v��  K��  � � K��    O@z  Z��  ��Z��  ��~Z÷  ��~ZϷ  ��~M۷  L H X�  M��  � � M�  � � M�  � � ;��A     ̸  k�  9U 9T��~9Q��~9R��9X��~ 8i�A     ~�  9Uu 9Ty 9Qq 9Rr 9Xx    J��  ��A       ��A            ۉ  K��  ^ \ Kſ  � �  J�  ��A      ��A            �  K��  � � K��  � �  Jc�  ��A      ��A            _�  Kq�  � � Kq�  � �  J-�  ܋A       ܋A            
��  K;�  � � K;�  � � KH�     NC�  ��A       �z  �  K^�  > : KQ�  x t  Nl�  ��A       �z  �  K��  � � Kz�  � �  N��  �A       �z  �P�  K��  & " K��  ` \  N��  x�A       {  ���  Kٻ  � � K̻  � �  N��  ΍A      @{  V{�  K��   
 K��  v n O@{  M��  � � M��  = 7 M��  � � [�  x�A     ^�  �{  �  M�  u q  YD�  ��A      �{  �Kp�  � � Kc�    � KV�  : 6 O�{  X}�  8��A     �c 9U 9Tt 9Qq      V}�  �A     ;       ь  W��  L�A     ;       M��  v p 8	�A     ��  9Uu    N3�  #�A      �{  �'�  KN�  � � KA�   � O�{  M[�  > 8 Mf�  � �   N��  ��A       |  �J�  K��  � � K��  ` X O |  Mε  � � M۵    M�  � � M��  � � M�  / % [�  W�A     :ΏA     Í  9U  : �A     ׍  9U  :8�A     �  9U 9Ts  :S�A     �  9U 9T� 9Q| 
��9Rs  ;F�A     =�  4�  9Us  8a�A     =�  9Us    J�  l�A      l�A     �       q)�  K)�  � � Ll�A     �       Z6�  ��ZB�  ��~ZO�  ��~Z[�  ��~Mg�  � � [t�  ��A     ;��A     ̸  �  9U 9T��~9Q��~9R��9X��~ 8$�A     ~�  9Uu 9Qq 9Rr 9Xx    J��  *�A      *�A     �       �Տ  K�  	  K�  . , L*�A     �       M�  W Q M'�  � � c��  {�A      {�A            9K��  � � K��  � �    Ji�  ��A      ��A            �
�  Kw�   
  N��  t�A      p|   3�  K��  1 /  J��  ܑA      ܑA     #       �h�  K��  V T  Jӿ  ��A      ��A            ���  K�  { y K�  � �  J��  �A      �A            ��  K
�  � � K�  � �  J%�  !�A      !�A            �.�  K3�    K@�  4 2  J��  2�A      2�A     #       �c�  K��  Y W  J��  U�A      U�A     #       ���  K��  ~ |  N��  x�A      �|  ���  K��  � �  J��  ��A      ��A            ���  K�  � �  J�  ��A      ��A            �+�  K!�  � �  N��  ��A      �|  �q�  K��    K��  N J S$�A     9U   J��  ԒA      ԒA            �Ò  K��  � � K��  � � SޒA     9U   Jg�  �A      �A     (       6 �  K��  � � Ku�  � � S�A     9U   J��  �A      �A     !       / J�  K��       J��  4�A      4�A            + �  K��  ?  =   JV�  J�A      J�A     +       � �  Kd�  d  b  LJ�A     +       Mq�  �  �  M|�  �  �  M��  �  �    J�  u�A      u�A            l /�  K�  �  �  K�  �  �   J+�  ��A      ��A            h q�  K9�  ! ! K9�  ! !  J��  ��A      ��A     u       � �  K�  C! A! K�  h! f! L��A     u       M �  �! �! M+�  �! �! M6�  �! �!   J�   �A       �A            ` .�  K�  w" u" K�  w" u"  J!�  ;�A      ;�A            X p�  K<�  �" �" K/�  �" �"  J��  K�A      K�A     0       T ͕  K��  �" �" K��  # 	# 8\�A     ��  9U 9T
A-  J��  {�A      {�A            ' �  K �  0# .#  J�  ��A      ��A     %       # 7�  K�  U# S#  J*�  ��A      ��A             ��  K8�  z# x# 8ǔA     ~y 9Q@  NF�  ԔA       }   ʖ  KT�  �# �# Ka�  �# �# 8�A     �y 9T@  Jo�  �A      �A             ��  K}�  $ $  J��  �A      �A             4�  K��  8$ 6$  J��  )�A       )�A             ��  K��  ]$ [$ K��  ]$ [$ K��  �$ �$  Jľ  @�A      @�A             ŗ  KҾ  �$ �$ K߾  �$ �$  J"�  Q�A      Q�A            � ��  K0�  �$ �$  N�  ƘA      @}  � #�  K�  % %  J��  ~�A      ~�A            �X�  K��  ;% 9%  N��  ��A      p}  ���  K��  `% ^%  Jʦ  ��A      ��A            � ��  Kئ  �% �%  N��  וA      �}  � �  K��  �% �% K��  �% �% O�}  M��  9& 1& M��  �& �& 8��A     ��  9Uu    J��  ,�A      ,�A     %       �w�  K�  ' ' K	�  :' 8' S<�A     9U 9Q0  J$�  Q�A      Q�A     *       �Ι  K?�  _' ]' K2�  �' �' Sa�A     9U 9Q0  JM�  {�A      {�A            ��  K[�  �' �'  Nr�  ��A      �}  � m�  K��  �' �' K��  ( ( O�}  M��  Y( U( M��  �( �( 8D�A     ��  9Uu    Nb�  m�A       ~  ��  K}�  �( �( Kp�  ) ) O ~  M��  C) =) M��  �) �) :��A     ՚  9U  S�A     9U    N��  ��A      P~  �@�  K��  �) �) K��  * * OP~  M��  )* '* SҗA     9U    N�  ߗA      �~  | ��  K:�  P* L* K-�  �* �* O�~  MG�  �* �* MR�  �* �* M]�  + 
+   Ni�  >�A      �~  x �  Kw�  J+ D+ O�~  M��  �+ �+ [��  ��A       J��  ٘A      ٘A     �       JΜ  K��  �+ �+ K��  H, F, L٘A     �       M��  m, k, M��  �, �, M̱  �, �, :,�A     y�  9U  :W�A     ��  9U 9T�9Q| 
��9Rs  Sk�A     9U 9T� 9Qv 
��9Rs    J��  t�A      t�A     Q       A ��  K�  E- C- K��  j- h- Lt�A     Q       M�  �- �- Y�_ ��A      �~   K�_ �- �- K�_ �- �- O�~  M�_ . �- M�_ F. B.     Jʽ  řA      řA     0       P ޝ  K�  �. �. Kؽ  �. �. 8֙A     ��  9U 9T
 @  N>�  њA         = f�  KY�  �. �. KL�  	/ / Y�  �A       P  TKD�  G/ ?/ K7�  �/ �/ K*�  -0 )0 OP  MQ�  m0 c0    N�  ��A      �  � T�  K�  1 �0 K��  ~1 x1 O�  M�  �1 �1 M�  �2 �2 M%�  �3 �3 M0�  K4 C4 M<�  �4 �4 MH�  Z5 R5 ^U�  �  �  MZ�  �5 �5 Mf�  =6 56  N��  t�A       �  \��  K�  �6 �6 K�  �6 �6 K��  �7 ~7 K��  �7 �7 O �  X�  8]�A     �v 9Q�9R�d�  �   ^s�  @�  ��  Mt�  L8 F8 M��  �8 �8  N��  ��A      ��  t>�  K�  �8 �8 K�  �8 �8 K��  \9 T9 K��  �9 �9 O��  X�  8>�A     �v 9Q�9R�d�  �   8ћA     �  9Uu    J#�  D�A      D�A     }       ���  K>�  : : K1�  C: A: LD�A     }       MK�  h: f: MV�  �: �: :y�A     Ԡ  9U  S��A     9U 9T�9Qs 
��   J�  ��A      ��A     $       �h�  K9�  �: �: K,�  �: �: L��A     $       MF�  �: �: SܜA     9U    N��  �A       ��  Fˡ  K��  #; ; K��  ]; Y; O��  M��  �; �; M��  �; �; P��A     �y   J4�  ��A      ��A     �       � 9�  KO�  �; �; KB�  < < L��A     �       M\�  @< << Mg�  y< w<   J��  l�A       l�A            � {�  K��  �< �< K��  �< �<  Nչ  ��A      ��  � ޢ  K�  �< �< K�  &= "= O��  M��  ^= \= M�  �= �= M�  �= �=   Nĺ  �A       �  � '�  Kߺ  �= �= KҺ  > > O �  M�  X> T>   J��  ԟA      ԟA     D       � ��  K��  �> �> K��  �> �> LԟA     D       M��  �> �> M��  ? �>   Jv�  �A      �A     t       � A�  K��  ;? 9? K��  `? ^? L�A     t       M��  �? �? M��  �? �? c��  *�A      *�A            rK��  �? �? K��  �? �?    ;h~A     �  Y�  9Uu  ;KA     �  w�  9U 9Tv  ;��A     �  ��  9U  ;^�A     <�  ��  9U  ;�A     ��  Ť  9U 9Tv  8��A     %i 9U d�  v   UP�  ��  7def � 1O  &@ "@ 4�� � 1O  s@ o@ O��  4�{  � �  �@ �@ YD�  A      ��  � Kp�  A 	A Kc�  FA DA KV�  kA iA O��  X}�  8%A     �c 9U 9Tt 9Qq      N��  �zA      �s  Eѥ  K�  �A �A K�  B �A  8�zA     �  9Uu   7O  H�i  ��A     �       �ʦ  fexc � �<  U7def �1O  �C �C 4�� �1O  D D O�]  4�c ��  �D �D YD�  ?A      ^  �	Kp�  �D �D Kc�  E E KV�  UE OE O^  X}�  8PA     �c 9Uu 9Tt 9Qq      0�~  ~�  -��  ~�+   0�  `4�  gexc `%�<  -��  a%�+  /�m  c
	  /�  d�  .i f
	   0�c  �u�  gexc � �<  -��  � �+  .K �	  /K1 ��J   0�h  &�  gexc &�<  -��  '�+  /mv  )"	  .k )"	  .A *"	  .C *"	  .P *"	  .B +	  1�0  h H��  ��@     �      ��  bexc �<  �E �E 3��  ��+  :F 2F 4mv  �"	  �F �F 7k �"	  �F �F 7A ��  �G xG 7C �"	  �G �G 7P �"	  �H vH 7B �	  I �H 5�0  W�@     :��@     ͨ  9Us  S��@     9Us 9Ts�   H�s  � GA           ���  bexc ��<  EJ 7J hV �W  ��4� �  �J �J 4c+  
	  GK CK 4�k  
	  �K }K 44w  
	  �K �K 4�  
	  �K �K 4oI 

	  LL @L 4� �  �L �L N��  !IA       @k  Vf�  KȬ  9M 3M K��  �M �M K��  �M �M K��  =N 9N K��  {N sN O@k  Xլ  X�  X�  X��  X�  X�  X!�  X.�  X;�  8�HA     �n 9U��9X|    J��  =IA       =IA     7       e?�  KȬ  �N �N K��  O O K��  ,O *O K��  SO OO K��  �O �O L=IA     7       Xլ  X�  X�  X��  X�  X�  X!�  X.�  X;�  8jIA     �n 9U��9T
��9Qv 9R 9Xs    J��  {IA       {IA     *       l�  KȬ  �O �O K��  P 	P K��  2P .P K��  lP jP K��  �P �P L{IA     *       Xլ  X�  X�  X��  X�  X�  X!�  X.�  X;�  8�IA     �n 9U��9Qs9R 9Xs    Y��  �IA       pk  bK��  �P �P K��  �P �P K֭  (Q $Q Kʭ  bQ ^Q K��  �Q �Q Opk  M�  �Q �Q M�  nR hR    0�r  ���  -Հ  �(�W  gp1 �(
	  gp2 �(
	  -1v  �(
	  -zf  �(
	  .i �
	  /�  �;	  /
�  �;	  /�  �;	  //�  �%;	  /'j  �+;	  /,j  �1;	  /؊  �7;	  /�k  �?;	  Rh�  /A  �;	  /#�  �
	   Ry�  .x �;	   E/�� �H	  /jw  ��  E.x �;	     09�  ~��  -Հ  ~"�W  gp1 "
	  gp2 �"
	  gp �"
	  .i �
	  .dx �;	   0�z  V<�  gexc V�<  -��  W�+  /oI Y�  /� Z�   H�n  � �@           ���  bexc ��<  �R �R 4�a  �;	  ^S TS 4)c  �;	  �S �S 4�  �T  ,T &T 4Bw  �T  {T uT 4�~  ��  �T �T 5�0  I	�@     U�V  ��  7vec ��  6U ,U N�_ ��@      �V  �^�  K�_ @W <W K�_ ~W xW O�V  M�_ �W �W M�_ (X $X   N�_ ��@      �W  ���  W�_ W�_ O�W  M�_ gX cX M�_ �X �X   S�@     9Us   UpU  S�  4oI 
	  �X �X 4|�  ;	  HY >Y 4�j  ;	  �Y �Y /��  ';	  6��@     _       �  7vec �  Z Z N�_ ��@      �U  ��  K�_ �[ �[ K�_ �[ �[ O�U  M�_  \ �[ M�_ C\ ?\   N�_ �@      @V  а  W�_ W�_ O@V  M�_ �\ ~\ M�_ �\ �\   S<�@     9Us   :J�@     ��  9Us  :q�@     	�  9Us  :��@     .�  9Us 9Ts�9Q 
�� 8w�@     ~y 9U~ 9T��9Q��  :��@     g�  9Us  :��@     {�  9Us  S&�@     9Us   0�  �ڱ  gexc �!�<  -��  �!�+  .p1 ��  .p2 ��  /3{  �;	   0Yv  6��  gexc 6�<  -��  7�+  /oI 9�  .a0 :�  .a1 :�  .b0 ;�  .b1 ;�  /�f  =;	  /�i  =;	  .dx ?;	  .dy ?;	  .dax @;	  .day @;	  .dbx A;	  .dby A;	  .val C;	  .R E�   0��  ���  gexc � �<  /oI ��  /3{  �;	  1�0  ) H��  ��@     �      ���  bexc �<  ]  ] 3��  �+  k] g] 4oI �  �] �] 4�q  "	  ^ �] 4�  ;	  �^ �^ 43{  ;	  T_ P_ 4�j  ;	  �_ �_ 4|�  ;	  ` ` 4g  ;	  V` T` 4+{  ;	  }` {` 5�0  ���@     N�  P�@      �T  �M�  KD�  �` �` K7�  a �` K*�  wa sa O�T  XQ�    :�@     a�  9Us  ;��@     =�  y�  9U  ;��@     =�  ��  9U  :��@     ��  9Us  :	�@     ��  9Us  :��@     Ӵ  9Us 9T  S��@     9Us 9Ts�9Q} 
��  0Cm  }��  gexc }�<  -��  ~�+  /oI ��  /|�  �;	  /3{  �;	  /+{  �%;	  1�0  �Rz�  /�(  �T  /�(  �T   E/�(  �T  /�(  �T  E.vec ��     0�  �  gexc �<  -��  �+  /�q  "	  /oI �  /3{  ;	  /|�  ;	  /g  ;	  1�0  p 0��  �i�  gexc ��<  -��  ��+  /oI ��  /�j  �;	  /3{  �;	   0Sp  ���  gexc ��<  -��  ��+  /oI ��  /3{  �;	   0؋  ��  gexc ��<  -��  ��+  .dx �;	  .dy �;	  /oI ��  /�~  ��  1�0  � 0;g  ���  gexc ��<  -��  ��+  .zp �v<  /Hg  ��  .dx �;	  .dy �;	  /�� ��  .i ��   0g  ��  gexc ��<  -��  ��+  .zp �v<  /Hg  ��  .dx �;	  .dy �;	  /� ��  /�! ��  /�S ��  /�� ��  .i �$�   0a  Q~�  gexc Q�<  .zp Sv<  /Hg  T�  .dx V;	  .dy V;	  /oI W�  1�0  } 0f~  (̸  gexc (#�<  -oI )#�  gdx *#;	  gdy +#;	  -Mu  ,#�   26d  ��  P�@     �      �Ϲ  bexc �/�<  �a �a bx �/Ϲ  b b by �/Ϲ  qb eb 3Xc  �/�<  �b �b 3Hg   /\1  Qc Kc 7zp v<  �c �c 7p �  ff `f 7d ;	  �f �f :0�@     ��  9Us  ;J�@     ~y ��  9U}  8i�@     ~y 9U}   ;	  0
h  ��  gexc �"�<  -��  �"�+  .I ��  .K ��  .L ��   0��  �i�  gexc �!�<  -��  �!�+  .I ��  .K ��  .L ��   0ņ  ���  gexc ��<  /oI ��  1�0  � 0n�  jĺ  gexc j!�<  -��  k!�+   0�i  ;��  gexc ;!�<  -��  <!�+  .A >�   0�e  �C�  gexc �!�<  -��  �!�+  .K  "	  .L  "	  .Kf  "	   0;|  �l�  gexc ��<  -��  ��+   0lr  ���  gexc ��<  -��  ��+   0cr  ���  gexc ��<  -��  ��+   0Zr  ��  gexc ��<  -��  ��+   0>�  -��  gexc -�<  -��  .�+  .A 0	  .B 0	  .C 0	  .p1 1�  .p2 1�  /6f  3�  Rs�  .v1 BT  .v2 CT   E.v1 _T  .v2 `T    0�|  �#�  gexc ��<  -��  ��+  .K ��  .L ��  .D �;	  R��  /�(  �T  /�(  �T   E/�(  T  /�(  T  E.vec �     0i�  �b�  gexc ��<  -��  ��+  .K �	  .L ��   0^�  ���  gexc ��<  -��  ��+  .L �"	  .R �;	   0�d  zʽ  gexc z!�<  -��  {!�+   0J{  i�  gexc i�<  -��  j�+   0A�  [�  gexc [�<   0��  M+�  gexc M�<   0�  ?G�  gexc ?�<   0�x  2c�  gexc 2�<   0j  %�  gexc %�<   0�h  ��  gexc �<   0*�  ľ  gexc �<  -��  �+   0��  ��  gexc ��<  -��  ��+   i4k  �0 }  ��  gexc � �<   0�h  �/�  gexc ��<   0>p  �X�  gexc ��<  -��  ��+   0Z�  ���  gexc ��<  -��  ��+   0��  ���  gexc ��<  -��  ��+   0�j  �ӿ  gexc ��<  -��  ��+   0r}  ���  gexc ��<  -��  ��+   0i}  |%�  gexc |�<  -��  }�+   0`}  nN�  gexc n�<  -��  o�+   0�  _w�  gexc _�<  -��  `�+   0�e  P��  gexc P�<  -��  Q�+   0�  7��  gexc 7�<  -��  8�+  .S :�  .X ;	  .Y ;	   0P�  4�  gexc �<  -��  �+  .S �  .X  	  .Y  	   0�d  P�  gexc �<   0�i  �y�  gexc ��<  -��  ��+   0�x  ���  gexc ��<  -��  ��+   0�}  ���  gexc ��<  .AA ��  .BB ��  /6f  ��   ,w�  ��  p�  gexc ��<  -/e  ��  -5e  ��  gVec �p�  .A �	  .B �	  .C �	  .p1 �T  .p2 �T  /6f  ��   �	  0�f  a��  gexc a�<  -��  b�+  .L d�  .K d�   0Of  G��  gexc G�<  -��  H�+  .L J�  .K J�   0�g  (3�  gexc (�<  -��  )�+  .L +�  .K +�   0�g  r�  gexc �<  -��  �+  .L �  .K �   08u  ���  gexc ��<  -��  ��+  .def �1O  /�� �1O   0�  ]�  gexc ]!�<  -��  ^!�+  .F `"	  /�  a�  .def b1O  1�0  �E/�� w1O    0��  ��  gexc �<  -��  �+  .F "	  /�  �  .def 	1O  1�0  QE/�� 1O    0Lm  ���  gexc ��<  /��  ��   0E�  ���  gexc ��<  -��  ��+  .n �"	  .rec �1O  /�� �1O   0ky  �!�  gexc ��<  -��  ��+   0e�  J�  gexc �<  -��  ��+   0&e  \s�  gexc \�<  -��  ]�+   i�o  O0��  .��  gexc .�<  /Ca  0�   0ot  ��  gexc �<  -��  �+  /Ca  �  .Out �   2K�  ��  �@     �       �-�  fexc ��<  U5}  �^�@      0��  �V�  gexc ��<  -��  ��+   0І  ���  -��  ��+  .A �	  .B �	  .C �	   05�  ���  gexc ��<  -��  ��+  .L �	   0�  ~�  gexc ~�<  -��  �+  .L �	  .K �	   0�|  p"�  -��  p�+   0�~  b>�  -��  b�+   0�h  Qg�  gexc Q�<  -��  R�+   0	�  @��  gexc @�<  -��  A�+   0Ef  3��  gexc 3�<   i�s  $0$�  ��  gexc �<  -��  �+  .I "	   0p  ��  gexc ��<  -��  ��+  .I �"	   04x  �R�  gexc ��<  -��  ��+  .I �"	   0d�  ���  gexc ��<  -��  ��+  .I �"	   0�  ���  gexc ��<  -��  ��+  .I �"	   0Au  ���  -��  ��+   0"s  ~��  -��  ~�+   0.~  q�  -��  q�+   0go  c*�  -��  c�+   0S�  VF�  -��  V�+   0�f  Eo�  gexc E�<  -��  F�+   0�q  8��  -��  8�+   0�p  +��  -��  +�+   0�m  ��  -��  �+   0�~  ��  -��  �+   0'y  ��  -��  �+   0@t  �
$�  gexc �
�<  -��  �
�+   0�d  �
M�  gexc �
�<  -��  �
�+   0�}  �
i�  -��  �
�+   0n  �
��  -��  �
�+   0��  �
��  -��  �
�+   0Qq  �
��  -��  �
�+   0�k  �
��  -��  �
�+   0�|  �
��  -��  �
�+   0�w  �
�  gexc �
�<  -��  �
�+   0
t  z
E�  -��  z
�+  .L |
	   0�g  m
a�  gexc m
�<   i��  `
0��  S
��  -��  S
�+   0e  8
��  gexc 8
�<  -��  9
�+   0~  *
��  gexc *
�<  -��  +
�+   ,nj  �	�  �  gVx �	;	  gVy �	;	  gR �	p�  .V �	�   H�x  �	@�@     �      �I�  fexc �	"�<  U 2�  �	;	  0�@            ���  fexc �	�<  Ufdx �	�  Tfdy �	�  Q 2�q  }	;	   �@            ���  fexc }	�<  Ufdx ~	�  Tfdy 	�  Q 2��  b	;	  ��@     8       ���  fexc b	!�<  Ubdx c	!�  �f �f bdy d	!�  +g 'g c��  ��@      ��@     5       f	K�  fg dg K
�  �g �g K��  �g �g K��  h h L��@     5       M"�  ,h &h M/�  �h }h    2��  G	;	  ��@     8       ���  fexc G	�<  Ubdx H	�  �h �h bdy I	�  �h �h c��  ��@      ��@     5       K	K�  8i 6i K
�  hi fi K��  �i �i K��  �i �i L��@     5       M"�  �i �i M/�  Sj Oj    HKv  �@�@     \      ���  fexc �"�<  U3 �   	".	  �j �j 3�N 	"	  �k |k  0�e  �'�  gexc �"�<  -dt  �"�   ,�y  �;	  n�  gexc �#�<  -3{  �#;	  -r�  �#;	  .val �;	   ,�i  l;	  ��  gexc l �<  -3{  m ;	  -r�  n ;	  .val p;	   ,i  :;	  ��  gexc :)�<  -3{  ;);	  -r�  <);	  .val >;	   ,vl  ;	  C�  gexc %�<  -3{  %;	  -r�  %;	  .val ;	   ,Fj  �;	  ��  gexc �'�<  -3{  �';	  -r�  �';	  .val �;	   ,K�  �;	  ��  gexc �'�<  -3{  �';	  -r�  �';	  .val �;	   ,cq  �;	  �  gexc �"�<  -3{  �";	  -r�  �";	  .val �;	   ,�d  _;	  _�  gexc _�<  -3{  `;	  -r�  a;	  .val c;	   H�{  = �@            ���  fexc ='�<  UIXc  >'�<  T3oI ?'�  Yl Ul I3{  @';	  R H�  1��@            �#�  fexc 1'�<  UIXc  2'�<  T3oI 3'�  �l �l I3{  4';	  R H<{  ��@     M       ���  fexc "�<  UIXc  "�<  T3oI "�  �l �l I3{  ";	  R H�n  �P�@     G       ���  fexc �"�<  UIXc  �"�<  T3oI �"�  m m I3{  �";	  R Hч  �`�@     �       ���  bexc �%�<  Um Im 3Xc  �%�<  �m �m 3oI �%�  hn \n 33{  �%;	  �n �n 7v �;	  �o �o ;��@     ~y ��  9U}  8��@     ~y 9U}   H{  � �@     +      �D�  bexc � �<  �o �o 3Xc  � �<  Bp :p 3oI � �  �p �p 33{  � ;	  'q q 7v �;	  �q �q P��@     ~y 8�@     ~y 9U��  ,�x  E�  ��  gexc E'�<  -�  F'�  gaIP G'	  /�a  I��   �L  ,Mg  +�  ��  gexc + �<   H�i  ��@     -       �<�  bexc '�<  r r bidx '"	  Zr Tr 3�\ ';	  �r �r ;��@     1�  '�  9Uv  8��@     �x 9U|   H �  
@�@            ���  fexc 
�<  Ufidx "	  TI�\ ;	  Q Hd�  ��@     0       ��  bexc (�<  �r �r bidx ("	  Ps Js 3�\ (;	  �s �s ;��@     1�  ��  9Us  8��@     �x 9Uv   H�  �0�@            �a�  fexc ��<  Ufidx �"	  TI�\ �;	  Q 22�  �;	  ��@     9       ��  bexc �'�<  �s �s bidx �'"	  Ft @t N�_ ��@       �Y  ��  K�_ �t �t K�_ �t �t O�Y  M�_ /u +u M�_ ru nu   8��@     1�  9Us   2֐  �;	   �@            �[�  fexc ��<  Ufidx �"	  T 2��  �	   �@     &       ���  bexc �+�<  �u �u N�_ )�@       �Y  ���  K�_ v �u K�_ *v $v O�Y  M�_ �v �v M�_ �v �v   8)�@     1�  9Us   2Sh  �	  �@            �1�  fexc �!�<  U 2��  �	   �@     �       ���  bexc �"�<  w w LT�@     *       7x �;	  fw bw 7y �;	  �w �w P_�@     =�  ;l�@     =�  ��  9Uq 9Tr 0$0& Pw�@     �y   ,b  b[  =�  gax b$[  gay c$[  gbx d$�  gby e$�  /  j.  /Bo  k.   2��  [  ��@            ���  fa $[  Ubb $�  �w �w 7ret .  3x +x 7tmp .  �x �x  a?�  G�<  ��A     �       ���  3K1 G�J  �x �x 4R�  Iu  <y 8y )� JU	  �X4�6  L�<  |y ry 1�0  _N��  �A       �  Y��  K�  �y �y K�  ,z &z O �  Z)�  �\[6�  h�A     ;�A     �x ��  9Uv 9T 9Q09R 9X09Y�\ 8p�A     @�  9Us    8թA     �y 9Uv 9T
P9Q�X  ,~  U	  �  -�6  #�<   0ہ  �5�  -�6  �$�<  -�  �$�@  .i ��   2�h  �U	  ��@     T      �(�  3�6  �$�<  z uz 3�  �$�4  �z �z 3�  �$�@  y{ s{ 7i ��  �{ �{ htmp �"	  �X4'I ��a  8| .| 4� �U	  �| �| ;=�@     (�  �  9T�X9Q89Rs0 8��@     (�  9T�X9Q19Rs�  2b  UU	  `�@     W       ���  3R�  Uu  �| �| 3�  V�-  9} 3} 3�z  W"	  �} �} 3;o  Xa   �} �} 3�:  Y"	  ~ ~ )� [U	  �\4<o  \�   l~ f~ 8��@     �x 9T19Rv �Q9Y�\  ,Su  U	  @�  -�6  !�<  -R�  !u  /� U	  1�v  4 `��  �0�@     �       ���  >�6  �$�<  �~ �~ ?R�  �u  #  ;S�@     �x ��  9Uv  ;r�@     �x ��  9Uv  ;��@     �x ��  9Uv  j��@     �x 9T�U  k�h  �
�  B�6  �'�<  B�a  �'�   k��  �H�  B�6  �%�<  B�a  �%�  B2�  �%a   Bss  �%	   k�w  }��  B�6  }&�<  B�a  ~&�  _IP &	  Cpn  ���   Hٌ  cP�@     	      ���  3�  c�4  a Y 4R�  eu  � � 4�  f�2  � � O X  7i k
	  O� M� 4�m  k
	  u� s� ;��@     �x (�  9U|  ;��@     �x @�  9U|  ;��@     �x X�  9U|  ;��@     �x p�  9U|  ;��@     �x ��  9U|  ;�@     �x ��  9U|  ;,�@     ��  ��  9U~  ;<�@     �x ��  9U|  ;T�@     �x ��  9U|  ;h�@     �x  �  9U|  ;��@     ��  �  9U~  ;��@     �x 0�  9U|  ;��@     �x H�  9U|  ;��@     �x `�  9U|  ;��@     ��  x�  9U~  ;��@     �x ��  9U|  ;��@     �x ��  9U|  ;�@     �x ��  9U|  ;)�@     �x ��  9U|  GG�@     �x   H��  >p�@     �       ���  3�  >6�4  �� �� 3�{  ?6�P  ۀ Հ 4R�  Au  )� '� 7i B
	  \� L� ;��@     �x p�  9U}  ;��@     �x ��  9U}  ;��@     �x ��  9U}  ;"�@     �x ��  9U}  8;�@     �x 9U}   ,�e  U	  !�  -�  "�4  -�u  "�;  -�   "�G  -�  !"�G  -2�  ""G   2M�  �U	  P!A     �      �l�  3�  �,�4  � 
� 3�^ �,
	  �� �� 3�S  �,l�  (� � 3Z�  �,
	  �� �� 4Jy  �A  *� � 4R�  �u  �� �� 4�  ��2  �� � 4�  �T  � � 4,q  �T  �� �� 4�y  �r�  *�  � )� �U	  ��4��  �"	  �� �� 4�u  �
	  E� ?� 4C�  �"	  ň �� 4�  �"	  � � 7i �
	  �� |� 7j �
	  *� �� 4:�  ��  � � 4h  ��  �� �� 4
�  ��  e� Y� )�  �
	  ��)�  �
	  ��4oo  �\1  � � 4f  �\1  � � 4�  �\1  -� %� 4�u  ��;  �� �� 4~  ��;  u� c� 5��  
"A     5lE  �(A     Up`  ��  4V�  
	  E� ;� 4Sn  
	  � ޓ 4�� H	  �� x� U�`  ��  4Um  _�  � ޔ 4]m  `�  �� �� N�_ �,A      a  _V�  W�_ K�_ �� �� Oa  M�_  �� M�_ � �   Y�_ �,A      @a  `W�_ K�_ �� �� O@a  M�_ ї ˗ M�_ )� #�    Upa  P�  7idx ��  �� �� N�_ l&A      �a  � �  W�_ K�_ ʘ Ƙ O�a  M�_ (� $� M�_ k� g�   Y�_ �&A      �a  � W�_ W�_ O�a  M�_ �� �� M�_ � �    U�b  ��  4Um  ��  2� (� 4]m  ��  �� ��  Nx�  �&A      0b  �	U�  K��  a� Y� K��  a� Y� K��  ՛ ś K��  �� � K��  � � O0b  M��  a� W� M��  �� ҝ M��  {� u� M��  Ҟ Ğ M��  �� i� M��  �� y� N	�  d)A       �b  \��  KV�  �� �� KI�  8� 4� K<�  v� r� K/�  �� �� K#�  � �� K�  R� N� O�b  Xc�  Xn�  Xy�  X��  X��  X��  X��  X��  X��  8I)A     �k 9Rv 9X��}9Y��}   J	�  **A       **A     J       s��  KV�  �� �� KI�  �� �� K<�  آ ֢ K/�  �� �� K#�  7� 5� K�  ^� Z� L**A     J       Xc�  Xn�  Xy�  X��  X��  X��  X��  X��  X��  8\*A     �k 9U9Ts 9Q 9R} 9X��}9Y��}   J	�  �*A       �*A     9       {��  KV�  �� �� KI�  �� �� K<�  � � K/�  � 	� K#�  2� .� K�  l� j� L�*A     9       Xc�  Xn�  Xy�  X��  X��  X��  X��  X��  X��  8�*A     �k 9U~ 9T}9Q 9R} 9X��}9Y��}   c��  �+A      �+A     �       jK"�  �� �� K�  �� �� K�  ߤ ݤ K��  � � K��  +� '� L�+A     �       M/�  i� c� X:�      ;�$A     �x m�  9U}  ;�$A     �x ��  9U}  ; %A     �y ��  9U��~ ;#%A     � ��  9U~ 9Ts 
��9Q��~9R��~9X��~ ;�%A     
# ��  9U}  ;�%A     
# 	�  9U}  ;#(A     �x +�  9U��~9T��~ ;>(A     �x K�  9Us 9T��~ ;K(A     �x k�  9Us 9T��~ ;�)A     �x ��  9U}  ;�)A     �x ��  9U}  ;+A     �$ ��  9U} 9Q�� 8X+A     �x 9U}   ;�!A     �x �  9U 9T@9Q09R| 9X09Y�� ;"A     �x #�  9U 9T��} ;!"A     �x C�  9U 9T��} ;-"A     �x b�  9U 9Tw  ;}"A     �x ��  9U 9T@9Q09R| 9X09Y�� ;�"A     �x ��  9U 9T19Qw 9R| 9Xw 9Y�� ;�"A     qy ��  9U}  ;#A     �x ��  9U}  ;:#A     �x ,�  9U 9T89Q09X09Y�� ;k#A     �x Z�  9U 9T89Q09X09Y�� ;�#A     �x ��  9U 9T89Q09X09Y�� ;�#A     �x ��  9U}  ;�#A     �x ��  9U}  ;�(A     �x ��  9U 9T��~ ;�(A     �x ��  9U 9T��~ ;�(A     �x �  9U 9T��~ ;�(A     �x 0�  9U}  ;�(A     �x P�  9U 9T��~ 8�-A     �$ 9U} 9Q��  `  �  0�o  0	�  -�S  0'l�  -�  1'T  -�q  2'T  -�y  3'r�  /c+  5�  /�k  6�  /yu  8�  /u~  9�  /oI ;�  /� <�   0��  ���  gp1 �%S   gp2 �%S   -1v  �%S   -zf  �%S   -�q  �%T  -�  �%T  .p �
S   .i �S   .out ��  .in1 ��  .in2 ��  /�a  ��  /�a  �"�  .d1 �(�  .d2 �,�  E/�� H	    0  �H�  gp1 �S   gp2 �S   gref �S   -�q  �T  -�  �T  .p �S   /� ��   2�h  �U	  @A     �      ���  3�  � �4  ʥ �� 3Jy  � A  �� �� )� �U	  ��4R�  �u  �� t� 4�q  �"	  #� � )>k  �"	  ��4�u  �
	  �� �� 4C�  �"	  -� � 4�  �"	  �� �� 7i �
	  =� 1� 7j �
	  � ǫ 4:�  ��  �� � 4h  ��  �� �� 4
�  ��  � � 4�  ��2  }� y� )�  �
	  ��)�  �
	  ��4oo  �\1  Ǯ �� 4f  �\1  �� �� 4�  �\1  ð �� 4�o  ��;  @� 4� 5�u  ��A     5�u  �tA     U[  ��  4V�  
	  ͱ ñ 4Sn  
	  t� f� 4�� H	  >� 6� U�[  ��  4(�  j	  �� �� c�_ �A      �A            n&W�_ K�_ ҳ г L�A            M�_ � � M�_ K� G�    UP[  y�  4{}  �S   �� �� 4(�  �	  �� �� Y�_ �A      �[  �+W�_ K�_ � � O�[  M�_ $�  � M�_ g� c�    ;�A     �x ��  9U|  ;�A     �x ��  9U|  ;�A     �y ��  9U~  ;�A     � ��  9U} 9Ts 
��9Q~ 9Rw 9X  ;A     
# �  9U|  ;A     �x 0�  9U��9T��~ ;*A     �x P�  9U��9Tv  ;�A     �x h�  9U|  ;A     �x ��  9U|  ;\A     �$ ��  9U| 9Q�� 8�A     �x 9U|   :�A     ��  9Uv 9Travc9Q| 9R�� ;�A     �x ��  9Us  ;�A     �x �  9Us 9T~  ;�A     �x 3�  9Us 9Tw  ;�A     �x Q�  9Us 9T  ;�A     �x i�  9U|  ; A     y ��  9U|  ;>A     �x ��  9U|  ;kA     �x ��  9Us 9T89Q09X09Y�� ;�A     �x ��  9U|  ;�A     �x �  9Us 9T89Q09X09Y�� ;�A     �x %�  9U|  ;�A     �x S�  9Us 9T89Q09X09Y�� ;
A     �x k�  9U|  ;A     �x ��  9U|  ;�A     �x ��  9U|  PBA     �x ;j	A     �$ ��  9U| 9Q�� 8�	A     �x 9U|   2ty  EU	  `cA     �       �c�  3�  E#�4  �� �� 3� F#
	  F� 6� 4� HU	  � �� 4�  I�2  �� �� 46~  JG  ݷ ׷ 4�|  L
	  +� '� 5�u  ��cA     Un  -�  4R�  `u  q� m� 4$S  a�F  �� �� 4��  cx-  Ҹ θ )A  d�  �H:�cA      �  9Us 9Q�H ;dA     �x �  9U|  84dA     Q�  9Us   ;�cA     Q�  O�  9Us 9T09Q0 8GdA     � 9T0  2i�  �
U	  `dA           �Q�  3�  �
!�4  � � 3�u  �
!
	  �� �� 3�   !�  #� � 4� U	  �� �� 4�  �2  � � 7i 
	  i� ]� 7nc 
	  �� � ;/eA     � -�  9T0 8YeA     �  9U} 9T09Q09R1  2�o  v
U	  �`A     c      ���  3�  v
!�4  L� @� 3�u  w
!
	  ׼ Ѽ 3�  x
!�  2�  � )� z
U	  ��4�  {
�2  �� �� 46~  |
G  <� 4� 7i }

	  �� �� 4R�  ~
u  E� A� 7c �
�  �� {� 7n �
�  �� �� 4cj  �
�  �� �� 4(�  �
�  -� � 5�u  �
UbA     6�aA     L       ��  4� �

	  R� N� 4��  �
x-  �� ��  6xbA     P       ��  7a �
r-  �� ��  ;�aA     �x �  9U| 9T89Q09X09Y�� ;&bA     �q 4�  9Ts 9R d8 }  ;6bA     �  W�  9U} 9Q 9R0 ;`bA     �x u�  9U| 9T  ;�bA     �  ��  9U}  ;�bA     � ��  9T0 8cA     �x 9U| 9T89Q09X09Y��  2�  (
U	  peA           ���  3�  (
�4  #� � 3�u  )

	  �� �� 3�  *
�  2� &� 4� ,
U	  �� �� 4�  -
�2  #� � 7i .

	  x� l� 7nc .

	  �  � ;?fA     � ��  9T0 8ifA     �  9U} 9T09Q09R1  ,�n  �	U	  �  -�  �	�4  -�u  �	
	  -�  �	�  /�  
U	   2�  &	U	  @XA     �      �� 3�  &	�4  c� O� 3�u  '	
	  O� 7� 3�  (	�  [� C� 3'�  )	�  e� ]� )� +	U	  ��4�  ,	�2  �� �� 46~  -	G  &� � 7i .	
	  �� �� 4�d  0	�  j� R� 4R�  2	u  �� p� lZ   5	�  Bz   m�  ��   4cv  :	��  :� 0� 5�u  �	�[A     U�l  ��  4(�  {	�  �� �� .j |	
	  7c }	�  K� C� 7n ~	�  �� �� LwYA     N       7idx �	
	  3� -�   N� @ZA        m  �	.  K� �� �� K� �� �� K� V� N� K� �� �� O m  M� � � M� �� �� M� �� �� M� B� (� M ^� T� M �� �� ^ pm  |�  M f� `� P�[A     ~y  N�_ F[A      �m  T��  K�_ �� �� K�_ �� �� O�m  M�_ �  � M�_ G� C�   c�_ �[A      �[A             QK�_ �� �� K�_ �� �� L�[A             X�_ X�_     N� �]A      �m  b	� K� �� �� O�m  M� R� L� M� �� �� M� �� �� Z� ��M� �� �� M� D� <� Z� ��M �� �� M �� �� Z" ��[F M_A     :�]A     
 9U| 9Travg9Q��~9R�� ;�]A     Wy $ 9U��~ ;^A     �y R 9U��~9T	�6H     9Q�� ;�^A     �x � 9U��~9T89Q09X09Y�� ;�^A     �x � 9U��~ ;_A     y � 9U��~ ;A_A     �x � 9U��~ ;�_A     �x � 9U��~ ;�_A     �x  9U��~ ;#`A     �x 4 9U��~9T89Q09X09Y�� ;G`A     qy N 9U��~ ;j`A     �x h 9U��~ ;�`A     �x � 9U��~ 8�`A     �x 9U��~   ;ZA     �y � 9T~ 9Q
s ����3$ ;)\A     �x � 9Uw  ;E\A     �Y  � 9U|  ;Z\A     �x 
 9Uw  ;�\A     � ! 9T0 ;(]A     H�  9 9U|  ;K]A     �x h 9Uw 9T89Q09X09Y�� 8�]A     �x 9Uw 9T89Q09X09Y��  2�  �U	   MA     ?      �h 3�  ��4  � �� 3��  �G  � � 4Jy  �A  �� z� 4R�  �u  �� �� )>k  �"	  ��~)� �U	  ��~4�  �"	  i� [� 7i �
	  �  � 7j �
	  �� �� 46~  �G  !� � 4a�  ��  �� �� 7nsc ��  � � 4dk  ��  �� �� 7a �r-  `� R� 7c ��  � �� 7ns �x-  �� �� )��  �gV  ��~4��  ��  s� g� 4�|  �
	  � � 4�m  �
	  �� �� 4�  �\1   � � 4��  �o	  �� �� 4e�  �o	  � � 4$~  �o	  g� a� 4�l  �o	  �� �� 4;e  �o	  � � 42�  �o	  �� �� 4bs  ��  � � )�u  �"x 	 7H     )�t  �"� 	 7H     5�u   	�WA     6�QA     �       { )X�  _�V  ��8�QA     �y 9Uv 9T	 7H     9Q~   6WWA     -       � 4x  �"	  t� p� ;_WA     Wy � 9Uv  ;jWA     �  � 9U}  8uWA     qy 9Uv 9T~   U`l  � 4$S  ��F  �� �� 4;�  ��  �� �� )vw  ��  ��~)�c  �!�  ��4c  �
	  b� \� :�RA     � 9U} 9TA9Q��~9R~  :SA     � 9U} 9T29Q��~9R~  S)SA     9U} 9T69Q��~9R��~  U0l   7n �
	  �� �� ;�MA     �y  9U��}9Q��~ P�MA     �y  N6 xSA      �l  � KD �� �� O�l  MQ )� %� M^ a� _� Mk �� �� Mx �� �� M� � � M� j� b� Z� ��~M� �� �� Z� ��M� �� �� M� /� -� M� V� T� ]� XA            	 M� }� {� 8XA     � 9U} 9Tt   :�SA     C	 9U} 9TRAVM9Qv 9R��~ ;�SA     Wy [	 9Uv  ;�SA     �y z	 9Uv 9T��~ ;�SA     �y �	 9Uv 9T2 ;!TA     �y �	 9U~ 9T09Q��~ ;@TA     �y �	 9Uv 9T4 ;hTA     �y �	 9Uv 9T��~ ;�TA     �y 
 9Uv 9T��~ ;�TA     Wy /
 9Uv  ;�TA     = Y
 9U} 9T��~�
����~" ;�TA     �x �
 9U~ 9T@9Q09X09Y��~ ;"UA     qy �
 9Uv 9T��~ ;FUA     �x �
 9Uv  ;~UA     y �
 9Uv  ;�UA     �x �
 9Uv  ;�UA     �x  9Uv  8�WA     �x 9Uv    :OA     A 9Travg9Qv 9R��~ :3OA     k 9U} 9T2FFC9Qv 9R��~ :XOA     � 9U} 9Travf9Qv 9R��~ ;oOA     Wy � 9Uv  ;�OA     �y � 9Uv 9T	 7H     9Q��~ ;�OA     �y   9U��}9T�9Q��~ ;WPA     �y H 9U��}9T#| 2$| "������~"��~"��}"��~"# 9Q��~ ;BQA     qy ` 9Uv  ;�RA     �x � 9U��}9T89Q09X09Y��~ ;]VA     �x � 9Uv 9T��~ ;tVA     �x � 9Uv  ;�VA     �x � 9Uv  ;�VA     y � 9Uv  ;�VA     �q # 9T��~�9R| d8 ��~ ;�VA     �x ; 9Uv  ;(WA     �x S 9Uv  8>WA     qy 9Uv   �#  x L    	h �#  � L    	} 07�  * -�   �4  -�u   
	  -�   �  -�v   �  /�  �2  /6~  G  .a r-  .i 
	  .j 
	  .nc 
	  E.av 0�O    0Yj  �� -�  �$�4  -�u  �$
	  -�  �$�  -cj  �$�  /�  ��2  /6~  �G  .i �
	  .j �
	  .a �r-  .av ��O  E/�a �H	    2x  >H	  P�@           �� 3�  >"�2  �� �� 3Sn  ?"�  :� 4� 3:�  @"�  �� �� 3h  A"�  &� � 3
�  B"�  �� �� 7i D
	  � �� 4�� EH	  �� �� P��@     ~y P�@     ~y  ,^{  �U	  P -�  ��4  /Jy  �A  /R�  �u  /�  ��2  /� �U	  .i �
	  .j �
	  />k  �"	  /��  �"	  /C�  �"	  /��  ��U  ) �  �"x 	�6H     1�u   0v   � -�   �4  /�  "�2  /�\ #�Q  /�� #�Q  R� .p .�;  /� /�   E/�� KT    2�  U	  0�@            �6 3D� (�
  *� &� 3R   (a   g� c� 4�  	�@  �� �� 8B�@     �]  9T1  0�u  �� -�  ��4  /Jy  �A  /R�  �u  /�  ��2  /�{  ��P  /�\ ��Q  /�� ��Q  /� �U	  /�y  ��  />k  �"	  /� �"	  /B�  ��  /��  �"	  E.p ��;    2�l  I�;  @�@     �      �V 3�  I'�4  � �� I�l  J'"	  T7p L�;  �� ��  2Os  .U	  PkA     
       �� 3�  . �4  �� �� 3n�  / 
	  � � 3"c  0 yD  I� E� jZkA     l 9U�U9T�T9Q�Q9R1  2�x  %U	  `kA            �l 3�  % �4  �� �� 3n�  & 
	  �� �� 3"c  ' yD   � �� jgkA     l 9U�U9T�T9Q�Q9R0  2u  �U	  0jA           � 3�  �!�4  C� 9� 3n�  �!
	  �� �� 3"c  �!yD  �� �� 3�(  �!�  e� U� 4� �U	  %� � 4]c  �
	  �� �� 4�n  �
	  �� �� 4� ��  "�  � 4>) ��Q  I� E� 5�u  �jA     6�jA            � 7idx �
	  �� �  6�jA            � 4k  P  �� ��  ;�jA     � � 9T0 ;�jA     Qm � 9Us�	9Rv d s  8:kA     � 9T1  ,<~  T�  � -�  T+�4  -�{  U+�P  -�n  V+
	  -]c  W+
	  /k  YP  /~  Z�;  /��  \
	  .j \
	  /\d  ]H	  /[�  ^H	  /� _H	  E/sf  kH	  /(�  l
	  /dh  n_P  E/�{  tH	     2�  �U	  �fA     l      �D 3�  ��4  �� �� 3�(  ��  y� q� 4Jy  �A  �� �� 4R�  �u  !� � 4�  ��2  �� �� 4>) ��Q  �� �� 4� �U	  � � 4�y  ��  @� <� )>k  �"	  ��4� �"	  �� v� 4B�  �"	  �� �� 4�p  �"	  L� B� 1�u  6ND �hA      @n  *	 K} �� �� K} �� �� Kp �� �� Kc &� � KV �� �� O@n  M� �� �� M� � � M� s� q� M� �� �� M� �� �� M� <� 8� M� �� �� M� �� �� M�     [� jA     ^ �n  K M m  g  M �  �  M �  �  m, �n  M-   8�iA     �y 9U 9T��   ;�hA     qy m 9U 9Tw s " ;�hA     �y � 9U 9T�� ;�hA     �y � 9U 9T�� ;iA     �x � 9U��9T49Q09X09Y�� 8<iA     �x 9U��9T49Q09X09Y��   :gA     3 9U~ 9TRAVV9Qs 9R�� :;gA     W 9TRAVH9Qs 9R�� ;OgA     Wy o 9Us  ;`gA     �y � 9Us 9T�� ;zgA     �y � 9Us 9T2 ;�gA     �y � 9Us 9T�� ;�gA     �y � 9Us 9T�� ;�gA     �y  9U} 9T89Q�� ;hA     = 6 9U~ 9Tw  "9Q}  P`hA     �y  ,��  gU	  = -�  g;�4  -x  h;"	  gmap i;LQ  -�{  j;�P  /Jy  lA  /R�  mu  /� oU	  /ߣ  q�  /��  r
	  /�q  s
	  /�  t
	  .i u
	  .j u
	  1�u  �E/nl  �
	  /�n  �
	  /]c  �
	  E/�U  ��     2��  �U	  �A     
      ��  3�  �6�4  F B 3x  �6"	  �  3�{  �6�P  � � 4Jy  �A  Q M 4R�  �u  � � )� �U	  ��4ߣ  ��  � � 4t�  �"	   � 7i �
	  ` N 7j �
	  @ $ 7k �
	  d b 43c  �
	  � � 4�  ��2  � � 4k  �P   � 4|�  ��-  . $ 5�u  _)A     6�A     �       � 4�k  �_P  � � U \  n 4�S ��  � � 4T�  ��  � � 7end � �    ;IA     �y 3 9Us 9T�� ;gA     �y R 9Us 9T�� 8�A     �y 9Us 9T��  8A     �x 9Uv 9TH9Q09X09Y��  UP\  � 4� H�  9 7 8wA     �y 9Us 9T��  U�\   4� T�  ^ \ 8�A     �y 9Us 9T��  ;A     qy + 9Us 9T|  ;4A     �x I 9Uv 9T  ;]A     �y h 9Us 9T�� ;�A     �y � 9Us 9T�� ;�A     �y � 9Us 9T�� ;�A     �x � 9Uv 9T89Q09X09Y�� ;A     �y � 9Us 9T�� ;=A     qy  9Us 9T��| " ;VA     �y 5 9Us 9T�� ;vA     �y T 9Us 9T�� ;�A     �x � 9Uv 9T89Q09X09Y�� ;�A     �x � 9Uv 9TH9Q09X09Y�� ;3A     qy � 9Us  ;LA     �y � 9Us 9T�� ;jA     �y   9Us 9T�� ;�A     �y %  9Us 9T�� ;�A     �x S  9Uv 9T49Q09X09Y�� ;�A     �y r  9Us 9T�� 8;A     �x 9Uv 9T29Q09X09Y��  H��  5�
A           �
# 3�  5�4  � � 4Jy  7A  � � 4R�  8u    4�  9�2  b \ 4zx  :�O  � � )� ;U	  ��4��  <	  � � 4�q  =	  B	 4	 7i >�  �	 �	 7j >�  T
 J
 )>k  ?"	  ��5�u  �iA     :A     �! 9U�U9Trava9Qs 9R�� ;=A     �x �! 9Us  ;MA     y " 9Us  ;XA     y " 9Us  ;qA     �x 3" 9Us  ;�A     �x g" 9U} 9T@9Q09R~ 9X09Y�� ;�A     �x " 9Us  ;A     �x �" 9U} 9T@9Q09X09Y�� ;7A     �x �" 9Us  ;QA     �x �" 9Us  ;�A     �x �" 9U}  8�A     �x 9U}   <@�  ��;  ��@     X      ��$ >Jy  �'A  �
 �
 >�  �'"	  I E >Cc  �'
	  � � ?�o  ��;    ?|  �
	  � � @cnt �
	  � � @i �
	  9 ) @j �
	  � � ?R�  �u  � � (� �U	  ��;��@     �x ($ 9U��9T29Q09Rv ����9X09Y�� ;�@     %y @$ 9U~  ;<�@     %y X$ 9U~  ;��@     �x p$ 9U~  8��@     �x 9U��  <�  �\1  ��@     �      �Z& >Jy  �'A    >�  �'"	  z n >In  �'�;    ?�  �\1  � � @n �
	    ?|  �
	  � � @i �
	  S 7 @j �
	  � z ?N� ��    � ?R�  �u  P J (� �U	  ��;��@     %y �% 9U|  ;?�@     �x �% 9U} 9T29Q09R~����9X09Y�� ;h�@     %y �% 9U|  ;��@     %y �% 9U|  ;��@     %y & 9U|  ;,�@     �x -& 9U|  ;d�@     �x E& 9U|  8�@     %y 9U|   2�s  
U	  P�A     �      ��- 3�  
 �@  � � 3)�  �
 K     3�^ �
 
	  o g 3:1  �
 [  � � 4� �
U	    )��  �
BB  ��|1�u  I6�A     �       ( 4�  �
�4  � � )R0  �
�  ��{)C  �
(�  ��|)�  �
�  ��|)  �
)�  ��|NZ �A      ��  �
�' K6Z %  K*Z z t KZ � � KZ � � S:�A     9U��{9Ts 9Q} 9R��{9X��|  8T�A     �Y 9U��{9T} 9Qs 9R��|9X|   NI7 ��A       �  �
�( K[7   K�7 � x Ku7 � � Kh7 F @ O �  M�7 � � M�7 � � M�7 � � M�7   Z�7 ��|SзA     9Q} 9R 9Yv�   J�- ϸA      ϸA             �
) K�- } { 8�A     	z 9U|�9T09R0  N�_ �A      `�  �
t) K�_ � � K�_ � � O`�  M�_ � � M�_ : 6   N�_ E�A      ��  �
�) K�_ w u K�_ � � O��  M�_ � � M�_     N�7 ��A      ��  <~, K�7 V J K�7 � � O��  M�7 r f M
8 � � Z8 ��|M$8 S E M18 � � M>8 N  H  ^K8 0�  �* MP8 �  �  Y�W  ��A       `�  iKX  �  �  KX  /! +! KX  u! q! O`�  M,X  �! �! M8X  " �! MEX  X" T" MRX  �" �"    ^^8 ��  \, M_8 �" �" Ml8 a# S# ^y8 ��  :+ M~8 �# �# 8 �A     �x 9T��{  ^�8 �  �+ M�8 8$ 4$ Z�8 ��|M�8 w$ s$ S��A     9T} 9Q19R��|  N�_ ̼A      @�  ��+ K�_ �$ �$ K�_ �$ �$ O@�  M�_ �$ �$ M�_ @% <%   N�_ �A      ��  �+, K�_ }% {% W�_ O��  M�_ �% �% M�_ �% �%   ;z�A     �x E, 9T��{ 8��A     �x 9T��{  8(�A     z 9U��{#�9T��|   J�- /�A      /�A             ?�, K�- & & 8O�A     	z 9U|�9T09R0  ;��A     �- - 9U| 9T~ 9Qv 9R 9X1 ;ϸA     �8 )- 9U| 9T} 9Q09R1 ;ڹA     �- X- 9U| 9T~ 9Qv 9R 9X0 ;�A     �8 �- 9U| 9T} 9Q09R0 8پA     "z 9Uv�9Q0  0�  Z
�- -��  Z
9   2��  0	U	  ��A     �      �I7 3��  0	!9  .& && 3�  1	!�@  �& �& 3)�  2	!K  s' ]' 3:1  3	![  p( b( 3��  4	!�  +) ) 4�  6	�4  x* t* 4Jy  7	A  �* �* 4� :	U	  �* �* 4�  ;	�  2+ "+ 4K1 >	�J  , , U`�  7 4�6  M	�<  �, �, 4�g  N	�  - �, 4�m  P	�  . . 4y�  Q	�  s. k. 4�p  b	�  �. �. 6�A     �       �/ 7i  

	  �/ �/ J�_ @�A      @�A     '       $
�/ K�_ �/ �/ K�_ 0 0 L@�A     '       M�_ D0 @0 M�_ �0 �0   8��A     �b  9Uv 9T����  N�`  ��A      ��  g	�6 K�`  �0 �0 K�`  >1 <1 O��  M�`  o1 a1 [�`  ��A     N�`  ��A      ��  jD6 K a  2 2 W�`  O��  Za  ��Xa  M'a  �2 �2 M4a  �2 �2 XAa  MNa  +3 %3 e[a  ^da  0�  �0 Mia  �3 }3  N�r  m�A      p�  <72 K�r  �3 �3 K�r  4 4 W�r  K�r  U4 O4 Op�  Z�r  ��;w�A     �x B1 9U��9T@9Q09R��9X09Y�� ;��A     �x z1 9U��9T@9Q09R��9X09Y�� ;�A     �r  �1 9U�� ;��A     �x �1 9U��9T@9Q09R��9X09Y�� ;¶A     �x 2 9U��9T19Q09R��9X09Y�� 8�A     �x 9U��9T29Q09R09X09Y��   ^wa  ��  R2 Mxa  �4 �4  N�d  �A      ��  W�4 K�d  �4 �4 K�d  C5 =5 O��  M�d  �5 �5 M�d  �5 �5 M�d  6 6 ]�d  w�A     ?       �2 M�d  q6 i6 M�d  �6 �6  J
�  ��A      ��A            SC3 K;�  [7 Y7 K/�  �7 ~7 K#�  �7 �7 K�  �7 �7  J��  ĲA      ĲA            Y�3 K��  �7 �7 K��  8 8  J��  ڲA      ڲA            Z�3 K��  ;8 98 K��  a8 _8  J�   �A       �A     ]       n(4 K�  �8 �8 K�  �8 �8 L �A     ]       M)�  �8 �8   JH�  �A      �A     #       ^�4 Km�  89 69 Ka�  ^9 \9 KU�  �9 �9 L�A     #       Mx�  �9 �9   ;��A     5�  �4 9U��9T 9Qv  SH�A     9U��   ;ȭA     �x �4 9U�� ;�A     �x 5 9U�� ; �A     �x 5 9U�� ;�A     �x 85 9U�� PL�A     @�  ;t�A     �r  _5 9U�� P��A     ��  ;;�A     �x �5 9U��9T(9Q09X09Y�� ;w�A     �x �5 9U��9T(9Q09X09Y�� ;��A     �x �5 9U��9T89Q09X09Y�� ;�A     �x .6 9U��9T89Q09X09Y�� 82�A     �a  9Uv    m�`  ��  M�`  �9 �9 M�`  k: g: J�_ ��A      ��A     '       {�6 K�_ �: �: K�_ �: �: L��A     '       M�_ ; �: M�_ D; @;   8�A     �b  9Uv     8ݫA     5�  9U 9T| 9Qv   L%�A     3       4�V  D
�  �; ; 8A�A     /z 9U}    ,Z �U	  �7 -�  �"�@  -)�  �"K  -�^ �"
	  -:1  �"[  /�  ��4  /$S  ��F  /Jy  �A  /� �U	  /�  ��0   ,��  9U	  �8 -��  9%9  -�^ :%
	  /�  <�4  /K1 ?�J  /�!  B  /�� CH	  /)�  DK  /�  E�@  R^8 /Ą  f�.   E.top ��  /�  ��  R�8 /�  ��   E/�i  �'�"  /f  �'�!  /� �'U	     2R~  �U	  �-A     �      ��K 3��  �#9  �; �; 3�^ �#
	  = �< 3Q�  �#
	  �> U> 3bl  �#�  w@ o@ )� �U	  ��}4�� �H	  �@ �@ 4�� �H	  �A �A 4x  �"	  �B �B 4�  ��4  2C C 4�V  ��  rD XD 4'  ��  �E �E )Fy  �{  ��~)��  �=
  ��}4�z  ��  �F �F 5�u  &03A     5Ii  �<A     6�3A     �      �: )�  ��K ��~)s  ��K ��})[  ��K ��})�S  �`  ��~8�4A     !�  9Ts 9Q��~9R4  U�d  �E 4R�  �u  �H pH 4-1 �
	  @I 6I 4�e  �
	  �I �I 4�8  �"	  �J �J 4D� ��
  K K 4�i  ��
  :K 6K U�h  �< 7i 0A  �K pK 4�� 0A  YL SL 4�l  1�  �L �L )�S  3`  ��~4�  4T  >M 6M 4s  5�   �M �M 4[  6Z  
N N ;j9A     �x �; 9U��}9T@9Q09X09Y��} ;�9A     �x < 9U��}9T19Q09X09Y��} ;�9A     �x =< 9U��}9T29Q09X09Y��} ;';A     !�  b< 9U~ 9Ts 9Q��~ ;(<A     �x z< 9Us  ;D<A     �x �< 9Us  8`<A     �x 9Us   U@e  �B 7n �
	  XN TN 4ŀ  �
	  �N �N 4�l  ��  O �N 42]  �
	  �O �O 44  �
	  Q Q 4o�  �
	  IQ EQ 4�}  �A  �Q Q 4
�  ��  9R -R U�f  �@ 7pp ��K �R �R 4g�  ��  �T �T 4��  ��  �T �T NWM ~?A       g  �@ K�M �T �T K�M ?U 5U KvM �U �U KiM @V 6V O g  M�M �V �V Z�M ��~M�M W W M�M iW WW M�M @X .X ]�M >A     E       �> M�M Y Y M�M �Y �Y M�M �Y �Y MN DZ BZ MN iZ gZ  ];N �?A     |       �? M<N �Z �Z MIN �Z �Z N�_ �?A      `g  �? K�_ �Z �Z K�_  [ �Z O`g  M�_ '[ #[ M�_ j[ f[   N�_ @A      �g  �`? K�_ �[ �[ W�_ O�g  M�_ �[ �[ M�_ \ \   nVN =@A     .       MWN O\ M\ MdN u\ s\   ]N �BA     n       k@ M N �\ �\ M-N �\ �\ N�_ �BA      �g  �@ K�_ �\ �\ K�_ ] ] O�g  M�_ 9] 5] M�_ |] x]   N�_ �BA      @h  �P@ W�_ W�_ O@h  X�_ X�_   P�BA     �y P�BA     �y  ;�@A     ;z �@ 9U��~9T��|# 8�@A     "z 9U��~9T| 9Q}    8�>A     �8 9Us 9Q��}�9R0  N�L �AA      �e  yB K�L �] �] K�L O^ G^ K�L �^ �^ O�e  Z�L ��~MM T_ P_ MM �_ �_ ^ M f  �A M!M �_ �_ M.M 1` -` M;M m` g` ZHM ��~;�6A     �y �A 9Us 9T��~ ;<7A     (�  �A 9T��~9Q19Xv  ;r7A     Hz �A 9Us 9Qv  8xBA     qy 9Us   N�P �7A       `f  6AB KQ �` �` KQ �` �` K�P &a "a K�P ea ca  ;\8A     O ^B 9U} 9T1 8-CA     Uz 9Us 9Q0   8�=A     az 9U��|  NL ]5A       e  �B K$L �a �a KL �a �a O e  M1L %c c   N�_ �<A      �h  �/C K�_ �c �c K�_ �c �c O�h  M�_ �c �c M�_ d d   N�_ =A       i  ��C K�_ Ud Sd K�_ |d zd O i  M�_ �d �d M�_ �d �d   J�_ �<A      �<A            ��C K�_ %e #e K�_ Le Je L�<A            M�_ ue qe M�_ �e �e   J�_ �<A      �<A            �aD K�_ �e �e K�_ f f L�<A            M�_ Ef Af M�_ �f �f   J�_ +=A      +=A     !       ��D K�_ �f �f K�_ �f �f L+=A     !       M�_ g g M�_ Xg Tg   J�_ V=A      V=A     !       �=E K�_ �g �g K�_ �g �g LV=A     !       M�_ �g �g M�_ (h $h   ;�5A     mz ]E 9U��}9T|  ;�8A     mz |E 9U}�9T|  :�8A     �E 9U}  :�8A     �E 9U}  ;AA     �y �E 9U��}9TH9Q��} ;0AA     yz �E 9U��} 8?AA     az 9U��|  NtN &/A      c  ��G K�N kh ch Oc  M�N �h �h M�N 7i +i M�N �i �i M�N 0j .j ^�N `c  SG M�N [j Sj M�N �j �j M�N pk jk M�N �k �k M�N l l N�_ @0A      �c  �F W�_ K�_ Ll Hl O�c  M�_ �l �l M�_ �l �l   c�_ e0A      e0A            W�_ W�_ Le0A            M�_ 
m m M�_ Mm Im    N�P 6A      d  ��G KQ �m �m KQ �m �m K�P �m �m K�P �m �m  ;�/A     !�  �G 9Q|�  ;�0A     O �G 9U} 9T0 P~6A     �y   J�_ >2A      >2A            �VH K�_  n �m K�_ 'n %n L>2A            M�_ Pn Ln M�_ �n �n   J�_ _2A      _2A            ��H K�_ �n �n K�_ �n �n L_2A            M�_  o o M�_ co _o   N�_ �2A      @d  �I K�_ �o �o K�_ �o �o O@d  M�_ �o �o M�_ 3p /p   N�_ �2A      pd  �pI K�_ pp np K�_ �p �p Opd  M�_ �p �p M�_ q �p   J�_ �2A      �2A            ��I K�_ @q >q K�_ gq eq L�2A            M�_ �q �q M�_ �q �q   J�_ �2A      �2A            �LJ K�_ r r K�_ 7r 5r L�2A            M�_ `r \r M�_ �r �r   :n.A     gJ 9Ts 9Q��} ;�.A     �[  �J 9Uu 9Ts 9Qq  ;�.A     ?L �J 9Uu  ;�.A     !W �J 9Ts  :/A     �J 9U}  :&/A     �J 9U}  ;�0A     az �J 9U��| ;01A     �z K 9U  :g1A     /K 9U} 9Ts  :|1A     CK 9U}  :�1A     WK 9U}  :�1A     lK 9T��} ;�1A     X �K 9U} 9Ts  ;2A     ?L �K 9U}  ;2A     !W �K 9Ts  8r3A     X 9U} 9Ts   �  �K L    �   �K L    A  L L    ,b�  ��
  ?L -�$ �!�
  gidx �!
	  .cur ��
   He  �`�@     �       ��L I��  � 9  U4�x  ��  �r �r 4�g  ��  7s 1s 4�~  ��  �s �s 4K1 ��J  �s �s  ,��  �U	  WM -��  �*9  --1 �*
	  -�e  �*
	  /� �U	  /�S  �l�  .i �
	  E/Jy  A  /s  �  /�v  �  .tmp "	    ,5�  <U	  tN -��  <09  -�l  =0�  --1 >0
	  -ŀ  ?0
	  /�V  A�  /�� B`  /�  C�  .x D�  .y D�  RN /2]  W
	  .k X
	  .l Y
	  .p1 ZT  .p2 [T   R;N /��  �H	  /P|  �H	   E/�� �H	  /�� �H	  E/�  ��4  /K1 ��J     ,f  �U	  O -��  �'9  /�V  ��  /� �U	  /�S  �l�  /Z�  ��  E.vec �T  /�� �T  /�� �H	  /�� �H	  /�n  ��    o�  U	   �@     Y      ��P 3��  9  Yt Mt 3aa  �  �t �t 4�  �4   u u 4K1 �J  Ju Du 4Xc  �<  �u �u 4s  	  ?v 9v 6��@     `      �P 4� MU	  �v �v 4�V  O�  �v �v 4Rl  P`  �v �v N
�  ��@       �X  SPP K;�  w w K/�  :w 8w K#�  _w ]w K�  �w �w  Y��  �@       Y  YK��  �w �w YH�  �@      PY  Km�  �w �w Ka�  �w �w KU�  x x OPY  Mx�  @x >x     PF�@     �y PM�@     �y  0Mc  �&Q -Xc  �"�<  -��  �"'  --1 �"
	  -�e  �"
	   0ih  �BQ -�  �#�4   2�  /U	   A     4      ��R 3��  /'9  nx fx 4� 1U	  �x �x 7p 2�.  �y ]y 4�� 3�.  �{ �{ 4�V  4�  �{ �{ 4�l  5�  
| | 44  6
	  a| S| 5�0  � A     1Г  �U�\  �R 7xx =H	  	} �| 7xy =H	  �} �} 7yy =H	  x~ d~ 7yx =H	  a S 4.� >
	  � � 8�A     �z 9Us 9T   O ]  4Jy  �A  �� �� PA     Wy   2�p  FU	  P�@     �      ��U 3��  F$9  � ր 4� HU	  �� �� 7p I�.  �� M� 4�� J�.  �� �� 4�V  K�  � � 4�  L�  (� $� 4�S  Ml�  d� ^� 4s  N�  �� �� 4Z�  O�  �� �� 4&| Q�.  r� X� 4Xq  Q�.  �� � 7c R�  ܇ · 4.� R�  x� t� 7vec ST  �� �� 4Es  ST  � �� 7x T�  �� u� 4�t  U�;  � � 4-i  U�;  �� �� 4�t  U)�  C� ;� QE�  V�   1�0  %1��  (U�Y  �T htmp �"	  ��;
�@     (�  �T 9T��9Q19Xw  8_�@     �y 9Tw 9Q��  U0Z  U 7y ��  �� �� 7f ��  �� ��  UpZ  KU 7y �  �� � 7f �  �� ��  ;� A     Uz nU 9U| 9T09Q~  8� A     Uz 9U| 9T9Q0  2�  *U	  ��@     �       ��U I��  *$9  U7p ,�.  ?� 1� 4�� -�.  �� ގ  H�t   ��@     	       �@V 3��   %9  	� � 4Jy  "A  F� B� G��@     �x  2ur  U	  `�@     R       �!W 3��  %9  �� }� 3�^ %
	   � �� 3x  %"	  =� 9� 3�  	%
	  �� v� 4� U	  �� �� 4Jy  A  3� /� ;y�@     qy  W 9Us 9T�Q 8��@     �x 9Us 9T| ����  `�s  � �@     �       �X >��  �-9  q� i� >�^ �-
	  ֑ Б ?�  ��4  &� "� ?R0  ��  d� ^� pC  �"�   ?�  ��  �� �� p  �#�   q�u  ���@     O�T  (f  �"�!  �P?� �"U	  � � Sv�@     9T�T9Q09Rw    <_�  zU	  �A     �       ��Y >��  z9  -� '� >�^ {
	  � y� ?�  }�4  ͓ ˓ ?� �U	  � � ?Jy  �A  � � (R0  ��  �H(C  �"�  �J(�  ��  �L(  �#�  �N@pos �"	  >� :� rZ :A      p]  �_Y K6Z x� t� K*Z �� �� KZ � � KZ *� (� SOA     9Uv 9T09Q} 9R�H9X�L  ;-A     Wy wY 9U|  ;hA     �Y �Y 9Uv 9T} 9R�J9X�N 8sA     qy 9U| 9T~   k6y  ]Z B�  ] �4  _idx ^ 
	  B/  _ �  _tsb ` �;  _ah a \1   k�~  KBZ B�  K �4  _idx L 
	  _lsb M �;  _aw N \1   ,�}  8�  �Z -K1 8"*  -[x  9"  /k  ;h  /E  <�  /�|  =*  /$S  >�F   2,s  �U	  @�A     �       ��[ 3�q  � �  [� M� 3�k  � (  � �� 3�^ � 
	  � �� 3:1  � [  �� {� 4 �K  I� ;� 4�  ��@  �� � 4�  �T  �� � )� �U	  Ps��A     Z& �[ 9U�T9T�U j��A     Z& 9U�T9T�U  ,!z  IU	  (\ -�  I%(  greq J%Q  /�k  L�@  /� MU	  R\ /e5  T�4  /$S  U�F  /-U V"	   E/��  m
	    2p  $U	  ��@     S       �2] 3�  $(  ܚ Қ 3-U %"	  Y� Q� 4e5  '�4  �� �� 4�k  (�@  �� �� 4� )U	  e� _� 6��@     !       ] 4$S  7�F  �� �� 44  8�C  ߜ ל S��@     9T�T9Qs  P�@     �z 8�@     �]  9Us 9T0  Az  �U	  �] Be5  �T  B�S �
	  B.� �
	  B?1  �[  B\-  ��  Fnn �
	  C�  ��4  R�] Ftsb ��  Fah ��   E.lsb �  .aw �    <�n  �U	  ��@     3       ��^ >e5  �T  J� D� >�U  �
	  �� �� >B7  �
	  � � >Y�  �T  B� :� ?�  ��4  �� �� ?$S  ��F  �� � S�@     9U�U9T�T9Q�Q  <Zw  xU	  @A     /       �=_ >~ x!*  H� D� >n  y!  �� ~� =�\ z!9  Qp� |U	   ?K1 }�J  �� �� ?Nz  
	  � ݟ LlA            @val ��;  � �   A  ?U	  �_ B~ ?!*  Bn  @!  B�\ A!9  B�R  B!�  C� DU	  CK1 E�J  ECNz  N
	  R�_ Fs T   EFiv \�;     A�6  �[   ` _a �[  _b �[  Fret �.  Ftmp �.   t�  �@     (       �J` u*�  UK7�  F� @� KD�  �� �� MQ�  �� ��  t�Y pA     |       �!a K�Y (� � K�Y �� �� K�Y O� I� K�Y �� �� K�Y  � � ^�Y @]  �` K�Y p� l� K�Y �� �� K�Y У Σ K�Y �� � K�Y � �  v�A     9U�U9T19Q�T9R�R9X�X  t2] �A           ��b KC] I� =� KO] ؤ Τ K[] W� M� Kg] Х ̥ Ks] � 	� M] �� �� M�] Ц Ħ 6A     "       �a Z�] ��Z�] ��8)A     �Y 9U| 9Ts9Q09R} 9X~   m2] �]  Kg] Y� U� Ks] �� �� K[] � � KO] ?� 9� KC] �� �� O�]  M] ި ڨ X�] n�] �A     +       Z�] ��Z�] ��cZ �A      �A     "       	K6Z � � K*Z =� ;� KZ f� `� KZ �� �� S�A     9U| 9T09Qs9R} 9X~       t��  �A     f       ��c K��  ܩ ֩ K��  .� (� K��  �� z� u�  Ru�  Xn��   A     #       K��  Ϊ ̪ K�  � � K�  � � K��  =� ;� K��  b� `�   tD�  PA     ]       ��c uV�  Uuc�  Tup�  QM}�  �� ��  t��  �A     7       �{d u��  Uu��  TK��  ë �� M
�  1� %� n��  �A            K��  ݬ ۬ K��  �  � K��  ?� =� L�A            M
�  l� b�    t��  �A     <       �e u��  Uu��  TK��  � � M��  w� q� n��  �A            K��  Ϯ ͮ K��  �� � K��  1� /� L�A            M��  X� T�    tC�   A     :       ��e uU�  Uub�  TKo�  �� �� M|�  � � nC�   A            KU�  �� �� Ko�  а ʰ Kb�  � � L A            M|�  K� A�    t��  @A     7       �[f u�  Uu�  TK(�  � � M5�  V� J� n��  `A            K�  �  � K(�  )� %� K�  d� b� L`A            M5�  �� ��    t��  �A     7       ��f u��  Uu��  TK��  4� ,� M��  �� �� n��  �A            K��  N� L� K��  u� q� K��  �� �� L�A            M��  ݵ ӵ    tn�  �A     R       ��g u��  Uu��  TK��  |� x� M��  �� �� nn�  �A            K��  � � K��  >� <� K��  c� a� L�A            M��  �� ��    t'�   A     U       �;h u9�  UuF�  TKS�  ӷ ˷ M`�  =� 5� n'�  XA            KS�  �� �� KF�  �� � K9�  � � LXA            M`�  @� <�    tJ�  �A     �       ��h uX�  Uue�  TnJ�  �A     "       Ke�  �� �� KX�  �� ��   t~�  A     �       �%i u��  UK��  � ܹ u��  Qu��  Ru��  Xm~�  @^  K��  2� .� K��  l� h� K��  �� �� K��  � ܺ K��  � �   t��  �A     �      ��k K�  X� P� W�  M�  �� �� M*�  *� � M7�  Ǽ �� MD�  %� #� [Q�  A     ]Z�  #A     $       �i M_�  N� J� Ml�  �� �� SDA     9Us   N�  hA      p^  �-j KD�  �� �� K7�  6� 2� K*�  p� l� Op^  MQ�  �� ��   ^z�  �^  �k M{�  � � M��  w� q� ]��  �A     ]       'k M��  ڿ п N�_ �A      �^  ��j K�_ �� �� K�_ �� �� O�^  M�_ � � M�_ \� X�   N�_ �A      `_  �k W�_ W�_ O`_  M�_ �� �� M�_ �� ��   SA     9Us   J�_ [A      [A            ��k K�_ � � K�_ B� @� L[A            M�_ i� e� M�_ �� ��   S[A     9Us   :�A     �k 9Us 9T  :�A     �k 9Us  SA     9Us 9Ts�9Q} 
��  t	�  �A     �      �Qm K�  �� �� K#�  R� N� K/�  �� �� K<�  R� D� KI�  �� �� KV�  B� 8� Mc�  �� �� Mn�  � � My�  6� ,� M��  �� �� M��  C� 7� M��  �� �� M��  �� {� M��  �� �� M��  �� �� m��  �_  M��  �� �� N�_  !A      0`  !8m W�_ K�_ �� �� O0`  M�_ � � M�_ O� K�   8 A     �x 9Ts |    t pCA     �      ��n K$ �� �� K1 � � K> ^� X� W MK �� �� MX �� �� Me 8� ,� Mr �� �� M} Z� P� M� �� �� M� 0� *� m� Pi  M� �� �� M� a� [� M� �� �� ^� �i  Kn M� �� �� P�DA     �x  Y�_ RDA      �i  �K�_ #� � K�_ �� �� O�i  M�_ �� �� M�_ &� "�     t��  `EA     �      �Dp K��  i� a� K��  �� �� K��  O� G� K��  �� �� KȬ  �� �� Mլ  ,� (� M�  j� b� M�  �� �� M��  2� .� M�  p� h� M�  �� �� M!�  '� � M.�  �� �� M;�  �� �� ^y�   j  ,p Mz�  _� W� M��  �� �� m��  Pj  M��  U� M� N�_ �FA      �j  �p K�_ �� �� K�_ �� �� O�j  M�_ 	� � M�_ L� H�   8�FA     �x 9Uw ��9T	����   mh�   k  Mm�  �� ��   t�[ @JA     �       ��q K�[ �� �� K�[ h� X� M�[ '� � M�[ �� �� U�k  �p M�[ l� j� M�[ �� �� Z
\ �X:iJA     �p 9T| 9Q�X 8KA     (\ 9Us   ]�[ �JA     P       �q K�[ �� �� K�[ �� �� L�JA     P       X�[ M�[ 6� 0� ]\ �JA     @       q M\ �� � 8�JA     ~y 9T
   8�JA     �]  9Us 9T0   8�JA     �z 9T|   t* 0KA     �      ��r KE �� �� KR � � K_ �� �� W8 Ml �� �� My 3� /� M� �� i� M� �� �� M� � � M� ~� t� ^� �k  yr M� �� �� P�KA     �x P�LA     �x  P�LA     ~y  t��  �fA     7       �Us K��  y� s� K��  �� �� K��  � � M��  V� T� ]��  �fA            .s K��  {� y� K��  �� �� K��  �� �� L�fA            X��    8�fA     �  9Us 9Tv 9Q�Q9R1  tP pkA     k      �|t K^ �� �� Mk �� � Mx �� �� M� �� �� 6�kA     /       t M� 7� 1� M� �� �� ;�kA     � �s 9U~ 9Tt  8�kA     Qm 9U} d ~   mP  o  K^ �� �� O o  Xk Xx X� m�  o  M� � � j�lA     �z 9U�U#�9T	0�@     9Q0     tBZ pwA     b       ��u KTZ �� y� KaZ � � XnZ M{Z �� �� X�Z X�Z ^BZ �r  ^u KaZ � � KTZ ]� W� O�r  MnZ �� �� X{Z M�Z �� �� M�Z �� �� ;�wA     �z Du 9T	�1H      v�wA     9U�U9T�T   8�wA     �z 9U	@AH     9Tv   t=_ �wA     ~       ��v KN_ (� � KZ_ �� �� Kf_ � �� Kr_ �� }� w~_  M�_ �� �� m=_  s  KZ_ }� {� Kr_ �� �� Kf_ �� �� KN_ {� q� O s  X~_ X�_ m�_  s  M�_ �� �� ]�_ xA            kv M�_ q� o�  n�_ PxA            M�_ �� �� 8\xA     �z 9U�Q9T09Q:      t��  `xA     R       �w K��  �� �� K��  =� 9� W�  W�  Z�  �P8}xA     �z 9Uw   t��  �xA     �       ��x K��  �� v� K�  � � K�  �� �� K�  C� ;� M)�  �� �� M4�  Q� E� M?�  �� �� MJ�  � � MV�  ?� /� Mb�  ]� Q� N��  yA      @s  �,x K�  �� �� K�  z� p� K��  �� �� K��  Z� P� O@s  X�  8UyA     �v 9Q�R9R�R#d�  �R   n��  (yA            K�  �� �� K�  � � K�  A� =� K��  {� w� L(yA            X)�  X4�  X?�  XJ�  XV�  Xb�     x?  ?  �y�6  �6  &�x�3  �3  �xxL  xL  �yg?  g?  Tx5<  5<  ?yF\  F\  &�x�J  �J  �y�+  �+  '(xRH  RH  �xiD  iD  �x�*  �*  �x�H  �H  �zBi  8i  ( xF  F  mx!,  !,  Ux9  9  cxjO  jO  x�=  �=  y�Z �Z 'x@:  @:  uy�K  �K  &vz�D  �D  ( x�N  �N  �x>Q  >Q  �x _   _  hx?U  ?U  �x�F  �F  �x�9  �9  )y�,  �,  *�xcL  cL  *yC  C  `x�-  �-  *BxE1  E1  ry],  ],  eyo+  o+  �y�]  �]  )^y�H  �H  )ox�X  �X  XyaG  aG  �xP  P  �x�=  �=  �y7  7  )�x�R  �R  x�*  �*  [y�\  �\  +.x02  02  7 V�   �  �  ��  $"  @�A     p^      	� X  ^� 	�@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  .�  
�5  -  �[  
�H  �  	H  >   
G   �	  
	N   �  B"z  �     ��  R   �U    �� ��  �N ��  �6  �
   �  Y�  �  U   �  n  -      n�  �  
  n  U    �  �    U   :  n  -   -   U    �  �"F  L  �   PJ�  2�  LI   �  M@   pos N@   �  P  SF  Q   �1 R  (=9 SV  0R�  Un  8y�  VI  @�� WI  H �  �  �\ �-   m  �U    o  ��  �  �%  +  @   I  :  @   I  @    O  �  2  c  i  t  :     :-   �  J�  x Lt   y Mt   )  O�  	�  B   s�  M   ut   }  ut  V  vt  /  vt   t
  x�  k	  (�  �  N    ��  N   �  	G   B� 
I  L  H    O  s  O  v	  U     �    	�  �  (N�  �  P5   Z�  Q5  �  S�  s  T�   [  U�  ?1  WG     �  5    Y�  �  =  N   �T  �   M
  pmoc5  stib	  ltuo|  tolp 	  �  b   "n  t  �  %  <�  x >5   len ?H  *� @O   %  By  	�    `�  �  �  G   G   �  U    �  �  q    G   !  G   G   U    �  .  4  I  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  �!  0R   �U   8�  ��  @ �  �  �  �I  	�  �       G     U      a  �  /  5  @  a   �  ?M  S  h  a  I  @    �  Yu  {  G   �  a  @   U    s  ��  �  G   �  a  �   �  W  0�$  �  �T   e� ��  �� �@  �� �h  �� ��   �� �"  ( �'  ��  �!  lO  �  �I  �  -  �O  	P  \  �L  �a  �  ��   	s  �
  �5  �  �H  �  �G   
  �N   	�  �  �-   \#  �@   �   -   �  ,G   \&  7U   �0  D4   b   �H	  xx ��   xy ��  yx ��  yy ��   a  �	  	H	  z'  ��	  m  �a   ss  ��   �  �Z	    ��	  �	  �	  U    �  ��	  �U  �U      ��	   %  ��	  �  $�	  �	  �   4
  �� "�	   �@ #�	  �U  $U    �  7_
  �; 9�	   ��  :�	   L  <4
  N   #��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=.  ��  ?t   �  @t  ~  Bt  �  Ct  �  Dt   5  Ft  (B  Gt  0�  Ht  8 �	  J�  
   s�  �  u�   ��  v�  �  xt  �
  zt  (  {t   �  };  �  �#�  �  k  `�_  R�  �n   (  ��  |  ��  �  ��  �  ��  �  �C$  v  �_
  �  �  (�%  �_  07&  �S$  8G   ��  X �  �"l  r  h  �  �M $   k  �  R�  n   �  �"�  �  %  8;  �� =#$   �M >�    ?_
   r$  @�  0 5  �$    %  ��  �� #$   �M 0$  �  T   �    (�� 
a  h�� �  p�� �  x K  � �  �  �  �,]  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9�  8  :�  @�  <�  H�  =�  PE-  ?�	  X�!  D�  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R]  ��� S  �K1 W�  �R�  Xn  �Jy  Y:  �%  [_
  ��	  ]�	  �    ^U   ��8  `M  � L   j  p    X��  �  ��   E-  ��	  N ��  �8  ��  P �  *%�  �  �  0t  k  v�   �  w�  �@ x�  ݖ y�  E-  z�	   N |.  0�  }�  pR  ~�  x�  �  �ߣ  �T  ��I ��  ��  ��  �h  ��  ��S  �  �4  ��  �8  ��  �  �U    �  �-   �  �t  o  �t  �L �U    �8  �E  ( �
  L#!  '  W  Hn  �  J�   = K3    L�  d  M�   �  N   �3  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  n  (0  O'  #   g)Z  `  �   ���  =  �H	   L  ��   $  ��  0�  �Y   8m  �#�!  h�  �=  pآ  �T  tG   ��  x s  �    �?  d�  �
  �)    �   H�J  �  �U    "  ��  �!  ��   ~	  8f�  �
  h�   (  i�  �� k�  �� l�    nt  �  ot   �  pt  (�  qt  0 y  sJ  �a  �p    �$�  �  �  0'E  �N  )�   ?1  *�  }0  +�  i/  ,�  � -H	   �  �)R  X     H��  ��  ��   ?1  ��  (  �1  4  �H	  \  ��  0  �U   @ ��  ��  +!  �  tag �   �U  �   �  �  �  `  N   
>  w%   }#  �&  h  �  &     
  E   9
�  � ;
>   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  K  �  N   ��  :   �   ^$  1  �!  �!   :  ��  �  ��  �#  �    �  %  _   I$  �1  7  B  _   �&  �N  T  �  h  _  h   �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  �  0�   �%  8��  �B  @   R  �n  x  =�	  H  E#!  	  �  @J�  �  L�   �  MT  �� O�  .� P  �  Q�   �  R4  (�!  Sa  08'  T�  8   W!�  �  -  (l�  k  n�   �M o�  ߣ  pT  �  q�     k  )�    �    �  �   w   .#  )  4  �   �  1@  F  [  �  [     U	  K  6m  s  �  �  �   �  �  :�  �  �  �  �  �   �  >�  "  Y�  �  �  �    �  �     �  _�  �  �      �  [     $  f'  -  B    �  �   �  lN  T  �  m    �  �   #  x��  �� � �   �  � T  H  � �  P�  � �  X9!  �   `l� � B  h  � �  p $    �m  P  �  @    �  H2G  �S  4   �  5�  (  6�  04  7�  88  8�  @ �  :�  �  �=�  R�  ?n   �  @�  n  A�  �  B�  1$  C1  2�  EG  �� FG  `�L HU   � �  J�  S  P   �  �  �    :  �  �  �      �  &  "  -  �   �%  *9  ?  �  N  ]   �%  -Z  `  k  ]   {  1w  }  �  �  �   �  4�  �  �  �   l  8�  �  �  �  ]  �   �  <�  �  �  �  ]  �   �  @    �  %  �  ]  �  T   �  G1  7  �  U  �  �  �  �   �'  Na  g  �  {  �  :   �  S�  �  �  �  �  �  �  T  �   �  &  ���  �� ��   i'  ��  H   ��  P  ��  X�A ��  `Y �  h�#  �-  p�  �N  x�  �k  �  ��  ���  ��  �U�  �%  ��!  �U  ���  �{  ��  ��  �&  ��  �   ��  	�  �&  ��  �  U   �>  ��  'O  �h   xC  ��   s/  ��  	�  �  0tY   �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�  �  U'r   x   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {}   �  ��   �   �  �   f   �  �    �	  �  �!  !  !  f   �    �'  �*!  0!  �  N!  f   �  1  N!   �   �!  �!  ��  )�    ��  )�   �  )!   }  T!  	�!  O  ;�!  _� =%�!   ݰ  >%f    �!  �  @�!  �!  cA  �,�!  �!  /  �"  �� �@   �M �"   ?<  �,)"  �"  �5  P��"  �  ��   �� ��"  �Y ��"  �H �#  U@ �9#   �9 �#e#  (�A  �#�#  0�^  �#�#  8�^  �#�#  @N7  �#$  H 	/"  ��  ��!  (Z  ��"  �"  �  �"  �!  �   17  �#  #  #  �!   �G  �#  %#  �  9#  �!  a   %G  �E#  K#  �  _#  �!  _#   a  �@  �q#  w#  �  �#  �!  �!  a  a   �;  ��#  �#  1  �#  �!  a  a   �W  ��#  �#  _#  �#  �!  n   *;  ��#  �#  _#  $  �!  n  a   �T  ��#  �  �  r  �  -1  B�  _  S$  @      c$  @    i$  h  x$  �   ~$  �  �$  �  �  �  �   �$  �  �$  �  �   �  �%$  �  8YF%  ��  [�   Ǧ  \�  ��  ]�  d> ^�  ��  _�   I�  `�  (�  a1  0U  b�  2�  c�  4 ��  e�$  ��  p$^%  �$  ��  ���&  ֤  ��   Ğ  ��  ��  �P  �  �P  	��  �P  
�  �P  ��  ��&  �  ��&  (��  ��&  <�  ��&  X��  ��  p��  ��  x��  ��  |��  ��&  ��  ��&  �R�  �P  ���  �P  ���  �1  �F�  �1  �V�  ��&  ���  ��&  ���  ��  �"�  ��  ��  ��  �@�  ��&  � �  �&  @    �  �&  @   	 �  �&  @     �  �&  @    �  '  @    ��  �d%  o�  �#'  d%  �  �'  ��  j'  2]   P   U�  !j'  5�  "�   �  �  $1'  ʭ  $�'  1'  ��   *^(  m�  ,�   `h  -�  �  /^(  #�  0n(  (��  1~(  ��  3�  z�  4�  ��  6�(  ��  7�(  ��  9�  (Ԯ  ;�(  0��  C�(  ���  D�  � �  n(  @    �  ~(  @    p'  �(  @    R%  �(  @    '  �(  @    �  �(  @    �  �(  @    3�  F�'  ��  F�(  �'  �  N   0 )  ��   r�  �  E�  Ϊ   H�  8�(  �  N   w[*  U�   ��  ��  �  ��  ��  ޟ  $�  ��  �  	t�  
�  ܖ  �  ��  ��  d�  {�  ך  ʕ  �  ��  ��  m�  ,�  �  ^�  ׭  ~�  @�  �  ��  N�   ��  !��  "��  #ݴ  $��  %�  &�  ',�  (a�  )��  *x�  +��  ,"�  -"�  - a�  �-)  ��  )$t*  z*  H�  ��  ,�*  �*  �  �*  n  �*  �*   %'  h*  ��  1�*  �*  �*  h*  �  �  �  �   ��  8�*  �*  +  h*   �  ;9+  M� =*   �� >�*  Յ ?�*   ��  AE+  +  �  h!W+  ]+  ��  ��  u-n+  �+  ��  8V�+    XK+   j�  Y�+  =9 Z\,  �� [,  Q� \.,   �� ]:,  (�� ^�,  0 	t+  ��  ��+  �+  ,  K+   ��  �,  ,  .,  K+  �  �   K�  �,  å  �F,  L,  \,  K+  �   ��  
i,  o,  �  �,  K+  �   ?�  1�,  �,  �  �,  K+  �,  h*  �     1�  �!�,  �,  $�  ��  �-�,  V-  .�  8�V-    ��,   j�  �[-  =9 ��-  �� �y-  +�  ��-   �� ��-  (�� �".  0 	�,  ǡ  �h-  n-  y-  �,   ��  ��-  �-  �-  �,  �  �  �   ��  ��-  �-  �-  �,  �  �  a   !�  &�-  �-  �-  �,  �  a   K�  D.  .  �  ".  �,  �   	�  k/.  5.  �  S.  �,  �,  h*  �   ��  ��.  ��  ��.   X� ��.  l� ��.   9+  �.  _   �.  b+  �.  _   �.  �,  �.  _   �.  $�  �S.  �  � �.  �.  �3  5/   num 7�   str 8h   +P  :�.  �J  =E/  key ?/   �U  @4    �7  D$Q/  /  O  Hc/  i/  �  x/  x/   /  �Z  K�/  �/  1  �/  x/  x/   �S  (O 0  �� Q�   �  R�  �6 S�  �B  UW/  3  V~/  >) X 0    E/  e-  \ 0  �/  ��  #$0  *0  a  90  h   d�  )E0  K0  h  Z0  �   0�  /E0  K�  6�0  �> 8a   �^ 9�   �  ;f0  Ѽ  >$�0  �0  ў  (@�0  
H B�"   ��  C�  XT D�0    �0  ��  N�0  �0  h  1  �  �   B�  V1  1  /1  �  h   ��  Z;1  A1  �  i1  n  �0  �  �0  1  �   ��  bu1  {1  �  �1  �0  a   ��  f�1  �1  a  �1  �0  _#   ��  @j+2  �\ l 0   8` n /1  �\ o i1  �_ p �1  �T r 90   }�  s Z0  (ʬ  t B2  0�  u B2  8 	�1  ��  j<2  +2  O  7�   F�2  ~�  H�   ̰  I�  V�  J�  �H L�2  �  M�2   �  �  b�  OH2  �  O�2  H2  ��  W�2  ��  Y�    ��  [�2  !�  ^D4  �  `F%   8�  a�2  8-�  b'  @"�  c�   "E�  e )  ("= f�2  0"�  hD4  P"
�  iD4  X"��  jD4  `"��  l�  h"��  mJ4  p"h�  nP4  x"��  o0  �"�  q�  �"V r�2  �"� sJ4  �"'�  tP4  �"��  vP  �"�  wP  �"��  xH	  �"w�  y�  �";�  z�  �"* {�   "ܲ  }�   P  D4  �  �  �2  �  n4  �2  ��  (��4  �9  ��   ��  ��  ɲ  ��  �  ��  �  ��    T�  ��4  t4  ��  �5  ��  ��   ��  ��  x ��  y ��   �  �5  �4  z�  X��5  ��  �1   ��  ��  �Z  ��  (%?  ��  0L�  ��4  8)�  ��  @W�  �5  HѺ  ��  P b�  ��5  %5  �  �!�5  �5  !6�  x��6  �� ��   �6  �V4  �"s  ��  "Q  ��  "Y�  ��  "B�  ��6   "�  ��6  @"�  ��(  P"�  ��  X"�  ��  \"�  ��  `"�  �j'  h"2�  ��  p @  �6  @      �6  @    x�  ��5  �  - �6  �6  W�  XZ�6  �� \�    �  8%�6  �6  !u�  Pt]7  �� v�   "�� x1  0"��  y1  1"�� {�  8"�� |�  @"�  ~�  H"n  �  L �6  `SH8  �<  U�   �Q  V�  a(  X�  VA  Y�  Q) [�   nX  \�  "�D  ^H8  (�5  _H8  8M   a�  H}  b�  JV  c�  L/  d�  N7K  f�  P>D  g�  R�:  i�  T�3  j�  V=]  k�  X �  X8  @    �5  m]7  �Q  8�B9  �  ��   �Z  ��  %?  ��  
L/  ��  �<  ��  �Y  ��  �7  ��  �)  ��  �O  ��  �H  ��  vH  ��  ^  �B9  �>  ��  $�7  ��  &0>  �U   (�+  �U   0 �  R9  @    �H  �d8  �?  8AM:  �  C�   �Z  D�  %?  E�  
L/  F�  S.  H�  �W  J�  �W  K�  C  L�  �O  M�  �H  N�  vH  O�  ^  QB9  �>  S�  $�B  T�  &0>  ZU   (�+  [U   0 �]  ]^9  �B  �|�<  ��  ~�   �)  �  �)  ��  �.  ��  U  ��  �V  ��  
�0  ��  �6  ��  �C  ��  U?  ��  6P  ��  �C  ��  &L  ��  *J  ��  �L  ��  HP  ��  N*  ��<   [2  ��  0k2  ��  8.  ��  @{2  ��  HQ2  ��<  P�0  ��  Tp4  ��  VmU  ��  X�Z  ��  Z ?  ��  \:  ��  ^�I  ��  `E8  ��  b�;  ��  h�;  ��  p�O  ��  xDF  ��  zfV  ��  |�9  ��  ~[9  ��  ��G  ��  �zQ  ��  � P  �<  @   	 =  �<  @    {D  �Z:  �1  @�E=  �I  ��   6Y  ��  �^  ��  S  ��  )  ��  @3  ��   �0  ��  (4C  ��  0�C  ��  8 aM  ��<  �I  @�3>  �  ��   _7  ��  )  ��  �O  ��  �n ��  �T  ��  EF  ��  I  ��  �K  �3>  N:  �C>  ,L  �S>  4�E  �=  :�Z  �=  ;�Z  �P  <^  �P  = =  C>  @    =  S>  @    =  c>  @    eU  �R=  �9  (7Q?  ��  9�   a@  :�  b<  ;�  
8  <�  .  =�  �H  >�  �Q  ?�  X  @�  �.  A�  �;  B�  ))  C�  eH  D�  I_  E�  �B  F�   !3  G�  " �)  Ip>  �  I�?  F@ K�   I�  L�  K�  M�   ԃ  O^?  �b  hh�?  `h  j�   m�  k�  dh  l�?   �?  �?  @    ��  n�?  �j  0�L@  F@ ��   I�  ��  def ��  K�  ��  tag ��   c  ��  ( )�  ��?  �  ��@  �  ��   c  ��  Cg  ��   �~  �X@  z�   ��@  `h  ��   m�  ��  L�  ��  dh  ��@  e  ��@   L@  �@  J�  ��@  �R   FBA  tag H�   ��  I�  .� J�  �P  KBA   �  DG  M A  f3   ��A  Tag ��   Q  ��  .*  ��  �K  ��   gW  ��A  TA  �^   B  k@  �   aE  �  p0  �  �>  �  H  �  �/  �  �� D4   �F  �A  �<  0_B  H  2�   �/  3�  �� 8D4   qS  :&B  A9  0U�B  ߣ  W�   �E  X�  �^  Y�  =Y Z�B  <  [�  �=  \�B   Jy  ]:  ( B  _B  rY  _lB  �1  ~!C  �.  ��   �L  ��   Z  �.C  �B  �V  �mC  ��  ��   f>  ��  Y  �!C   �)  �4C  �A  /#D    1=   �  2=  �N  3P  o=  4=  D4  5=  �^  6=  `*  7=  �0  8=  �G  9=  �D  :=  	I:  ;#D  
 =  3D  @    �@  =zC  �\  ��D  +  �3D   Y�  �3D  �
  �P  (  �P  �F  �P  �C  �P   <)  ��D  @D  �,  �D  �  �   AK  �  z8  �2  V �D   E  =  �R  �D  	F  .AE  �  0�   �P  1E   ">  3E  #IsE  $�K K	E  $`B LAE   �[   E�E  �z  G1   =Y NNE   �6  PsE  O]  a!�E  �E  �(  7N  (�&F  >) �D4   -N  �D4  V` �D4  TE  ��  �/  ��   �z  �1  $ G  ��E  &8  � @F  FF  eS  po�J  �� q�   ^  sHA  ��^  u�  [>  v�   �W  w�A  (� yX8  0�=  zR9  ��,  |Q?  ���  ~1  ��(  M:  �AK  ��  0XL  ��B  8%os2 ��<  hp�  �E=  �T  �D4  0#9  ��  8!H ��L  @�+  ��L  H@.  �M  P�E  ��L  X�P  ��L  `@  ��L  h$S  �U   ps  �U   x%mm �U   �%var �U   �Q  �U   �<B �mC  �2Y �c>  �=  ��  �=  ��D  �UV  ��E  ��(  ��  =  �D4   /:  ��  (�?  �D4  0�]  ��  8%cvt �aM  @�R  ��J  H5$  ��	  P��  �h  `HT  ��  h�*  ��  p�J  �1  x�+  �1  y�  ��E  ��C  �a  ��-  �h  �j7  ��  �kN  ��  ��F  ��  �#7  ��  ��(  �D4  �rE  �D4  �QZ  ��  �4  ��  ��@  ��  �:L  �D4  ��G  �D4  ��]  ��  ��W  �TM  ��/  ��  ��B   P4   �I  D4  s-  �  �*  �  ,  a  ,  a   %bdf 	&F  (�T  �  P#F  �  X�U  �  `�K  �  h �=  ��J  �J  �  �J  U    �Q  �"�J  �J  �\  xc�L  �  e3F   �  f5N  )�  g�  �V  h�  :1  j�   �^ k�  (Jy  m:  0�  n�  8�  p�  <�!  q�  @R0  r�  `�  s�  duN t�  h6  u1  lpp1 v�  ppp2 w�  �2�  zN  �Xc  {N  ��6  }N  )  ~D4  �8  �   �L �U   (C  ��  0��  ��  4%pp3 ��  8%pp4 ��  Hy�  �D4  X�� �D4  `U  �_
  h �I  ��L  �L  �  �L  3F  �  :  BA    1  �L  �L  �  �L  �J  �  �  �   �M  +�L  �L  �  M  �J   �<  :M  M  "M  �J   y*  N   =TM  4   �^  J  b8  �T   lK  H"M  �  |T  @?N  R�  An   �  B�  n  C�  
Z�  D�  �  E�  org G�  cur H�  ��  I�   s  KD4  ([  L�2  0c+  N�  8 R8  PgM  RG  T'*N  0N  [  O  _ BN  HN  LL  ͳ  @ @�N  Jy   B:   �S  C�  ܱ   D�  .�  E�  ��   FP  ��   G�   
�   H�  (�P   JBA  0Ӏ  KD4  8 ,�   MMN  !
�   P-O  ߣ   R�   x   S�  .�  U�  ē   V-O  " �  W-O   �  =O  @   � ��   Y�N  ��  ( \�O  ߣ   _�   x   `�  ē   b�2  ��   c�2  Ӷ   e�   �   f�  $ r�   hIO  W�   m�O  Kw   t�   7�   uP4   0�   w�O  j�   {P  ��   }�   �   ~�  �w   �   J�   ��O  1�   �AP  �{   �AP    P  �   �&P  �    ��P  ��   ��   k   ��P  �q   ��   q   ��  y|   ��P   �O  GP  �   �SP  %�   �!�P  �P  �  � MS  k   O�   Jy   P:  R�   Qn  ��   R�  �    S�   �   T�  $(   VP  (|   WP  )x�   XP  *п   Z�  ,�J   \1  0i�   ^�N  8�   _�N  xC�   `�N  �=  b=O  ���   c�O  p�   e�N  8��   f�N  x=�   g�N  ���   h�N  ��   j�  8��   mJ4  @V�   p�  HV`  qJ4  P��   rD4  X��   s�  `/�   uY  h��   v�  0��   wY  8j�   y�X  82�   |�.  Xs   02  `��   ��  h�   �%Y  pd�   ��  x|�   ��  �˽   ��	  �ʞ   ��P  �8�   �+Y  � ֥  0 ��S  ��   �1   �   �1  v�   ��P  �   ��  ݺ   ��  ��   ��  c�   ��   BV  ��S  ( T  �   �S  !��  H ��U  ��   ��   Ǧ   ��  @�   ��  ��   ��  d>  ��  ��   ��  �   �1  I�   ��   U   ��  (�   ��  0��   ��  8�&  ��  <��   �H	  @?�   �1  `U�   ��  hw�   ��  p֤   ��  �;�   ��  �ܲ   �t  �w�   ��  ���   ��  ��   ��  ���   ��  �ٛ   ��  ��   ��  �g�   ��  �`�   ��  �x�   ��  ��   ��  �|�   ��  �"��   ��   "�   ��  "n�   ��  "��   ��  "��   ��   "`�   ��  ("�   ��  0"m�   ��  4"�m   ��  6"A�   ��  8"��   ��  @ ��   ��S  S�   �$�U  �U  ��  � *�V  Ҳ   ,�U   -�   -}X  H�   0�S   ݺ   1�  P%NDV  2�  X�   <D4  `K�   =D4  h�   >�  p��   ?�  t��   A�N  xZ�   BJ4  �l�   Ea  � !E�  � �MX  ��   �P   �   �P  ��   �P  �   �P  ��   �MX  �   �]X  x��   �MX  �"�   �]X  8"��   ��  �"��   �t  �"��   �t  �"��   �t  ��    t  �R�   P  ���   P  �V�   mX  ���   mX   ��   1  �6�   �  �Ğ   �  �"�   	�  ���   
�  �Т   �  �P�   �  �W�   t  ���   t  ���   �  ���   �U  � t  ]X  @    t  mX  @   	 t  }X  @    ��   �V  a�    �X  ߣ   P   �   �  �U   D4  
�   �  w�   !�  .�   "�  �   #P   �   %�X  9�   G�U  �U  %Y  @   � F%  �2  8�  `!,YY  �� !.�   -U !/�  X `�  !1eY  1Y  !~�  H!<�Y  �� !>�   "�� !@1  0"��  !A1  1"�� !C�  8"�� !D�  @ Z�  !F�Y  kY  �C  h"* Z  �� ",6$   �Z  ".�  8�  "/1  <X;  "0 Z  @آ  "1T  ` �  0Z  @    �D  "3<Z  �Y  ��  "?-NZ  TZ  ۳  `"��Z  ��  "�D4   y�  "��  �� "��  �� "��  ��  "��   Ǩ  "��  $(2 "�J4  (Ϛ  "�P4  0R�  "�n  8_� "�z[  @ ��   "T&[  �� "W?[   �Y "\P[  add "_t[  �x "eP[   �  ?[  BZ  �  n   &[  P[  BZ   E[  �  t[  BZ  �  U   �   V[  r�  "g�Z  	z[  �  "�TZ  �  "�"�[  �[  ��  �"�\  y�  "�D4   2�  "�D4  �� "�D4  � "��  R�  "�n   _� "�/`  ( ��  "�"\  \  ��  "�S\  �S "�D4   �� "�D4  � "�%]   ��  "�"d\  	S\  j\  ��  0"��\  9�  "�h   �{  "��]  � "��]  ��  "�^  x  "��  �  "�P  m�  "��   �  "��  $��  "�  ( &��  N   "�%]  ˟   .�  ��  ��  ��  ��   ��  "��\  ��  "�\  &L�  N   "��]  ��   ��  Ʊ  ��  ��  g�  �  ��  W�  �  	|�  
K�  ��   8�  "�=]  &��  N   "��]  c�   ��  p�  �  �  ��  �  ��  ��  }�  	 ��  "��]  ��  "�^  ^  '^  �  �   [�  "j\  	'^  �  h"k�^  �� "n_   �Y "t)_  �? "w)_  �2 "y)_  �! "|>_   �$ "~X_  (�* "��_  0�3 "��_  8k! "��_  @�A "��_  HV- "� `  P�F "�)`  X  "�)`  ` _  �[  D4  D4  n   �^  )_  �[   _  �  >_  �[   /_  �  X_  �[  �   D_  �  �_  �[  D4  �  BA  1   ^_  �  �_  �[  �  aM   �_  �  �_  �[  �  �  �   �_  �_  �[  \   �_  �_  �[  \  �  �_   �  �_  �  )`  �[  _\  �  �  BA   `  �  "�9^  	/`  �  "��[  ~�  "�[`  l�  p"Xa  R�  "n   �  "�  )�  "�Y  ��  "�  2�  "�,   �� "�,  (��  "�a  0��  "�a  8R0  " �  @�  "!�  H�!  "#�  P��  "$1  X�� "%1  Yb�  "&1  Z��  "(1  [�  ")1  \_� "+�a  ` ګ  "��a  �� "��a   �Y "��a   �a  �a  U   1   N`  �a  �a  �a   �a  �  "�Xa  t  î  "Bb  2�  "DD4   �� "ED4  y�  "FD4   {�  "H�a  ��  "Lb  !b  �  ?b  3F  �  J4  BA   l�  "RLb  Rb  gb  3F  J4  �   ��  �"W�d  <0 "YN`   4� "[�d  p%top "\�  �O� "^�d   Xc  "_�d  ���  "a�  ��  "b�  ��  "c�d  �%cff "e�P  �  "f�U   ˽  "g�d  (
�  "i�a  0�  "j1  8��  "k�  <z�  "m�  @�  "n�  D��  "p�  H�  "q�  L~�  "sJ4  P9� "tJ4  XV "vJ4  `�  "w�  h&  "y�  l�J "{1  p�  "}&b  x��  "~&?b  �s  "�02  �Ğ  "��  ���  "�P4  �q�  "�0  ���  "�H	  �w�  "��  ��  "��(  ��  "�j'  ��  "��  � �  �d  @   0 b  �d  @    b  �  �d  @    �	  x�  "�gb  ջ  "�#�d  �d  �  �"�e  R�  "n   �  "�  )�  "�  ��  "�  2�  "�,   �� "�,  (��  "t  0��  "t  8R0  "�  @�  "�  P�!  "�  `��  "�g  ��� "1  �b�  "1  ���  " 1  ��  ""U   �L�  "#U   �_� "%Zg  � ��  "��e  �e  �  f  �d  �   q�  "�f  #f  =f  �d  t  t  P   j�  "�Jf  Pf  �  if  �d  t  t   ��  "�vf  |f  �  �f  �d   *�  "�Jf  �  "��f  �f  �f  �d   �  @"�5g  �� "�Tg   �Y "��f  �? "�$�e  kI "�$f  rL "�$=f   � "�$if  (-1 "�$�f  0��  "�$�f  8 Tg  �d  �  ]  �  1   5g  T�  "��f  	Zg  a�  N   "��g  ��   J�  �  ,�   ה  "�lg  ��  "'�d   �  "F�g  y�  "HD4   2�  "ID4  �� "JD4   ɠ  "L�g  ݬ  "Lh  �g  �  "O/h  h  ��  �"}�i  <0 "�g   4� "��j  �%top "�j'  �O� "��j  �Xc  "��g  x
s  "�02  �
�  "��  �
V "�J4  �
Ğ  "��  �
��  "��  �
��  "�J4  �
h�  "�P4  �
��  "�0  �
��  "�H	  �
w�  "��  �
��  "��  �
�  "��  �
�  "��d  �
�  "��(  `&  "��  h�  "�j  p_� "��j  x�  "�j'  ��  "��  ��J "�1  �˽  "��	  � ��  "P/�i  	�i  j  �   "Xj  �� "[tj   �Y "f�j  �; "o�j  � "u�j   	�i  �  "T#j  )j  �  =j  h  �   �  tj  h  �  ]  �  J4  �(  1  �  j   =j  �j  h   zj  �  �j  h  D4  �   �j  �  �j  �j  D4  �   �d  �j  X�  "z�i  	�j  �  �j  @   � �g  k  @    �  "�h  <�  "� k  ��  �"&l  R�  "n   �  "3F  )�  "�Y  ��  "�  2�  "�,   �� "�,  (��  "t  0��  "t  8R0  "�  @�  " �  P�!  ""�  `��  "$1  ��� "%1  �b�  "&1  ���  "(1  ��  "*U   �L�  "+U   �_� "-�m  � c�  "�3l  9l  �  Ml  Ml  �   k  ˯  "�`l  fl  �l  Ml  t  t  P   N�  "��l  �l  �  �l  Ml  t  t   Ԝ  "��l  h�  "��l  �l  �l  Ml   8�  "��l  �l  �  �l  Ml   p�  @"�xm  �� "��m   �Y "��l  �? "�%&l  kI "�%Sl  rL "�%�l   � "�%�l  (-1 "�%�l  0��  "�%�l  8 �m  Ml  3F  YY  �Y  1   xm  +�  "��l  !�  "E�m  2�  "GD4   �� "HD4  y�  "ID4   ��  "K�m  j�  �"N�o  <0 "Pk   cff "Q�P  �4� "S�d  �%top "T�  hO� "V�o  pXc  "W�o  ��  "Y�  �  "Z�  �  "[�d  
�  "]t  ���  "^t  ���  "`1  ��  "a1  ���  "b�  ��  "c�o  �z�  "e�  ��  "f�  ���  "h�  ��  "i�  �~�  "kJ4  �9� "lJ4  �V "nJ4  ��  "o�  �&  "q�  ��J "s1  ��  "u�U  ��  "w&b  ���  "x&?b  � �m  �o  @    �m  �  �o  @    1�  "z�m  l�  "p  �� "�Ap   >'  "�`p  � "��j   ;p  ;p  3F  YY  �Y  1  �  b  ?b   �o  p  �  `p  ;p  YY  �   Gp  U�  "��o  	fp  :�  "�#�p  �p  ,�  ("��p  R�  "�n   Jy  "�uq  � "��5  p�  "��q  o�  "�U     4�  "�q  �� "�7q   �Y "�Hq  gP "�]q   �  7q  xp  n  D4  D4   q  Hq  xp   =q  �  ]q  xp   Nq  \�  "��p  	cq  ١  "�#�q  �q  ��  �  �q  h  �  U    �q  C�  "��p  �  "�.�q  r  0�   "�r  ��  "�"   �0 "�"  ک  "�"  �> "�"   	�q  �  X"��r  b�  "!�r   �  "!�r  E�  "!�r  b�  "!�r  ,�  "�r   h�  "s  (�  "s  0��  "9s  8c�  "�q  @:�  "!?s  Hs�  ""Es  P �[  <`  gg  �j  �r  D4  �  �   �r  a  s  a   �r  s  �j  U   1   	s  9s  �  '  �U   $s  pq  sp  ��  "Xs  r  N   #��u  +�   ��  ʵ  ݒ  �  b�  ��  ׾  �  ݘ  	7�  
=�  ��  I�  p�  �  ��  ��  ɓ  Q�  ��  4�   R�  !�  "�  #ŧ  $�  %��  &�  '�  (V�  0ݕ  1��  @��  A��  Qt�  R  SO�  T��  Uݼ  V��  W�  Xn�  `�  aͷ  b�  c��  pV�  ��  �Φ  ��  �X�  ���  ���  �ɴ  �(�  ���  �^�  �i�  �Z�  �ĸ  �7�  �F�  �۹  �B�  �;�  �c�  �A�  �S�  ���  �Ѩ  ��  �E�  �ř  �k�  ���  ��  ���  ���  �/�  �.�  �!�  � �  ���  �=�  ���  �"�  ��  ���  ���  ��  �i�  �6�  ���  � 
;  $".�  ��  �%=0v  �� %?A`   Jy  %@:  ���  %BD4  ���  %C�  �-�  %ED4  �Ȝ  %F�  ��  %H1  �O�  %I1  ���  %J1  � �  %L�u  ��  %LHv  �u  !I�  �&"w  �  &$0v   ~�  &&�  ���  &'�[  �"�  &*�  ("V &+�[  0"� &,�[  �"V�  &-�[  �"��  &/�  P"��  &0�[  X"��  &10  �"��  &21  �"B�  &4�  � ܠ  &6Nv  �  &6w  Nv  ��  '',w  2w  �  Fw  �  Fw   �?  jd  '+Xw  ^w  �  rw  �  rw   xw  �@  �g  '/�w  �w  �  �w  �  �  j'   �{  '6�w  �w  �  �w  �  �  �    l  '=�w  �n  'B�w  �x  'G�w  �w  �  x  �  �   1j  'K�w  �}  'P*x  0x  �  Sx  �  P4  Sx  Sx  rw   �  ��  'W  ��  'Zvx  	ex  �b  P'Zy  h  '\ w   �v  ']~w  ��  '^�w  ��  '_x  .�  '`Lw   �  'a�w  (V�  'b�w  0��  'c�w  88�  'fx  @��  'gYx  H f.  (&x$  <B  (,�$  %�  (0/y  	y  �3  (0Wy  tW (2!y   i�  (3!y   FO  ))c$  ��  ),ty  	cy  Y  ),�y  6 ).Wy    =�  *!�y  �y  �  �y  �  %Y   T�  *%�y  �y  �  �y  �  +Y   ��  *)�y  �y  �  �y  �   �  *,z  z  �  "z  �  "z   '  ��  *04z  :z  �  ]z  �  [*  �  U   �   �  *7nz  	]z  ,�  (*7�z  ۽  *9�y   1�  *:�y  G�  *;�y  #�  *<�y  )�  *=(z    n)  +�z  �z  �  �z  _  h  �  1   �)  +$�z  �z  �  {  _  h  U    nk  +)){  	{  �;  +)Q{  �=  ++�z   z+ +,�z   �N  , ]{  c{  �  �{  �  �  �  �   /�  ,%�{  	�{  �I  ,%�{  �2  ,'Q{    '�  \)*y  	`QH     '�  o*oy  	PQH     '��  {,qx  	 QH     (E�  Z&iz  	�PH     (N�  e'�{  	�PH     ('�  q${  	�PH     �  D|  @    	4|  (�  }#D|  	 PH     )�u  �	`OH     4^  �|  @   . 	s|  (J�  ��|  	�FH     *a�  �  �}  +�  '<v  +Q  'Ks  ,Jy  :  ,R�  	n  ,� 
�  ,�  �  -�0  -��  U-�u  -�Y �.C}  ,��  �  /tag �   0/cur OD4  ,�� PD4  ,1�  Q�  ,Y�  R1  0/len ��     1�  ��}  2�  �"<v  3R�  �n   4?�  ��  ~  2�  �!<v  2Jy  �!:  2R�  �!n  2Q  �!Ks  3� ��  5tag ��  3�  ��  6�u  � 4ӣ  b�  �~  2Jy  b$:  2ϒ  c$h  2n�  d$4   3� f�  5tag g�  3��  h�  7�u  �tB      8�  F�  @�A     n       �U  9Jy  F:  �� �� 9��  G�2   � � 9�Y  HBA  �� � '� J�  �L:tag K�  �� �� ;�  L�  9� 5� <i�A     p�  :  =Uv =T�L >��A     }�  =Uv =T�L  ?z�  {p�A            ��  @K1 {_  U A
�  F�  ��A     x       ��  @~ F_  UBK1 H0Z  q� o� (ߢ  Ja  �t A��  -�  �B     �      ��  CJy  - :  �� �� C�  . �  �� �� C�  / �  �� �� CG  0 �  � � CG  1    R� N� B�  3�5  �� �� B� 4�  h� L� Bs  502  �� �� BQ  6Ks  #� � B�6  7b4  �� �� B��  8R%  �  �  D�u  2B     E��  K�  B~ A_  s o B�O  A�  � � >�B     ��  =T	�BH     =Q1  E�  ��  B�� j�  A 9 E@�  ��  Bs�  ��   � � Br? ��   J D F��  B�  �1  � �   F��  (�  �t  �@<OB     ��  �  =Us =Tw  G)B     ��    E�  ��  B�� ��  � � FP�  (�� �@  �@Bf�  ��q  $  B�M �"  } m <�B     ��  y�  =T0=Qw =R0 >B     ��  =T0=Qw =R0   <B     ��  ��  =T	�BH      <EB     ��  ׂ  =T	`BH      >TB     a�  =Us   H��  �p�A     Q      �i�  9�  ��  1 ) ;�  ��5  � � ;R�  �n  � � ;�6  �b4  "  E��  �  ;��  �R%  { w <��A     ��  ��  =Uv  <��A     ��  ��  =Uv  <�A     ��  ��  =Uv  <"�A     ��  ׃  =Uv  ><�A     ��  =Uv   <��A     ��  �  =Uv  <��A     ٫  �  =Us  <V�A     ��  4�  =Uv  <p�A     ��  L�  =Uv  <��A     ��  d�  =Uv  <��A     ��  |�  =Uv  <��A     ��  ��  =Uv  <��A     ��  ��  =Tv  <��A     ��  Ą  =Uv  <�A     ��  ܄  =Uv  <�A     ��  �  =Uv  <5�A     ��  �  =Uv  <O�A     ��  $�  =Uv  <i�A     ��  <�  =Uv  <��A     ��  T�  =Uv  >��A     ��  =Uv   IX�  ��  ��A     M       �3�  9 �$�  � � ;�  ��5    ;2�  ��.  _ ] J��A     .       ;~ �_  � � K��A            �  ;_� �b+  � �  >��A     ��  =T	`BH        Hȩ  ���A            �`�  L �$�  U 8��  u�   B     C       ��  9�  u%]  � � Mreq v%�  $  ;�  x�6  v p ;_� y9+  � � <2B     ��  �  N0�  s  <@B     ��  �  =T|  O\B     =R0=X0  8��  ]�  pB     H       ��  9�  ]]  	 � ;�  _�6  T	 N	 ;� `�  �	 �	 ;_� a9+  �	 �	 K�B     (       ԇ  '9� fh*  �h;�  g�5  
 
 O�B     =Q�h  >�B     ��  N0�  s   1ι  I�  2�  I]  3�  K�6  03_� P9+    4��  99+  a�  2�  9'�6  3�  ;�5  32�  <�.  3~ =_   A�  ��  �B           ���  C�  ��5  T
 :
 (��  �w  ��yB�   	<v  p j B�6  	b4  � � B��  	'  3  (� 	�  ��yBQ  	Ks  � v D�u  �	�B     E�  Q�  Pi F	�  I G >�B     ٫  =U~   KPB     @       ��  BR�  U	n  o m >kB     ��  =T8=Q0=X0=Y��y  E �  H�  B�j �	�  � � Pidx �	�  j b B��  �	 �  � � Bb�  �	*�  = 3 Bla �	D4  � � Fp�  B�  �	D4    >HB     ��  =U} =Tv    Q�  �B      ��  	~�  R�  � g R�  � �  Q�}  2B      �  	6�  R�}  � � R�}  � � R�}  = 3 R�}  � � F�  S�}  ��yS�}  ��yS~  ��yT~  >B     UCB     �  =Us =T0=Q0=R  <�B     ~  H�  =U| =T	�BH     =Q> <�B     ~  r�  =U| =T	�BH     =Q: <�B     �  ��  =U| =T0 <	B     �~  ��  =U| =T��y=Q}  <,B     �  ы  =U| =T0 <�B     ��  �  =U  <�B     �  �  =U =Q��y <�B     !�   �  =U|  >�B     .�  =U|    Q��  �B      ��  �	��  Rː  ) % F��  Vؐ  c _ V�  � � Q�}  }B      ��  ���  R�}  � � F��  V�}  � � <�B     ��  ό  =Uv  U�B     �  =Us  >XB     ��  =Uv    U�B     �  =Us� U�B     #�  =Us� UB     8�  =Us� U+B     M�  =Us� UAB     b�  =Us� <QB     ��  z�  =Tv  >aB     ��  =Uv    Q�|  UB       �  "	l�  R�|  > 2 R�|  > 2 R�|  � � F �  V�|  0 ( V�|  � � S�|  ��yS�|  ��yT�|  �B     W}  T}  �B     T}  QB     XC}  ��  j�  VD}    VQ}  � � V^}  k e Vk}  � � Yx}  �B     P       ��  Sy}  ��yO�B     =Us =R��y=X0  UB     Î  =Us  UB     ׎  =Us  UsB     �  =Us  <�B     ;�  �  =U} =T:=Q��y <�B     ;�  6�  =U} =T==Q| }  <�B     G�  N�  =T}  >�B     �  =U =Q��y  X#}  ��  Y�  V(}  � � S5}  ��y<�B     S�  ��  =U|  < B     .�  ��  =U|  <:B     �~  �  =U| =T} =Qv  <�B     �  �  =U| =T��y <�B     �   �  =U =Q��y <B     !�  8�  =U|  >(B     �~  =U| =T} =Q   O)B     =Q
q�   <IB     �  ��  =U~ =Ts  <�B     �  ��  =U~ =Ts  >�B     ٫  =U~   Z��  ��  +��  �w  ,�  �<v  ,R�  �n   Z��  ��  +��  �w  +�  ��5   [� �  @�A     �      �^�  C�  �5  2 . C��  w  z j C2�  D4  ) % C�  �  f b B�  <v  � � B�� D4  ` Z Bם  D4  � � Ba�  1  6 * D�u  �T�A     E �  M�  Pcur +D4  � � .2�  /s R�  /b SD4   K-�A     C       ��  \s _�  ��\b `D4  ��>X�A     �  =U =T��=Q��  Ep�  �  Plen l�  � � E��  �  B��  {S\  � � F��  BF@ �D4  m  i  EP�  Ó  B��  ��  �  �  ]B�  ��A      ��  �&Rn�  �! ~! Ra�  /" !" RT�  �" �" F��  V{�  # # S��  ��V��  �# h# V��  �$ �$ V��  �% �% T��  �A     U�A     ��  =U��=T  Of�A     =U =T~ =X0    <'�A     `�  ݓ  =U�� >C�A     l�  =U| =T��=Q��   O��A     =U   U��A     (�  =U  U��A     <�  =U  O��A     =U   On�A     =U   ?� ���A     �      ���  C�  �!�5  �& �& C��  �!w  F' :' B�  �<v  �' �' B�  �BZ  v( b( BXL  �BZ  v) b) BV�  �BZ  x* b* BR�  �n  }+ w+ B� ��  �+ �+ BQ  �Ks  , , Pcur �D4  V, @, B�� �D4  D- >- Pn ��  �- �- B�  ��  �- �- B#�  ��  L. @. B4�  �P  �. �. D�0  �e�A     E �  X�  (�  ��  ��(2�  �D4  ��E0�  3�  Plen (�  _/ Y/ K�A     �       ǖ  B/� PD4  �/ �/ <'�A     �  [�  =U��~=Q�� <H�A     w�  s�  =U  U]�A     ��  =U =Q
� U��A     ��  =U��=T}  >��A     ��  =U��~=T   <C�A     �  �  =U~ =T��=Q�� U~�A     �  =U��=T} =Q=R��~�# O�A     =U��=T}   U��A     G�  =U~  O��A     =U~   K��A           F�  (�  ��  ��Bf�  ��   '0 %0 U��A     ��  =Us =T0 U*�A     ŗ  =Us =T1 UQ�A     �  =Us =T0=Q	�1H     =R8 Ux�A     �  =U =T0=Q��=R5 U��A     /�  =Us =T}  O��A     =U =T}   U�A     Z�  =U~  U��A     }�  =U~�=T} =Q��~ U��A     ��  =U~�=T} =Q��~ U��A       =U~�=T4=Q��~ U�A     ۘ  =U =T0 UI�A     ��  =U =T1 U~�A     �  =U =T2 U��A     &�  =U =T3 U��A     @�  =U =Ts  U�A     ]�  =Us =T��� U=�A     v�  =U =T0 Oj�A     =Us =T0  ^�  ���A     :      ���  C�  ��5  c0 S0 C��  �w  &1 1 B�  �<v  �1 �1 B>) �BZ  �2 �2 BR�  �n  �3 �3 (� ��  ��B��  ��  #4 4 B.� ��  �4 �4 BQ  �Ks  5 5 D�0  �m�A     E`�  1�  Pidx O�  \5 R5 (�  P�  ��(2�  QD4  ��E��  \�  B/� �D4  �5 �5 <��A     �  �  =U~ =Q�� <��A     w�  
�  =U}  U��A     %�  =U} =Q
� U��A     A�  =U��=Ts  >��A     ��  =U~ =T}   U1�A     p�  =U  U8�A     ��  =U  <^�A     �  ��  =U =T��=Q�� Um�A     ��  =U  U��A     қ  =U  U��A     �  =U  U��A     ��  =U  <��A     ��  �  =Ts =R~  O�A     =U��=Ts   U��A     E�  =U  U�A     Y�  =U  U!�A     m�  =U  UD�A     ��  =U��=T���=Q~  UC�A     ��  =U  <��A     �  ˜  =U~ =T(=Q�� >��A     ��  =T~   ?� ��A     �      �_�  C�  �5  e6 G6 C��  w  �7 �7 B�  <v  �8 �8 Pcur D4  �9 �9 B�� D4  e; W; BQ  Ks  < �; E��  N�  BН  '�2  �< �< B.� (�  o= k= B.�  (�  �= �= Pn ('�  > k> BI5 )BZ  ]? U? BR�  *n  �? �? (� +�  ��B�  ,1  G@ A@ E0�  o�  B^�  [�   �@ �@ OY�A     =U} =Ts=Q	�1H     =R8  E`�  �  B�j ��  �@ �@ K��A     n       �  Plen ��  ,A &A U��A     ˞  =U  O��A     =U��=T| =Q} =Rv  U��A     �  =U  O��A     =U   Ue�A     )�  =U  U~�A     =�  =U  <��A     ��  V�  =Uw  <��A     ��  o�  =Uw  U��A     ��  =U�� <�A     ��  ��  =Uw =T2=Q0=R��=X0=Y�� <��A     ��  �  =Uw =T8=Q0=R��=X0=Y�� U�A     �  =U�=T| =Qw  Ui�A     )�  =U  U��A     =�  =U  O�A     =U   O��A     =U   ?��  ���A     3      ��  C�  �$�5  �A zA C��  �$w  B B B�  �<v  �B �B B:  ��  C C Bx  ��  �C �C B�� ��  dD XD (/� ���  ��B��  ��  �D �D BE  ��  0E ,E U��A     [�  =Uv =T6=Qw =R3 <}�A     ��  z�  =U
�=Tv  <��A     ��  ��  =Tv  <��A     ��  ��  =Tv  <��A     ��  ¡  =Tv  <��A     ��  ڡ  =Tv  >��A     ��  =Tv   H	  �  �  @    A��  �G   @�A     �       ��  C�  � <v  pE fE C�  � BA  �E �E C2�  � J4  nF dF C�  � 1  �F �F Pcur �D4  $G  G B�� �D4  ]G [G Kt�A     ;       �  Ps ��  �G �G Uz�A     �  =Us  O��A     =Us   Oa�A     =Us   ?;�  �0�A            �B�  @�  ��5  U@��  �w  T *��  !�  ƣ  +�  !$�5  +��  "$w  +�F #$_\  ,� %�  ,װ  &U   ,>�  '�  ,:�  (�  ,�  )�(  -�u  � ?�  
�A            �0�  C�  
�5  �G �G C��  w  H H O#�A     =U�T=T0=Q0=R0  ?�  �p�A           ���  C�  �#�5  jH ^H C��  �#w  �H �H (w�  ���  ��|(m�  ��  ��|B� ��  cI YI B�  �<v  �I �I B�  ��(  @J <J B�2 �\  zJ vJ Pn ��  �J �J Bu�  �D4  K K B��  �D4  \K TK D�u  ��A     U��A     d�  =Us =T��|=Q@=R��| <��A     �  ��  =Uv =Q0 OG�A     =Us =T0  1]  ��  @    ?��  b@�A           ��  C�  b&�5  �K �K C��  c&w  L L (� e�  ��zB�  f<v  �L �L B�  g�(  	M M (��  h�  ��{Pn i�  GM AM (`h  i�  ��zBu�  jD4  �M �M B��  kD4  �M �M BR�  ln  %N !N D�u  �%�A     K �A     �       ħ  /map �}'  B��  �\  _N ]N (��  ��  ��{Pp ��  �N �N (2]  ��  ��zK��A     H       p�  B�  �\  �N �N U��A     Z�  =U  O��A     =U =T0  U,�A     ��  =U =T��{=QD=R��z >e�A     ��  =U��z=T8=Q0=X0=Y��z  U��A     �  =U =T��{=Q4=R��z >��A     �  =Us =T0  1]  �  @    1]  %�  @    ?��  ���A     �      �*�  C�  �,�5  O O C��   ,w  mO cO (w�  ��  ��|(m�  �  ��{B`h  �  �O �O B�  <v  =P 3P B� �  �P �P B�  �(  /Q +Q D�u  \�A     E �  �  Bu�  D4  oQ gQ B��  D4  �Q �Q Pn �  ER 9R FP�  (��  '�  ��{B�2 (\  �R �R Bdh  )�  S S (+�  )�  ��{E��  ��  B�  O\  LS HS O��A     =U =T0  UI�A     �  =U =T��{=Q4=R��{ >z�A     �  =Us =Q��{�   O��A     =U =T��|=Q@=R��{  ?��  ���A     &      �٫  C�  �&�5  �S �S C��  �&w  �S �S (��  ��  ��~Pn ��  XT RT (`h  ��  ��~B� ��  �T �T B�  ��(  �T �T BR�  �n  U U D�u  ���A     EЌ  ��  B�2 �\  DU <U BF@ �D4  �U �U Plen ��  �U �U <R�A     ��  X�  =U~  <b�A     �  ��  =U~ =Ts����=Q��~ >��A     w�  =Qs   U��A     ��  =U} =T��~=Q4=R��~ >�A     �  =Us =T0  ?e�  }��A           ���  C�  }�5  5V -V BR�  n  �V �V B�  ��(  �V �V F��  Bm�  ��  �V �V B`h  ��  3W /W Pn ��  wW iW K��A            ��  Bim �}'  X X >�A     ��  =U|   <��A     ��  Ь  =U|  <�A     ��  �  =U|  <9�A     ��   �  =U|  <S�A     ��  �  =U|  <��A     ��  0�  =U|  <��A     ��  H�  =U|  <"�A     ��  `�  =U|  <O�A     ��  x�  =U|  <i�A     ��  ��  =U|  >��A     ��  =U|    A0�  Y�  � B     �       ���  C�  Y!�5  WX QX C�u  Z!�  �X �X C�  [!�  )Y !Y B�  ]�(  �Y �Y (��  _��  ��Pi `�  �Y �Y Pnc `�  \Z XZ <� B     ��  y�  =Uu =Tt =Qq  >� B     �  =Uvh  �  ��  @    A��  F�   B     c       �R�  C�  F!�5  �Z �Z C�u  G!�  �Z �Z C�  H!�  M[ G[ (9�  JR�  ��Pi K�  �[ �[ GYB     ��  >vB     ϯ  =U} =Tv =Qw   �  b�  @    A(�  7�  �B            �ϯ  C�  7�5  �[ �[ C� 8�  ,\ (\ _�B     ��  =U�U=T0=Q0  As�  ��  pB     �      ���  C�  ��5  s\ e\ C�u  ��  ] ] C�  �j'  �] u] B� ��  ^ ^ B�  ��(  Y^ U^ Pn ��  �^ �^ Pp ��  _ _ (ͫ  ���  ��~D�Y #/B     Ep�  l�  B�v  ��  �_ �_ B��  ��  �_ �_ Pmap �}'  ?` 9` Bq�  �j'  �` �` Bӫ  ��  �` �` BAT  ��  7a )a B;  �#�  �a �a E��  ^�  B��  �  Hb <b  G�B     ��   <VB     �  ��  =Qq N�  s  >�B     �  =U~ =T0=Qq N�  ��~  �  Ʊ  @    AS�  ��  ��A     �       ���  C�  ��5  �b �b C�u  ��  .c $c C�  ��  �c �c B�  ��(  d 	d (��  ���  �@Pi ��  bd Zd Pnc ��  �d �d > B     ��  =Uu =Tt =Qq   *�  ��  ܲ  +�  ��5  +�u  ��  +�  ��  ,� ��   *��  r�  d�  +�  r�5  +�u  s�  +�  t�  ,�  v�(  /n w�  /m w�  ,(�  y1  0,E  ��  0,��  ��     A7�  .�  `B     �      ���  C�  .�5  .e *e C��  /rw  se ge BR�  1n  �e �e B6~  2xw  Af 5f (��  3�?  ��~(� 4�  ��~Pi 5�  �f �f (��  6��  ��~B�  7�(   g g D�u  l�B     <�B     X�  f�  =U�U=Tt  <�B     �  �  =Q��~ <B     ��  ��  =Uu =Tt =Qq  >HB     �  =Ush  Z��  �  +r�  �  +��   �  +$�   �   8��  ��   �A     �       �X�  9��  � }'  �g g Mncv � �  h �g :j �
G   ih eh G��A     ��   8�  ��  ��A     n       �
�  9�  �*�5  �h �h L��  �*Fw  T;�  ��(  �h �h :n ��  i i `� ��  J��A     5       ;dh  �
�  Wi Si :map �}'  �i �i   �?  8��  h�  ��A     �      �N�  9�  h�5  �i �i 9m�  i�  �j �j 9`h  j�  _k Ok ;�  l�(  l l ;R�  mn  �l �l ;� n�  �l �l 7�u  ��A     7�0  ��A     K(�A     P      ʷ  :nn ��  �l �l <E�A     ��  '�  =U =T8=Q0=R~ =X0=Y�� <r�A     ��  \�  =U =T�=Q0=R~ =X0=Y�� <��A     ��  ��  =U =T =Q0=R~ =X0=Y�� >��A     ��  =U =T8=Q0=R
| 1$����=X0=Y��  K�A     a       +�  :n ��  "m  m >%�A     ��  =U =T8=Q0=R| v ����=X0=Y��  >��A     �  =U =T
 =Q��  A��  J�  ��A     �      �?�  C'�  J �  Nm Fm C�  K ]  �m �m C�^ L �  �n �n C:1  M T  �o �o B)�  O�6  1p )p B� P�  �p �p (�3 Qk  ��hB�  R�5  bq ^q BZy  S1  �q �q B��  T1  }r sr (=�  U1  ��gB�6  Vb4  	s s BQ  WKs  Ks Es Be�  X�i  �s �s (��  ZH	  ��gBw�  [�  Zt Rt (��  \�	  ��gB<�  ]1  �t �t B�z  _1  Su Gu -�u  7K��A     Y       >�  B�8  �E  �u �u G��A     ��  G��A     ��   E��  ��  (C!  ��  ��gBN �?�  v  v E0�  R�  Pn �  @v >v Pcur �,  ov kv Pvec �  �v �v B�� �  2w .w B�� �  pw lw a}�  ��A      ��A            "C�  b��  R��  �w �w J��A            V��  �w �w V��  x x   a}�  	�A      	�A            "��  b��  R��  Ux Sx J	�A            V��  ~x zx V��  �x �x   Q}�  ��A      `�  ��  b��  R��   y �x F`�  V��  <y 8y V��  y {y   c}�  ��A      ��A            b��  b��  J��A            V��  �y �y V��  z �y    Q}�  L�A      Љ  �"��  R��  >z <z R��  ez cz FЉ  V��  �z �z V��  �z �z   Q}�  q�A       �  �"��  R��  { { R��  5{ 3{ F �  V��  ^{ Z{ V��  �{ �{   G��A     ��  G��A     ��  <L�A     ��  7�  =U} =T��g <��A     ��  ]�  =U} =T��g=Q~  <7�A     ��  |�  =U} =T��g <z�A     ��  ��  =Us0 G%�A     ��  G:�A     ��   U��A     ֽ  =U��h=Tv =Q} =Rs  <)�A     w�  �  =U��h=T~ =Q��g=R��g U��A     �  =U��h U@�A     -�  =T��g O��A     =U��h  .  A_�  �  `�A     T      ���  C�  �  �{ �{ CN� �  `| X| C.� �  �| �| C:1  T  *} &} C\-  �  m} c} B�  �5  �} �} (�3 k  ��hB�6  b4  e~ [~ BQ  Ks  �~ �~ Pnn �    B� �  � � U��A     o�  =U��h=T} =Q0=R0 <U�A     ��  ��  =Uw =Tv  Gj�A     ��   8;�  ��  @�A           ���  9�  �$�5  � � 9�  �$�a  G� A� ;� ��  �� �� '�3 �k  ��h;�^ ��  � � ;�6  �b4  %� � ;Q  �Ks  �� �� U��A     j�  =U��h=Tv =Q0=R0 <"�A     ��  ��  =Uw =Ts  OJ�A     =Uw   8۶  ��  ��A     Q       �w�  9�3 �h  �� �� 9�^ ��  � � '��  ��	  �`'=�  �1  �_;� ��  H� D� K �A     +       O�  ;�  ��5  �� � O'�A     =T�`  >��A     w�  =Us =T�T=Q�`=R�_  8�  +�  ��A           ���  9�3 +3h  �� �� 9�^ ,3�  � � 9�  -3�   �� �� 9=�  .3��  � � ;�  0�5  n� j� ;�6  1b4  �� �� ;� 2�  � � ;Q  4Ks  �� �� ;e�  5�i  ˅ Å 'A�  6�d  ��u:inc 9"�!  /� +� Kc�A     }       ��  '��  hY  ��lUw�A     ��  =U��u=Ts =Q1 U��A     ��  =Uv =Tv�=Q��l U��A     ��  =U��u O��A     =U��u  K��A     |       h�  'N �"�   ��lG�A     ��  G �A     ��  G2�A     ��  OQ�A     =T} =Q0=R��l  UN�A     ��  =T} =Q  O��A     =Us   1  AB�  ��   �A     �       ���  C�  ��  i� e� C�U  ��  �� �� CB7  ��  � ߆ @Y�  ��  RB�  ��5   � � ]F�  ?�A       ��  �RT�  a� Y� RT�  ч ɇ Rz�  =� 9� Rz�  =� 9� Rm�  y� s� R`�  Έ Ȉ F��  V��  !� � V��  ]� W� V��  �� �� V��   � �� d��  Ў  V��  d� ^�     A ��  ��A     
       �G�  C~ �$_  �� �� CM�  �$�  � � _��A     ��  =U	 PH     =T�T  8&�  ��  ��A     J	      �;�  9�  �'�  =� '� Mkey �'[*  .� *� Midx �'�  }� g� 9�\ �'U   �� h� 9³  �'�  �� ~� ;ʼ  ��  � W� ;;�  ��  � �� ;�  ��5  ՗ �� ;�6  �b4  ؘ  Ep�  ;�  :val ��  �� �  E@�  Y�  :val ��  �� ��  E�  ��  Pok W1  d� ^� K��A            ��  Pval ];�  �� �� >��A     ��  =U�Q  G��A     w�   <��A     `�  ��  =U|  <��A     w�  �  =U�H=T| =Qv  <k�A     `�  �  =U}  >��A     w�  =U�H=T} =Q|   4   8 �  ��  ��A     �       ���  L�  �+�  ULۮ  �+"z  T 8D�  ��  ��A            ���  L�  �#�  U 8.�  ��  ��A            ���  L�  �+�  UL��  �++Y  T 8ؽ  ��  ��A     1       �/�  L�  �)�  ULù  �)%Y  T 8��  ih  p�A            �`�  L�  i�5  U 8b�  I�  ��A     p       ���  9�  I"�5  ۛ ՛ 9la J"�  3� '� :i L�  ǜ �� FЊ  ;��  Q�  Q� O� >�A     ��  =Uv    8��  =�  ��A     %       ���  9�  ="�5  ~� z� 9�^ >"�  �� �� 9B� ?"�  �� �� 9(5  @"�  L� F� >�A      �  =U�Q=Q	�R����  A7�  s�  ��A     �       �F�  C�  s$�  �� �� C��  t$�  �� � C�9  u$�  p� f� CY�  v$�  � � Pfi x�5  d� ^� Pi y�  �� �� FЍ  Ptk ��4  � �� Gz�A     ��    Z?�  J��  efi J!�5  +Z�  K!�  +2�  L!�  +Y�  M!�  /min O5  /mid O5  /max O5  /idx P�  0,y�  Y�    8�  ��  �B     Y      �V�  9v�  ��  V� N� 9Jy  �:  �� �� ;Q  �Ks  $� � ;R�  �n  �� �� '�  ��q  ��:fi ��5  Ȣ �� '� ��  ��;�  ��5  g� _� ;s�  �b4  Σ ƣ D�u  @	B     E �  w�  B�S D4  A� 9� ]V�  �
B      `�  %R�  �� �� R�  �� �� Rs�  Τ Ȥ Rg�  � � F`�  S��  ��V��  r� f� V��  � �� V��  Y� O� V��  ܦ ʦ V��  �� �� V��  :� 2� V��  �� � V��  }� s� V��  � � T��  �B     <�B     ��  ��  =U��~=T@=Q0=X0=Y�� <$B     �  ��  =Us  <8B     �  �  =Us  <zB     �  "�  =Us =T��~ <�B     '�  F�  =Q@=R	@�A      <�B     ��  `�  =U��~ >�B     �  =Us     <�B     ��  ��  =U|  <	B     �  ��  =U| =TX=Q�� <<	B     3�  ��  =U  U�	B     ��  =U�� <�	B     @�  ��  =U  <�	B     ��  �  =U| =Tv  U
B     ,�  =U�� U
B     A�  =U�� >�
B     @�  =U   4K�  m�  �  2v�  m�  2Jy  n:  ffi o�5  3� q�  3R�  rn  3�S sD4  3�� tD4  5p uD4  5kp v5  3ї  w�  3�  x  3�� y  5n z�  6�u  � 8�% XG   @�A     )       ���  ga X$�  Ugb Y$�  T;�  [5  � � ;ǫ  \5  ;� 9� ;��  ^�  `� ^� ;��  _�  �� ��  4m�  7�  ��  2F@ 7h  flen 8�  2o�  9U   3�6  ;b4  5n <�  03��  E�     HP�  (P�A     P       �}�  9R�  ("n  ܪ Ԫ Mfi )"�5  C� ;� <e�A     ��  H�  =Uv  <��A     ��  `�  =Uv  _��A     ��  =U�U=T�T  4�6  �T  ��  fa �T  fb �T  5ret �"  5tmp �"   h��  ��A           ��  iƴ  UiӴ  Ti�  Qd��  �  R�  �� �� RӴ  � ܫ Rƴ  � �   hܲ  `B           �*�  R��  Z� P� i�  Qb�  V�  Ь ̬ V"�  � � V-�  �� �� V8�  � � jE�  �B     �       VF�  �� �� dS�  @�  VT�  � �� c}�  B      B            �R��  @� >� R��  e� c� JB            V��  �� �� V��  ݯ ۯ      h��  �B     1       ���  R��  � � R��  Y� S� R��  �� �� Vβ  � � Y��  �B            ��  R��  � � R��  F� D� R��  k� i� J�B            kβ    >�B     �  =Tv =Qq N�  s   l�  �B     <       �W�  b0�  V<�  �� �� VH�  �� �� VT�  � � >�B     ��  =T	`BH       m�  �B     9       � �  R��  /� '� V�  �� �� j�  �B     "       R��  �� �� J�B     "       k�  j�  �B     "       V�  I� G� >�B     ��  N0�  s      h��   B     �       ���  R��  t� l� R��  ۳ ӳ R��  B� >� V��  � {� k��  j��  B     k       b��  b��  b��  JB     k       k��  V��  �� �� d��  ��  V��  '� !� <jB     `�  ��  =Uv  >�B     M�  =Uv =T~ =Q��     h~  B     �       �p�  R.~  z� p� R:~  �� � RF~  x� n� VR~  �� � S^~  �VSj~  �XY~  tB     )       ��  RF~  h� f� R:~  �� �� R.~  �� �� JtB     )       VR~  ݷ շ k^~  kj~  Tv~  �B     <�B     l�  ��  =T| =Qv  >�B     @�  =Us    <(B     �  �  =Us =T0 <JB     �~  8�  =Us =T�V=Q�X <aB     �  U�  =Us =T0 >pB     3�  =Us =Tv   n>Q  >Q  -�n�P  �P  -�nKM  KM  Yn\  \  Vn�3  �3  1n!,  !,  UoF\  F\  .�oUP  UP  hn�R  �R  n�=  �=  �o�6  �6  .�oBi  Bi  /n9  9  -co�K  �K  .vnE1  E1  -rn _   _  -ho�[ �[ /"o�Z �Z /nF  F  -mo�O  �O  /2p�  �  0 p�D  �D  0 o�4  �4  to�-  �-  dn5<  5<  ?njO  jO  n�-  �-  1BncL  cL  1o�,  �,  1�n�D  �D  �n�*  �*  [o�X  �X  ~nq]  q]  .zn)=  )=  gnB2  B2  /o_T  _T  2Xn�3  �3  -�nxL  xL  -�o��  ��  /   3"  �  )�  $"  �B     �o      �� :G  �9   X  ^� �L   �i int �i {S @	�   g
  	�      	 	@   v  	#	@   �  	&	@   |
  	)	@    h  	,	@   (�  	-	@   0�	  	2S   8�  	5S   < �   �  	�   �
  	8"c   
  	K  �   
�  	L  
�  	M  S  .�  
�A  -  �[  
�T  �  	T  >   
S   	`  �	  
	Z   �  B"�  �     ��  R   �a    �� ��  �N ��  �6  �   �  Y�  �  a   �    9      n        a    �  �'  -  a   K    9   9   a    �  �"W  ]  �   PJ�  2�  LZ   �  ML   pos NL   �  P  SF  Q   �1 R*  (=9 Sg  0R�  U  8y�  VZ  @�� WZ  H �  �  �\ �9   m  �a    o  ��  �  �6  <  L   Z  K  L   Z  L    `  �  2  t  z  �  K     :9   �  J�  x L�   y M�   )  O�  	�  B   s  M   u�   }  u�  V  v�  /  v�   t
  x�  k	  (�  �  Z    ��  Z   �  	S   B� 
Z  L  T    `  s  `  v	  a     �    	�  �  (N  �  PA   Z�  QA  �  S  s  T�   [  U  ?1  WS     �  A    Y�  �  =  Z   �e  �   M
  pmoc5  stib	  ltuo|  tolp 	  �'  b   "  �  �  %  <�  x >A   len ?T  *� @`   %  B�  	�    `�  �     S   S      a    �  �  q    S   2  S   S   a    �  ?  E  Z  S   S   a    �  `��  �  ��   �% ��  ?1  �S   �&  ��  !  ��   I  �  ()  �2  0R   �a   8�  �  @ �  �  �  �Z  	�  �       S   -  a   -   r  �  @  F  Q  r   �  ?^  d  y  r  Z  L    �  Y�  �  S   �  r  L   a    s  ��  �  S   �  r  �     W  0�5  �  �e   e� �  �� �Q  �� �y  �� ��   �� �3  ( �'  ��  �!  l`  �  �Z  �  -  �`  	a  m  �L  �r  �  ��   	�  �
  �A  �  �T  	�  �  �S   
  �Z   �  �9   	�  \#  �L   �   9   �  ,S   \&  7a   �0  D@   �H  Q-   b   �k	  xx ��   xy ��  yx ��  yy ��   a  �(	  	k	  z'  ��	  m  �r   ss  ��   �  �}	    ��	  �	  �	  a    �  ��	  �U  �a      ��	   %  ��	  �  $
  
  �   W
  �� "
   �@ #
  �U  $a    �  7�
  �; 9
   ��  :
   L  <W
  Z   #��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=Q  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  J�  
   s�  �  u�   ��  v�  �  x�  �
  z�  (  {�   �  }^  �  �#�  �  k  `��  R�  �   (  ��  |  ��  �  ��  �  ��  �  �g$  v  ��
  �  �(  (�%  ��  07&  �w$  8G   ��  X �  �"�  �  h  �  �M A$   k  �  R�     �  �"�  �  %  8;(  �� =G$   �M >�    ?�
   r$  @�  0 5  �$5  ;  %  ��  �� G$   �M T$  �  e   �  3  (�� 
r  h�� �  p�� �  x K  � �  �  �  �,�  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6  (A  7  0T  9�  8  :  @�  <�  H�  =  PE-  ?�	  X�!  D  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R�  ��� S7  �K1 W�  �R�  X  �Jy  YK  �%  [�
  ��	  ]�	  �    ^a   ��8  `p  � L   �  �    X��  �  ��   E-  ��	  N ��  �8  �!  P �  *%�  �  �  0t7  k  v�   �  w�  �@ x�  ݖ y�  E-  z�	   N |Q  0�  }�  pR  ~�  x�  �  �ߣ  �e  ��I ��  ��  ��  �h  ��  ��S  �  �4  ��  �8  �  �  �a    �  �9   �  ��  o  ��  �L �a    �8  �h  ( �
  L#D  J  W  H�  �  J�   = KV    L�  d  M�   �  Z   �V  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  (0  OJ  #   g)}  �  �   ��  =  �k	   L  ��   $  ��  0�  �l   8m  �#�!  h�  �N  pآ  �`  tG   ��  x �  �  7  �?  d�  �
  �).  4  �   H�m  �  �a    "  �  �!  ��   ~	  8f�  �
  h�   (  i�  �� k�  �� l�    n�  �  o�   �  p�  (�  q�  0 y  sm  �a  ��    �$    �  0'h  �N  )�   ?1  *�  }0  +�  i/  ,�  � -k	   �  �)u  {     H��  ��  ��   ?1  ��  (  �B  4  �k	  \  ��  0  �a   @ ��  ��  +!    tag �   �U  	   �  �    `  Z   
a  w%   }#  �&  h  �  &     
)  E   9
�  � ;
a   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  n  �  Z   �  :   �   ^$  1  �!  �!   :  ��  �  �	  �#  �3  9  �  H  �   I$  �T  Z  e  �   �&  �q  w    �  �  �   �   �!  H�  �  ��   S"  ��     �  �"  ��  �  ��   ;  ��  (%  �'  0�   �H  8��  �e  @ �  R  ��  x  =�	  H  E#D  	3  �  @J�  �  L�   �  Me  �� O  .� P:  �  Q�   �  RW  (�!  S�  08'  T�  8   W!�  �  -  (l  k  n�   �M o  ߣ  pe  �  q�   ?  k  )   &  �  :  �  �   w   .F  L  W  �   �  1c  i  ~  �  ~  !   x	  K  6�  �  �  �  �     �  :�  �  �  �  �  �   �  >   "  Y�  �  �    (  �    !   �  _     �  >  (  �  ~  !   $  fJ  P  e  (  �  �   �  lq  w  �  �  (  �  	   #  x��  �� �    �  � e  H  � �  P�  �   X9!  � >  `l� � e  h  � �  p 5    ��  �  H2Z  �S  4   �  5  (  6  04  7�  88  8  @ �  :  �  �=�  R�  ?   �  @�  n  A�  �  B�  1$  CB  2�  EZ  �� FZ  `�L Ha   � �  J�  f  P   �     �  #  K  �  �  �  #   �  &/  5  @  �   �%  *L  R  �  a  �   �%  -m  s  ~  �   {  1�  �  �  �  �   �  4�  �  �  �   l  8�  �  �  �  �  �   �  <�  �  �    �  �   �  @    �  8  �  �  �  `   �  GD  J  �  h  �  �  �     �'  Nt  z  �  �  �  K   �  S�  �  �  �  �  �  �  `  �   �  &  ���  �� �   i'  ��  H   ��  P  ��  X�A ��  `Y �#  h�#  �@  p�  �a  x�  �~  �  ��  ���  �  �U�  �8  ��!  �h  ���  ��  ��  ��  �&  ��  �   ��  	�  �&  ��  �  a   �>  ��  'O  ��   xC  ��   s/  ��  	�  �  0tl   �  v	   a   w	  �'  x	  !  y	  �#  z	   �  {	  ( �  }	   �  U'�   �   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {�   �  ��   �   �  	!  y   �  	!   �	  �  �!  !!  1!  y   	!   �'  �=!  C!  �  a!  y   �  B  a!   �   �!  �!  ��  )�    ��  )!  �  )1!   }  g!  	�!  O  ;�!  _� =%�!   ݰ  >%y    �!  �  @�!  �!  cA  �,"  "  /  �0"  �� �c   �M �0"   ?<  �,<"  �"  �5  P��"  �  ��   �� ��"  �Y �	#  �H �&#  U@ �L#   �9 �#x#  (�A  �#�#  0�^  �#�#  8�^  �#�#  @N7  �#$$  H 	B"  ��  �"  (Z  ��"  �"  �  	#  �!  	   17  �#  #  &#  �!   �G  �2#  8#  �  L#  �!  r   %G  �X#  ^#  �  r#  �!  r#   r  �@  ��#  �#  �  �#  �!  �!  r  r   �;  ��#  �#  B  �#  �!  r  r   �W  ��#  �#  r#  �#  �!     *;  �$  $  r#  $$  �!    r   �T  �$  g�  �B"  	0$    �  �  �  -1  B�  �  w$  L    &  �$  L    �$  �  �$  �   �$  �  �$  �  �  	  �   �$  �  �$  �     �  �%5  �  8Yj%  ��  [   Ǧ  \  ��  ]  d> ^  ��  _   I�  `�  (�  aB  0U  b�  2�  c�  4 ��  e�$  ��  p$�%  �$  ��  ���&  ֤  ��   Ğ  ��  ��  �a  �  �a  	��  �a  
�  �a  ��  ��&  �  ��&  (��  ��&  <�  ��&  X��  ��  p��  ��  x��  ��  |��  ��&  ��  ��&  �R�  �a  ���  �a  ���  �B  �F�  �B  �V�  �'  ���  �'  ���  ��  �"�  ��  ��  ��  �@�  �'  � �  �&  L    �  �&  L   	 �  '  L     �  '  L    �  +'  L    ��  ��%  o�  �#C'  �%  �  �+'  ��  �'  2]   a   U�  !�'  5�  "�   �  �  $U'  ��   *o(  m�  ,�   `h  -�  �  /o(  #�  0(  (��  1�(  ��  3�  z�  4�  ��  6�(  ��  7�(  ��  9�  (Ԯ  ;�(  0��  C�(  ���  D�  �   (  L    �  �(  L    �'  �(  L    v%  �(  L    7'  �(  L    �  �(  L    �  �(  L    ��  F�(  �'  �  Z   w *  U�   ��  ��  �  ��  ��  ޟ  $�  ��  �  	t�  
�  ܖ  �  ��  ��  d�  {�  ך  ʕ  �  ��  ��  m�  ,�  �  ^�  ׭  ~�  @�  �  ��  N�   ��  !��  "��  #ݴ  $��  %�  &�  ',�  (a�  )��  *x�  +��  ,"�  -"�  - a�  ��(  ��  #9*  ?*  r  N*  �   d�  )Z*  `*  �  o*  �   0�  /Z*  K�  6�*  �> 8r   �^ 9�   �  ;{*  Ѽ  >$�*  �*  ў  (@�*  
H B�"   ��  C�  XT D�*    �*  ��  N+  +  �  "+  	  �   B�  V.+  4+  D+  	  �   ��  ZP+  V+  �  ~+    �*  �  �*  "+  	   ��  b�+  �+  �  �+  �*  r   ��  f�+  �+  r  �+  �*  r#   ��  @j@,  �\ l -*   8` n D+  �\ o ~+  �_ p �+  �T r N*   }�  s o*  (ʬ  t W,  0�  u W,  8 	�+  ��  jQ,  @,  [  ��  )$i,  o,  H�  ��  ,�,  �,  �  �,    �,  �,   I'  ],  ��  1�,  �,  �,  ],  �  �  �  �   ��  8�,  �,  �,  ],   �  ;.-  M� =t,   �� >�,  Յ ?�,   ��  A:-  �,  �  h!L-  R-  ��  ��  u-c-  �-  ��  8V�-    X@-   j�  Y�-  =9 ZQ.  �� [�-  Q� \#.   �� ]/.  (�� ^x.  0 	i-  ��  ��-  �-  �-  @-   ��  �.  .  #.  @-  �  �   K�  �.  å  �;.  A.  Q.  @-  �   ��  
^.  d.  �  x.  @-  �   ?�  1�.  �.  �  �.  @-  �.  ],       1�  �!�.  �.  $�  ��  �-�.  K/  .�  8�K/    ��.   j�  �P/  =9 ��/  �� �n/  +�  ��/   �� ��/  (�� �0  0 	�.  ǡ  �]/  c/  n/  �.   ��  �{/  �/  �/  �.  �  �  �   ��  ��/  �/  �/  �.  �  �  r   !�  &�/  �/  �/  �.  �  r   K�  D�/  0  �  0  �.  �   	�  k$0  *0  �  H0  �.  �.  ],     ��  ��0  ��  ��0   X� ��0  l� ��0   .-  �0  �   �0  W-  �0  �   �0  �.  �0  �   �0  $�  �H0  �  � �0  �0  �3  51   num 7�   str 8�   +P  :�0  �J  =:1  key ?1   �U  @@    �7  D$F1  1  O  HX1  ^1  �  m1  m1   1  �Z  K1  �1  B  �1  m1  m1   �S  (O�1  �� Q�   �  R�  �6 S�  �B  UL1  3  Vs1  >) X�1    :1  e-  \ 2  �1  �    ��  W42  ��  Y�    ��  [2  a  @2  �  ��  (��2  �9  ��   ��  ��  ɲ  ��  �  ��  �  ��    T�  ��2  R2  ��  ��2  ��  ��   ��  ��  x ��  y ��   �  ��2  �2  z�  X�y3  ��  �B   ��  �  �Z  ��  (%?  ��  0L�  ��2  8)�  ��  @W�  ��2  HѺ  ��  P b�  ��3  3  ͳ  @@4  Jy  BK   �S C�  ܱ  D�  .� E�  ��  Fa  ��  G�   
�  H�  (�P  J4  0Ӏ K@2  8 �  ,�  M�3  ��  M,4  �3  !
�  P�4  ߣ  R�   x  S�  .� U�  ē  V�4  " � W�4   �  �4  L   � ��  Y24  ��  Y�4  24  ��  (\5  ߣ  _�   x  `�  ē  b2  ��  c2  Ӷ  e�   �  f�  $ r�  h�4  ��  h%5  �4  W�  mS5  Kw  t�   7�  uL2   0�  w+5  j�  {�5  ��  }�   �  ~�  �w  �   J�  �_5  1�  ��5  �{  ��5    �5  �  ��5  �   �6  ��  ��   k  �6  �q  ��   q  ��  y|  �"6   S5  �5  �  ��5  ��  �@6  �5  %�  �!R6  X6  �  �M�8  k  O�   Jy  PK  R�  Q  ��  R�  �   S�   �  T�  $(  Va  (|  Wa  )x�  Xa  *п  Z�  ,�J  \B  0i�  ^4  8�  _4  xC�  `4  �= b�4  ���  c5  p�  e4  8��  f4  x=�  g4  ���  h4  ��  j  8��  mF2  @V�  p�  HV` qF2  P��  r@2  X��  s�  `/�  u�>  h��  v�  0��  w�>  8j�  y�>  82�  |�0  Xs  E,  `��  ��  h�  ��>  pd�  �  x|�  �  �˽  ��	  �ʞ  �(6  �8�  �?  � ֥  0�9  ��  �B   �  �B  v�  �F6  �  ��  ݺ  ��  ��  ��  c�  ��   BV �9  ( `  �  ��8  ��  �59  �8  !��  H�j;  ��  ��   Ǧ  ��  @�  ��  ��  ��  d> ��  ��  ��  �  �B  I�  ��   U  ��  (�  ��  0��  ��  8�& ��  <��  �k	  @?�  �B  `U�  ��  hw�  ��  p֤  ��  �;�  �  �ܲ  ��  �w�  ��  ���  ��  ��  ��  ���  ��  �ٛ  ��  ��  ��  �g�  ��  �`�  ��  �x�  ��  ��  ��  �|�  ��  �"��  ��   "�  ��  "n�  ��  "��  ��  "��  ��   "`�  ��  ("�  ��  0"m�  ��  4"�m  ��  6"A�  ��  8"��  ��  @ ��  �;9  ~�  ��;  ;9  S�  �$�;  �;  ��  �*]<  Ҳ  ,j;   -�  -->  H�  09   ݺ  1�  P#NDV 2�  X�  <@2  `K�  =@2  h�  >�  p��  ?�  t��  A4  xZ�  BF2  �l�  Er  � !E�  ���=  ��  �a   �  �a  ��  �a  �  �a  ��  ��=  �  �>  x��  ��=  �"�  �>  8"��  ��  �"��  ��  �"��  ��  �"��  ��  ��   �  �R�  a  ���  a  �V�  >  ���  >   ��  B  �6�  �  �Ğ  �  �"�  	�  ���  
�  �Т  �  �P�  �  �W�  �  ���  �  ���  �  ���  �;  � �  >  L    �  >  L   	 �  ->  L    ��  ]<  ��  G>  ]<  a�   �>  ߣ  a   �  �  �U  @2  
�  �  w�  !�  .�  "�  �  #a   �  %M>  �  %�>  M>  9�  G�;  �;  �>  L   � j%  42  d�  �X6  �6  `S�?  �<  U�   �Q  V�  a(  X�  VA  Y�  Q) [�   nX  \�  "�D  ^�?  (�5  _�?  8M   a�  H}  b�  JV  c�  L/  d�  N7K  f�  P>D  g�  R�:  i�  T�3  j�  V=]  k�  X �  @  L    �5  m?  �Q  8��@  �  ��   �Z  ��  %?  ��  
L/  ��  �<  ��  �Y  ��  �7  ��  �)  ��  �O  ��  �H  ��  vH  ��  ^  ��@  �>  ��  $�7  ��  &0>  �a   (�+  �a   0 �  	A  L    �H  �@  �?  8AB  �  C�   �Z  D�  %?  E�  
L/  F�  S.  H�  �W  J�  �W  K�  C  L�  �O  M�  �H  N�  vH  O�  ^  Q�@  �>  S�  $�B  T�  &0>  Za   (�+  [a   0 �]  ]A  �B  �|BD  ��  ~�   �)  �  �)  ��  �.  ��  U  ��  �V  ��  
�0  ��  �6  ��  �C  ��  U?  ��  6P  ��  �C  ��  &L  ��  *J  ��  �L  ��  HP  ��  N*  �BD   [2  ��  0k2  ��  8.  ��  @{2  ��  HQ2  �RD  P�0  ��  Tp4  ��  VmU  ��  X�Z  ��  Z ?  ��  \:  ��  ^�I  ��  `E8  ��  b�;  ��  h�;  ��  p�O  ��  xDF  ��  zfV  ��  |�9  ��  ~[9  ��  ��G  ��  �zQ  ��  � a  RD  L   	 N  bD  L    {D  �B  �1  @��D  �I  ��   6Y  ��  �^  ��  S  ��  )  ��  @3  ��   �0  ��  (4C  ��  0�C  ��  8 aM  �oD  �I  @��E  �  ��   _7  ��  )  ��  �O  ��  �n ��  �T  ��  EF  ��  I  ��  �K  ��E  N:  ��E  ,L  �
F  4�E  �N  :�Z  �N  ;�Z  �a  <^  �a  = N  �E  L    N  
F  L    N  F  L    eU  �	E  �9  (7G  ��  9�   a@  :�  b<  ;�  
8  <�  .  =�  �H  >�  �Q  ?�  X  @�  �.  A�  �;  B�  ))  C�  eH  D�  I_  E�  �B  F�   !3  G�  " �)  I'F  �  IJG  F@ K   I�  L�  K�  M�   ԃ  OG  �b  hh�G  `h  j�   m�  k�  dh  l�G   JG  �G  L    ��  nVG  �j  0�H  F@ �   I�  ��  def ��  K�  ��  tag ��   c  ��  ( )�  ��G  �  �DH  �  ��   c  ��  Cg  ��   �~  �H  z�   ��H  `h  ��   m�  ��  L�  ��  dh  ��H  e  ��H   H  DH  J�  �PH  �R   F�H  tag H�   ��  I�  .� J�  �P  K4   DG  M�H  f3   �GI  Tag ��   Q  ��  .*  ��  �K  ��   gW  �SI  I  �^   �I  k@  �   aE  �  p0  �  �>  �  H  �  �/  �  �� @2   �F  YI  �<  0J  H  2�   �/  3�  �� 8@2   qS  :�I  A9  0U�J  ߣ  W�   �E  X�  �^  Y�  =Y Z�J  <  [�  �=  \�J   Jy  ]K  ( �I  J  rY  _J  �1  ~�J  �.  ��   �L  ��   Z  ��J  �J  �V  �K  ��  ��   f>  ��  Y  ��J   �)  ��J  ��  ��K  �  ��   ��  ��  ~  ��  �  ��  �  ��  5  ��  
B  ��  �  ��   �w  �+K  �A  /`L    1N   �  2N  �N  3a  o=  4N  D4  5N  �^  6N  `*  7N  �0  8N  �G  9N  �D  :N  	I:  ;`L  
 N  pL  L    �@  =�K  �\  ��L  +  �pL   Y�  �pL  �
  �a  (  �a  �F  �a  �C  �a   <)  ��L  }L  �,  :M  �  �   AK  �  z8  2  V :M   @M  N  �R  �L  	F  .~M  �  0�   �P  1@M   ">  3SM  $I�M  %�K KFM  %`B L~M   �[   E�M  �z  GB   =Y N�M   �6  P�M  O]  a!�M  �M  �(  7N  (�cN  >) �@2   -N  �@2  V` �@2  TE  ��  �/  ��   �z  �B  $ G  � N  &8  � }N  �N  eS  po�R  �� q   ^  s�H  ��^  u�  [>  v�   �W  wGI  (� y@  0�=  z	A  ��,  |G  ���  ~B  ��(  B  �AK  ��  0XL  ��J  8#os2 �bD  hp�  ��D  �T  �@2  0#9  ��  8!H ��T  @�+  ��T  H@.  �AU  P�E  �U  X�P  �U  `@  �U  h$S  �a   ps  �a   x#mm �a   �#var �a   �Q  �a   �<B �K  �2Y �F  �=  ��  �=  ��L  �UV  ��M  ��(  ��  =  �@2   /:  ��  (�?  �@2  0�]  ��  8#cvt ��U  @�R  ��R  H5$  ��	  P��  ��  `HT  ��  h�*  ��  p�J  �B  x�+  �B  y�  ��M  ��C  �r  ��-  ��  �j7  ��  �kN  ��  ��F  ��  �#7  ��  ��(  �@2  �rE  �@2  �QZ  ��  �4  ��  ��@  ��  �:L  �@2  ��G  �@2  ��]  ��  ��W  ��U  ��/  ��  ��B   L2   �I  @2  s-  �  �*  �  ,  r  ,  r   #bdf 	cN  (�T  �  P#F  �  X�U  �  `�K  �  h �=  ��R  �R  �  �R  a    �Q  �"S  S  �\  xc�T  �  epN   �  frV  )�  g�  �V  h�  :1  j�   �^ k�  (Jy  mK  0�  n�  8�  p�  <�!  q  @R0  r�  `�  s�  duN t�  h6  uB  lpp1 v�  ppp2 w�  �2�  zMV  �Xc  {MV  ��6  }ZV  )  ~@2  �8  �   �L �a   (C  ��  0��  ��  4#pp3 ��  8#pp4 ��  Hy�  �@2  X�� �@2  `U  ��
  h �I  ��T  �T  �  �T  pN  �  K  4    1  �T  U  �  U  �R  �  �  �   �M  +,U  2U  �  AU  �R   �<  :NU  TU  _U  �R   y*  Z   =�U  4   �^  J  b8  �T   lK  H_U  �  |T  @?MV  R�  A   �  B�  n  C�  
Z�  D�  �  E�  org G  cur H  ��  I   s  K@2  ([  L2  0c+  N�  8 R8  P�U  RG  T'gV  mV  [  O  _ V  �V  LL  @�   !pN  8�  ` ,�V  ��  .�   -U  /�  X `�   1�V  �V  !~�  H <$W  ��  >�   "��  @B  0"��   AB  1"��  C�  8"��  D�  @ Z�   F0W  �V  !@�   Q_W  �   S],   ��   T_W   ],  oW  L   � ��   V{W  6W  ��  !$$�W  �W  ��   !&�W  
H !(�"   �  !)2   
��  !.<$  
e�  !;<$  ��  H"4pX  k  "6�   �S "7@2  �� "8@2  y�  "9@2  4� ";F2   top "<F2  (�m  "=�  0s�  "?�  4ݰ  "@a   8m�  "B�  @�m  "C�  B ��  "E�W  ��  "E�X  �W  Z   "_�X  >�   u�  �  ��  ��  d�  ��  �  �  T�  	 S�  "o�X  �X  �  �X  |X   a�   "qcY  ��  "sS    � "tS   x  "u�  �  "va  ��  "w�X  m�  "x�  �  "y�   F�  "�X  	cY  Z   #��[  ��   ��  G�  ��  ��  ��  \�  W�  ��  l�  	��  
 �  ��  �  F�  ��  �  <�  ��  ��  ��  4�   v�  !�  ":�  #�  $ �  %�  &��  '9�  (y�  0"�  1��  @��  A7�  Q��  R��  S��  T!�  UX�  V�  W��  XI�  `�  aJ�  b��  c�  p��  ���  ���  �(�  ���  �w�  �%�  �P�  ���  ���  ���  �Q�  �$�  ���  �l�  ���  �_�  �e�  ���  ���  ���  �>�  �E�  ��  �(�  ���  ���  ���  ��  ���  ��  �)�  ��  ���  �*�  ���  ���  ���  ���  ���  �&�  ��  ���  ���  ���  �}�  �t�  � &�W  k	�gH     &�W  �	@gH     '�(  Z   $9X\  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  $V�\  �\ $Xa   �  $Ya  x  $Z�   �7  $\X\  	�\  Y�  %E�\  �\  �  �\  K  pN  �  �  #   ��  %k�\  �y  %��\  �\  �\  pN   �m  %�]  ]  �  1]  pN  �  �  @2  4   t�  %">]  D]  �  q]  pN  �  �  �  K  q]  w]   �  �K  ن  %@�]  �]  �  �]  pN  �  4   �}  %Z�]  �]  �  �]  pN  �  �]   �  kp  %s�]  �]  �  ^  pN  �  2   T�  %�^  ^  �  3^  pN  K  B   �m  %�@^  F^  e^  pN  B  �  �U  2   1z  %�r^  x^  �  �^  pN  �  2   �a  %��^  �^  B  �^  pN  �  �^  �^   �  sz  %��^  �^  �  �^  pN  K   �w  %�\  �m  %!	_  _  �  (_  pN  �  �   3b  �%2�`  !H %4"�T   �A %6"�\  �M %7"�\  Y %8"�\  ��  %9"e   K %;"�\  (�; %?"�^  0|G %@"^  8H %A"�^  @"I %B"�^  H�Y %C"�^  P�Z %D"�^  X�S %F"�^  `�< %G"�^  h�9 %J"�^  p7B %L"�^  x-Y %M"�^  �(K %Q"�^  �Z %S"1]  ��i  %V"�]  �s  %W"�^  �U�  %\"�^  ��@ %b"�^  �x> %c"^  ��j  %e"�^  ��w  %f"�^  ��V %h"}]  ��= %i"�]  ��D %k"3^  �tW %m"e^  ��9 %n"�^  � ��  %p(_  ~c  %ta  �`  �C  h&*Xa  �� &,Z$   �Z  &.�  8�  &/B  <X;  &0Xa  @آ  &1`  ` �  ha  L    �D  &3ta  	a  ��  &?-�a  �a  ۳  `&�b  ��  &�@2   y�  &�	  �� &�	  �� &��  ��  &��   Ǩ  &��  $(2 &�F2  (Ϛ  &�L2  0R�  &�  8_� &��b  @ ��   &T^b  �� &Wwb   �Y &\�b  add &_�b  �x &e�b   �  wb  za  �     ^b  �b  za   }b  �  �b  za  �  a   �   �b  r�  &gb  	�b  �  &�"�b  �b  ��  �&�8c  y�  &�@2   2�  &�@2  �� &�@2  � &��  R�  &�   _� &�7g  ( ��  &�"Dc  Jc  ��  &�c  �S &�@2   �� &�@2  � &�Qd   ��  &�"�c  	c  �c  ��  0&�d  9�  &��   �{  &�e  � &��d  ��  &�%e  x  &��  �  &�a  m�  &��   �  &��  $��  &�  ( '��  Z   &�Qd  ˟   .�  ��  ��  ��  ��   ��  &�d  'L�  Z   &��d  ��   ��  Ʊ  ��  ��  g�  �  ��  W�  �  	|�  
K�  ��   8�  &�]d  '��  Z   &�e  c�   ��  p�  �  �  ��  �  ��  ��  }�  	 ��  &��d  ��  &�1e  7e  Ge  �  	   �  h&kf  �� &n&f   �Y &t7f  �? &w7f  �2 &y7f  �! &|Lf   �$ &~ff  (�* &��f  0�3 &��f  8k! &��f  @�A &��f  HV- &�g  P�F &�1g  X  &�1g  ` &f  �b  @2  @2     f  7f  �b   ,f  �  Lf  �b   =f  �  ff  �b  �   Rf  �  �f  �b  @2  	  4  B   lf  �  �f  �b  �  �U   �f  �  �f  �b  �  �  �   �f  �f  �b  8c   �f  g  �b  8c  �  �^   �f  �  1g  �b  �c  �  �  4   g  �  &�Ge  	7g  ~�  &�Vg  l�  p&Sh  R�  &   �  &�  )�  &$W  ��  &�  2�  &�.   �� &�.  (��  &�h  0��  &�h  8R0  &   @�  &!  H�!  &#�  P��  &$B  X�� &%B  Yb�  &&B  Z��  &(B  [�  &)B  \_� &+�h  ` ګ  &�~h  �� &��h   �Y &��h   �h  �h  a   B   Ig  ~h  �h  �h   �h  �  &�Sh  �  î  &B�h  2�  &D@2   �� &E@2  y�  &F@2   {�  &H�h  ��  &Li  i  �  :i  pN  �  F2  4   l�  &RGi  Mi  bi  pN  F2  �   ��  �&W}k  <0 &YIg   4� &[}k  p#top &\�  �O� &^�k   Xc  &_�k  ���  &a�  ��  &b�  ��  &c�k  �#cff &eF6  �  &f�;   ˽  &g�k  (
�  &i�h  0�  &jB  8��  &k�  <z�  &m�  @�  &n�  D��  &p�  H�  &q�  L~�  &sF2  P9� &tF2  XV &vF2  `�  &w�  h&  &y  l�J &{B  p�  &}&	i  x��  &~&:i  �s  &�E,  �Ğ  &��  ���  &�L2  �q�  &��1  ���  &�k	  �w�  &��  ��  &��(  ��  &��'  ��  &��  � �  �k  L   0 �h  �k  L    �h  �  �k  L    �	  x�  &�bi  ջ  &�#�k  �k  �  �&�l  R�  &   �  &�  )�  &�  ��  &�  2�  &�.   �� &�.  (��  &�  0��  &�  8R0  &�  @�  &�  P�!  &  `��  &�n  ��� &B  �b�  &B  ���  & B  ��  &"a   �L�  &#a   �_� &%Un  � ��  &��l  �l  �  m  �k  �   q�  &�m  m  8m  �k  �  �  a   j�  &�Em  Km  �  dm  �k  �  �   ��  &�qm  wm  �  �m  �k   *�  &�Em  �  &��m  �m  �m  �k   �  @&�0n  �� &�On   �Y &��m  �? &�$�l  kI &�$m  rL &�$8m   � &�$dm  (-1 &�$�m  0��  &�$�m  8 On  �k  �  �  �  B   0n  T�  &��m  	Un  a�  Z   &��n  ��   J�  �  ,�   ה  &�gn  ��  &'�k   �  &F�n  y�  &H@2   2�  &I@2  �� &J@2   ɠ  &L�n  ݬ  &L o  �n  �  &O/o  o  ��  �&}�p  <0 &�n   4� &��q  �#top &��'  �O� &��q  �Xc  &��n  x
s  &�E,  �
�  &��  �
V &�F2  �
Ğ  &��  �
��  &��  �
��  &�F2  �
h�  &�L2  �
��  &��1  �
��  &�k	  �
w�  &��  �
��  &��  �
�  &��  �
�  &��k  �
�  &��(  `&  &�  h�  &��p  p_� &��q  x�  &��'  ��  &��  ��J &�B  �˽  &��	  � �   &X�p  �� &[Rq   �Y &fcq  �; &o�q  � &u�q   �  &Tq  q  �  q  o  �   �  Rq  o  �  �  �  F2  �(  B    �p   q  cq  o   Xq  �  �q  o  @2  �   iq  �  �q  �q  @2  �   �k  �q  X�  &z�p  	�q  �  �q  L   � �n  �q  L    <�  &� �q  ��  �&�r  R�  &   �  &pN  )�  &$W  ��  &�  2�  &�.   �� &�.  (��  &�  0��  &�  8R0  &�  @�  & �  P�!  &"  `��  &$B  ��� &%B  �b�  &&B  ���  &(B  ��  &*a   �L�  &+a   �_� &-nt  � c�  &�s  
s  �  s  s  �   �q  ˯  &�1s  7s  Qs  s  �  �  a   N�  &�^s  ds  �  }s  s  �  �   Ԝ  &�^s  h�  &��s  �s  �s  s   8�  &��s  �s  �  �s  s   p�  @&�It  �� &�ht   �Y &��s  �? &�%�r  kI &�%$s  rL &�%Qs   � &�%�s  (-1 &�%}s  0��  &�%�s  8 ht  s  pN  �V  $W  B   It  +�  &��s  !�  &E�t  2�  &G@2   �� &H@2  y�  &I@2   ��  &K{t  j�  �&Nrv  <0 &P�q   cff &QF6  �4� &S}k  �#top &T�  hO� &Vrv  pXc  &W�v  ��  &Y�  �  &Z�  �  &[�k  
�  &]�  ���  &^�  ���  &`B  ��  &aB  ���  &b�  ��  &c�v  �z�  &e�  ��  &f�  ���  &h�  ��  &i�  �~�  &kF2  �9� &lF2  �V &nF2  ��  &o�  �&  &q  ��J &sB  ��  &u�;  ��  &w&	i  ���  &x&:i  � �t  �v  L    �t  �  �v  L    1�  &z�t  ��  &}0�v  	�v  �v  l�  &�v  �� &�/w   >'  &�Nw  � &��q   	�v  )w  )w  pN  �V  $W  B    	i  :i   �v  �v  �  Nw  )w  �V  �   5w  U�  &��v  	Tw  :�  &�#sw  yw  ,�  (&��w  R�  &�   Jy  &�cx  � &�y3  p�  &��x  o�  &�a     4�  &�x  �� &�%x   �Y &�6x  gP &�Kx   �  %x  fw    @2  @2   x  6x  fw   +x  �  Kx  fw   <x  \�  &��w  	Qx  ١  &�#px  vx  ��  �  �x  �  	  a    {x  �  &�.�x  �x  0�   &��x  ��  &�0"   �0 &�0"  ک  &�0"  �> &�0"   	�x  �  X&��y  b�  &!�y   �  &!�y  E�  &!�y  b�  &!�y  ,�  &�y   h�  &�y  (�  &�y  0��  &z  8c�  &�x  @:�  &! z  Hs�  &"&z  P �b  Dg  bn  �q  �y  @2  	  �   �y  r  �y  r   �y  �y  �q  a   B   �y  z  �  7'  �;   z  ^x  aw  ��  &9z  �x  ��  'Kz  Qz  �  oz  �  oz  oz  �^   �  ��  '$�z  �z  �  �z  �  �z   B  �  ''�z  �z  �  �z  �  �  L2   d�  '+�z  	�z  ��  '+{  �  '-/?z   N�  './uz  ��  '//�z   =�  (!{  ${  �  8{  �  �>   T�  (%D{  J{  �  ^{  �  ?   ��  ()j{  p{  �  {  �   �  (,�{  �{  �  �{  �  �{   +'  ��  (0�{  �{  �  �{  �   *  �  a   �   �  (7�{  	�{  ,�  ((7@|  ۽  (9{   1�  (:8{  G�  (;^{  #�  (<{  )�  (=�{    FO  ))�$  ��  ),]|  	L|  Y  ),x|  6 ).@|    	]|  �O  ),�|  x|  &I  *:�|  �8  *<�   ߣ  *=�   `K  *?�|  'B  *C�|  �|  �  �|  7  �|   �|  �  *G }  	�|  b:  *G}  '�  *I�|    	 }  SQ  *G,}  }  "�  +!>}  D}  �  S}  �   �  +$_}  e}  �  �}  F6  �;  �  �   �  +*�}  �}  a  �}  �>  �   ��  +.�}  �}  B  �}  )9  �  �  �   ��  +4�}  �}  �  	~  )9  �  �  �   ��  +:~  		~  9�  (+:i~  i�  +<$2}   (�  +=$S}  Z�  +>$�}  ��  +?$�}  ��  +@$�}    	~  R�  +:z~  i~  
�  ,�  ��  -'�~  �~  �  �~  �  �~   �G  jd  -+�~  �~  �  �~  �  �~   �~  �H  �g  -/�~  �~  �    �  �  �'   �{  -6!  '  �  @  �  �  �    l  -=�~  �n  -B!  �x  -Gd  j  �  ~  �  �   1j  -K�~  �}  -P�  �  �  �  �  L2  �  �  �~   �  ��  -W/  ��  -Z�  	�  �b  P-Zr�  h  -\�~   �v  -]�~  ��  -^@  ��  -_~  .�  -`�~   �  -a  (V�  -bL  0��  -cX  88�  -f�  @��  -g�  H 	�  h�  -Z��  r�  i  .'��  ��  �  ��  �  �  �^   4�  .,��  \�  .1��  �l  .8��  ~�  .=��  ŋ  .B��  �w  .G��  H�  .N/  �r  .Q�  	�  ȅ  @.Q��  ��  .S��   ��  .T��  �n  .U��  Rs  .W̀  ��  .X؀   F}  .Y�  (�|  .Z��  0��  .\��  8 	�  w�  .Q��  ��  f.  /&�$  <B  /,�$  %�  /0ρ  	��  �3  /0��  tW /2!��   i�  /3!��   	ρ  �?  /0�  ��  n)  0�   �  �  >�  �  �  �  B   �)  0$J�  P�  �  i�  �  �  a    nk  0)z�  	i�  �;  0)��  �=  0+�   z+ 0,>�   (��  �ʁ  	0gH     (��  F�{  	 gH     (��  uX|  	�fH     (�  ��|  	�fH     (��  (�z  	�fH     (��  9u�  	�fH     ("�  ��  	`fH     (f�  ��  	 fH     (��  �~  	�eH        ��  L   
 	q�  (��  ���  	 eH     )�~  N	`dH     �  ��  L   	 	��  *��  ���  	 dH     *��  ���  	�cH     oY   �  L   L 	��  (p�  # �  	 ZH     �  ,�  L   � 	�  *��  +,�  	 XH     �  W�  L   � 	G�  *�  LW�  	�VH     �  ��  L   V 	r�  *��  e��  	 VH     �  ��  L   � 	��  *^�  t��  	 TH     *��  ���  	 RH     +��  ��#B            ��  ,~ ��  U -B�  ��  `#B     x       �e�  ,~ ��  U.K1 �ha  =� ;� (ߢ  �r  �t /��  c�PB     �      ��  0��  c�  h� `� .�  e�V  ϸ Ǹ .R�  f  0� .� .$S  g�`  U� S� 1�PB     D      m�  2cff tF6  z� x� 3�  
QB       �  y	X�  4��  �� �� 5 �  6�  Ĺ ¹ 6�  � � 7o�  XQB       XQB            �		��  4��  %� #� 4}�  J� H� 8eQB     
 9U|   3w�  �QB      P�  �	Ȇ  4��  o� m�  3I�  �QB       ��  �	|�  4d�  �� �� 4W�  �� �� 5��  6q�  � � 3�  �QB      П  }f�  4��  	� � 4��  	� � 4��  1� /� 8�QB     " 9U}   8�QB     " 9U}    3o�  RB      �  �	͇  4��  Z� T� 4}�  �� �� 8$RB     
 9U| 9Ts�  3`�  $RB      @�  �	�  4{�  л λ 4n�  �� �� 8>RB     . 9Ts�&  :QB     �  1�  9Us� :&QB     �  J�  9Us�
 :/QB     �  b�  9Us8 :;QB     �  {�  9Us�
 :�QB     " ��  9U|  :RB     ��  ��  9Us�'9T|  :hRB     " ʈ  9U|  :�RB     " �  9U|  :�RB     " ��  9U|  :�RB     " �  9U|  :�RB     " *�  9U|  :�RB     " B�  9U|  8SB     " 9U|    83SB     " 9U~   7��  >SB      >SB            щ  4��  � � ;>SB            6��  C� A� <PSB     9Uv    <�PB     9Uv   -��  ��   iB     E&      �=�  0Jy  �!K  �� f� 0��  �!�  0� �� 0�  �!�  r� @� 0G  �!�  �� �� 0G  �!#  C� 1� .�  ��V  D� � .� ��  X� T� .$S  ��`  �� �� .s  �E,  � � .2�  ��0  �� �� .Q  �,z  � 
� .��  �n~  9� /� .��  �B  �� �� .�J  �B  �� Z� .K�  �B  e� Y� .k  ��  �� �� =�u  ]�xB     =��  <HxB     > �  ˋ  .~ �  i� g� .�O  	  �� �� 8|iB     ; 9T	�BH     9Q1  >`�  �  .~ �  � � .�O  	  >� 4� 8�iB     ; 9T	xQH     9Q1  >��  ��  2cff ]F6  �� �� .��  ^v;  L� H� .R�  _  �� �� .?1  ``  �� �� 2i a�  {� u� 1�qB     ]       �  2mm �'w�  �� �� 2var �'��  �� �� .� ��  .� *� ?rB     ��  9U} 9T~  <6rB     9U}   >P�  �  .:  �=�  r� h� .x  �  �� �� 2upm �4  �� |� ./� ��  � � :{B     H ��  9Ts  :{B     H ��  9Ts  ::{B     H ��  9Ts  :U{B     H ʍ  9Ts  :p{B     H �  9Ts  :�{B     H ��  9Ts  8�{B     H 9Ts   >��  ď  2sub v;  W� Q� 2top v;  �� �� .:  =�  �� �� .x  	  V� P� 2upm 
4  �� �� ./� �  �  � 1�rB     k       �  .C�  �  Q� O� :"sB     U �  9Uv 9T|� 9Q~  :2sB     b 
�  9U|� 9Tv 9Q~  8FsB     o 9Q~   :tB     H 7�  9T~  :'tB     H O�  9T~  :9tB     H g�  9T~  :KtB     H �  9T~  :]tB     H ��  9T~  :otB     H ��  9T~  8�tB     H 9T~   >��  ��  .A  M�   ~� t� 1|B     F       ��  .d> r�   �� �� 3ا  2|B      ��  w$z�  4��  � � 4�  >� :� 5��  @�  ��6�  x� v� 8:|B     | 9U��}9Q    8|B     ��  9U��}  > �  ��  .s�  ��   �� �� .X�  ��   �� �� .r? ��   �� |� 3ا  �}B      `�  �G�  4��  �� �� 4�  	� � 5`�  @�  ��6�  C� A� 8�}B     | 9U��}9Q    3C�  �}B      ��  ��  4^�  j� f� 4Q�  �� �� 5��  6k�  �� �� 6x�  �� �� A��  Ы  ��  6��  !� �  :�}B     � Α  9Us  8�}B     � 9U|    8%vB     ��  9U��}  >��  ��  .�  ��   �� �� 7ا  L}B      L}B            �$��  4��  � � 4�  5� 3� ;L}B            @�  ��6�  \� Z� 8\}B     | 9U��}9Q    8>}B     ��  9U��}  >0�  �  .��  ��   �� � 8�vB     ��  9U��}  3ا  �vB       �  �!f�  4��  �� �� 4�  �� �� 5 �  @�  ��6�  � � 8�vB     | 9U��}9T	�BH     9Q    7��  �|B      �|B     �       �ԓ  4��  =� 3� ;�|B     �       6��  �� �� 6��  X� V� 6ʧ  �� {�   8w|B     ��  9U��}9T��}�  >�  Ĕ  (��  c  ��.
H 7  � � 2nn �  �� v� .= �4  �� �� >@�  ��  .�M ?0"  7� 1� 8�xB     � 9U	�gH     9T09Q��9R0  8xB     � 9U	@gH     9T09Q��9R0  3&�  3kB      �  h��  4��  �� �� 4y�  .� ,� 4l�  t� R� 4_�  �� �� 4R�  y� W� 4E�  � �� 48�  �� �� 5�  @��  ��~6��  � � 6ı  Q� 3� 6ѱ  �� �� @ޱ  ��~6�  �� �� B��  ]qB     B�  �pB     A�  ��  �  @"�  ��6/�  ;� /� 6<�  �� �� 3��  nB       �  J	U�  4��  \� X� 4��  �� �� 4��  3� � 4��  f� `� 5�  6
�  �� �� @�  ��6$�  �� i� 61�  �� �� 6<�  �� �� BG�  BnB     AP�  P�  �  6Q�  � � 6^�  m� k� 6k�  �� �� Cx�  r�B     �       ��  6}�  �� �� C��  ��B     �       k�  6��  %� #� 6��  J� H� 6��  q� o� 6��  �� �� :͌B     � 2�  9Us 9T  :�B     � P�  9Us 9T  8�B     � 9Us 9T   8��B     � 9U��}9TH9Q09X09Y   C��  6�B           Z�  6��  �� �� :`�B     � ՗  9Us  :|�B     � �  9Us 9T4 :��B     � �  9Us 9T  :͎B     � ?�  9U��}9T49Q09X09Y  8��B     � 9U| 9T   :}B     � r�  9Us  :�B     � ��  9Us 9T2 :�B     � ��  9Us  :�B     � Ř  9Us 9T  :��B     � �  9Us 9T  :ۊB     � �  9Us 9T  :�B     � 6�  9U��}9T89Q��}9X��}9Y  :W�B     � T�  9U} 9T  :��B     � y�  9Us 9T	��~��~" :ЋB     � ��  9Us 9T  :��B     � ��  9Us 9T  :-�B     � �  9U��}9T89Q09X09Y  8��B     � 9U��}9T@9Q09X09Y   :VnB     " 2�  9U��}9T��} 8GB     ��  9U��}#�'9T��}   3��  �oB       ��  �	]�  4�  �� �� 4�  � � 4��  a� ]� 4��  �� �� 5��  @&�  ��~63�  �� �� 6@�  � � BM�  �pB     BV�  {pB     :�oB     � ��  9Us  :
pB     � �  9Us 9T��~ :TpB     � <�  9Us 9T��~ 8�pB     � 9Us 9Q��}#�&   :�nB     � u�  9Us  :�nB     ��  ��  9U 9Ts 9Q09R��~� :oB     � ԛ  9U��}9T
�9Q09X09Y��} :�oB     ��   �  9T 9R| 9X��}9Y~  8�pB     �  9U   C
�   yB     R       X�  6�  [� Y� 8yB     � 9Us 9T��}  AJ�  Ш  [�  6K�  �� ~� 3��  x�B        �  �	g�  4��  �� �� 4��  �� �� 4��  >� 0� 4��  �� �� 4��  w� o� 4��  �� �� 5 �  6��  �� �� @��  ��6�  �� �� B�  ^�B     A!�  `�  o�  6"�  =� 3� C-�  ͇B     �       ��  6.�  �� �� 6;�  � � :�B     � {�  9Us 9T  :�B     � ��  9Us 9T  Dh�B     �  :3�B     � ��  9Us  :Z�B     � ݝ  9Us 9T  :��B     � �  9U��}9T29Q09R| ����9X09Y  :ՉB     	 B�  9Us 9T|����1$���� :�B      Z�  9U}  84�B     # 9Us   :߀B     � ��  9U��}9T29Q09Rv 9X09Y�� :R�B     ��  ͞  9U��}9T| 9Q��} :��B     � �  9U��}9T29Q09Rv 9X09Y�� :��B     " �  9U  :��B     " 3�  9U  8~�B     � 9U��}9T29Q09Rv 9X09Y��   E\�  ��B       ��  �	4��  Y� O� 4��  �� �� 4��  W� O� 4��  �� �� F{�  4n�  !� � 5��  @��  ��6ɺ  �� �� 6ֺ  �  �  6�  � � 6�  � � B��  /�B     B�  D�B     AZ�  �  ��  6[�  � � 6h�     G��  ��B      ��B            'F��  F��  4��  w q ;��B            6��  � �    C�  '�B           �  6#�    60�  > 6 6;�  � � :_�B     �  �  9Us 9T  8�B     � 9Us 9T   AG�   �  ��  6L�  � � :I�B     � S�  9Us 9T  :��B     � q�  9Us 9T  8��B     � 9Us 9T   C�  �B     ~       �  6�    :�B     	 ӡ  9Us 9Tv � 8i�B     # 9Us   :e�B     ��  �  9U��}9T|  :��B     �  �  9Us  :ЃB     � >�  9Us 9T  8��B     � 9Us 9T     :�kB     � s�  9Us  :�kB     0 ��  9Us 9T	�QH     9Q��} :lB     � ��  9Us 9T��} :HlB     � آ  9Us  :�lB     � �  9Us  :�lB     � �  9Us  :�lB     ��  2�  9U��~9Ts 9Q19R1 :�mB     ��  ��  9U��}#�9Tv 9Q��~�9Rs 9X 9Y	�0| �0)(  �#�` :�mB     � ��  9Us  :�mB     ��  ͣ  9U��}#�
9Ts 9Q09R��~� :�pB     �  �  9U��} :lqB     �  �  9U��} :�xB     �  �  9U��} :hyB     � 3�  9Us  :�yB     ��  _�  9U��}#89Ts 9Q09R0 :�yB     ��  ��  9Uv 9Ts 9Q09R0 :zB     ��  ��  9U��}9Ts 9Q19R0 :@zB     ��  ۤ  9U��~9Ts 9Q19R0 :szB     h�  �  9U��}9T��}#�9Q��}#�9R��}#� :�~B     �  0�  9U��} :,�B     h�  _�  9U��~9T��}#�9Q09R0 8��B     ��  9U��}9T��~�   8kB     = 9U��}9T
�9Q��~  :ZiB     I ʥ  9Uv 9T	�1H      :�iB     I �  9Uv 9T	`BH      :�iB     I �  9Uv 9T	�BH      :�iB     � 1�  9Us 9T0 ?�iB     a�  9Us 9T} 9Q~ 9Rw �9X��} ?=jB     ��  9U} 9Tdaeh9Qs 9R0 ?WjB     ��  9U} 9Ts  ?}jB     ˦  9U} 9T2FFC9Qs 9R0 :�jB     � �  9Us 9T0 ?&qB     �  9Us 9T} 9Q~ 9Rw �9X��} <�tB     9U} 9T FFC9Qs 9R0  k	  H��  ���  Id> �#  IA  �#  J��  �`  J�  �#`  KLidx ��    Hy�  �ا  IF@ �%  Lidx �`  Jss  �`  J��  �B   M7�  �  �  IR�  �!  I�% �!  J� ��  JE  �   N��  f�  �$B     T       ��  0 f �  � � .�  h�V  � � .v�  iF6  J F .2�  j�0  � � ;�$B     .       .~ o�  � � 1%B            �  ._� v�.  � �  8%B     V 9T	`BH        +��  _P#B            �3�  , _ �  U -�  �  @;B     D      ���  0�  &�  � � Oreq &�  z p .V�  �V  � � ._� .-  r n >��  �  .��  �V  � � .$S  �`  � � (-U  �  ��?o;B     	�  9Ts 9Q�� 8u<B     ��  9Uv   1�;B     �       a�  .��  1�V  � � .v�  2F6  	 	 .�8  3oW  A	 ?	 .S�  5�  f	 d	 2i 6�  �	 �	 >��  L�  2sub ?�;  �	 �	 .�  @�  �	 �	 .�� A�  H
 @
 .�� A�  �
 �
 :�;B     o �  9T| 9Q�� :<B     o 7�  9T| 9Q�� </<B     9R09X0  <�;B     9R09X0  :�;B     c y�  9Ts  8�;B     � P��  v   QA�  ��  �9B     �       �l�  R�  ��  �
 �
 R-U ��  5 1 SV�  ��V  t n S_� �.-  � � 1�9B     �       <�  S�  ��V  � � Sv�  �F6  "   S�8  �oW  G E SS�  ��  l j Ti ��  � � >�  '�  Tsub ��;  � � S�  ��  � � S�� ��  N F S�� ��  � � :;:B     o �  9T| 9Q�� :S:B     o �  9T| 9Q�� <o:B     9R09X0  <:B     9R09X0  :�9B     p U�  9T�T 8�9B     � P��  v   Q)�  ��  �<B     >      �&�  RV�  ��  � � S�  ��V  T L *� ��  ��}S_� �.-  � � U�u  ��=B     >��  �  S�  ��V  . , Sv�  �F6  W Q S�8  �oW  � � *��  �+'  ��}SR�  �  5 3 Ti ��  Z X 1j=B     C       ��  Tsub ��;   } :|=B     &�  ��  9Tt  <�=B     9T��}9Q s "  :�<B     = �  9T
9Q��} :!=B     &�   �  9U}�9Tt  <8=B     9T��}9Q   D�<B     �  V��  v@%B     �      ���  R��  v'�;  � � W��  w'7'  TS��  y:>  � � Tn z�  G # S.� z�  � �  X��  S�:B     �       ���  RV�  S�  S M SR�  U  � � S�  V�V  � � S�  W�V    Sv�  XF6  C A S�8  YoW  s k 5@�  S_� ^.-  � � 1�:B     -       x�  Ti d�   
  :�:B     � ��  P��  �U Y&;B     "   Z/�  B.-  �  [�  B)�V  \�  D�V  \v�  EF6  \2�  F�0  \~ G�   H��  �	&�  Iv�  �	F6  JR�  �	  Lidx �	�   M��  g�  Z�  Ik  g�  IJy  hK  I�  i�  Iv�  jF6  I�  k�V  I��  lB  I�J  mB  (R�  o"j�  	�QH     J� {�  JR�  |  J��  }�  J��  ~v;  J��  4  J��  ��  ]�u  �	]��  �	^�  Jc�  �a   ^J�  Jn�  C	4  Lsub D	�;  Lidx E	�   KJ��  �	B    �\  j�  L    	Z�  H��  W��  IR�  W"  I��  X"�;   N'�  ��   eB     �      �f�  0��  �"�;  N F Oidx �" 4  � � 0��  �"�  � � 0Jy  �"K  S K 0��  �"�  � � 0� �"�  ; 5 0v�  �"F6  � � 0�  �"�V  � � .� ��  +  (�  �pX  ��~(��  �@2  ��~(��  ��  ��~2top �v;  � � .��  �:>  < 4 .Q  �,z  � � .�J  �B    .�m  ��  f \ =�u  OgB     1�hB     A       P�  .K1 ha     3 �  �eB       ��  �K�  4y�  = 9 4m�  = 9 4a�  { u 4U�  � � 4I�    4=�  k c 41�  � � 5��  6��    @��  ��~B��  gB     :�eB     � 5�  9U} 9T89Q09R	�0s  $0)( 
�#`9X09Y��~ 8gB     " 9U}    3��  �fB      �  �ŵ  4��  M I 4��  M I 4��  � � _��  �hB            6��  � � 8�hB     . 9T}    7��  gB      gB            P3�  4�  � � 4�  � � ;gB            6�      D)gB     "   :�fB     ��  a�  9Uv 9T��~�9Q} 9R��~ :LgB     � y�  9U|  :ggB     � ��  9U| 9Q}  :�gB     *�  ��  9U��~ :�gB     . ζ  9U| 9T}  :�gB     f�  ��  9U� 9T~ 9Q09R0 :YhB     � �  9U|  :�hB     ��  @�  9Uv 9T| 9Q19R
s  $0)� 8�hB     h�  9Uv 9T~�	9Q09R0  -$�  I�  �XB     �      �\�  0v�  I'F6  =  3  0��  J'�;  �  �  0ݺ  K'�  R! D! ONDV L'�  " �! .� N�  �" �" (�  OpX  ��2top Pv;  �# �# .��  Q:>  :$ .$ .Jy  RK  �$ �$ .�m  S�  (% $% =w\  ��XB     =�u  �IZB     3 �  �YB      P�  p
[�  4y�  d% `% 4m�  �% �% 4a�  �% �% 4U�  & & 4I�  X& P& 4=�  �& �& 41�  '  ' 5��  6��  D' @' @��  ��~B��  �ZB     :�YB     � E�  9U~ 9T89Q09X09Y��~ 8�ZB     " 9U~    7��  IZB      IZB            ���  4��  |' z'  7��  eZB      eZB            ���  4�  �' �' 4�  �' �' ;eZB            6�  �' �' DrZB     "   :$ZB     � �  9Us  ::ZB     	 .�  9Us  :�ZB     *�  G�  9U�� 8�ZB     # 9Us   M�  R�  w�  I= R$�4  I��  S$5  I�  T$�  IJy  U$K  I��  V$�  Ix  W$�  J� Y�  J.� Z�  Lj [�  J�  \�  J[�  ]�  ]�u  =]x�  ^�  Lp �@2   ^G�  J��  ��  Li ��  Lk ��   ^Z�  Jn�  ��   KLsid "�  Lgid #�    H��  I��  I= I$�4   H��  <��  I�  <�V  Lmm >w�   -4�  *�   #B     
       ���  0�  *#�V  �' �' 0�u  +#L2  0( ,( 0�  ,#�  m( i( 0�  -#�  �( �( 02�  .#�~  �( �( 2mm 0w�  ")  ) `*#B     9U�U9T�T9Q�Q9R�R9X�X  -��  B   .B     ;       �%�  0�  &)9  K) G) 0��  &�  �) �) 0ݺ  &�  �) �) ONDV &�  * �) 8Q.B     } 9U�R9Q�Q����3$  -��  k�  `.B     �      ���  0�  k&)9  G* ;* 0��  l&�  �* �* 0ݺ  m&�  @+ 8+ ONDV n&�  �+ �+ .� p�  , 
, .R�  q  4, 0, 2len s�  t, l, 2vs t46  �, �, .k  u6  "- - .��  v�  f- Z- =�u  
�/B     >@�  �  2j ��  �- �- 2idx ��  . . .i�  �"6  Q. M. 5��  .dh  ��5  �. �. .�{  ��  / / 7� d0B       d0B     $       ��  F� 4� B/ @/ ;d0B     $       6� j/ f/ 6� �/ �/   D�0B     H   :/B     � B�  9U��9T19Rs 2$9Y�� :1B     � n�  9U��9T19Rs 9Y�� 8+1B     � 9T��9Qs   M��   �  ��  I��   #�;  I�  #|X  I��  #�  J� �  J2�  �  Li �  Lj �  J�  �  J�  	)9  JR�    J� �  J��  �  J.� �  ]�u  a^��  J��  !@2  Jo�  "@2  KJx  4	  Lp 5F2    KJ��  F��  Lsum Gr    m  H��  ���  I��  �!�;   M��  a�  ��  Iʞ  a$��  IJy  b$K  I��  c$�  Ix  d$�  JR�  f  J� g�  J|�  i4  Li j�  Lj j�  ]�u  �KJ��  p�  Jߣ  q�  J^�  r�  ^��  J1�  �"6  KJdh  ��5  J�  �5  J��  �5  Ja�  �&5    KJ�U  �6     (6  +��  D $B     �       ���  0ʞ  D$��  �/ �/ 0R�  E$  @0 :0 2i G�  �0 �0 :Z$B     " L�  9U}  :s$B     " d�  9U}  :�$B     " |�  9U}  8�$B     " 9U}   M��  ��  I�  I��  �"5  I�  �"�  IJy  �"K  I��  �"�  Ix  �"�  I��  �"B  JR�  �  J� ��  J�  ��  ]�u  4KLj ��  KJ��  ��  Li ��     H��  w�  I��  w"5  IJy  x"K  JR�  z   H��  n��  I��  n'5  IR�  o'   M[�  `�  ��  I��  `+5  acid a+�  JE  c�   -E�  ;�  0-B     �       ��  0��  ;*5  T1 J1 0�  <*�  �1 �1 0R�  =*  N2 B2 (� ?�  �\2i @�  �2 �2 2j A�  3 3 .Ӷ  B�  =3 73 =�u  Z0-B     :�-B     � ��  9U�Q9T29Q09Rs 
��#9X09Y�\ 8.B     � 9U�Q9T29Qs 9R19Xs 9Y�\  -V�  �a  @"B     �       ���  ,��  �$�>  U,�^ �$�  T2fd �a  �3 �3 =�u  -X"B     5�  2p 
@2  '4 4 .3o  @2  �4 �4 2fd2 a  5 �4 .N� �  k5 a5 .�� �  �5 �5   M?�  ��  `�  I��  �%�>  I�  �%�  IJy  �%K  Ix  �%�  J� ��  Jߣ  �a  J5�  ��  ]�u  �]��  � H��  ���  I��  �%�>  IJy  �%K   M��  �  ��  Iv�  �'F6  asid �'�   Mu�  �  ��  Iv�  �#F6  I��  �#�   -��  c  0@B     �       ���  0v�  c!F6  c6 S6 0��  d!�  7 7 2idx f 4  c7 Q7 .R�  g  98 78 (Ӏ h@2  �P(�  i�  �X(� j�  �L.F@ k  l8 \8 =�u  �@B     3��  �@B      `�  }*�  4��  9 9 4��  �9 �9 4��  : �9 _��  �@B            6��  f: d: 8�@B     . 9T�P   :Y@B     ��  U�  9Us89T�T9Q�P9R�X :w@B     = s�  9Uv 9Q�L 8�@B     � 9Uv   H�  T��  aidx T( 4  IqI  U(F2  KJJy  YK    -��  ��  0>B     �      �h�  Oidx �( 4  �: �: 0��  �(�  (; ; 0qI  �(F2  �; �; 0Q�  �(4  M< C< .� ��  �< �< =�u  NT>B     5 �  .Jy  �K  �< �< .ti ��  @= 8= .Ϭ ��  �= �= 1H?B     �       .�  2pos �  n> l> :i?B     � ��  9U  :�?B      
�  9T} 9Q��P��  s  8�?B      9T} 9Q��P��  s   :�?B     � F�  9U  8@B     � 9U 9Tv 9Q~    -<�  ��  01B           �u�  Oidx �' 4  �> �> 0>) �'u�  ? ? 0�� �'F2  �? �? 0��  �'4  j@ ^@ (� ��  ��.R�  �  �@ �@ 2t �F2  gA UA .W�  �@2  =B -B .6^  ��  �B �B =�u  �3B     >��  ��  2n ��  JC <C .T�  ��  �C �C .5$  ��  �D �D .��  �@2  YE SE 5 �  .��  ��  �E �E Dr2B     �   3{�  3B      p�  ��  4��  #F F 5p�  @��  ��6��  �F F 6��  �F �F B��  >4B     A��  И  �  6��  QG GG 6��  �G �G 6��  �H �H 6��  �I �I 6��  aJ IJ :L3B     � ��  9U| 9T89Q09Rv 9X09Y�� :�3B     � ��  9U  :�3B     	 ��  9U 9Tv  8>4B     # 9U   8u3B     " 9U|    :�1B     � Q�  9U| 9T89Q09R}����9X09Y�� 8�1B     = 9U| 9T��9Q��  F2  M�  V�  �  aidx V& 4  J� X�  JJy  YK  JR�  Z  ]�u  �KJ��  _a  J
�  `�  Lp a@2  J��  b@2  J	�  c4    +�  D�&B     Q       ���  Oidx D 4  |K tK 5 �  .Jy  HK  �K �K .R�  I  L  L :�&B     . ��  9Ts8 8'B     " 9Uv    Q��  ��  �@B     �      �v�  bidx � 4  5L %L RJy  �K  �L �L R��  �B  �M �M R�J  �B  �M �M *� ��  ��SR�  �  >N 6N S.� ��  �N �N =�u  ;aBB     >��  �  .��  	a  2O .O .�  
�  sO iO :�AB     � ��  9Uv 9T  :BB     � ��  9Uv  :/BB      ��  9Ts9Q P��  s  :]BB     � �  9Uv 9Qs8 8�BB     � 9Uv   :6AB     � 2�  9Uv  :JAB     � P�  9Uv 9T  :�AB     " h�  9U}  D�AB     �  Z��  ��  ��  cidx �% 4  [��  �%��  \� ��  \Jy  �K  dtmp ���  \E  ��  Kdnn ��    �  a  ��  L    Qe�  ��   "B            �*�  R�j �'�  �O �O  -��  �  0UB     �      �	�  0�  |X  :P .P 0�S @2  �P �P 0�� @2  Q �P 2p @2  �Q PQ .� �  �S ~S .k  �  �S �S =զ  �VVB     =�u  �VVB     ]��  �]��  �=��  �VB     =�Y ��VB     5P�  2v *�  'T T 5��  .� �#�  �U �U .��  �#�  PV @V .�F �#	�  EW 7W 5 �  2val ��  �W �W 2q �@2  �X {X 1pWB     �       �  .��  I@2  �X �X .�U  LF2  5Y 1Y 8�WB     > 9U��P[�  | Ph�  }   7��  �VB      �VB            x�  4��  nY lY 4��  �Y �Y 4��  �Y �Y 8�VB     �
 9Q3P�  |   7��  �VB      �VB            ��  4��  �Y �Y 4��  Z Z 8 WB     �
 9Q0P�  |   ?WB     ��  9U|  8;WB     > 9U|P[�  |      oY  -��  ��  �[B     7       ���  0�  �#|X  0Z (Z .��  �v;  �Z �Z .�U  �F2  �Z �Z .� ��  R[ N[ =�u  ��[B     8�[B     > 9U�U#P[�  �U  -s�  ��  @]B     ^      ���  0�  � |X  �[ �[ .��  �:>  9\ 3\ .��  ��;  �\ �\ .�  �)9  �\ �\ .��  ��  A] ?] .� ��  j] d] =�u  ��_B     3��  �]B      `�  �(�  4��  �] �] 4��  �] �] 4��  D^ >^ 5`�  6Ŀ  �^ �^ 6ѿ  b_ `_ 6޿  �_ �_ 6�  �_ �_ 6��  1` )` 6�  �` �` 6�  �` �` @�  ��6(�  ,a (a 65�  fa ba BB�  �_B     A��  ��  ��  6��  �a �a 6��  
b b :n^B     > ��  9U| P[�    8�^B     > 9U| P[�     _K�  �_B     �       6P�  lb hb 6]�  �b �b Cj�  S`B     E       �  6k�  �b �b 6x�  	c c  8`B     � 9T19X��9Y��    :�]B     ��  R�  9Us 9Tv 9Q| 9R}  :�]B     %�  |�  9Us 9Tv 9Q| 9R}  8�]B     > 9U| P[�     -��  l�  @[B     G       �W�  0�  l"|X  Hc @c .��  o:>  �c �c .�U  pF2  d �c .�  q)9  hd fd .� r�  �d �d =�u  �V[B     8t[B     > 9U�U#P[�  �U  -e�  L�  �[B     b       �C�  0�  L"|X  �d �d .��  Nv;  
e e .�U  OF2  4e .e .� P�  �e �e :�[B     > ��  9Us P[�  spPh�  v  :\B     > �  9Us P[�  spPh�  v 8#\B     > 9Us P[�  spPh�  v  -��  �  @\B     q       ���  0�  *|X  �e �e .��  v;  f f .�  �  8f 6f 5�  .m�  2�  af ]f 8q\B     > 9Us   -g�  ��  �\B     r       ���  0�  �'|X  �f �f .��  �v;  �f �f .�U  �F2  g g .� ��  �g �g =�0  �\B     5 �  2tmp ��  �g �g :�\B     > ��  9Us P[�  spPh�  v  8]B     > 9Us P[�  spPh�  v   -1�  ��  TB     �       ���  0�  �$|X  Oh Ih .��  �v;  �h �h .�!  ��  �h �h .�U  �F2  �h �h .� ��  Zi Vi 7��  /TB      /TB            ���  4��  �i �i 4��  j �i 8ATB     �
 9Q0P�  s P�  v   3��  [TB      ��  ��  4��  =j 7j 4��  �j �j 8`TB     �
 9Q0P�  s P�  v  3��  zTB      �  �h�  4��  �j �j 4��  �j �j 8TB     �
 9Q0P�  s P�  v  3��  �TB       �  ���  4��  k k 4��  =k ;k 8�TB     �
 9Q0P�  s P�  v  DITB     � DhTB     � D�TB     � D�TB     �  -B�  Y�  �`B     U      �"�  0�  Y&|X  lk `k .��  [v;  �k �k .:  \=�  l l .x  ]  Fl Dl 2upm ^4  pl nl .�U  _F2  �l �l .� `�  �m �m =�u  ��`B     5У  (�D e"�  ��~(0�  f2�  ��.��  h�  �m �m .G�  h�  _n Un 2i iS   �n �n >��  j�  .�\ ��  o  o .��  ��  �o �o .��  ��  3p #p  EB�  �aB      �  {4T�  �p �p Fl�  4a�  oq gq Ay�  `�   �  6z�  �q �q 6��  jr Xr DbaB     H :�aB     ��  ��  9Uu 9Tt  D�aB     H  8dcB     t�  9Q09R� ~ "p    �  2�  L    �  B�  L    M��  .�  ��  I�  .(|X  ad /(F2  IC�  0(�'  KJ��  8�  Jf�  9�    M��  "�  ��  I�  "'|X  ad #'F2  IC�  $'�   M�  �  ��  I�   |X  ad  F2   M��  ��  I�  I�  �|X  ad �F2  IC�  ��  ](�  KLval ��    M�  ��  t�  I�  �|X  ad �F2   Qr�  ��   (B     �      ���  R�S �@2  2s .s R�� �@2  �s ks Rb�  ��  �t �t RC�  ��'  (u  u Tp �@2  �u �u Tnib ��  !v v S t  ��  �v �v SE  ��  �w �w S��  ��  y �x ST�  ��  �z �z S�b ��  �{ �{ e��  ��   S��  �,�  j| \| S��  ��  } } Sf�  ��  �} �} S��  �-�  ~ �} fBad ��(B     =�u  ��(B     =��  ��(B     =(�  ��(B     1c)B     R       Q�  .��  Y�  �  .�� Y+�  � �  D+B     H D�+B     H :�+B     H ��  9T: D�+B     H  Z�  \�  ��  [�S \ @2  [�� ] @2  dp _@2  dv `�  dval a�  gBad ��5B     U�u  ��5B      h��  Q �  [�  Q |X  \R�  S   Z^�  *�  ��  [�  * |X  [� + �  [ݰ  , a   [k  - �  [�m  . �  [m�  / �  [�m  0 �  \R�  2  \� 3�  i�u  K Q	�  ��  PCB     �
      ���  R)�  �!$W  � � R�  �!�V  J� 0� R�^ �!�  m� ]� R:1  �!`  -� � S� ��  �� �� *�3 ��v  ��s*A�  ��k  ��iS�  �pN  :� 0� SZy  �B  �� �� S��  �B  _� W� S=�  �#B  � ц Tcff �F6  � � SQ  �,z  p� h� Se�  ��v  ܈ Ԉ *��  �k	  ��iSw�  ��  \� L� ] �  �> �  �  S�  ��V  G� A� S$S  ��`  �� �� SJy  �K  � � 5 �  (N �K  ��s>`�  ��  .��  B  N� H� (�  �  ��i(��  �  ��i?�HB     ��  9U~ 9T09Q} 9R��i9X��i <MIB     9U~ 9T19Q} 9R��i9X��i  <	HB     9U~ 9Q} 9Rv 9Ys�   >p�  ��  .S�  d�  �� �� .�  d�  ڋ ֋ .n�  ea  � � :/GB     �  ��  9Uu 9T}  :�GB     o ��  9T��h9Q��i 8�GB     o 9T��h9Q��i  >��  �  (ٶ �@2  ��i(��  ��  ��i1�MB     6       �  .��  � 4  P� N�  ?EB     J�  9U��s9T~ 9Q| 9Rs 9Yv @&? :DEB     "�  v�  9U~ 9T} 9Q��i9R��i ?eEB     ��  9U��s9T| 9Q}  ?�EB     ��  9U��i9T��s9Q0 ?�EB     ��  9U��i :�EB     ��  ��  9U~ 9T��i ?FB     �  9U��s <�IB     9U��i  >@�  J�  (N �"�   ��i<�FB     9T} 9Q09R��i  1�FB     I       u�  .�8  h  x� v�  1�IB     �      x�  (C!  #  ��i.N $��  �� �� .��  %B  Ȍ  >��  �  (~  *�  ��i(�  +�  ��i<�IB     9U~ 9T09Q} 9R��i9X��i  >Н  p�  (B  E�  ��i(�  F�  ��i<pJB     9U~ 9T 9Q} 9R��i9X��i  >��  U�  2n ~�  � � 2cur �.  E� A� 2vec �  �� �� .�� ��  �  � .�� ��  B� >� 7� �KB      �KB            �"F�  F� 4� ~� |� ;�KB            6� �� �� 6� � �   7� �KB      �KB            �"��  F� 4� '� %� ;�KB            6� P� L� 6� �� ��   3� �LB      ��  ���  F� 4� ҏ Ώ 5��  6� � 
� 6� Q� M�   G� �LB      �LB            �F� F� ;�LB            6� �� �� 6� Ӑ ϐ    3� �JB       �  k"��  4� � � 4� 7� 5� 5 �  6� `� \� 6� �� ��   3� KB      `�  m"�  4� �� ޑ 4� � � 5`�  6� 0� ,� 6� s� o�   :�JB     �  �  9U| 9T��i :`KB     � D�  9U| 9T~ 9Q}  :�KB     � c�  9U| 9T��i 8;MB     � 9Us0  j��  �CB      Л  �4��  �� �� 4��  �� �� 4��  �� � 5Л  6��  C� =�    Q  h��  Q"�  [�  Q#pN  [m  R#F2  [ss  S#�  ^�  \�U  ^�	   Kdcff kF6    Z��  -�  ��  [�  -"pN  [�^ ."�  [m  /"F2  [ss  0"4  ^��  \�U  7�	  \� 8�   Kdcff GF6    M��  !  ��  IK1 !#�  I;  "#�  Jk  $�  J$S  %�  JE  &   +��  �"B     
       �?�  0�  �!�V  �� �� 2var �#��  ͓ ˓ `"B     9U�U  -��  ��   "B     	       ���  0�  �"�V  �� � 0n�  �"�  3� /� 0"c  �"�^  p� l� 2var �#��  �� �� `	"B     9U�U9T�T9Q�Q  -��  ��  �!B     
       �P�  0�  ��V  Ԕ Д 0� ��  � � 2mm �w�  L� J� `�!B     9U�U9T�T  -R�  w�  �!B     
       ���  0�  w"�V  u� q� 0�u  x"�  �� �� 0�  y"�  � � 2mm {w�  *� (� `�!B     9U�U9T�T9Q�Q  -��  k�  �!B     
       �|�  0�  k"�V  S� O� 0�u  l"�  �� �� 0�  m"�  ͖ ɖ 2mm ow�  � � `�!B     9U�U9T�T9Q�Q  -*�  `�  �!B     
       ���  0�  ` �V  1� -� 0��  a �~  n� j� 2mm cw�  �� �� `�!B     9U�U9T�T  -��  T�  �!B     
       ���  0�  T �V  җ Η 0�u  U �  � � 0�  V �  L� H� 2mm Xw�  �� �� `�!B     9U�U9T�T9Q�Q  -C�  H�  �!B     
       �"�  0�  H �V  �� �� 0�u  I �  � � 0�  J �  *� &� 2mm Lw�  e� c� `�!B     9U�U9T�T9Q�Q  -u�  �  P!B     A       ���  ,�  +�V  U,�^ +�  Tkcid +L2  Ql� �   2cff F6  �� �� =�0  #t!B     5��  2c �  � ۙ .��  v;  �� ��   -8�  ��   !B     !       �a�  ,�  ��V  U,R�  ��z  Tl� ��   2cff �F6  ͚ ˚ ;/!B            .��  �v;  � �   -��  ��  `6B     �       �[�  0�  ��V  � � 0d�  �oz  _� U� 0|�  �oz  ۛ ћ 0�  ��^  W� M� .� ��  Ϝ ɜ 2cff �F6  � � =�0  ��6B     5p�  .��  �v;  Y� U� :�6B     ��  E�  9Us  87B     ��  9Us    -��  ��  0'B     ~       ���  0�� �$7  �� �� 0+�  �$�|  L� >� .
H ��!  �� � l� ��   .�  ��  �� �� .k  ��  П ̟ 5P�  .$S  ��  � � .YM  � }  =� ;� :h'B     V C�  9T	�1H      :w'B     ; g�  9T	v.H     9Q0 `�'B     9U�U9T�T   -��  Y�  �'B     o       �}�  0�  Y�V  l� `� 2cff [F6  �� �� .$S  \�`  4� .� 5��  .k  d�  �� �� .�  e�  �� �� .YM  f}|  С Ρ :�'B     V F�  9T	�1H      :(B     ; j�  9T	V.H     9Q0 `(B     9U�U   -��  ��  @8B            �)�  0�  �,�V  �� � 0��  �,?  g� ]� 2cff �F6  ݢ ٢ (� ��  �L=�0  A@8B     ;�8B     �       .��  v;  � � .8�  ?  A� ;� .R�    �� �� .g�    ɣ ǣ >��  ��  .�    � � .��    ,� (� >��  ��  2s   f� b�  :�8B     � ��  9T	pQH      8�8B     � 9U} 9T	�1H       :�8B     = �  9T29Q�L 8�8B     ��  9U|    -��  ��  7B     &      ���  0�  �*�V  �� �� 0ù  �*�>  � � 2cff �F6  q� m� (� ��  �\=�0  �7B     ;p7B     �       .��  �v;  �� �� .�  ��>  ե ϥ .R�  �  #� � :�7B     = �  9T89Q�\ :�7B     ��  2�  9U|  :�7B     ��  J�  9U|  :�7B     ��  b�  9U|  :�7B     ��  z�  9U|  8�7B     ��  9U|    -��  ��  !B     
       ���  ,�  �$�  U Nu�  y�   ,B     
      ���  0�  y#�V  k� [� 0la z#  (� � 2cff |F6  �� �� .��  }5  � � .s  ~E,  .� *� .F@   h� d� 2sid ��  �� �� 2i ��  � � >�  0�  .k  ��  S� O� .�  ��  �� �� .YM  ���  �� �� :�,B     V ��  9T	�1H      :�,B     ; �  9T	K.H     9Q0 `*-B     9U�U9T�T  1I,B            ��  .~ ��  ֩ ԩ .�O  �	  �� �� 8X,B     ; 9T	�BH     9Q1  7��  ~,B       ~,B            ���  4��  7� 5� 4��  7� 5� 4��  \� Z�  8�,B     � 9Us   M4�  6�  ��  I�  6#�V  I�^ 7#�  IB� 8#	  I(5  9#�  Jv�  ;F6  J��  <  Lsid =�  J� >�  ]�u  sKJk  E�  J�  F�  JYM  G��    Q��  ��  �NB     �      �W�  R�  � �  �� � R�S � �  K� =� R.� � �  �� � R?1  � `  �� �� R\-  � �  7� )� Tnn ��  � խ S� ��  �� � S ��  � �� =�  XOB     >�  6�  Se5  �pN  �� x� *��  ��  ��1OB     .       ��  mah ��  ��<-OB     9U| 9T19Qs9R} 9X~   ; PB     +       naw 
�  ��<"PB     9U| 9T09Qs9R} 9X~    8�OB     W�  9U 9Qs 9R}   Q��  ��  0NB     V       �\�  R��  �!�  � ܯ RV�  �!�  �� �� R�^ �!�  B� 4� R:1  �!`  � � *� ��  PS �$W  �� �� S�  ��V  H� :� oMNB     ��  -�  9U�U9T�T9Q�Q9R�R oWNB     ��  D�  9T0 phNB     ��  9R�R3!  Qx�  m�  � B     3       �  Re5  m �  � � R�U  n �  >� 8� RB7  o �  �� �� RY�  p   � ܴ S�  rpN  I� C� S$S  s�`  �� �� <� B     9U�U9T�T9Q�Q  Q��  �r  � B            ��  RyW �,�*  � � R��  �,r#  '� #� S�  �pN  b� `� Tcff �F6  �� �� Ss  �E,  �� �� `� B     9U�U9T�T  Q]�  ��  � B            �T RyW �-�*  � ޶ R��  �-r  � � S�  �pN  Z� X� Tcff �F6  �� ~� Ss  �E,  �� �� `� B     9U�U9T�T  V@�  ��#B     (       �� RyW �'�*  ܷ ַ S�  ��  *� (� SR�  �  P� N� D$B     "  Qt�  ��  @ B     F       �� RyW �'�*  �� x� Rm  �'	  � ߸ S�  �pN   � � SR�  �  Z� V� Tcff �F6  �� �� S��  �5   � �� Ss  �E,  v� p� `v B     9T�U9R	@6B     9X0  Q��  ��  @6B            �" R�  �#pN  ɺ ź bidx �#�  � � Tcff �F6  A� ?� S��  �5  f� d� Tsid ��  �� �� YV6B     ��   Q8�  Jr    B     ;       �� W
H J.�W  UW��  K.r#  TSE  M�  � � S��  Nr  }� {� 5��  S� U�  �� ��   Q�  <�  �B            �� W
H <.�W  UR��  =.r  � � SE  ?�  G� E�  V�  5�B     	       �) W
H 5(�W  U Q��  $�  �B            �� W
H $(�W  UWm  %(	  TS�  'pN  m� k� Tcff (F6  �� �� S= )�4  �� ��  Z�6  �`  � ca �`  cb �`  dret �.  dtmp �.   q��  0#B            �) 4��  � � 6��  @� <� `?#B     9U�U  q��  @5B     �       �� r��  Ur��  T6��  z� v� 6��  ľ �� 6��  �� �� _��  k5B            4��  G� E� 4��  l� j� ;k5B            s��  s��  6��  �� �� t��  B��  r5B        q��  �5B     K       �� 4��  �� �� 4��  � � A��  �  � 4��  �� �� 4��  �� �� E��  6B       @�  �4��  � �� 4��  � �� 4��  &� $�   `6B     9U�T  u��  `9B     D       � F��  6��  K� I� 6˰  p� n� 6װ  �� �� 6�  �� �� 8�9B     V 9T	`BH       qv�  �=B     Q       �� 4��  � 	� F��  F��  6��  a� [� 6��  �� �� @��  �\6��  �� �� C��  �=B     %       � 6��  &� "�  8�=B     � 9T�\  q"�  �BB     Z       �� 43�  e� ]� 4?�  �� �� 4K�  =� 1� 4W�  �� �� 1�BB            1 @h�  �P6t�  [� Y� <�BB     9T�T9Qw   _"�  �BB            4W�  �� ~� 4K�  �� �� 4?�  �� �� 43�  3� /� _��  �BB            6��  r� l� 8�BB     ��  9T�T9Qs 9Rv     q��  �BB     W       �
 4��  �� �� 4��  2� *� 4��  �� �� 1CB            0	 @�  �`<CB     9Tw   _��  (CB            4��  � �� 4��  ?� ;� 4��  |� x� _�  (CB            6�  �� �� v��  /CB      /CB            n4��  �� �� 4��  �� �� 4��  � � _��  9CB            6��  A� ?� 8ECB     . 9T�T      qo�  @PB     �       ��
 4}�  l� f� 4��  �� �� :XPB     �  a
 9Us� :gPB     " y
 9Uv  :�PB     " �
 9Uv  :�PB     " �
 9Uv  8�PB     " 9Uv   q��  pSB     �       �> 4#�  � 
� F�  F�  t0�  A9�  p�  * 6:�  �� �� 8�SB     ��  9Uu 9Tt   p�SB     t�  9R0  qI�  �TB     g       �� Fh�  F[�  o�TB     ��  � 9Uu 9Tt  8UB     t�  9Q09R0  q��   dB     Y       �� 4��  	� �� 4��  �� ~� s��  s��  6��  � � A��  �  c 4��  |� v� 4��  �� �� 5�  6��  � � 6��  ,� *� s��  :AdB     V P 9T	�1H      `YdB     9T�T   8dB     � 9U	 eH     9Tv   q��  `dB     �       �" 4�  _� O� 4�  � � 4 �  �� �� 4-�  �� z� 6:�  V� P� 6G�  �� �� 6T�  �� �� sa�  A��  0�  � 4-�  '� � 4 �  �� �� 4�  � � 4�  l� d� 50�  s:�  sG�  sT�  sa�  tn�  ww�  0�  6x�  �� �� 6��  �� �� 6��  � � :�dB     V � 9T	�1H      :�dB     ; � 9T	K.H     9Q0 `eB     9U�U9Q�Q9R�R    D�dB     ��  8�dB      9U} 9Q| ����  xF\  F\  1�y�J  �J  $�yKM  KM  Yy5<  5<  ?y)S  )S  y]  ]  )yjO  jO  y�?  �?  1^x�O  �O  22y�3  �3  1y>Q  >Q  $�x�6  �6  1�y9  9  $cy _   _  $hyF  F  $my�F  �F  $�y?U  ?U  $�y�*  �*  $�y�3  �3  $�y?  ?  $�yxL  xL  $�y�N  �N  $�x�K  �K  1vy!,  !,  Uy�R  �R  y�=  �=  �yP  P  �z�  �  3 z�D  �D  3 y\  \  Vy�-  �-  4BycL  cL  4x�,  �,  4�y�D  �D  �x�+  �+  2(xBi  Bi  2yE1  E1  $ry�*  �*  [yq]  q]  1z ��   |)  �  <�  $"  p�B     �$      �' �  B"9   ?      ��   R   ��    �� ��   �N ��   �6  ��    �  Y�   �   �   �   -   �    	X    n�   �   
�   -   �    �  ��   �   �     -   �   �   �    �  �"    �   PJ�  2�  L   �  M  pos N  �  P�  SF  Q�   �1 R�  (=9 S%  0R�  U-   8y�  V  @�� W  H �  ��  �\ ��   m  ��    o  ��  �  ��  �               	�i   	�  2  2  8  
C     ^� �  int 	�i {S @	�  g
  	�     	 	C  v  	#	C  �  	&	C  |
  	)	C   h  	,	C  (�  	-	C  0�	  	2O  8�  	5O  < �  	�  �  �
  	8"]    	K
  �  �  	L
  �  	M
  	S  	-  	�  6  >   
O  �	  
	V    :�   �  J�  x L\   y M\   )  Oh  �  B   s�  M   u\   }  u\  V  v\  /  v\   t
  x�  k	  (j  �  V   ��  V  �  	O  B� 
  L  6      s    v	  �     �  �  j  �  (N�  �  P/   Z�  Q/  �  S�  s  T�  [  U�  ?1  WO    �  /    Y|  �  =  V  �<  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "V  \  �  %  <�  x >/   len ?6  *� @   %  Ba  �    `�  �  
�  O  O  �  �    �  �  q�  �  O  	  O  O  �    �      
1  O  O  �    �  `��  �  ��   �% ��  ?1  �O  �&  ��  !  ��   I  ��  ()  �	  0R   ��   8�  ��  @ w  �  �  �1  �  �   �  �  O    �      I  �      
(  I   �  ?5  ;  
P  I       �  Y]  c  O  |  I    �    s  ��  �  O  �  I  �   �  W  0�  �  �<   e� ��  �� �(  �� �P  �� �|   �� �
  ( �'  ��  �!  l  �  �1  	�  -  �  8  D  �  ��  O  �
  �/  �  �6  �  �O  
  �V  �  ��   \#  �  �   �   �  ,O  \&  7�   �0  DC  b   �	  xx ��   xy ��  yx ��  yy ��   a  ��  	  z'  �\	  m  �I   ss  �x   �  �1	    �v	  |	  
�	  �    �  ��	  �U  ��      �i	   %  ��	  �  $�	  �	  �   
  �� "�	   �@ #�	  �U  $�    �  76
  �; 9�	   ��  :�	   L  <
  V  #��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=  ��  ?\   �  @\  ~  B\  �  C\  �  D\   5  F\  (B  G\  0�  H\  8 �	  J�  
   sg  �  u`   ��  v`  �  x\  �
  z\  (  {\   �  }  �  �#�  �  k  `�6  R�  �-    (  �x  |  �x  �  �x  �  ��  �  �
$  v  �6
  �  ��  (�%  �6  07&  �$  8G   �x  X �  �"C  I  h  �  �M �#   k  t  R�  -    �  �"�  �  %  8;�  �� =�#   �M >l    ?6
   r$  @�  0 5  �$�  �  %  �`  �� �#   �M �#  �  <   �  �  (�� 
I  h�� |  p�� �  x K  � m  s  �  �,4  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9x  8  :�  @�  <x  H�  =�  PE-  ?�	  X�!  D�  h:  Fl  �  G`  ��  H`  ��  I`  ��  K`  �  L`  �U  N`  ��  O`  �)�  Q�  ��  R4  ��� S�  �K1 W�  �R�  X-   �Jy  Y  �%  [6
  ��	  ]�	  �    ^�   ��8  `$  � L   A  G    X��  �  �`   E-  ��	  N ��  �8  ��  P �  *%�  �  �  0t�  k  vt   �  w`  �@ x�  ݖ y�  E-  z�	   N |  0�  }�  pR  ~�  x�  �  �ߣ  �<  ��I �j  ��  �x  �h  �x  ��S  ��  �4  ��  �8  ��  �  ��    �  ��   �  �\  o  �\  �L ��    �8  �  ( �
  L#�  �  W  HE  �  J`   = K
    Ll  d  Ml   �  V  �
  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  E  (0  O�  #   g)1  7  �   ���  =  �	   L  ��   $  �x  0�  �    8m  �#�!  h�  �%  pآ  �B  tG   �x  x O  g  �  �?  ds  �
  �)�  �  �   H�!  �  ��    "  ��  �!  ��   ~	  8f�  �
  hl   (  il  �� k�  �� l�    n\  �  o\   �  p\  (�  q\  0 y  s!  �a  �G    �$�  �  �  0'  �N  )x   ?1  *l  }0  +x  i/  ,x  � -	   �  �))  /     H��  ��  ��   ?1  ��  (  �  4  �	  \  ��  0  ��   @ ��  ��  +!  �  tag �   �U  �   �  �  �  `  V  
  w%   }#  �&  h  �  &     
�  E   9
w  � ;
   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  "  �  V  ��  :   �   ^$  1  �!  �!   :  ��  �  ��  �#  ��  �  �  �  6   I$  �    
  6   �&  �%  +  �  ?  6  ?   �  �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  �  @ [  R  �E  x  =v	  H  E#�  �  �  @Jn  �  L�   �  M<  �� O�  .� P�  �  Q`   �  R  (�!  S8  08'  T�  8   W!z  �  -  (l�  k  nt   �M o�  ߣ  p<  �  q�   �  k  )�  �  �  �  n  �   w   .�     
  n   �  1    
2  n  2  �   ,	  K  6D  J  
Z  n  Z   �  �  :l  r  �  �  n  n   �  >�  "  Y�  �  �  �  �  �  �  �   �  _�  �  �  �  �  �  2  �   $  f�    
  �  �  Z   �  l%  +  �  D  �  �  �   #  x��  �� � �   �  � <  H  � �  P�  � �  X9!  � �  `l� �   h  � �  p     �D  �  H2  �S  4�   �  5�  (  6�  04  7�  88  8�  @ �  :�  �  �=�  R�  ?-    �  @�  n  A�  �  B�  1$  C  2�  E  �� F  `�L H�   � �  J�    P   �  �  �  �    `  x  x  �   �  &�  �  
�  `   �%  *     �    4   �%  -!  '  
2  4   {  1>  D  �  S  �   �  4_  e  
p  �   l  8|  �  �  �  4  w   �  <�  �  �  �  4  �   �  @�  �  �  �  �  4  �  B   �  G�  �  �    `  �  �  �   �'  N(  .  �  B  `     �  SN  T  �  w  `  �  �  B  w   �  &  ��[  �� ��   i'  ��  H   ��  P  ��  X�A ��  `Y ��  h�#  ��  p�  �  x�  �2  �  �S  ���  ��  �U�  ��  ��!  �  ���  �B  ��  �p  �&  ��  �   �}  [  �&  �x  }  �   �>  ��  'O  �?   xC  ��   s/  ��  �  �  0t    �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�  �  U'9   ?   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {D   �  ��   �   �  �   -   �  �    \	  �  ��   �   
�   -   �    �'  ��   �   �  !  -   �    !   �   �!  T!  ��  )�    ��  )�   �  )�    }  !  T!  O  ;�!  _� =%�!   ݰ  >%-    a!  �  @f!  �!  cA  �,�!  �!  /  ��!  �� �   �M ��!   ?<  �,�!  �"  �5  P��"  �  ��   �� ��"  �Y ��"  �H ��"  U@ � #   �9 �#,#  (�A  �#\#  0�^  �#�#  8�^  �#�#  @N7  �#�#  H �!  ��  ��!  (Z  ��"  �"  �  �"  �!  �   17  ��"  �"  
�"  �!   �G  ��"  �"  �   #  �!  O   %G  �#  #  �  &#  �!  &#   O  �@  �8#  >#  �  \#  �!  �!  O  O   �;  �h#  n#    �#  �!  O  O   �W  ��#  �#  &#  �#  �!  -    *;  ��#  �#  &#  �#  �!  -   O   �T  ��#  �  �  I  �  -1  B�  6  $     �  *$     0$  ?  ?$  `   �  �%  �  8Y�$  ��  [�   Ǧ  \�  ��  ]�  d> ^�  ��  _�   I�  `�  (�  a  0U  b`  2�  cl  4 ��  eL$  ��  p$�$  L$  ��  ��@&  ֤  �x   Ğ  �x  ��  �8  �  �8  	��  �8  
�  �8  ��  �@&  �  �P&  (��  �@&  <�  �P&  X��  ��  p��  �x  x��  �x  |��  �`&  ��  �`&  �R�  �8  ���  �8  ���  �  �F�  �  �V�  �p&  ���  �p&  ���  ��  �"�  ��  ��  ��  �@�  ��&  � `  P&     `  `&    	 l  p&      `  �&     `  �&     ��  ��$  o�  �#�&  �$  �  ��&  ��  �&  2]   8   U�  !�&  5�  "w   �  �  $�&  ��   *�'  m�  ,�   `h  -�  �  /�'  #�  0�'  (��  1�'  ��  3w  z�  4w  ��  6(  ��  7(  ��  9�  (Ԯ  ;$(  0��  C4(  ���  D�  � �  �'     w  �'     �&  (     �$  (     �&  $(     Z  4(     �  D(     ��  FQ(  '  ��  PU)  -�  W�&   �  Y�  ��  Z�  �ܲ  [\  ���  \�  ���  ^8   �  _8  ��  `	  w�  a�  (��  c�  8�  d�  @��  ex  H T�  gW(  ��  r%0)  W(  ��  H�I*  �  ��   ��  ��  �  �x  d�  ��  |�  ��   �  �x  (�  ��$  0;�  ��  h��  ��  ���  �x  ���  �I*  ���  ��  L�  �x   ��  �x  $n�  ��  (��  �x  0��  �#)  8��  ��  @ �  Y*     M�  �6)  ��  �%s*  6)  �  V  w�+  U�   ��  ��  �  ��  ��  ޟ  $�  ��  �  	t�  
�  ܖ  �  ��  ��  d�  {�  ך  ʕ  �  ��  ��  m�  ,�  �  ^�  ׭  ~�  @�  �  ��  N�   ��  !��  "��  #ݴ  $��  %�  &�  ',�  (a�  )��  *x�  +��  ,"�  -"�  - a�  �y*  ��  )$�+  �+  H�  ��  ,�+  �+  �  �+  -   �+  �+   �&  �+  ��  1,  ,  
3,  �+  �  �  �  �   ��  8?,  E,  
P,  �+   �  ;�,  M� =�+   �� >,  Յ ?3,   ��  A�,  P,  �  h!�,  �,  ��  ��  u-�,  1-  ��  8V1-    X�,   j�  Y6-  =9 Z�-  �� [S-  Q� \z-   �� ]�-  (�� ^�-  0 �,  ��  �B-  H-  
S-  �,   ��  �_-  e-  
z-  �,  �  w   K�  �_-  å  ��-  �-  
�-  �,  �   ��  
�-  �-  �  �-  �,  �   ?�  1�-  �-  �   .  �,   .  �+  �   �  1�  �!.  .  $�  ��  �-+.  �.  .�  8��.    �.   j�  ��.  =9 �G/  �� ��.  +�  ��.   �� �/  (�� �n/  0 1.  ǡ  ��.  �.  
�.  .   ��  ��.  �.  
�.  .  �  x  w   ��  ��.  /  
/  .  �  �  I   !�  &,/  2/  
G/  .  �  I   K�  DT/  Z/  �  n/  .  �   	�  k{/  �/  �  �/  .   .  �+  �   ��  ��/  ��  ��/   X� ��/  l� �0   �,  �/  6   �/  �,  �/  6   �/  .  0  6   0  $�  ��/  �  � 10  0  �3  5]0   num 7x   str 8?   +P  :70  �J  =�0  key ?]0   �U  @C   �7  D$�0  i0  O  H�0  �0  �  �0  �0   ]0  �Z  K�0  �0    �0  �0  �0   �S  (OL1  �� Q�   �  R�  �6 S�  �B  U�0  3  V�0  >) XL1    �0  e-  \ ^1  �0  ��  #p1  v1  O  �1  ?   d�  )�1  �1  ?  �1  �   0�  /�1  K�  6�1  �> 8O   �^ 9�   �  ;�1  Ѽ  >$�1  �1  ў  (@-2  
H B�"   ��  C�  XT D-2    �1  ��  N?2  E2  ?  Y2  �  �   B�  Ve2  k2  
{2  �  ?   ��  Z�2  �2  �  �2  -   �1  �  32  Y2  �   ��  b�2  �2  �  �2  �1  O   ��  f�2  �2  O  3  �1  &#   ��  @jw3  �\ l d1   8` n {2  �\ o �2  �_ p �2  �T r �1   }�  s �1  (ʬ  t �3  0�  u �3  8 3  ��  j�3  w3  =  l  ��  W�3  ��  Yl    ��  [�3  8  �3  �  ��  ��3  ��  �x   � ��3   �  �4  �3  ��  (�\4  �9  �x   ��  ��  ɲ  ��  �  ��  �  ��    T�  �h4  4  ��  ��4  ��  ��   ��  ��  x �x  y �x   �  ��4  n4  z�  X�45  ��  �   ��  ��  �Z  ��  (%?  ��  0L�  �\4  8)�  ��  @W�  ��4  HѺ  ��  P b�  �@5  �4  ��  �!R5  X5  !(�  x��5  �� ��   s  ��   �"Q  ��    #cid �Y*  "8�  ��3  P"��  ��3  X"2�  ��   `"��  ��3  h"��  �  p �6  `S�6  �<  U�   �Q  V�  a(  X�  VA  Y�  Q) [l   nX  \l  "�D  ^�6  (�5  _�6  8M   a`  H}  b`  JV  c`  L/  d`  N7K  fl  P>D  gl  R�:  i`  T�3  j`  V=]  k`  X �  �6     �5  m�5  �Q  8��7  �  ��   �Z  �`  %?  �`  
L/  �`  �<  �l  �Y  �`  �7  �`  �)  �`  �O  �`  �H  �`  vH  �`  ^  ��7  �>  �`  $�7  �l  &0>  ��   (�+  ��   0 `  �7     �H  ��6  �?  8A�8  �  C�   �Z  D`  %?  E`  
L/  F`  S.  Hl  �W  J`  �W  K`  C  L`  �O  M`  �H  N`  vH  O`  ^  Q�7  �>  S`  $�B  Tl  &0>  Z�   (�+  [�   0 �]  ]�7  �B  �|;  ��  ~l   �)  `  �)  �l  �.  �l  U  �l  �V  �`  
�0  �`  �6  �`  �C  �`  U?  �`  6P  �`  �C  �`  &L  �`  *J  �`  �L  �`  HP  �`  N*  �;   [2  ��  0k2  ��  8.  ��  @{2  ��  HQ2  �!;  P�0  �l  Tp4  �l  VmU  �l  X�Z  �`  Z ?  �`  \:  �`  ^�I  �l  `E8  �l  b�;  ��  h�;  ��  p�O  �`  xDF  �`  zfV  �l  |�9  �l  ~[9  �l  ��G  �l  �zQ  �l  � 8  !;    	 %  1;     {D  ��8  �1  @��;  �I  ��   6Y  ��  �^  �`  S  �`  )  ��  @3  ��   �0  ��  (4C  ��  0�C  ��  8 aM  �>;  �I  @��<  �  ��   _7  ��  )  �l  �O  �l  �n �l  �T  �l  EF  �l  I  �l  �K  ��<  N:  ��<  ,L  ��<  4�E  �%  :�Z  �%  ;�Z  �8  <^  �8  = %  �<     %  �<     %  �<     eU  ��;  �9  (7�=  ��  9�   a@  :l  b<  ;l  
8  <l  .  =l  �H  >l  �Q  ?l  X  @l  �.  Al  �;  Bl  ))  Cl  eH  Dl  I_  El  �B  Fl   !3  Gl  " �)  I�<  �R   F&>  tag H�   ��  I�  .� J�  �P  K&>   �  DG  M�=  f3   �z>  Tag ��   Q  ��  .*  ��  �K  ��   gW  ��>  8>  �^   �>  k@  l   aE  l  p0  l  �>  l  H  l  �/  �  �� �3   �F  �>  �<  0C?  H  2l   �/  3�  �� 8�3   qS  :
?  A9  0U�?  ߣ  Wl   �E  X�  �^  Y�  =Y Z�?  <  [�  �=  \�?   Jy  ]  ( �>  C?  rY  _P?  �1  ~@  �.  �l   �L  �l   Z  �@  �?  �V  �Q@  ��  �l   f>  �l  Y  �@   �)  �@  �A  /A    1%   �  2%  �N  38  o=  4%  D4  5%  �^  6%  `*  7%  �0  8%  �G  9%  �D  :%  	I:  ;A  
 %  A     �@  =^@  �\  ��A  +  �A   Y�  �A  �
  �8  (  �8  �F  �8  �C  �8   <)  ��A  $A  �,  �A  �  l   AK  l  z8  �3  V �A   �A  %  �R  �A  	F  .%B  �  0l   �P  1�A   ">  3�A  $IWB  %�K K�A  %`B L%B   �[   E�B  �z  G   =Y N2B   �6  PWB  O]  a!�B  �B  �(  7N  (�
C  >) ��3   -N  ��3  V` ��3  TE  ��  �/  ��   �z  �  $ G  ��B  &8  � $C  *C  eS  po~G  �� q�   ^  s,>  ��^  u�  [>  vl   �W  wz>  (� y�6  0�=  z�7  ��,  |�=  ���  ~  ��(  �8  �AK  �l  0XL  ��?  8&os2 �1;  hp�  ��;  �T  ��3  0#9  ��  8!H �dI  @�+  ��I  H@.  ��I  P�E  ��I  X�P  ��I  `@  ��I  h$S  ��   ps  ��   x&mm ��   �&var ��   �Q  ��   �<B �Q@  �2Y ��<  �=  ��  �=  ��A  �UV  ��B  ��(  ��  =  ��3   /:  ��  (�?  ��3  0�]  ��  8&cvt �EJ  @�R  �~G  H5$  ��	  P��  �?  `HT  ��  h�*  ��  p�J  �  x�+  �  y�  ��B  ��C  �O  ��-  �?  �j7  ��  �kN  ��  ��F  ��  �#7  ��  ��(  ��3  �rE  ��3  �QZ  ��  �4  ��  ��@  ��  �:L  ��3  ��G  ��3  ��]  ��  ��W  �8J  ��/  ��  ��B   �3   �I  �3  s-  �  �*  �  ,  O  ,  O   &bdf 	
C  (�T  �  P#F  �  X�U  �  `�K  �  h �=  ��G  �G  �  �G  �    �Q  �"�G  �G  �\  xcdI  �  eC   �  fK  )�  g�  �V  h�  :1  j�   �^ k�  (Jy  m  0�  nx  8�  p`  <�!  q�  @R0  rx  `�  sx  duN tx  h6  u  lpp1 v�  ppp2 w�  �2�  z�J  �Xc  {�J  ��6  }K  )  ~�3  �8  �   �L ��   (C  �x  0��  �x  4&pp3 ��  8&pp4 ��  Hy�  ��3  X�� ��3  `U  �6
  h �I  �qI  wI  �  �I  C  �    &>    1  �I  �I  �  �I  �G  �  �  �   �M  +�I  �I  �  �I  �G   �<  :�I  �I  
J  �G   y*  V  =8J  4   �^  J  b8  �T   lK  HJ  `  |T  @?�J  R�  A-    �  Bl  n  C`  
Z�  Dl  �  E`  org G�  cur H�  ��  I�   s  K�3  ([  L�3  0c+  Nl  8 R8  PKJ  RG  T'K  K  [  O  _ &K  ,K  LL  ͳ  @@�K  Jy  B   �S C�  ܱ  D�  .� E�  ��  F8  ��  G�   
�  H�  (�P  J&>  0Ӏ K�3  8 ,�  M1K  !
�  PL  ߣ  R�   x  S�  .� U�  ē  VL  " � WL   l  !L    � ��  Y�K  ��  (\�L  ߣ  _�   x  `�  ē  b�3  ��  c�3  Ӷ  e�   �  f�  $ r�  h-L  W�  m�L  Kw  t�   7�  u�3   0�  w�L  j�  {�L  ��  }�   �  ~�  �w  �   J�  ��L  1�  �%M  �{  �%M    �L  �  �
M  �   ��M  ��  ��   k  ��M  �q  �l   q  ��  y|  ��M   �L  +M  �  �7M  %�  �!�M  �M  �  �M�O  k  Ot   Jy  P  R�  Q-   ��  R�  �   S�   �  T�  $(  V8  (|  W8  )x�  X8  *п  Z�  ,�J  \  0i�  ^�K  8�  _�K  xC�  `�K  �= b!L  ���  c�L  p�  e�K  8��  f�K  x=�  g�K  ���  h�K  ��  j�  8��  m�3  @V�  p�  HV` q�3  P��  r�3  X��  s�  `/�  u�U  h��  v�  0��  w�U  8j�  y�U  82�  |$0  Xs  |3  `��  ��  h�  �	V  pd�  ��  x|�  ��  �˽  ��	  �ʞ  ��M  �8�  �V  � ֥  0�oP  ��  �   �  �  v�  ��M  �  ��  ݺ  ��  ��  �w  c�  ��   BV �oP  ( B  �  ��O  !��  H��R  ��  ��   Ǧ  ��  @�  ��  ��  ��  d> ��  ��  ��  �  �  I�  ��   U  ��  (�  ��  0��  �x  8�& �x  <��  �	  @?�  �  `U�  ��  hw�  ��  p֤  ��  �;�  ��  �ܲ  �\  �w�  ��  ���  ��  ��  ��  ���  ��  �ٛ  ��  ��  ��  �g�  ��  �`�  ��  �x�  ��  ��  ��  �|�  ��  �"��  ��   "�  ��  "n�  ��  "��  ��  "��  ��   "`�  ��  ("�  ��  0"m�  �l  4"�m  �l  6"A�  ��  8"��  ��  @ ��  ��P  S�  �$�R  �R  ��  �*�S  Ҳ  ,�R   -�  -aU  H�  0uP   ݺ  1�  P&NDV 2w  X�  <�3  `K�  =�3  h�  >�  p��  ?�  t��  A�K  xZ�  B�3  �l�  EO  � !E�  ��1U  ��  �8   �  �8  ��  �8  �  �8  ��  �1U  �  �AU  x��  �1U  �"�  �AU  8"��  ��  �"��  �\  �"��  �\  �"��  �\  ��   \  �R�  8  ���  8  �V�  QU  ���  QU   ��    �6�  �  �Ğ  x  �"�  	x  ���  
�  �Т  �  �P�  �  �W�  \  ���  \  ���  �  ���  �R  � \  AU     \  QU    	 \  aU     ��  �S  a�   �U  ߣ  8   �  �  �U  �3  
�  �  w�  !�  .�  "�  �  #8   �  %nU  9�  G�R  �R  	V    � �$  �3  8�  `,=V  �� .�   -U /�  X `�  1IV  V  !~�  H<�V  �� >�   "�� @  0"��  A  1"�� C�  8"�� D�  @ Z�  F�V  OV  �C  h*W  �� ,�#   �Z  .�  8�  /  <X;  0W  @آ  1B  ` x  W     �D  3 W  �V  ��  ?-2W  8W  ۳  `��W  ��  ��3   y�  ��  �� ��  �� ��  ��  �x   Ǩ  �x  $(2 ��3  (Ϛ  ��3  0R�  �-   8_� �^X  @ ��   T
X  �� W#X   �Y \4X  add _XX  �x e4X   �  #X  &W  x  -    
X  
4X  &W   )X  �  XX  &W  x  �   �   :X  r�  g�W  ^X  �  �"{X  �X  ��  ���X  y�  ��3   2�  ��3  �� ��3  � ��  R�  �-    _� ��\  ( ��  �"�X  �X  ��  �+Y  �S ��3   �� ��3  � ��Y   ��  �"<Y  +Y  BY  ��  0��Y  9�  �?   �{  ��Z  � �jZ  ��  ��Z  x  ��  �  �8  m�  ��   �  ��  $��  �  ( '��  V  ��Y  ˟   .�  ��  ��  ��  ��   ��  ��Y  'L�  V  �jZ  ��   ��  Ʊ  ��  ��  g�  �  ��  W�  �  	|�  
K�  ��   8�  �	Z  '��  V  ��Z  c�   ��  p�  �  �  ��  �  ��  ��  }�  	 ��  �vZ  ��  ��Z  �Z  
�Z  `  �   [�  BY  �Z  �  hk�[  �� n�[   �Y t�[  �? w�[  �2 y�[  �! |
\   �$ ~$\  (�* �M\  0�3 �l\  8k! ��\  @�A ��\  HV- ��\  P�F ��\  X  ��\  ` 
�[  oX  �3  �3  -    �[  
�[  oX   �[  �  
\  oX   �[  �  $\  oX  x   \  �  M\  oX  �3  �  &>     *\  x  l\  oX  x  EJ   S\  x  �\  oX  x  w  x   r\  
�\  oX  �X   �\  
�\  oX  �X  �  �\   x  �\  �  �\  oX  7Y  ~  �  &>   �\  �  �[  �\  �  ��X  ~�  �']  l�  p$^  R�  -    �  `  )�  �V  ��  �  2�   .   ��  .  (��  �^  0��  �^  8R0   �  @�  !�  H�!  #Z  P��  $  X�� %  Yb�  &  Z��  (  [�  )  \_� +�^  ` ګ  �O^  �� �j^   �Y �{^   
d^  d^  �      ]  O^  
{^  d^   p^  �  �$^  \  î  B�^  2�  D�3   �� E�3  y�  F�3   {�  H�^  ��  L�^  �^  �  _  C  �  �3  &>   l�  R_  _  
3_  C  �3  �   ��  �WNa  <0 Y]   4� [Na  p&top \w  �O� ^^a   Xc  _na  ���  ax  ��  bx  ��  cta  �&cff e�M  �  f�R   ˽  g�a  (
�  i�^  0�  j  8��  kx  <z�  m�  @�  n�  D��  px  H�  qx  L~�  s�3  P9� t�3  XV v�3  `�  w�  h&  y�  l�J {  p�  }&�^  x��  ~&_  �s  �|3  �Ğ  �x  ���  ��3  �q�  �R1  ���  �	  �w�  ��  ��  �D(  ��  ��&  ��  ��  � �  ^a    0 �^  na     �^  �  �a     �	  x�  �3_  ջ  �#�a  �a  �  ��b  R�  -    �  `  )�  �  ��  �  2�   .   ��  .  (��  \  0��  \  8R0  �  @�  �  P�!  �  `��  dd  ���   �b�    ���     ��  "�   �L�  #�   �_� %&d  � ��  ��b  �b  �  �b  �a  x   q�  ��b  �b  
	c  �a  \  \  8   j�  �c  c  �  5c  �a  \  \   ��  �Bc  Hc  �  Wc  �a   *�  �c  �  �qc  wc  
�c  �a   �  @�d  �� � d   �Y �qc  �? �$�b  kI �$�b  rL �$	c   � �$5c  (-1 �$Wc  0��  �$dc  8 
 d  �a  `  4  �     d  T�  ��c  &d  a�  V  �dd  ��   J�  �  ,�   ה  �8d  ��  '�a   �  F�d  y�  H�3   2�  I�3  �� J�3   ɠ  L~d  ݬ  L�d  ~d  �  O/�d  �d  ��  �}~f  <0 qd   4� ��g  �&top ��&  �O� ��g  �Xc  ��d  x
s  �|3  �
�  ��  �
V ��3  �
Ğ  �x  �
��  �x  �
��  ��3  �
h�  ��3  �
��  �R1  �
��  �	  �
w�  ��  �
��  �x  �
�  �x  �
�  �ta  �
�  �D(  `&  ��  h�  ��f  p_� �~g  x�  ��&  ��  ��  ��J �  �˽  ��	  � �   X�f  �� [#g   �Y f4g  �; oSg  � uxg   �  T�f  �f  �  �f  �d  �   �  #g  �d  `  4  �  �3  D(    �  �f   �f  
4g  �d   )g  �  Sg  �d  �3  �   :g  �  rg  rg  �3  �   �a  Yg  X�  z~f  ~g  �  �g    � �d  �g     �  ��d  <�  � �g  ��  ��h  R�  -    �  C  )�  �V  ��  �  2�   .   ��  .  (��  \  0��  \  8R0  �  @�   �  P�!  "�  `��  $  ��� %  �b�  &  ���  (  ��  *�   �L�  +�   �_� -Lj  � c�  ��h  �h  �  �h  �h  x   �g  ˯  �i  i  
/i  �h  \  \  8   N�  �<i  Bi  �  [i  �h  \  \   Ԝ  �<i  h�  �ui  {i  
�i  �h   8�  ��i  �i  �  �i  �h   p�  @�'j  �� �Fj   �Y �ui  �? �%�h  kI �%i  rL �%/i   � �%�i  (-1 �%[i  0��  �%hi  8 
Fj  �h  C  =V  �V     'j  +�  ��i  !�  E�j  2�  G�3   �� H�3  y�  I�3   ��  KYj  j�  �NPl  <0 P�g   cff Q�M  �4� SNa  �&top Tw  hO� VPl  pXc  W`l  ��  Yx  �  Zx  �  [ta  
�  ]\  ���  ^\  ���  `  ��  a  ���  bx  ��  cfl  �z�  e�  ��  f�  ���  hx  ��  ix  �~�  k�3  �9� l�3  �V n�3  ��  o�  �&  q�  ��J s  ��  u�R  ��  w&�^  ���  x&_  � �j  `l     �j  �  vl     1�  z�j  l�  �l  �� ��l   >'  �m  � �xg   
�l  �l  C  =V  �V    �  �^  _   vl  �l  �  m  �l  =V  �   �l  U�  ��l  m  :�  �#4m  :m  ,�  (��m  R�  �-    Jy  �$n  � �45  p�  �Un  o�  ��     4�  ��m  �� ��m   �Y ��m  gP �n   �  �m  'm  -   �3  �3   �m  
�m  'm   �m  �  n  'm   �m  \�  ��m  n  ١  �#1n  7n  ��  x  Un  ?  �  �    <n  �  �.hn  �n  0�   ��n  ��  ��!   �0 ��!  ک  ��!  �> ��!   nn  �  X�co  b�  !co   �  !io  E�  !oo  b�  !uo  ,�  �o   h�  �o  (�  �o  0��  �o  8c�  [n  @:�  !�o  Hs�  "�o  P jX  ]  3d  �g  
�o  �3  �  l   {o  O  �o  O   �o  
�o  rg  �      �o  
�o  `  �&  �R   �o  n  "m  ��  �o  �n  -�  � =vp  ��  ?]   Jy   @  �p�   B�3  ���   C�  ���   E�  �'�   G�  �cid  If*  �l�   Jx  � ��   L p  ]�  �!�p  �  !!vp   ~�  !"x  � I�  !$�p  ;�  "8!�p  �p  �  `"]�p  �� "_�   pw  "`  X ��  "C&�p  q  !��  H"eVq  �� "g�   "�� "i  0"��  "j  1"�� "l�  8"�� "m�  @ V  #��s  p�   �  ��  (�  �  
�  ��  @�  ��  M�  	��  
F�  u�  �  ��  �  ;�  ��  ��  ��  �  G�   {�  !��  "��  #�  $�  %��  &t�  '��  (��  0��  1�  @��  Av�  Qd�  RF�  S��  T��  U��  VD�  Wn�  X��  `��  a��  bn�  c5�  p�  ���  �6�  ���  ���  ���  ���  ���  �o�  �o�  ��  �b�  ���  �]�  �^�  ��  ���  ���  ���  �5�  �%�  �t�  ���  �Y�  �W�  ���  �}�  �g�  ���  ���  ���  ���  �D�  ���  ��  ���  ��  ���  ���  �P�  �5�  ���  �"�  �2�  ���  �(�  �d�  �  [  �s    2 �s  (8�  2�s  	�jH     V'  $#g  FO  %)*$  ��  %,�s  �s  Y  %,	t  6 %.�s    =�  &!t  t  �  /t  `  	V   T�  &%;t  At  �  Ut  `  V   ��  &)at  gt  x  vt  `   �  &,�t  �t  �  �t  `  �t   �&  ��  &0�t  �t  �  �t  `  �+  �  �   �   �  &7�t  �t  ,�  (&77u  ۽  &9	t   1�  &:/t  G�  &;Ut  #�  &<vt  )�  &=�t    ��  'Cu  Iu  �  gu  `  gu  gu  �\   ?  ��  '$yu  u  �  �u  `  �u     �  ''�u  �u  �  �u  `  �  �3   d�  '+�u  �u  ��  '+
v  �  '-/7u   N�  './mu  ��  '//�u   n)  (v  v  �  :v  6  ?  �     �)  ($Fv  Lv  �  ev  6  ?  �    nk  ()vv  ev  �;  ()�v  �=  (+
v   z+ (,:v   )S�  A*�s  	�jH     )��  ^&�t  	�jH     )��  �#�u  	PjH     )_�  �qv  	@jH     �  w     �v  ).�  �#w  	�iH     *�s  �	 iH     +��  ��  �B     
       ��w  ,~ �#6  X� T� ,�  �#?  �� �� -�B     Z�  .U	�iH     .T�T  +��  ��  �B     
       ��w  /�  �+F5  U/�^ �+�  T0cid �+�3  Q1� ��    +J�  ��   �B            �Ex  /�  �F5  U/R�  ��u  T1� ��    +�  p�  АB     .       ��x  /�  pF5  U/d�  qgu  T/|�  rgu  Q/�  s�\  R2cid uf*  �� ��  +i�  V�  ��B            ��x  /�  V+`  U/��  W+V  T +��  M�  ��B     1       �2y  /�  M*`  U/ù  N*	V  T +��  5?  `�B            �wy  /�  5&F5  U3E  7?  �� ��  4��  �y  5�  !�y  67Jy      vp  8�  9�  �z  9�  9"�y  9Jy  :"  9R�  ;"-   9Q  <"�o  :� >�  :��  ?�  :x  ?�  :�  ?$�  ;cur @�3  :�� @�3  :}0  A�3  :i/  A�3  <�u  �<��  Z<�Y �=�z  :B� o�z  :2�  r�  :��  s�  ;p t�3  6:��  y�    6;tmp ��    8  �z  >  	 ?(�  P�B            ��z  @K1 6  U A^�  ��  ЏB     x       �J{  @~ �6  UBK1 �W  4� 2� (ߢ  �O  �t C��  �  |  5Jy  !  58�  !`  5�  !x  5G  !x  5G  !�  7�  F5  7� �  7Q  �o  72�   $0  D�u  ���B     6Ecid _f*  7��  `�$  67s�  x�  7r? y�     F�  ���B     �      �4~  ,8�  �`  _� W� 3�  �F5  �� �� 3R�  �-   '� %� 2cid �f*  P� J� 3��  ��$  �� �� G�B     w       /}  2n �x  �  � G �B     D       }  3�8 ��3  T� R� H�B     g�  }  .U}  I1�B     g�  .U}   IU�B     g�  .U}   Ho�B     g�  G}  .U}  H��B     g�  _}  .U}  H��B     g�  w}  .U}  H��B     g�  �}  .U}  HלB     g�  �}  .U}  H�B     g�  �}  .U}  H�B     g�  �}  .U}  H/�B     g�  �}  .U}  HI�B     g�  ~  .U}  Hs�B     g�  ~  .U}  I��B     g�  .U}   +��  ��  `�B     4       ��~  ,�  �&4  }� w� Jreq �&w  �� �� 3_� ��,  � � Hl�B     s�  �~  .T�T Ht�B     ��  �~  K�  s  L��B     .R0.X0  +��  ��  ��B     Y       ��  ,g�  �4  1� +� 3�  ��p  �� }� 3� ��  �� �� 3_� ��,  � 
� G��B     9       �  )9� ��+  �h3�  �F5  H� D� 3��  �#)  �� � 3��  ��&  �� �� L�B     .Q�h  I��B     ��  K�  s   M��  p�  9g�  p4  :�  r�p  6:_� w�,    8��  `�,  J�  9�  `)�p  :�  bF5  :2�  c$0  :~ d6   N��  :�   �B     M       ��  , : �  -� '� 3�  <F5  � y� 32�  =$0  �� �� O6�B     .       3~ E6  �� �� GS�B            ��  3_� L�,  � �  IN�B     ��  .T	`BH        F��  3��B            �A�  / 3 �  U Ca�  ��  �  5�  �F5  5�  �x  7��  ��p  7�  ��y  7R�  �-   7� ��  En �x  Ecid �f*  7'�  ��  7U�  ��  P�u  H67��  #)    C��  P�  ւ  5�U  P �3  5)  Q �  5x  R �  5�  S F5  7Jy  U  7� V�  7B� Xւ  Ep Y�3  7`�  Y�3  Ed Z�3  7@�  Z�3  Eval [8  7��  ]  7�Y ]  P�u  �67�  o�  7�  p�    8  �    � 49�  E�  5��  E!�  7�  G�y   �p  4��  ;>�  5��  ;!�  5�  <!F5   C��  ��  f�  5�  �F5  Ecid �f*  7R�  �-   7Jy  �  7� ��  En �x  7�8 ��3  7U�  ��  7�P  �&>  7Q  ��o  P�u  &P�0  *67��  �#)  7Ğ  �x  7.� ��  7��  ��  7)  ��  Ep ��3  =B�  7�:  ��   =U�  Elen �   6Elen �     C��  @�  �  5�  @ F5  5��  A �  52�  B �3  5�  C �  7�  E�y  6Ecur M�3  7�� N�3  67�  S�3  6Elen w�  67��  �+Y  67F@ ��3  6En ��         A��  �  p�B     K       ���  Q�  (F5  ?� 9� Q�   (�y  �� �� B��  "#)  �� �� L��B     .U�T.T0  +)�  ��   �B     �       ��  ,�  � F5  � � ,�  � �y  �� ~� 2cid �f*  �� �� 3R�  �-   2� .� 3Jy  �  l� h� )� ��  �L3��  ��  �� �� D�u   �B     G��B     j       ׆  Rn x  �� �� G�B            ��  B��  #)  � �  I��B     ��  .Uv .T
P.Q0.Rs .X0.Y�L  LI�B     .U�T  +��  ��  ��B     c      �z�  ,�  �'F5  ^� V� ,�  �'�y  �� �� 3��  �#)  � � 3�� �`  o� g� )/� �z�  ��3��  ��  �� �� S�  3:  ���  � � 3x  ��  j� f� 3E  �x  �� �� T��B     �  .U�T.T6.Qw .R3 H��B     ��  �  .U
�.T}  H��B     ��  �  .T}  H��B     ��  4�  .T}  HӞB     ��  L�  .T}  H�B     ��  d�  .T}  I��B     ��  .T}    �  ��     	  8�  F�  �  9�  F%F5  9��  G%�  9��  H%7Y  :� J�  :�  K�y  :ݰ  L�3  :װ  M�   ;cid Nf*  <�u  �6:��  n#)    8��  *�  X�  9�S *�3  9��  +8  :E  -�  ;p .�3   A��  Q�  @�B     u      ���  Q��  Q&�  � �� Qg�  R&4  s� e� Q�^ S&�  � � Q:1  T&B  �� �� B)�  V�p  �� �� B� W�  )� � (�3 X�g  ��hB�  YF5  �� �� BZy  Z  A� 3� B��  [  �� �� BQ  ]�o  �� �� (��  ^	  ��gBw�  _�  �� �� B<�  `  f� Z� P�u  
G��B     V       �  B�8  �  �� �� U�B     ��  U!�B     ��   V�  8�  (C!  ��  ��gBN ���  � � V��  ��  Rn �x  S� Q� Rcur � .  �� ~� Rvec ��  �� �� B�� ��  E� A� B�� ��  �� � W��   �B      ��  �ԋ  XՔ  Y˔  �� �� S��  Zߔ  �� �� Z�  @� <�   [��  %�B      %�B            �2�  XՔ  X˔  O%�B            Zߔ  � {� Z�  �� ��   [��  L�B      L�B            � ��  XՔ  Y˔  �� �� OL�B            Zߔ  (� $� Z�  k� g�   \��  m�B      m�B            � XՔ  Y˔  �� �� Om�B            Zߔ  �� �� Z�  � �    W��  L�B      0�  � Q�  YՔ  Q� O� Y˔  x� v� S0�  Zߔ  �� �� Z�  �� ��   W��  q�B      `�  � ��  YՔ  !� � Y˔  H� F� S`�  Zߔ  q� m� Z�  �� ��   U��B     ��  UӘB     ��  HL�B     ��  ��  .U| .T��g H��B     ��  �  .U| .T} .Q~  H��B     ͤ  #�  .U| .T��g I��B     ٤  .Us0  T�B     i�  .U��h.T| .Q} .Rs .X0.Y0 H1�B     ��  ��  .U��h.T~  T��B     ��  .U��h Lh�B     .U��h    +��  -�  p�B     �      ���  ,�3 -�d  �� �� ,�^ .�  �� �� 3�  0F5  �� �� 2cid 1f*  k� a� 2p 2�3  �� �� 3j�  3�  �� �� 3Jy  4  �� �� )� 5�  ��k3ٶ 6�3  Y� C� 3R�  7-   G� ?� 3��  8�  �� �� 3Q  9�o  �� �� 3=�  ;  $� � 2inc >#�!  �� �� ]�u  ��B     V��  ߐ  )��  K\	  ��u^�  �B      ��  Tg�  Y5�  �� �� Y)�  6� 2� S��  ZA�  |� v� ZM�  �� ��   TבB     ��  .T��k�.Q��u TQ�B     ��  .T��u H+�B     �    .Uw .T��k.Q��k IV�B     �  .U} .Q��k  V@�  ��  3U�  l�  � � 3ti m�  ?� ;� 3Ϭ m�  {� w� ^�  ЕB      ��  vy�  Y5�  �� �� Y)�  �� �� S��  ZA�  6� 0� ZM�  �� ��   _�  �B       �B     1       w�  Y5�  �� �� Y)�  <� 8� O�B     1       ZA�  �� |� ZM�  �� ��   ^�  ?�B      ��  y;�  Y5�  5� 3� Y)�  \� Z� S��  ZA�  �� �� ZM�  �� ��   H��B     ��  U�  .U��k H��B     
�  }�  .U��k.T
s 1$���� Hv�B     �  ��  .U��k H˖B     �  ��  .Uw .T��k.Q��k H��B     $�  �  .U��k.Q} .R��k I�B     �  .U��k  V�  2�  3��  �#)  � � 3��  ��3  c� _� 3-F  ��  �� �� GX�B     �       ��  )A�  ��a  ��u)��  ��U  ��lTu�B     ��  .U��u.Tv .Q1 T��B     ��  .Ts .Q��l T��B     ֓  .U��u.T��k.Qs  L��B     .U��u.T��k.Qs   T�B     �  .U} .T��k.Q
� LS�B     .Uv .T��k  Gv�B     �       ��  )N �"�   ��uU�B     ��  U��B     ��  U��B     ��  LٓB     .T��k�.Q0.R��u  I'�B     g�  .Uw .T}   8�6  �B  ��  `a �B  `b �B  ;ret �(  ;tmp �(   a�   �B     <       �[�  X�  Z%�  �� �� Z1�  � � Z=�  V� R� I=�B     ��  .T	`BH       b�   �B     9       ��  Y�  �� �� Z�  �� �� c�  �B     "       Y�  `� Z� O�B     "       d�  c�  �B     "       Z�  �� �� I�B     ��  K�  s      bJ{  @�B     �      �Z�  Y\{  �� �� Yi{  � �� Yv{  �� �� Y�{  L  D  Y�{  �  �  Z�{  D  Z�{  %  Z�{  � � Z�{    eJ{  0�  �  Y\{  ` T Y�{  � � Y�{  L F Yv{  � � Yi{   � S0�  d�{  Z�{  � w d�{  d�{  f�{  WA�  ��B      ��  H��  Y`�    YS�  � � S��  gm�  ��{Zz�  
 
 Z��  �
 �
 g��  ��{Z��  � � Z��  � � Z��  � � ZƁ  � � hӁ  G�B     W�  �B       �  ��  Y0�  f F Y#�  � �  W�y  �B      @�  �N�  Y�y  � � Y�y  ; + Y�y   � Y�y  � � S@�  Z�y  y a Z�y  � s Zz  Q 9 Zz  X L Zz   � Z%z  s a Z1z  D 8 Z=z  � � fIz  hQz  e�B     hYz  /�B     eaz   �  ��  gfz  ��}Zrz  K A Z~z  � � Z�z  d T e�z  @�  {�  Z�z    H��B     1�  /�  .Uv  H��B     >�  S�  .Uv .T| .Q  I?�B     K�  .U��}.T	�  "
Y.Q9  I��B     1�  .Uv   i�z  �B             ՙ  Z�z  S Q I�B     W�  .Us .T0.Q:  T�B     ��  .U~ .T0.Q0.R��{ H �B     1�  �  .Uv  H�B     
�  0�  .Uv .TO H?�B     �  H�  .Uv  Ue�B     �  HF�B     ��  u�  .Uv .T��{ H`�B     c�  ��  .Uv .Ts .Q~� T��B     ��  .U~  T��B       .U~  TťB     ֚  .U~  TϥB     �  .U~  T�B     ��  .U~  T�B     �  .U~  HG�B     p�  1�  .Uv .T~� IS�B     ��  .Uv .Tw    [�  G�B      G�B     )       I�  Y�  x v OG�B     )       Z�  � � \wy  G�B      G�B     )       KY�y  � � i�y  R�B            �  Z�y  � � If�B     p�  .T~�  Lp�B     .U~     Wf�  ��B       ��  �D�  Y��    Y��  5 3 Y��  j X Yx�  ' % S��  Z��  ^ J j��   �  Z��  H , ZǄ  ~ n jԄ  ��  ZՄ  M I e�  0�  �  Z�  � � j��  ��  Z�  /    j��  �  Z��  ! �  e�  p�  �  Z�  =! 7! k��  ͫB      е  �(Y��  �! �! Y��  O" ?" Y��  # �" Sе  Zň  x# p# Zш  �# �# Z݈  �$ �$ g�  ��}Z��  �$ �$ h�  9�B     e	�  @�  ��  Z
�  |% z%  T9�B     �  .U~ .T .Q��}.R0.X0 L��B     .U} .T~     I��B     }�  .U}     TϦB     0�  .U~  LڪB     .U~      W�  �B       p�  ���  Y%�  �% �% Y�  J& H& Y�  o& m& Y��  �& �& Sp�  Z2�  �& �& Z?�  b' Z' gL�  ��}ZY�  �' �' Zd�  ) �( Zq�  n) Z) Z|�  H* <* Z��  �* �* Z��  ++ + Z��  �+ �+ f��  e��  �  ��  Z��  �, �, Zǂ  - 
- H��B     1�  Z�  .Us  HجB     >�  y�  .Us .T��} I�B     1�  .Us   I$�B     ��  .Us    e܁   �  ��  Z݁  n- d-  W>�  ��B      P�  Fa�  YP�  �- �- SP�  Z]�  Q. K. Zj�  �. �. Zw�  (/  / g��  ��}Z��  �/ �/ Z��  �0 y0 Z��  �0 �0 Z��  �1 �1 ZÃ  �2 �2 hЃ  ��B     hك  ��B     e�  ��  ʢ  Z�  A3 73 Z��  �3 �3 Z��  �4 �4 Z
�  O5 C5 Z�  �5 �5 Z$�  6 �5 e/�   �  2�  Z4�  T6 N6 I��B     ��  .Uw .T8.Q��{�����.R��{�����.X| .Y��}  W�  �B       0�  ���  Y5�  �6 �6 Y)�  �6 �6 S0�  ZA�  '7 !7 ZM�  z7 r7   iB�  S�B            ��  ZG�  �7 �7  iU�  ��B            �  ZV�  8 8 L׳B     .Q
�  HðB     ��  ��  .U  H�B     
�  �  .U  HQ�B     �  /�  .U  HűB     ��  m�  .Uw .T8.Q0.R��{�����.X0.Y��} H��B     �  ��  .Uw .T��{.Q��} H�B     ��  ��  .U  ID�B     >�  .U .Q��{  H�B     ��  ��  .Uw .T@.Q0.X0.Y��} H:�B     g�  �  .Uw  H_�B     g�  +�  .Uw  H��B     g�  D�  .Uw  I��B     g�  .Uw .Ts    H��B     �  ��  .U��{.TP.Q��{ H�B     �  ��  .U��{.Q��{ U��B     ��    j�{  `�  Z�{  t8 j8 Z�{  �8 �8 j�{  ��  Z�{  �9 z9 Z|  ': !:     H��B     ��  �  .Us .T0 H�B     ��  >�  .T	�BH      I%�B     ��  .T	`BH       l�*  �*  [mF\  F\  )�l�=  �=  �l�R  �R  m�6  �6  )�l5<  5<  ?l\  \  Vl�-  �-  *BlcL  cL  *m�,  �,  *�l�D  �D  �m�K  �K  )vn�D  �D  . l9  9  +cl�3  �3  +�lxL  xL  +�l`I  `I  +xlF  F  +mlE1  E1  +rm�Z �Z ,m�\  �\  -.l�*  �*  +�l�J  �J  +�m�O  �O  ,2l�X  �X  +Xl!,  !,  U �t   �/  �  �  $"   �B     R5      �G X  ^� 	�@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  .�  
�5  -  �[  
�H  �  >   
G   �	  
	N   �  B"u  {     ��  R   �U    �� ��  �N ��  �6  �   �  Y�  �  U   �  i  -      n�  �    i  U    �  �    U   5  i  -   -   U    �  �"A  G  �   PJ�  2�  LD   �  M@   pos N@   �  P  SF  Q   �1 R  (=9 SQ  0R�  Ui  8y�  VD  @�� WD  H �  �  �\ �-   m  �U    o  ��  �  �   &  @   D  5  @   D  @    J  �  2  ^  d  o  5     :-   �  J�  x Lo   y Mo   )  O{  	�  B   s�  M   uo   }  uo  V  vo  /  vo   t
  x�  �J  N   �G  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  N    ��  N   �  	G   B� 
D  L  H    J  s  J  v	  U     �  G  	�  �  (N;  �  P5   Z�  Q5  �  S;  s  T�   [  UA  ?1  WG     �  5    Y�  �  =  N   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  �Z  b   "�  �  �  %  <�  x >5   len ?H  *� @J   %  B�  	�    `    3  G   G   3  U      �  qF  L  G   e  G   G   U    �  r  x  �  G   G   U    �  `�  �  �   �% �   ?1  �G   �&  �  !  �   I  �9  ()  �e  0R   �U   8�  ��  @ �  &  �  ��  	'  �   F  L  G   `  U   `   �  �  s  y  �  �   �  ?�  �  �  �  D  @    �  Y�  �  G   �  �  @   U    s  ��  �  G   �  �  �   4  W  0�h  �  ��   e� �9  �� ��  �� ��  �� ��   �� �f  ( �'  �  �!  lJ  �  ��  �  -  �J  	�  �  �  ��   	�  �
  �5  �  �H  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   �0  D4   b   �{	  xx �	   xy �	  yx �	  yy �	   a  �8	  	{	  z'  ��	  m  ��   ss  ��   �  ��	    ��	  �	  �	  U    �  �
  �U  �U      ��	   %  ��	  �  $(
  .
  �   g
  �� "
   �@ #
  �U  $U    �  7�
  �; 9
   ��  :
   L  <g
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=a  ��  ?o   �  @o  ~  Bo  �  Co  �  Do   5  Fo  (B  Go  0�  Ho  8 �	  J�  
   s�  �  u�   ��  v�  �  xo  �
  zo  (  {o   �  }n  �  �#�  �  k  `��  R�  �i   (  ��  |  ��  �  ��  �  ��  �  �d$  v  ��
  �  �8  (�%  ��  07&  �t$  8G   ��  X �  �"�  �  h  �  �M K$   k  �  R�  i   �  �"�  �  %  8;8  �� =Q$   �M >�    ?�
   r$  @�  0 5  �$E  K  %  ��  �� Q$   �M ^$  �  �   �  C  (�� 
�  h�� �  p�� �  x K  � �  �  �  �,�  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6  (A  7  0T  9�  8  :  @�  <�  H�  =  PE-  ?
  X�!  D�  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R�  ��� SG  �K1 W�  �R�  Xi  �Jy  Y5  �%  [�
  ��	  ]
  �    ^U   ��8  `�  � L   �  �    X��  �  ��   E-  �
  N ��  �8  �1  P �  *%�  �  �  0tG  k  v�   �  w�  �@ x�  ݖ y�  E-  z
   N |a  0�  }	  pR  ~	  x�  �  �ߣ  ��  ��I ��  ��  ��  �h  ��  ��S  �G  �4  ��  �8  �  �  �U    �  �-   �  �o  o  �o  �L �U    �8  �x  ( �
  L#T  Z  W  H�  �  J�   = Kf    L�  d  M�   �  N   �f  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  (0  OZ  #   g)�  �  �   ��  =  �{	   L  ��   $  ��  0�  �v   8m  �#�!  h�  ��  pآ  �O  tG   ��  x �  �  G  �?  d�  �
  �)>  D  �   H�}  �  �U    "  �  �!  ��   ~	  8f�  �
  h�   (  i�  �� k	  �� l	    no  �  oo   �  po  (�  qo  0 y  s}  �a  ��    �$#  )  �  0'x  �N  )�   ?1  *�  }0  +�  i/  ,�  � -{	   �  �)�  �     H��  ��  ��   ?1  ��  (  �u  4  �{	  \  ��  0  �U   @ ��  ��  +!  &  tag �   �U  	   �  �  &  `  N   
q  w%   }#  �&  h  �  &     
9  E   9
�  � ;
q   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  ~  �  N   �  :   �   ^$  1  �!  �!   :  ��  �  �	  �#  �C  I  	  X  �   I$  �d  j  u  �   �&  ��  �  +  �  �  �   �   �!  H�$  �  ��   S"  ��     �$  �"  �	  �  �	   ;  �   (%  �7  0�   �X  8��  �u  @ �  R  ��  x  =�	  H  E#T  	C  �  @J�  �  L�   �  M�  �� O$  .� PJ  �  Q�   �  Rg  (�!  S�  08'  T�  8   W!�  �  -  (l  k  n�   �M o  ߣ  p�  �  q�   O  k  )0  6  	  J  �  �   w   .V  \  g  �   �  1s  y  �  �  �  T   �	  K  6�  �  �  �  �   �  �  :�  �  	  �  �  �   �  >0  "  Y�     	    8  �    T   �  _*  0  	  N  8  �  �  T   $  fZ  `  u  8  �  �   �  l�  �  	  �  8  �  	   #  x�	  �� � *   �  � �  H  � �  P�  �   X9!  � N  `l� � u  h  � 	  p h    ��  �  H2j  �S  4G   �  5;  (  6;  04  7�  88  8  @ �  :  �  �=�  R�  ?i   �  @�  n  A�  �  B�  1$  Cu  2�  Ej  �� Fj  `�L HU   � �  J�  v  P   
    	  3  5  �  �  �  3   �  &?  E  P  �   �%  *\  b  	  q  �   �%  -}  �  �  �   {  1�  �  	  �  �   �  4�  �  �  �   l  8�  �  	  �  �  �   �  <�    	    �  �   �  @$  *  	  H  �  �  �  O   �  GT  Z  	  x  �  �  �  ;   �'  N�  �  	  �  �  5   �  S�  �  	  �  �  �  �  O  �   	  &  ���  �� �*   i'  ��  H   ��  P  ��  X�A ��  `Y �3  h�#  �P  p�  �q  x�  ��  �  ��  ���  �  �U�  �H  ��!  �x  ���  ��  ��  ��  �&  ��  �   ��  	�  �&  ��  �  �>  �   'O  ��   xC  �    s/  ��  	   �  0tv   �  v	   a   w	  �'  x	  !  y	  �#  z	   �  {	  ( �  }   �  U'�   �   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {�   �  ��   �   	  !  �   �  !   �	  �  �%!  +!  ;!  �   !   �'  �G!  M!  	  k!  �   �  u  k!   �   �!  �!  ��  )�    ��  )!  �  );!   }  q!  	�!  O  ;�!  _� =%�!   ݰ  >%�    �!  �  @�!  �!  cA  �,"  "  /  �:"  �� �s   �M �:"   ?<  �,F"  �"  �5  P��"  �  ��   �� ��"  �Y �#  �H �0#  U@ �V#   �9 �#�#  (�A  �#�#  0�^  �#�#  8�^  �#$  @N7  �#.$  H 	L"  ��  �"  (Z  ��"  �"  	  #   "  	   17  �#  %#  0#   "   �G  �<#  B#  �  V#   "  \   %G  �b#  h#  �  |#   "  |#   \  �@  ��#  �#  �  �#   "   "  \  \   �;  ��#  �#  u  �#   "  \  \   �W  ��#  �#  |#  $   "  i   *;  �$  $  |#  .$   "  i  \   �T  �$  g�  �L"  	:$  *  �  �    �  t$  @    6  �$  @     �  �%h  M�  l�%  ��   \   ��  !�  D�  "�  x�  #�  �  %�  �  &�  /�  (�  &�  )\  ��  *\   �  ,\  $h�  -\  (�  .\  ,Y�  0�  0=�  1\  4��  2\  8��  4�  <��  5�  @o�  6�  Da�  8�  H-�  9�  L��  ;\  PI�  <\  TE�  =\  X�  ?�  \v�  @�  `��  A�  d�  B�  h ��  D�$  ��  D&  �$  U�  0N�&  �  P\   x  Q\  :  S�&  ��  T�  ;�  U�  y  V�   ��  WO  $$�  Y\  (5�  Z\  , O  �&  @    F�  \&  '�  \�&  &  ��  v'  ��  x�   p  y�  ��  z\   t�  |'  �&  �  (��'  ��  ��   ��  ��  ?1  ��  p  �\  ��  �\  ��  �\  #�  �\  q�  ��  u�  �'    ��  �'  ��  ��'  '  �  ��'  ��  ��   �  ��  p  ��  ��  �\   3�  �(  �'  ��  �>(  ��  ��   .�  ��  ��  �>(   �  9�  �	(  <�  �%\(  b(  X�   ��(  �@ �P(   ��  ��  ?1  ��  	��  ��  
��  ��  x  �+	  �  �\  ǫ  �\   ��  ��y*  R�  �i   x  �\  ��  ��  ��  ��  ��  ��  �!  ��  ?1  ��  8��  ��  <�0 ��  @�1 ��  Dn ��  H�=  �D(  P�(  �D(  `* �  pd> �  xA  �  ��/  ��  ��  ��  ��/  �y*  ���  ��  ���  �>(  ���  ��  ���  ��  �~�  ��  ���  �+	  ��K ��'  ��  ��  ���  �P(  ���  �*  �#�  ��  �y�  ��*  � �'  P(  �  x�  ��(  N�  ��*  �(  �   +  ��  	   �� !	  ͩ "�  =�  #�  ��  $\  p  %�   -�  '�*  i�  '&+  �*  6�  80�+  ߣ  2�   ^�  8�  �  9�+  c�  :�+  ��  =�  ��  >�  ��  ?�+   ��  A�  (��  Bu  0 o  +  ��  D,+  m�  D�+  ,+  Z�  (,  
H �"   ~�   �  �K !�'    ��  #&,  �+  
��  &-F$  ��  !D,  J,  !k�  �"�,  �� $$   � %�%  �"�  &�&  d"�  '�*  � d�  !�,  �,  ��  X,�,  �� .	    ��  !�,  �,  !<�  h3�,  �� 5�   ")�  6�+  0 N   �;/  S�   ��  �  �  �  z�  �  �  ��  i�  	�  
��  H�  ��  L�  I�  D�  ��  #�  R�  3�  �     !��  "^�  #=�  $��  %�  &��  'Z�  (�  09�  1.�  @��  A��  Q��  R�  S6�  T��  U��  V��  W��  X��  `��  a��  b��  c�  p%�  ���  �+�  �m�  �J�  �<�  ���  ���  �g�  ��  ��  ��  ���  ���  �o�  �A�  ���  ���  ���  �(�  ���  ���  ���  �O�  �'�  ���  ��  ���  �T�  ���  ���  ���  �I�  ���  �n�  �a�  ���  �x�  ���  ���  �`�  ���  ���  ���  ���  �}�  ���  � #,,  �	�vH     �(  N   9�/  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  V0  �\ X�   �  Y�  x  Z�   �7  \�/  	0  0�  !0  $0  	  G0  �  G0  G0  �  �   �  ��  (T  e�  .e0  k0  	  �0  �  �  �+   w�  3�0  	�0  ��  3�0  �D 50   U�  6M0  �  7Y0   
6  ".�  $h�  �#�0  	�vH        �0  @    	�0  $��  �#�0  	�vH     #�0  �	�uH     l�  651  ;1  	  T1  �*  �*  	   ��  :|1  � <�   �  =)1   	T1  ��  ?T1  	�1  Q�  A,�1  |1  0  �1  @    	�1  $��  �!�1  	@uH     �1  �1  @    	�1  %��  �"�1  	�tH     ��  &J2  + (�*   �  )�  ��  *�  �  +�  y
 ,�   	�  .�1  �  .b2  �1  &7�  C	  �3  ')�  C#�,  '�  D#�,  '�^ E#�  '��  F#u  (� H	  (�  I8,  (Jy  J5  (L�  K�*  (��  L�  (p  M�  (Q  N�'  (�V O�'  )��  h)�u  #)Ii  *B3  +n W�   *U3  (f�  l�   ,(��  ��  (��  ��  (�  �%�  (�  ��  (�  ��  (ߣ  �'�  +p ��*  ,+len �     &[  	  ,4  -p %�*  '�� %�*  'ߣ  %�  '��  %u  '�  %,4  (� 	  (��  J2   �  &��  �	  =5  '	�  �'=5  '�� �'�*  '�  �'�  '��  �'C5  '��  �'C5  '�  �'G0  '�  �'G0  'D�  �'C5  '
�  �'G0  (� �	  (?1  ��  +b ��  +p ��*  (��  ��  (��  ��  (�  ��  (�  ��  (�  ��  )��  )�u  
 �*  �  .�  Z6  '2�  &�*  '�� &�*  '.� &�  '?1  &G0  '��  &�  '��  &Z6  '��  &Z6  +min �  +max �  (f�  �  +two u  (�� �*  )�0  w)��  }*=6  +p ,�*  +lim -�*  (� .�  (��  /�   ,+mid d�  (� d�    �  /x�  ��6  0��  �-V2  1p �-�*  0�� �-�*  2 t  ��  2.� ��  3n ��  29 ��  2�  ��  3cur ��*  2� ��  3c ��   /7  {�7  0��  {-V2  1p |-�*  0�� }-�*  2 t  �  2.� �  2�  �7  3n ��  29 ��  2�  ��  3cur ��*  2� ��  3c ��  ,3v ��    �  �7  @    /��  E 8  0��  E.V2  1p F.�*  0�� G.�*  3n I�  29 I�  2�  J�  3cur K�*  2� L�  3val M�  3c N�   /��  2R8  0��  2&V2  0�  3&,4  0��  4&u   4L�  �	  �B     #      ��:  5�  �%�  x: p: 5Z�  �%�  �: �: 52�  �%�  ; o; 5Y�  �%;  << .< 6�  �8,  �< �< 6� �	  J= >= 6�  ��*  �= �= 6n[ �\  M> E> 6%] �\  �> �> 6/< � \  :? 6? 7�u  S��B     7��  ϶B     7�Y F	��B     8��  6j �P(  t? p? 6Jy  �5  �? �? 9�  �:  6.� �  @ @ 6�  �  c@ _@ 6��  	�  �@ �@ 6��  
�  NA JA 65$  �  �A �A 62�  �*  �B ~B 6��  u  �B �B 6/�  u  $C  C :p �*  rC ZC 6N�  \  vD jD ;��B     %       6�\ C�  �D �D   <۶B     �s  �:  =U}  <�B     �s  �:  =U}  >�B     �s  =U}    4�  7	  `�B           ��F  5B�  7 �  5E E 5g�  8 �  HF 8F 5n�  9 �  G �F 5:1  : O  DH ,H 6 <�,  _I GI 6�  =�,  rJ bJ 6� >	  +K #K 6�  ?8,  �K �K 6��  @�'  �K �K 6�S  A�F  BL *L 6��  B�  oM iM 7�u  ���B     9 �  \>  %C!  n�  ��6N o�F  �M �M 6�  po   N �M 6S�  q�  KN IN 6�  q&�  pN nN 6C�  ru  �N �N ?��B     �       2>  :n ��  �N �N 6�� �	  O O 6�� �	  )O 'O :vec �;  SO MO @�o  �B      @�  �C=  A�o  B�o  �O �O 8@�  C�o  �O �O C�o  !P P   D�o  =�B      =�B            ��=  A�o  A�o  ;=�B            C�o  `P \P C�o  �P �P   @�o  d�B      p�  � �=  A�o  B�o  �P �P 8p�  C�o  Q Q C�o  JQ FQ   E�o  ��B      ��  � A�o  A�o  8��  C�o  �Q �Q C�o  �Q �Q    F��B     �s  >��B     �s  =Uv�=T��  @�[  ��B       ��  i�>  B\  R R B\  ER CR B \  lR hR B�[  �R �R B�[  �R �R F��B     �s  >%�B     (\  =Uv�=Tw =Q��=R| =X��~  Eh2   �B      ��  SB�2  DS 4S B�2  ST GT B�2  U �T Bz2  �U �U 8��  C�2  �V {V C�2  �W �W C�2  
X X C�2  5X /X C�2  �X �X C�2  �X �X C�2  7Y 5Y C	3  oY iY G3  O�B     H3  G(3  0�B     I13   �B     O       �?  C63  �Y �Y  JB3  0�  �A  CG3  �Y �Y @I5  ��B      ��  |FA  B�5  tZ nZ B�5  �Z �Z B�5  0[ *[ B~5  [ y[ Bq5  �[ �[ Ad5  BW5  \ \ 8��  C�5  e\ _\ C�5  �\ �\ C�5  /] '] C�5  �] �] C�5  �] �] G�5  ��B     G�5  M�B     J6  `�   A  C
6  �^ �^ C6  �^ �^ C"6  8_ 2_ C/6  �_ �_  K=6  ��  C>6  ` �_ CK6  �` �`    <��B     �s  _A  =Uw  <��B     �s  xA  =Uw  >��B     �s  =Uw   KU3  ��  CV3  �` �` Cc3  Wa Ma Cp3  �a �a C}3  �b �b C�3  Ec 9c C�3  �c �c C�3  �d �d @24  E�B       �  �C  B�4  Af =f B�4  �f �f B�4  �f �f B�4  g 	g Bx4  Qg Mg Bk4  �g �g B^4  �g �g BQ4  Qh Ah BD4  i 	i 8�  C�4  Qi Mi C�4  �i �i C�4  �j �j C�4  nk 6k C�4  �m �m C�4  �n }n C5  �o ~o C5  Pp <p C5  7q #q H*5  H35    J�3  @�  F  L�3  @�3  "�B      ��  �E  B4  r 
r B�3  �r �r B�3  8s 2s A�3  B�3  �s �s 8��  C4  Jt Dt C4  �t �t D 8  >�B      >�B     *       !�C  BE8  �v �v B98  �v �v B-8  �v �v  M`6   �  .	sD  A�6  By6  w w Am6  8 �  C�6  ?w ;w C�6  yw uw C�6  �w �w C�6  �w �w C�6  ^x Rx C�6  �x �x C�6  ?y 1y C�6  �y �y   D�7  $�B      $�B     �       &	'E  A�7  B�7  az [z B�7  �z �z ;$�B     �       C�7  �z �z C�7  { { C�7  A{ 5{ C�7  �{ �{ C�7  | �{ C	8  �| �| C8  }  }   N�6  ��  *	A7  B7  �} �} A�6  8��  C7  ~ �} C'7  �~ �~ C37  �~ �~ C?7  L J CI7  u o CU7  � � Ca7  B� >� Cm7  �� x� Cy7  1� '� O�7  /�B            C�7  �� ��      >�B     �s  =Uv   <9�B     �s  F  =Uw  F��B     �s  F��B     �s  <�B     �s  LF  =U|  <.�B     �s  lF  =U| =T�� >�B     �s  =Uw      G  a  Pf�  -��B     �       �?G  5B�  - �  "� � 6 /�,  t� n� E�j  ��B       �  2B�j  Ă �� 8 �  C�j  �  � <һB     �s  (G  =Uv  >�B     �s  =Uv     4��   	  0�B     H       ��G  5B�    �  +� %� 6 "�,  }� w� 6��  #�  ˃ Ƀ E�j  E�B      P�  &B�j  �� � B�j  � � Fq�B     �s    Q��  D	  0�B     B      ��Q  RJy  D!5  n� V� R�  E!�  �� w� R�  F!�  �� �� RG  G!�  H� D� RG  H!3  �� �� S�  J8,  և �� S� K	  � ߈ 7�u  �B     90�  cI  S�   a�  	� � TEZ  ��B      `�  dBqZ  D� @� BdZ  �� �� BWZ  ى Չ 8`�  U~Z  ��C�Z  � � C�Z  �� �� H�Z  <��B     �s  EI  =Uv =T}  >��B     �s  =Uv =T��    90�  �J  S�  ��*  �� ܊ 9p�  �I  Vnn ��   � �  ?"�B     �       FJ  Vn ��  Y� W� S.� ��  � }� S�  �  �� �� S�V ��'  �� � SR�  �i  F� D� >C�B     �s  =T =Q0=Rv ����=X0=Y��  9��  �J  Vmax ��  t� n� S.� ��  ǌ �� S��  ��'  +� '�  8��  %�� s  ��>��B     t  =U	�vH     =T0=Q��=R0   W�Z  C�B      ��  T]K  B�Z  g� a� B�Z  �� �� 8��  C[  � � <N�B     �s  3K  =Uv =T0 >|�B     t  =Uv =T	@uH     =Qs�   X�Z  ��B      ��B     /       X�K  B�Z  o� m� ;��B     /       C�Z  �� ��   WnY  k�B       ��  xnN  B�Y  �� �� B�Y  � � A�Y  B�Y  .� *� B�Y  h� d� 8��  C�Y  �� �� C�Y  ӏ Ϗ C�Y  � � C�Y  W� O� U�Y  ��GZ  C�B     GZ  3�B     GZ  ;�B     JZ  ��  �M  CZ  � Ő C)Z  |� x� C6Z  �� �� @�[  ��B      0�  ��M  B�[  H� F� B�[  m� k� Y[  ��B      ��B     8       �BF[  �� �� B:[  �� �� B.[  �� �� B#[  � �� ;��B     8       CR[  � 
� C^[  <� 0� Ch[   �� Ct[  � � C�[  1� -� H�[  H�[     <�B     �s  �M  =Uv  >(�B     �s  =Uv =T|   <p�B     �s  �M  =Uv  <��B     �s  �M  =Uv =T�� <��B     t  N  =Uv =T
 5���� <��B     �s  9N  =Uv =T�� <��B     *t  XN  =Uv =T�� >C�B     �s  =Uv    T�Q  u�B       `�  �BR  y� u� BR  �� �� BR  )� � B�Q  �� �� 8`�  U,R  ��C9R  � � CFR  �� }� CSR  )� � C`R  "� ޙ CkR  � � GxR  ��B     G�R  ��B     G�R  ��B     J�R  ��  �O  C�R  ڝ  C�R  ޞ ؞ K�R   �  C�R  5� '� C�R  � ܟ >��B     fS  =Qw    I�R  ;�B     �       �O  C�R  C� =� C�R  �� �� >��B     �s  =Uw =T4=Q0=R| =X0=Y��  J�R  @�  yP  C�R  Π ʠ C�R  � � CS  B� >� JS  p�  CP  CS  � y�  >��B     �s  =Uw =T@=Q0=R} 
��=X0=Y��  @[  ��B      ��  fGQ  B:[  ̡ ȡ BF[   � � B.[  Т Ƣ B#[  C� ?� 8��  CR[  �� �� C^[  � ԣ Ch[  �� �� Ct[  � ݤ C�[  9� 3� H�[  H�[  K�[   �  C�[  �� �� Z�B     =T} =Q|     <��B     �s  gQ  =Uv =T�� <��B     �s  �Q  =Uv =T|  <��B     �s  �Q  =Uv  >��B     7t  =Uv     /��  ,�Q  0�  ,�  2�  .8,  2R�  /i   &��  6	  !S  '�  6#�*  'Jy  7#5  'x  8#\  '�  9#\  (� ;	  (R�  <i  (?1  =�  (��  >�  +p ?�*  (�� @�*  )�u  )��  )�0  *�R  +q u�*  +q2 v�*  ,(ss  ~�  (� ~�    *�R  +n ��  (.� ��   ,+n ��  (.� ��  (�V  ��  ,+cur ��'     .��  
fS  '�  
#�*  'R�  #i  ,(j #P(  (�@ #P(    4��  �	  оB     �       ��T  [p �#�*  � �� [len �#�  �� �� 5R�  �#i  �� � 5~�  �#�T  �� �� %� �	  �L6E  �  &� � :n ��  ƨ �� :ok ��  (� $� 7�u  ��B     <��B     �s  PT  =U}  <U�B     Dt  zT  =U} =Ts����=Q�L >n�B     Pt  =Tv =Qs     4��  s	  ��B     �      ��U  [p s3�*  }� i� 5�� t3�*  a� U� 5�  u3�*  �� � 6j wP(  �� }� 6� x	  :� 8� 6R�  yi  d� ^� 7�u  ��B     7��  ��B     9��  �U  6��  ��  �� �� 6��  ��  j� T� :q ��*  R� 6�  <��B     Dt  �U  =U} =T =Q�L <�B     �s  �U  =U}  > �B     �s  =U}   4��  F	   �B     �       �W  [p F0�*  3� #� 5�� G0�*  � �� 5�  H0�*  l� d� 6.� J�  ٳ ˳ 6U�  J�  �� �� 6��  J!�  � � 6��  K>(  X� J� %� L	  �L6R�  Mi  � � 7�u  e^�B     7��  h^�B     >��B     �s  =T4=Q0=R} ����=X0=Y�L  4 ,	  P�B     u       �	X  [p ,-�*  d� Z� 5�� --�*  � ٶ 5�  .-�*  M� C� %� 0	  �\6R�  1i  ȷ · :len 2�   � � 7�u  ?P�B     <��B     Dt  �W  =Tv����=Q�\ >��B     Pt  =T| =Qv   4��  �	   �B     �      �nY  [p �1�*  � Ÿ 5�� �1�*  L� B� 5�  �1�*  ƺ �� 6R�  �i  )� %� 6�V ��'  o� _� 62�  ��  C� ?� :n ��  �� �� 6.� ��  �� �� 6��  ��  � � 6� �	   � � 7��  @�B     7�u  :�B     ;X�B     O       6�:  ��  H� D� >z�B     �s  =T(=R�������=Y��   &%�  G	  EZ  '�  G#�&  'Jy  H#5  -idx I#�  '��  J#\  '_�  K#u  (^�  M�  (?1  N�  (x  O\  (�  P\  (� Q	  )�u  �)��  �)�0  �,+p f�*  (�� g�*  (��  h�    &T�  !	  �Z  'Jy  !"5  '��  ""\  'A�  #"C5  (� %	  (.� &�  (E  '�  )�u  @ &��  u  �Z  '� !
&  (E  u   \<�  �	  [  0� � 
&  0Jy  � 5  2� �	   \��  �	  �[  1pp �*=5  0�� �*�*  0^�  �*�1  0��  �*	  2� �	  3p ��*  2��  ��  2J�  ��  2Y  �%�  ]��  �]�u  �,25$  ��1    \��  ~	  �[  1pp ~$=5  0�� $�*   &��  C	  (\  ')�  C�+  'Jy  D5  '��  E�  'x  F�  '�  G�   4��  �	   �B     2      �f  5)�  �"�+  �� �� 5Jy  �"5  � � 5��  �"�  v� N� 5x  �"�  5� 1� 5�  �"�  �� n� 6� �	  �� t� :p ��*  \� D� 6�� ��*  b� \� 7�u  =8�B     9�  <a  :n ��  �� �� 6��  ��  �� �� 6.� �%�  �� �� 6��  ��  *� $� 62�  ��F  |� v� 9 �  �^  :i ��  �� �� 6��  ��  � � 62]  �&�  �� �� 6�l   +  &� � ?o�B     v       �^  :vec ;  �� �� @�o  ��B      `�  =^  A�o  A�o  8`�  C�o  *� &� C�o  m� i�   E�o  ��B      ��  A�o  B�o  �� �� 8��  C�o  �� �� C�o  +� '�    ? �B     8       �^  :vec ";  h� f�  >-�B     (\  =U =T~ =Q��~  @f  ��B      ��  ��`  B�f  �� �� B�f  {� C� B�f  �� �� 8��  U�f  ��C�f  e� _� C�f  �� �� C�f  � � C�f  �� �� C�f  1� -� Cg  {� i� Cg  p� b� Cg  %� � C)g  �� �� H6g  H?g  GHg  ��B     JQg  @�  �_  CVg  �� �� >��B     �s  =T =R} ����=Y��  @�[  
�B      ��  H�`  B�[  !� � B�[  F� D� Y[  
�B      
�B     ^       �BF[  p� n� B:[  p� n� B.[  �� �� B#[  �� �� ;
�B     ^       CR[  �� �� C^[  !� 	� Ch[  4� .� Ct[  �� � C�[  1� %� H�[  H�[     Kdg  ��  Ceg  �� ��    <��B     �s  a  =U~  <��B     �s  'a  =U~  >@�B     �s  =U~   @tg  ��B      0�  8@f  B�g  o� a� B�g  R� � B�g  e� W� 80�  U�g  ��~C�g  � �� C�g  �� }� C�g  � � C�g  �� �� C�g  �� �� C�g  � � C�g  �� �� Ch  m� c� Gh  J�B     Gh  J�B     G"h  J�B     H+h  G4h  ��B     @�[  M�B      ��  U�b  B�[  �� �� B�[  � � T[  M�B      л  �BF[  a� ]� B:[  a� ]� B.[  �� �� B#[  �� �� 8л  CR[  � � C^[  i� S� Ch[  e� ]� Ct[  �� �� C�[  �� �� H�[  H�[     @j  ��B       �  Z(c  B*j  �� }�  JPh  0�  �e  UQh  ��C^h  �� �� Kkh  ��  Clh  q� c� Cyh  A� 3� C�h  �� �� C�h  �� �� C�h  F� 6� J�h   �  �c  C�h  �� �� C�h  �� ��  D�h  ��B      ��B            
%d  B�h  -� +� <��B     �o  d  =Uu =Tt ^Dj    F�B     [t   @�h  �B      @�  �d  Bi  X� P� Bi  �� �� 8@�  Ci  �� �� C(i  !� � < �B     �o  �d  =Uu =Tt ^Dj    <g�B     Tq  �d  =Q��^�i   ^�i  �� >��B     gt  =U��~=T1=Q1   @5i  ]�B      p�  �e  BFi  ]� W� BFi  ]� W� BRi  �� �� B^i  � �� Bji  \� V� 8p�  Cui  �� �� C�i  �  � C�i  f� ^� G�i  *�B     J�i  ��  �e  C�i  �� �� C�i  �� ��  >�B     gt  =U��~=T3=Q0   >��B     Tq  =Q��^�i   ^�i  ��   O=h  ��B     H       CBh  � � >��B     �s  =T8=R��~�����=Y��~    <K�B     �s  df  =U~ =T��~�R" >{�B     �s  =U~ =T}   &   /	  tg  ')�  /'�+  -p 0'�*  '�� 1'�*  (� 3	  (��  4�  (R�  5i  (�l  6+  (?1  7�  +i 7�  (.� 7�  ({�  7&�  (�s 8�  (��  8�  )��  �)��  �)�u  �*dg  (�:  Y�   ,(ߣ  p�    \g�  �	  �h  0)�  �%�+  1p �%�*  0�� �%�*  2� �	  2R�  �i  2?1  ��  2AX ��  2_�  � �  3i �)�  2.� �,�  2� �3�  +x  �  )��  &)��  %)�u  ")��  �	)"�  	*Ph  (�:  (�   ,+pos ^�h  +cur _;  ,(ߣ  g�  (��  g�  (\�  g&�  (A g7�  +n gC�  ,+idx ��  (� ��      �  �h  @    /��  ��h  0)�  ��+   \��  �	  5i  0)�  �"�+  1to �";  2��  ��  2� �	   \z�  �	  �i  0)�  �#�+  0*�  �#;  03�  �#;  1to �#;  2��  ��  2�S  ��F  2� �	  ]�u  �,3vec �;  3tag ��*    \��  	  j  0)�  "�+  1to �";  2��  ��  2�S  ��F  2� �	  ]�u  �,3n ��    /��  x7j  0)�  x�+   /}�  O�j  0)�  O'�+  2��  Q�  2�S  R�F  2k� S�  2N� S�  ,3p1 c;  3p2 d;    /��  5�j  0)�  5�+  2R�  7i   /��  (�j  0)�  (#�+  0��  )#�   Q�  �+  ��B     
       �Rk  R~ �&�  N� J� R�1  �&$  �� �� _ʿB     st  =U	�vH     =T�T  QC�  c	  пB     �       �Wl  R�  c�  �� �� R��  dG0  1� +� R��  eG0  �� }� R��  f�  �� �� R��  g�  >� 6� S�  i8,  �� �� SL�  j�*  � � S�� k	  � w� S�� k	  �� �� S�  l�  :� 6� F�B     �t  F4�B     �t   Q�  B	  ��B     5       �m  `�  B�  URn�  C�  v� p� `��  D�+  QS�  F8,  �� �� S� G	  �� �� a�u  ]ȵB     ;ȵB            SL�  S�*  '� %�   \�  	  bm  0�   �  0�    �  0�� ! �  0 �  " ;  2�  $8,  2L�  %�*   Q��  c\   �B     �       �?n  `
H c#,  U`��  d#|#  TSE  f�  a� M� S��  g\  >� 4� a��  j
�B     a�u  ���B     8`�  Vmin l�  �� �� Vmax m�  7� +� Vmid n�  �� �� S��  o�'  q� ]�   Q��  F�  ��B     h       ��n  `
H F#,  U`��  G#\  TVmin I�  �� �� Vmax J�  � �� 80�  S��  O�'  �� r� Vmid P�  ~� p�   b��  >��B            �o  `
H >,  U Q��  	   �B     V       ��o  `
H ,  URm  	  � � S� 	  T� P� S�   8,  �� �� a�u  8p�B     8 �  Vn +�  �� ��   \�6  �O  �o  1a �O  1b �O  3ret �"  3tmp �"   c7j  p�B     �       �Rp  ADj  ADj  CPj  �� �� C\j  � � Chj  @� :� Ctj  �� �� K�j  ��  C�j  �� �� C�j  � �   cm   �B     t       �Tq  Bm  [� O� B%m  �� �� B1m  $�  � B=m  i� ]� CIm  �� �� CUm  �  �  Jm  �  q  B%m  1 + B1m  � � B=m  � � Bm  J B 8�  LIm  LUm  Fq�B     �s    <1�B     R8  Fq  =Us =T�T=Q�Q=Rv  F��B     �s   c�i  ��B     q       ��q  A�i  A�i  A�i  C�i  � � C�i    C�i   } Gj  ��B     Ij  ��B     "       �q  Cj  � �  >�B     gt  =T1=Q0  c�Q  ��B     �      ��s  B�Q  � � C�Q  A 9 L�Q  K�Q  0�  B�Q  � � 80�  L�Q  C�Q  � � W!S  ��B      `�  <ns  B<S    B/S  @ < JIS  ��  �r  CJS  � | CWS  � � >��B     �s  =Uv   <��B     �s  �r  =Uv  <��B     �s  �r  =Uv  <��B     �s  s  =Uv  <�B     �s  )s  =Uv  <N�B     �s  As  =Uv  <s�B     �s  Ys  =Uv  >��B     �s  =Uv   >�B     �s  =U}     d9  9  cd�3  �3  �dxL  xL  �djO  jO  e�,  �,  �eC  C  `dT)  T)  �eF\  F\   �d>Q  >Q  �e�6  �6   �d�3  �3  1d�N  �N  �d _   _  hd*  *  �dF  F  me�K  �K   vf�D  �D  ! eo+  o+  �e],  ],  ed�*  �*  [d5<  5<  ? ��   �5  �  � $"  ��B     %      �x X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  	0  >   G   �	  	N   �  B"b  h     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  V  -      n�  �  �  V  U    �  ��    U   "  V  -   -   U    �  �".  4  �   PJ�  2�  L1   �  M@   pos N@   �  P�  SF  Q�   �1 R  (=9 S>  0R�  UV  8y�  V1  @�� W1  H �  ��  �\ �-   m  �U    o  ��  �  �    @   1  "  @   1  @    7  �  2  K  Q  \  "     :-   �  J�  x L\   y M\   )  Oh  	�  B   s�  M   u\   }  u\  V  v\  /  v\   t
  x�  k	  (j  �  N    ��  N   �  	G   B� 
1  L  0    7  s  7  v	  U     �  �  	j  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     �  )    Y|  �  =  N   �<  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "V  \  �  %  <�  x >)   len ?0  *� @7   %  Ba  	�    `�  �  �  G   G   �  U    �  �  q�  �  G   	  G   G   U    �      1  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  �	  0R   �U   8�  ��  @ w  �  �  �1  	�  �   �  �  G     U      I  �      (  I   �  ?5  ;  P  I  1  @    �  Y]  c  G   |  I  @   U    s  ��  �  G   �  I  �   �  W  0�  �  �<   e� ��  �� �(  �� �P  �� �|   �� �
  ( �'  ��  �!  	l7  �  	�1  �  -  	�7  	8  D  �  	��   	O  �
  	�)  �  	�0  �  	�G   
  	�N   �  	�-   \#  	�@   �  	 -   �  	,G   \&  	7U   �0  	D4   b   	�	  xx 	��   xy 	��  yx 	��  yy 	��   a  	��  		  z'  	�\	  m  	�I   ss  	�x   �  	�1	    	�v	  |	  �	  U    �  	��	  �U  	�U      	�i	   %  	��	  �  	$�	  �	  �  	 
  �� 	"�	   �@ 	#�	  �U  	$U    �  	76
  �; 	9�	   ��  	:�	   L  	<
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @
=  ��  
?\   �  
@\  ~  
B\  �  
C\  �  
D\   5  
F\  (B  
G\  0�  
H\  8 �	  
J�  
   
sg  �  
u`   ��  
v`  �  
x\  �
  
z\  (  
{\   �  
}  �  
�#�  �  k  `�6  R�  �V   (  �x  |  �x  �  �x  �  ��  �  ��/  v  �6
  �  ��  (�%  �6  07&  ��/  8G   �x  X �  
�"C  I  h  �  �M �/   k  t  R�  V   �  
�"�  �  %  8;�  �� =�/   �M >=    ?6
   r$  @�+  0 5  
�$�  �  %  �`  �� �/   �M �/  �  <   �  K(  (�� 
I  h�� |  p�� �)  x K  
� m  s  �  �
,4  �   
.�   �  
/�  O  
1�  C  
2�  �  
4�   d> 
6�  (A  
7�  0T  
9x  8  
:�  @�  
<x  H�  
=�  PE-  
?�	  X�!  
D�  h:  
Fl  �  
G`  ��  
H`  ��  
I`  ��  
K`  �  
L`  �U  
N`  ��  
O`  �)�  
Q�  ��  
R4  ��� 
S�  �K1 
W�  �R�  
XV  �Jy  
Y"  �%  
[6
  ��	  
]�	  �    
^U   ��8  
`$  � L  
 A  G    X
��  �  
�`   E-  
��	  N 
��  �8  
��  P �  
*%�  �  �  0
t�  k  
vt   �  
w`  �@ 
x�  ݖ 
y�  E-  
z�	   N 
|  0�  
}�  pR  
~�  x�  
�  �ߣ  
�<  ��I 
�j  ��  
�x  �h  
�x  ��S  
��  �4  
��  �8  
��  �  
�U    �  
�-   �  
�\  o  
�\  �L 
�U    �8  
�  ( �
  
L#�  �  W  
HE  �  
J`   = 
K
    
Ll  d  
Ml   �  N   
�
  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  
E  (0  
O�  #   
g)1  7  �   ���  =  �	   L  ��   $  �x  0�  �'  8m  �#}-  h�  �%  pآ  �<  tG   �x  x O  g  �  �?  
ds  �
  
�)�  �  �   H�!  �  �U    "  �N  �!  ��   ~	  8
f�  �
  
hl   (  
il  �� 
k�  �� 
l�    
n\  �  
o\   �  
p\  (�  
q\  0 y  
s!  �a  
�G    
�$�  �  �  0'  �N  )x   ?1  *l  }0  +x  i/  ,x  � -	   �  
�))  /     H��  ��  ��+   ?1  ��  (  �  4  �	  \  ��  0  �U   @ ��  
��  +!  
�  tag 
�   �U  
�   �  
�  �M  @
WV  ?1  
Y�   �I  
ZI  N  
[�  SF  
\�  Jy  
]"   K1 
^6  (G  
_x  0G  
`V  8 �  �O  
b�  `  N   

�  w%   }#  �&  h  �  &     

i  E   
9
  � 
;
�   ��  
<
�  �  
=
�  �  
>
�  �#  
?
�   �  
L
(  �  �  N   
�N  :   �   ^$  1  �!  �!   :  
�  �  ��  �#  �s  y  �  �  6   I$  ��  �  �  6   �&  ��  �  [  �  6  �   �   �!  H�T  �  ��   S"  ��     �T  �"  ��  �  ��   ;  ��  (%  �g  0�   ��  8��  ��  @ [  R  ��  x  =v	  P     �  �  �  "  `  x  x  V   �  &�  �  �  `   �%  *�  �  �  �  4   �%  -�  �    4   {  1    �  $  �   �  40  6  A  �   l  8M  S  �  g  4     �  <s  y  �  �  4  �   �  @�  �  �  �  �  4  �  <   �  G�  �  �  �  `  �  �  �   �'  N�  �  �    `  "   �  S  %  �  H  `  �  �  <  H   �  &  ��,  �� �Z   i'  ��  H   ��  P  ��  X�A �s  `Y ��  h�#  ��  p�  ��  x�  �  �  �$  ���  ��  �U�  ��  ��!  ��  ���  �  ��  �A  �&  �g  �   �N  	,  �&  �I  N  
   ".8  �  8Y�  ��  [�   Ǧ  \�  ��  ]�  d> ^�  ��  _�   I�  `�  (�  a  0U  b`  2�  cl  4 ��  e[  ��  p$�  [  � }�  ��  ��[  ֤  �x   Ğ  �x  ��  �8  �  �8  	��  �8  
�  �8  ��  �[  �  �k  (��  �[  <�  �k  X��  ��  p��  �x  x��  �x  |��  �{  ��  �{  �R�  �8  ���  �8  ���  �  �F�  �  �V�  ��  ���  ��  ���  ��  �"�  ��  ��  ��  �@�  ��  � `  k  @    `  {  @   	 l  �  @     `  �  @    `  �  @    ��  �  o�  �#�    �  ��  ��    2]   8   U�  !  5�  "H   �  �  $�  ��   *�  m�  ,�   `h  -�  �  /�  #�  0�  (��  1   ��  3H  z�  4H  ��  6   ��  7/   ��  9�  (Ԯ  ;?   0��  CU   ���  D�  � �  �  @    H     @         @    �  /   @    �  ?   @    O   O   @    �  �  e   @    ��  Fr   !  �  N   0�   ��   r�  �  E�  Ϊ   H�  8x   �  N   w�!  U�   ��  ��  �  ��  ��  ޟ  $�  ��  �  	t�  
�  ܖ  �  ��  ��  d�  {�  ך  ʕ  �  ��  ��  m�  ,�  �  ^�  ׭  ~�  @�  �  ��  N�   ��  !��  "��  #ݴ  $��  %�  &�  ',�  (a�  )��  *x�  +��  ,"�  -"�  - a�  ��   ��  )$�!  "  H�  ��  ,"  "  �  4"  V  4"  :"   �  �!  ��  1L"  R"  q"  �!  �  �  �  �   ��  8}"  �"  �"  �!   �  ;�"  M� =	"   �� >@"  Յ ?q"   ��  A�"  �"  �  h!�"  �"  ��  ��  u-�"  o#  ��  8Vo#    X�"   j�  Yt#  =9 Z�#  �� [�#  Q� \�#   �� ]�#  (�� ^$  0 	�"  ��  ��#  �#  �#  �"   ��  ��#  �#  �#  �"  �  H   K�  ��#  å  ��#  �#  �#  �"  �   ��  
�#  �#  �  $  �"  �   ?�  1$   $  �  >$  �"  >$  �!  N   �  1�  �!Q$  W$  $�  ��  �-i$  �$  .�  8��$    �D$   j�  ��$  =9 ��%  �� �%  +�  �0%   �� �]%  (�� ��%  0 	o$  ǡ  ��$  �$  %  D$   ��  �%  %  0%  D$  �  x  H   ��  �=%  C%  ]%  D$  �  �  I   !�  &j%  p%  �%  D$  �  I   K�  D�%  �%  �  �%  D$  �   	�  k�%  �%  �  �%  D$  >$  �!  N   ��  �&  ��  �%&   X� �:&  l� �O&   �"  %&  6   &  �"  :&  6   +&  \$  O&  6   @&  $�  ��%  �  � o&  U&  �>  ��&  'O  ��   xC  ��   s/  �u&  	�&  �  0t'  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�&  �3  5D'  num 7x  str 8�   +P  :'  �J  =x'  key ?D'   �U  @4    �7  D$�'  P'  O  H�'  �'  �  �'  �'   D'  �Z  K�'  �'    �'  �'  �'   �S  (O3(  �� Q�   �  R�  �6 S�  �B  U�'  3  V�'  >) X3(    x'  e-  \ E(  �'  H  E#\(  	K(  �  @J�(  �  L�   �  M<  �� O,)  .� PR)  �  Q�)   �  Ro)  (�!  S�)  08'  T�)  8   W!�(  �(  -  (l&)  k  nt   �M o&)  ߣ  p<  �  q�   W(  k  )8)  >)  �  R)  �(  �   w   .^)  d)  o)  �(   �  1{)  �)  �)  �(  �)  �   ,	  K  6�)  �)  �)  �(  O    �  :�)  �)  �  �)  �(  �(   �  >8)  "  Y�)  *  �   *  �  �  N  �   �  _,*  2*  �  P*  �  �  �)  �   $  f\*  b*  w*  �  �  O    �  l�*  �*  �  �*  �  �  �   #  x�+  �� � Z   �  � <  H  � �)  P�  �  *  X9!  � P*  `l� � w*  h  � +  p     ��*  �  H2l+  �S  4�   �  5�  (  6�  04  7�  88  8�  @ �  :+  �  �=�+  R�  ?V   �  @�  n  A�  �  B�  1$  C  2�  El+  �� Fl+  `�L HU   � �  J�+  x+  U   �  U',  ,  m  D   t_,  �  v�   A  w�  �  x�  &  y�   !  {,  �  �w,  },  �  �,  ,  �  �,   \	  �  ��,  �,  �,  ,  �,   �'  ��,  �,  �  �,  ,  �    �,   _,  �!  --  ��  )k,   ��  )�,  �  )�,   }  �,  	--  O  ;j-  _� =%j-   ݰ  >%,   :-  �  @?-  p-  cA  �,�-  �-  /  ��-  �� �   �M ��-   ?<  �,�-  _.  �5  P�_.  �  ��   �� �p.  �Y ��.  �H ��.  U@ ��.   �9 �#/  (�A  �#5/  0�^  �#`/  8�^  �#�/  @N7  �#�/  H 	�-  ��  ��-  (Z  �|.  �.  �  �.  �-  �   17  ��.  �.  �.  �-   �G  ��.  �.  �  �.  �-  I   %G  ��.  �.  �  �.  �-  �.   I  �@  �/  /  �  5/  �-  �-  I  I   �;  �A/  G/    `/  �-  I  I   �W  �l/  r/  �.  �/  �-  V   *;  ��/  �/  �.  �/  �-  V  I   �T  ��/  Z  �  I  +  -1  B�  6  �/  @    f  0  @    	0  �  0  `   0  �  <0  `  �  �  �   B0  �  V0  `  �    �  �%  ��  #o0  u0  I  �0  �   d�  )�0  �0  �  �0  �   0�  /�0  K�  6�0  �> 8I   �^ 9�   �  ;�0  Ѽ  >$�0  �0  ў  (@,1  
H Bd.   ��  C�  XT D,1    �0  6	 F�0  ��  NJ1  P1  �  d1  �  �   B�  Vp1  v1  �1  �  �   ��  Z�1  �1  �  �1  V  �0  �  >1  d1  �   ��  b�1  �1  �  �1  �0  I   ��  f�1  �1  I  2  �0  �.   ��  @j�2  �\ l c0   8` n �1  �\ o �1  �_ p �1  �T r �0   }�  s �0  (ʬ  t �2  0�  u �2  8 	2  ��  j�2  �2  7  7�   F�2  ~�  Hx   ̰  Ix  V�  Jx  �H L�2  �  M�2   l  �  b�  O�2  �  O3  �2  ��  W33  ��  Yl    ��  [3  !�  ^�4  �  `�   8�  a33  8-�  b�  @"�  c�   "E�  e�   ("= f�2  0"�  h�4  P"
�  i�4  X"��  j�4  `"��  lx  h"��  m�4  p"h�  n�4  x"��  o9(  �"�  qx  �"V r�2  �"� s�4  �"'�  t�4  �"��  v8  �"�  w8  �"��  x	  �"w�  y�  �";�  z�  �"* {�   "ܲ  }�   8  �4  �  �  ?3  �  �4  ?3  ��  (�5  �9  �x   ��  ��  ɲ  ��  �  ��  �  ��    T�  �&5  �4  ��  �j5  ��  ��   ��  ��  x �x  y �x   �  �v5  ,5  z�  X��5  ��  �   ��  ��  �Z  ��  (%?  ��  0L�  �5  8)�  ��  @W�  �j5  HѺ  ��  P b�  ��5  |5    6  @    �  $6  @    !*
 �!�6  �� #�   �6  $�4  �"s  %�  "Q  &�  "Q *�4  "� +�   "� ,`  ("B�  -6  0"�  .6  P"O /21  ` � 1�6  $6  �
 `%�6  �� '�   �k  (4  X D *7  �6  !� 8.37  �� 0�   "�q  1�  0 G 3?7  	7  0 @7m7  �� 9�/   � :=  8 �	 <y7  E7  N   ��9    
 � ] X �  | 9 � 	� 
� � z � � � � V � �
 t  u	 !o "n #P $� % &_ 'V (`
 0| 1~ @� A, Q R� S Ty
 U� V W� X� `� a� b c� pG �^ �� ��
 �Z �M �C �	 �� �� �< �y � �. �� � �� �� �d � �� �� �� �< �� �O �� ��	 �_ �x ��
 �� �� �� �J
 �E	 �l �= �� �� � �� ��	 ��	 � �� �p � f.  &0  <B  ,<0  %�  0�9  	�9  �3  0:  tW 2!�9   i�  3!�9   FO  )0  ��  ,0:  	:  Y  ,K:  6 .:    =�  !W:  ]:  �  q:  `  q:   �  T�  %�:  �:  �  �:  `  �:   33  ��  )�:  �:  x  �:  `   �  ,�:  �:  �  �:  `  �:   �  ��  0�:  ;  �  %;  `  �!  �  U   �   �  76;  	%;  ,�  (7�;  ۽  9K:   1�  :w:  G�  ;�:  #�  <�:  )�  =�:    #c \)�9  	�|H     #� p*+:  	�|H     ## �&1;  	`|H     �&  �;  @    	�;  #� �#�;  	 |H     $O  �	@{H     �6  `S�<  �<  U�   �Q  V�  a(  X�  VA  Y�  Q) [l   nX  \l  "�D  ^�<  (�5  _�<  8M   a`  H}  b`  JV  c`  L/  d`  N7K  fl  P>D  gl  R�:  i`  T�3  j`  V=]  k`  X �  �<  @    �5  m<  �Q  8��=  �  ��   �Z  �`  %?  �`  
L/  �`  �<  �l  �Y  �`  �7  �`  �)  �`  �O  �`  �H  �`  vH  �`  ^  ��=  �>  �`  $�7  �l  &0>  �U   (�+  �U   0 `  �=  @    �H  �=  �?  8A�>  �  C�   �Z  D`  %?  E`  
L/  F`  S.  Hl  �W  J`  �W  K`  C  L`  �O  M`  �H  N`  vH  O`  ^  Q�=  �>  S`  $�B  Tl  &0>  ZU   (�+  [U   0 �]  ]>  �B  �|2A  ��  ~l   �)  `  �)  �l  �.  �l  U  �l  �V  �`  
�0  �`  �6  �`  �C  �`  U?  �`  6P  �`  �C  �`  &L  �`  *J  �`  �L  �`  HP  �`  N*  �2A   [2  ��  0k2  ��  8.  ��  @{2  ��  HQ2  �BA  P�0  �l  Tp4  �l  VmU  �l  X�Z  �`  Z ?  �`  \:  �`  ^�I  �l  `E8  �l  b�;  ��  h�;  ��  p�O  �`  xDF  �`  zfV  �l  |�9  �l  ~[9  �l  ��G  �l  �zQ  �l  � 8  BA  @   	 %  RA  @    {D  �?  �1  @��A  �I  ��   6Y  ��  �^  �`  S  �`  )  ��  @3  ��   �0  ��  (4C  ��  0�C  ��  8 aM  �_A  �I  @��B  �  ��   _7  ��  )  �l  �O  �l  �n �l  �T  �l  EF  �l  I  �l  �K  ��B  N:  ��B  ,L  ��B  4�E  �%  :�Z  �%  ;�Z  �8  <^  �8  = %  �B  @    %  �B  @    %  
C  @    eU  ��A  �9  (7�C  ��  9�   a@  :l  b<  ;l  
8  <l  .  =l  �H  >l  �Q  ?l  X  @l  �.  Al  �;  Bl  ))  Cl  eH  Dl  I_  El  �B  Fl   !3  Gl  " �)  IC  �R    FGD  tag  H�   ��   I�  .�  J�  �P   KGD   �  DG   MD  f3    ��D  Tag  ��   Q   ��  .*   ��  �K   ��   gW   ��D  YD  �^    E  k@   l   aE   l  p0   l  �>   l  H   l  �/   �  ��  �4   �F   �D  �<   0dE  H   2l   �/   3�  ��  8�4   qS   :+E  A9  0 U�E  ߣ   Wl   �E   X�  �^   Y�  =Y  Z�E  <   [�  �=   \�E   Jy   ]"  ( E  dE  rY   _qE  �1   ~&F  �.   �l   �L   �l   Z   �3F  �E  �V   �rF  ��   �l   f>   �l  Y   �&F   �)   �9F  �A   /(G     1%   �   2%  �N   38  o=   4%  D4   5%  �^   6%  `*   7%  �0   8%  �G   9%  �D   :%  	I:   ;(G  
 %  8G  @    �@   =F  �\   ��G  +   �8G   Y�   �8G  �
   �8  (   �8  �F   �8  �C   �8   <)   ��G  EG  �,   H  �   l   AK   l  z8   �2  V  H   H  %  �R   �G  	F   .FH  �   0l   �P   1H   ">   3H  % IxH  &�K  KH  &`B  LFH   �[    E�H  �z   G   =Y  NSH   �6   PxH  O]   a!�H  �H  �(  7N  ( �+I  >)  ��4   -N   ��4  V`  ��4  TE   ��  �/   ��   �z   �  $ G   ��H  &8   � EI  KI  eS  p o�M  ��  q�   ^   sMD  ��^   u�  [>   vl   �W   w�D  (�  y�<  0�=   z�=  ��,   |�C  ���   ~  ��(   �>  �AK   �l  0XL   ��E  8'os2  �RA  hp�   ��A  �T   ��4  0#9   ��  8!H  ��O  @�+   ��O  H@.   �	P  P�E   ��O  X�P   ��O  `@   ��O  h$S   �U   ps   �U   x'mm  �U   �'var  �U   �Q   �U   �<B  �rF  �2Y  �
C  �=   ��  �=   ��G  �UV   ��H  ��(   ��  =   ��4   /:   ��  (�?   ��4  0�]   ��  8'cvt  �fP  @�R   ��M  H5$   ��	  P��   ��  `HT   ��  h�*   ��  p�J   �  x�+   �  y�   ��H  ��C   �I  ��-   ��  �j7   ��  �kN   ��  ��F   ��  �#7   ��  ��(   ��4  �rE   ��4  �QZ   ��  �4   ��  ��@   ��  �:L   ��4  ��G   ��4  ��]   ��  ��W   �YP  ��/   ��  ��B    �4   �I   �4  s-   �  �*   �  ,   I  ,   I   'bdf  	+I  (�T   �  P#F   �  X�U   �  `�K   �  h �=   ��M  �M  �  �M  U    �Q   �"�M  �M  �\  x c�O  �   e8I   �   f:Q  )�   g�  �V   h�+  :1   j�   �^  k�  (Jy   m"  0�   nx  8�   p`  <�!   q�  @R0   rx  `�   sx  duN  tx  h6   u  lpp1  v�  ppp2  w�  �2�   zQ  �Xc   {Q  ��6   }"Q  )   ~�4  �8   �   �L  �U   (C   �x  0��   �x  4'pp3  ��  8'pp4  ��  Hy�   ��4  X��  ��4  `U   �6
  h �I   ��O  �O  �  �O  8I  �  "  GD    1   �O  �O  �  �O  �M  �  �  �   �M   +�O  �O  �  	P  �M   �<   :P  P  'P  �M   y*  N    =YP  4   �^  J  b8  �T   lK   H'P  `  |T  @ ?Q  R�   AV   �   Bl  n   C`  
Z�   Dl  �   E`  org  G�  cur  H�  ��   I�   s   K�4  ([   L�2  0c+   Nl  8 R8   PlP  RG   T'/Q  5Q  [  O   _ GQ  MQ  LL  ͳ  @!@�Q  Jy  !B"   �S !C�  ܱ  !D�  .� !E�  ��  !F8  ��  !G�   
�  !H�  (�P  !JGD  0Ӏ !K�4  8 ,�  !MRQ  !
�  !P2R  ߣ  !R�   x  !S�  .� !U�  ē  !V2R  " � !W2R   l  BR  @   � ��  !Y�Q  ��  (!\�R  ߣ  !_�   x  !`�  ē  !b�2  ��  !c�2  Ӷ  !e�   �  !f�  $ r�  !hNR  W�  !m�R  Kw  !t�   7�  !u�4   0�  !w�R  j�  !{S  ��  !}�   �  !~�  �w  !�   J�  !��R  1�  !�FS  �{  !�FS    S  �  !�+S  �   !��S  ��  !��   k  !��S  �q  !�l   q  !��  y|  !��S   �R  LS  �  !�XS  %�  !�!�S  �S  �  �!MV  k  !Ot   Jy  !P"  R�  !QV  ��  !R�  �   !S�   �  !T�  $(  !V8  (|  !W8  )x�  !X8  *п  !Z�  ,�J  !\  0i�  !^�Q  8�  !_�Q  xC�  !`�Q  �= !bBR  ���  !c�R  p�  !e�Q  8��  !f�Q  x=�  !g�Q  ���  !h�Q  ��  !j�  8��  !m�4  @V�  !p�  HV` !q�4  P��  !r�4  X��  !s�  `/�  !u\  h��  !v�  0��  !w\  8j�  !y \  82�  !|b&  Xs  !�2  `��  !��  h�  !�q:  pd�  !��  x|�  !��  �˽  !��	  �ʞ  !��S  �8�  !��:  � ֥  0!��V  ��  !�   �  !�  v�  !��S  �  !��  ݺ  !��  ��  !�H  c�  !��   BV !��V  ( <  �  !�V  !��  H!��X  ��  !��   Ǧ  !��  @�  !��  ��  !��  d> !��  ��  !��  �  !�  I�  !��   U  !��  (�  !��  0��  !�x  8�& !�x  <��  !�	  @?�  !�  `U�  !��  hw�  !��  p֤  !��  �;�  !��  �ܲ  !�\  �w�  !��  ���  !��  ��  !��  ���  !��  �ٛ  !��  ��  !��  �g�  !��  �`�  !��  �x�  !��  ��  !��  �|�  !��  �"��  !��   "�  !��  "n�  !��  "��  !��  "��  !��   "`�  !��  ("�  !��  0"m�  !�l  4"�m  !�l  6"A�  !��  8"��  !��  @ ��  !��V  S�  !�$�X  �X  ��  �!*�Y  Ҳ  !,�X   -�  !-�[  H�  !0�V   ݺ  !1�  P'NDV !2H  X�  !<�4  `K�  !=�4  h�  !>�  p��  !?�  t��  !A�Q  xZ�  !B�4  �l�  !EI  � !E�  �!�R[  ��  !�8   �  !�8  ��  !�8  �  !�8  ��  !�R[  �  !�b[  x��  !�R[  �"�  !�b[  8"��  !��  �"��  !�\  �"��  !�\  �"��  !�\  ��  ! \  �R�  !8  ���  !8  �V�  !r[  ���  !r[   ��  !  �6�  !�  �Ğ  !x  �"�  !	x  ���  !
�  �Т  !�  �P�  !�  �W�  !\  ���  !\  ���  !�  ���  !�X  � \  b[  @    \  r[  @   	 \  �[  @    ��  !�Y  a�   ! \  ߣ  !8   �  !�  �U  !�4  
�  !�  w�  !!�  .�  !"�  �  !#8   �  !%�[  9�  !G�X  �X  *\  @   � 8�  `",R\  �� ".�   -U "/�  X `�  "1^\  *\  !~�  H"<�\  �� ">�   "�� "@  0"��  "A  1"�� "C�  8"�� "D�  @ Z�  "F�\  d\  ��  #?-�\  �\  ۳  `#�l]  ��  #��4   y�  #��  �� #��  �� #��  ��  #�x   Ǩ  #�x  $(2 #��4  (Ϛ  #��4  0R�  #�V  8_� #�^  @ ��   #T�]  �� #W�]   �Y #\�]  add #_�]  �x #e�]   �  �]  �\  x  V   �]  �]  �\   �]  �  �]  �\  x  U   �   �]  r�  #gl]  	^  �  #��\  �  #�"+^  1^  ��  �#��^  y�  #��4   2�  #��4  �� #��4  � #��  R�  #�V   _� #��b  ( ��  #�"�^  �^  ��  #��^  �S #��4   �� #��4  � #��_   ��  #�"�^  	�^  �^  ��  0#�v_  9�  #��   �{  #��`  � #�&`  ��  #��`  x  #��  �  #�8  m�  #��   �  #��  $��  #�  ( (��  N   #��_  ˟   .�  ��  ��  ��  ��   ��  #�v_  ��  #��^  (L�  N   #�&`  ��   ��  Ʊ  ��  ��  g�  �  ��  W�  �  	|�  
K�  ��   8�  #��_  (��  N   #��`  c�   ��  p�  �  �  ��  �  ��  ��  }�  	 ��  #�2`  ��  #��`  �`  �`  `  �   [�  #�^  	�`  �  h#k�a  �� #n�a   �Y #t�a  �? #w�a  �2 #y�a  �! #|�a   �$ #~�a  (�* #�	b  0�3 #�(b  8k! #�Lb  @�A #�bb  HV- #��b  P�F #��b  X  #��b  ` �a  ^  �4  �4  V   �a  �a  ^   �a  �  �a  ^   �a  �  �a  ^  x   �a  �  	b  ^  �4  �  GD     �a  x  (b  ^  x  fP   b  x  Lb  ^  x  H  x   .b  bb  ^  �^   Rb  �b  ^  �^  �  �b   x  hb  �  �b  ^  �^   ,  �  GD   �b  �  #��`  	�b  �  #�1^  ~�  #��b  l�  p#�c  R�  #V   �  #`  )�  #�\  ��  #�+  2�  #>$   �� #>$  (��  #Jd  0��  #Jd  8R0  # �  @�  #!�  H�!  ##O   P��  #$  X�� #%  Yb�  #&  Z��  #(  [�  #)  \_� #+=d  ` ګ  #�d  �� #�&d   �Y #�7d    d   d  U      �b  d  7d   d   ,d  �  #��c  \  î  #B�d  2�  #D�4   �� #E�4  y�  #F�4   {�  #HPd  ��  #L�d  �d  �  �d  8I  �  �4  GD   l�  #R�d  �d  �d  8I  �4  �   ��  �#W
g  <0 #Y�b   4� #[
g  p'top #\H  �O� #^g   Xc  #_*g  ���  #ax  ��  #bx  ��  #c0g  �'cff #e�S  �  #f�X   ˽  #g@g  (
�  #iJd  0�  #j  8��  #kx  <z�  #m�  @�  #n�  D��  #px  H�  #qx  L~�  #s�4  P9� #t�4  XV #v�4  `�  #w�  h&  #yN  l�J #{  p�  #}&�d  x��  #~&�d  �s  #��2  �Ğ  #�x  ���  #��4  �q�  #�9(  ���  #�	  �w�  #��  ��  #�e   ��  #�  ��  #��  � �  g  @   0 �d  *g  @    �d  �  @g  @    �	  x�  #��d  ջ  #�#`g  fg  �  �#qh  R�  #V   �  #`  )�  #�  ��  #�+  2�  #>$   �� #>$  (��  #\  0��  #\  8R0  #�  @�  #�  P�!  #�  `��  # j  ��� #  �b�  #  ���  #   ��  #"U   �L�  ##U   �_� #%�i  � ��  #�~h  �h  �  �h  Sg  x   q�  #��h  �h  �h  Sg  \  \  8   j�  #��h  �h  �  �h  Sg  \  \   ��  #��h  i  �  i  Sg   *�  #��h  �  #�-i  3i  >i  Sg   �  @#��i  �� #��i   �Y #�-i  �? #�$qh  kI #�$�h  rL #�$�h   � #�$�h  (-1 #�$i  0��  #�$ i  8 �i  Sg  `  4  �     �i  T�  #�>i  	�i  a�  N   #� j  ��   J�  �  ,�   ה  #��i  ��  #'fg   �  #Fsj  y�  #H�4   2�  #I�4  �� #J�4   ɠ  #L:j  ݬ  #L�j  :j  �  #O/�j  �j  ��  �#}:l  <0 #-j   4� #�Lm  �'top #�  �O� #�\m  �Xc  #��j  x
s  #��2  �
�  #��  �
V #��4  �
Ğ  #�x  �
��  #�x  �
��  #��4  �
h�  #��4  �
��  #�9(  �
��  #�	  �
w�  #��  �
��  #�x  �
�  #�x  �
�  #�0g  �
�  #�e   `&  #�N  h�  #��l  p_� #�:m  x�  #�  ��  #��  ��J #�  �˽  #��	  � �   #X�l  �� #[�l   �Y #f�l  �; #om  � #u4m   �  #T�l  �l  �  �l  �j  �   �  �l  �j  `  4  �  �4  e     N  �l   �l  �l  �j   �l  �  m  �j  �4  �   �l  �  .m  .m  �4  �   Fg  m  X�  #z:l  	:m  �  \m  @   � sj  lm  @    <�  #� ym  ��  �#�n  R�  #V   �  #8I  )�  #�\  ��  #�+  2�  #>$   �� #>$  (��  #\  0��  #\  8R0  #�  @�  # �  P�!  #"�  `��  #$  ��� #%  �b�  #&  ���  #(  ��  #*U   �L�  #+U   �_� #-�o  � c�  #��n  �n  �  �n  �n  x   lm  ˯  #��n  �n  �n  �n  \  \  8   N�  #��n  �n  �  
o  �n  \  \   Ԝ  #��n  h�  #�$o  *o  5o  �n   8�  #�Bo  Ho  �  Wo  �n   p�  @#��o  �� #��o   �Y #�$o  �? #�%�n  kI #�%�n  rL #�%�n   � #�%5o  (-1 #�%
o  0��  #�%o  8 �o  �n  8I  R\  �\     �o  +�  #�Wo  !�  #EAp  2�  #G�4   �� #H�4  y�  #I�4   ��  #Kp  j�  �#N�q  <0 #Plm   cff #Q�S  �4� #S
g  �'top #TH  hO� #V�q  pXc  #Wr  ��  #Yx  �  #Zx  �  #[0g  
�  #]\  ���  #^\  ���  #`  ��  #a  ���  #bx  ��  #cr  �z�  #e�  ��  #f�  ���  #hx  ��  #ix  �~�  #k�4  �9� #l�4  �V #n�4  ��  #o�  �&  #qN  ��J #s  ��  #u�X  ��  #w&�d  ���  #x&�d  � Ap  r  @    Ap  �  %r  @    1�  #zNp  l�  #kr  �� #��r   >'  #��r  � #�4m   �r  �r  8I  R\  �\    N  �d  �d   %r  kr  �  �r  �r  R\  �   �r  U�  #�2r  	�r  :�  #�#�r  �r  ,�  (#�>s  R�  #�V   Jy  #��s  � #��5  p�  #�t  o�  #�U     4�  #�ws  �� #��s   �Y #��s  gP #��s   �  �s  �r  V  �4  �4   ws  �s  �r   �s  �  �s  �r   �s  \�  #�>s  	�s  ١  #�#�s  �s  ��  x  t  �  �  U    �s  �  #�.t  dt  0�   #�dt  ��  #��-   �0 #��-  ک  #��-  �> #��-   	t  �  X#�u  b�  #!u   �  #!u  E�  #!u  b�  #!$u  ,�  #?u   h�  #Tu  (�  #ou  0��  #�u  8c�  #
t  @:�  #!�u  Hs�  #"�u  P ^  �b  �i  Gm  ?u  �4  �  l   *u  I  Tu  I   Eu  ou  .m  U      Zu  �u  `  �  �X   uu  �s  �r  ��  #�u  it   �$�u  �� $�b   Jy  $ "  ���  $"�4  ���  $#�  �O�  $%  �  $'�u  � $'v  �u  !� @$*�v  �  $,�u   ~�  $.x  ���  $/^  �"�  $2x  "V $3^   "� $4^  �"V�  $5^  � + $7v  , $7�v  v  �`  �v  @    	�v  #2 7�v  	�wH     E N   �v  7  M )	  �	 �v  )O /w  *��   �v  +�  
v   )� �Xw  *��  � �v  *�  � �6   ,� o�  8x  *�  o�6  *��  p�v  *2�  q�4  *�  r�  +�  t
v  +�� u�4  +� vx  -�u  �./cur ��4  0�w  +,j  ��4  .+�2 ��_    ./len ��  ./i �G   .+��  ��^  +F@ ��4       ,�
 8�  �x  *�  8!�6  *��  9!�v  *�F :!�^  +� <�  +װ  =U   +>�  > ,  +:�  ?�  -�u  i 1� P�B     "      ��|  2�  &�6  
  2��  &�v  K C 3�  	
v  � � 3�  
�\    3XL  �\  � � 3V�  �\  � � 3R�  V  p j 3� �  � � 3Q  �u  �	 �	 4cur �4  P
 >
 3�� �4    4n x  d \ 3#�  x  � � 34�  8  i ] 5�0  2z�B     6��B     j       zz  3.� =x  � � 7��B     Az  8U  7��B     Uz  8U  7��B     iz  8U  9��B     8U   6��B     s      :{  4len ��  = / 3� �  � � 77�B     �z  8U| 8T��� 7��B     �z  8U  7��B     �z  8U  7��B     {  8U  9�B     8Uv 8T���8Q��8R~  7v�B     N{  8U  7��B     b{  8U  7 �B     |{  8Uv 8Q}  7!�B     �{  8U| 8Q}  7B�B     �{  8U��8T48Q}  7{�B     �{  8U  7��B     �{  8U  :��B     =�  �{  8Uu  7F�B     |  8U~ 8T0 7p�B     )|  8U~ 8T1 7��B     B|  8U~ 8T2 7��B     [|  8U~ 8T3 7��B     u|  8U| 8Ts  7�B     �|  8Uv 8Ts  7B�B     �|  8U| 8T0 9g�B     8Uv 8T0  1? ��B     �      �>�  2�   �6  G ; 2��   �v  � � 3�  
v  o c 3R�  V  � � 4cur �4  \ H 3�� �4  : 2 ;� �  ��3[>  x  � � 3.� �  x \ 4n �  � � 3� �  � g 3� !�  � � ;U 2�  ��3�
 �4   k 30=   i Q 3%  �v  � p 5�0  ���B     5�u  ���B     <`�  �  3�  B�  t n <��  �~  4tmp h�  � � 7��B     �~  8U�� 9��B     8U��  < �  -  4i �G   � � 4len ��  9 3 <0�  �~  4p ��4  � �  =��B     ,�  8Uw 8T18Q���4$# $ &8Y��  7;�B     C  8U�� :��B     ,�  �  8Uw 8T18Q<8R���4$# $ &8Y�� 7��B     �  8U�� :J�B     ,�  �  8Uw 8T18Q��8R| 8X 8Y�� 9z�B     8U��8T 8Q| 8R��8X1  7�B     �  8Us  70�B     "�  8Us  =��B     8�  8Uw 8T   1� &��B     �      �ԃ  2�  &#�6   � 2��  '#�v  j V 3�  )
v  \ H 4cur *�4  ^ : 3�� +�4  � � 3Q  -�u  t  h  <`�  Ã  3Н  =3  ! �  3.� >x  �! �! 4n >x  >" *" 3I5 ?�\  # # 3R�  @V  �# �# ;� A�  ��3�  B  $ $ <��  ��  3^�  r�   j$ h$ 9i�B     8U} 8Ts8Q	�1H     8R8  <��  ^�  3�j �x  �$ �$ 6S�B     e       9�  4len ��  �$ �$ 7a�B     �  8U~  9��B     8U��8T| 8Q} 8Rv  7��B     M�  8U~  9��B     8U~   7�B     r�  8U~  79�B     ��  8U~  :_�B     8�  ��  8Uw  :z�B     8�  ��  8Uw  7��B     ΂  8U�� :��B     ,�  �  8Uw 8T28Q08R��8X08Y�� :��B     ,�  <�  8Uw 8T88Q08R��8X08Y�� 7%�B     ^�  8U~�8T| 8Qw  7y�B     r�  8U~  7��B     ��  8U~  7)�B     ��  8U~  7�B     ��  8U~  =��B     =�  8Uu   9��B     8U~   >� ���B           �'�  ?�  �&�6  A% 5% ?��  �&�v  �% �% @�  �
v  R& H& @:  �'�  �& �& @x  ��  y' m' #/� �-�  ��@��  ��  ( ( @E  �x  W( S( 7��B     ��  8Uv 8T68Qw 8R0 :��B     D�  ʄ  8Tv  :��B     D�  �  8Tv  :��B     D�  ��  8Tv  :��B     D�  �  8Tv  =��B     D�  8Tv   	  �  =�  @    A/ �G   Y�  Bc �8   Ce	 ��  D�  � 
v  ER�  �V   A� ��  �  D�  �#
v  DJy  �#"  DR�  �#V  DQ  �#�u  E� ��  E�  ��  F�u  � ,� ~�  i�  *)�  ~%�  *�  %4  *�^ �%�  *:1  �%<  +� ��  +	 �37  +[ ��6  +!	 ��6  +� �=   )o e��  * e&�   17
 [��B            �܆  2	 [%�  �( �( 3 ]37  �( �( G��B     Q�   H0 B�  ��B     Q       ���  2	 B%�  ) ) 3 D37  v) n) 3�  E`  �) �) 3!	 F�6  +* %* ;�q  G�  �h3� H�  {* u* =��B     ^�  8T�h  )� 0݇  *[ 04  +�  2�6  +�  3`  +!	 4�6  +D� 5�	   H� �  ��B     _       ���  2[ 4  �* �* 2-U �  + + 3�  �6  p+ j+ 3�   �6  �+ �+ 3� !�  �+ �+ I��B     k�  =��B     w�  8T|   H^ 	�   �B     _       �9�  2[ 	&4  , , Jreq 
&  ^, X, 3�  �6  �, �, 3�  �6  �, �, 3� �  #- !- I6�B     k�  =E�B     ��  8T|   H7 ��  ��B     6       ���  2�  �4  L- F- 3[ ��6  �- �- 3�  �`  �- �- 3!	 ��6  . . ;�k  �4  �X3� ��  <. 6. :�B     ��  �  8T�X I�B     k�   1� ���B            �*�  K~ �6  U H� ��  �B     /       ���  2~ �6  �. �. 3K1 �m7  / / 3� �6  �/ �/ ="�B     ��  8T	�.H       1? �0�B     �      ���  2!	 �`  �/ �/ 3�  ��6  ,0 $0 3�6  ��4  �0 �0 3��  ��  �0 �0 3R�  �V  C1 A1 IZ�B     ��  :i�B     8�  U�  8Uv  :��B     8�  m�  8Uv  :��B     8�  ��  8Uv  :��B     8�  ��  8Uv  :��B     8�  ��  8Uv  :��B     8�  ͋  8Uv  :�B     8�  �  8Uv  :�B     8�  ��  8Uv  :9�B     8�  �  8Uv  :S�B     8�  -�  8Uv  :m�B     8�  E�  8Uv  :��B     8�  ]�  8Uv  :��B     8�  u�  8Uv  :��B     8�  ��  8Uv  =��B     8�  8Uv   L� ��  �C     �      �-�  ?Jy  �!"  j1 f1 ?!	 �!`  �1 �1 ?�  �!x  3 {3 ?G  �!x  �3 �3 ?G  �!V  �3 �3 @�  ��6  W4 /4 @� ��  6 6 @s  ��2  7 7 @Q  ��u  W7 =7 @�� �`  �8 j8 @�6  ��4  j: B: @��  ��  �< b< 5�u  �	C     <��  �  @~ �6  �> �> @�O  ��  �> �> =�C     ��  8T	�BH     8Q1  <0�  I�  @s�  ��   �> �> @r? ��   �? �?  <p�  ��  ;��  !\  ��{:�C     ��  ��  8T	�.H      =5C     Ĝ  8Tv 8Q08Rs�  <��  (�  ;�� W  ��{3f�  X
t  �? �? 3�M Y�-  #@ @ :3C     ќ  	�  8T08Qv 8R0 =�C     ќ  8T08Qv 8R0  M-�  C      ��  � �  N>�  �@ �@ O��  PJ�  ��{QV�  �B zB Qb�  CC C Qn�  /E %E Pz�  ��zQ��  �E �E R��  PC     M/w  0C      p�  +܏  NJw  �F �F N=w  hH dH  Mw  PC      ��  �Đ  Nw  �H �H O��  Q!w  �H �H SY�  �C      ��  r�  Nf�  I I O��  Qr�  PI LI 7�C     c�  8Uv  IuC     8�    7fC     ��  8Uv� 7|C     ��  8Uv� 7�C     ��  8Uv� 9�C     8Uv�   M�  �C      �  8D�  N��  �I �I N��  �J xJ N��  �J �J N��  ]K UK O�  P��  ��zQ̅  �K �K R؅  �C     7�C     ^�  8Uv 8T08Q08R~  :/C     ޜ  {�  8U 8T0 :C     �  ��  8U 8TA :QC     ��  ��  8U  :lC     ޜ  ͑  8U 8T0 :�C     �  �  8U~ 8T| 8Q��z :�C     �  �  8U 8Q|  :0	C     8�  (�  8U~  =C     �  8U 8T|    MXw  �C      ��  ?^�  N�w  �K �K N�w  L L Nww  SL AL Njw  M M O��  Q�w  �M �M Q�w  �N �N Q�w  �N �N R�w  r
C     T�w  ��  L�  Q�w  9O #O T�w  P�  f�  Q�w  ,P "P Tx  ��  U�  Qx  �P �P Ux  ��  Qx  Q �P Q&x  �R �R S8x  C      0�  �$�  Ndx  �S �S NWx  �T �T NJx  }U wU O0�  Qqx  �U �U P~x  ��zQ�x  %V V Q�x  �V �V R�x  �C     7�C     ��  8Uv 8Ts  $ &34$�wH     "8Q��z8R08X0 9hC     8U��z8Tv    :�
C     +�  1�  8U}  =	C     7�  8U��z8T} 8Q    9fC     8Uv   V�w  �	C     �       '�  Q�w  �V �V V�w  $
C     4       ڔ  P�w  ��z7.
C       8Uv  9@
C     8Uv 8T��z  7�	C     �  8Uv  7�	C     �  8Uv  7�	C     �  8Uv  9�	C     8Uv   7�C     ;�  8Uv  9�C     8Uv   9C     8Uv    T��  ��  ޕ  Q��  $W W Q��  �W �W Q��  SX KX Q��  �X �X Q˖  :Y 4Y Uז  ��  Qؖ  �Y �Y =C     B�  8U| 8Ts    =;C     �  8U~ 8T<8Q��z   :�C     N�  �  8T	�BH      IPC     [�   A/  �  �  D�   �6  E��  "�v  E�  #
v  E�6  $�4  ER�  %V  E� &�  EQ  (�u  F�u  �.E�j ex  Widx ex  E��  e x  Eb�  e*x  Ela f�4  .E�  u�4     X �[  ��B     
       �T�  ?~ �(6  �Y �Y ?p �(T  (Z $Z Y��B     g�  8U	 |H     8T�T  X7 ��  ��B     �       ���  Z�  �,`  UZۮ  �,�:  T X| �x  ��B            �ė  Z�  �$`  U X� ��  ��B            ��  Z�  �,`  UZ��  �,�:  T X�	 }�  ��B     1       �B�  Z�  }*`  UZù  ~*q:  T X2 j�  ��B            �s�  Z�  j#�6  U X� H�  @�B     �       ��  ?�  H#�6  mZ aZ ?la I#�  [ �Z [i Kx  �[ �[ O �  @��  P�  �[ �[ :��B     B�   �  8U}  =��B     t�  8T08Q:   X <�   �B     %       ���  ?�  <#�6  �[ �[ ?�^ =#�  +\ '\ ?B� >#�  j\ d\ ?(5  ?#�  �\ �\ =�B     ��  8U�Q8Q	�R����  \=�  0�B            ���  ]N�  U^=�  0�B            NN�  
] ]   \�  0�B           �h�  N�  3] -] N �  �] ] N�  �] �] N�  )^ #^ Q'�  w^ u^ Q4�  �^ �^ QA�  �^ �^ QN�  @_ >_ Q[�  f_ d_ Si�  |�B      0�  �  Nw�  �_ �_ =��B     ��  8Us   V�  H C     �       3�  N �  �_ �_ _�  N�  �_ �_ N�  �_ �_ `H C     �       a'�  a4�  aA�  aN�  a[�    :r�B     t�  O�  8T08Q: 9@ C     8Q 8R| 8!  \��  PC     6       �,�  N��  #` ` Q��  u` o` Q��  �` �` Q  �` �` Qχ  a a V��  sC            �  N��  4a 2a `sC            a��  a��  a  aχ  I|C     [�    InC     ��   b�6  �6  %�bF\  F\  %�c5<  5<  
?c�M  �M  �c�D  �D  �bBX  BX  &�c�@  �@  
�	c�Z  �Z  
s
bU/  U/  &dc�R  �R  cA*  A*  
�	cKM  KM  Yc�?  �?  
<	c�3  �3  1c9  9  'cc�3  �3  '�cxL  xL  '�b�K  �K  %vcE1  E1  'rc _   _  'hb�O  �O  (2d�  �  + bBi  Bi  (c!,  !,  Ub�\  �\  &yc�*  �*  [b�\  �\  ).cq]  q]  %zc{X  {X  �b�]  �]  *^ E   �;  �  � $"  �C     a      �� X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �[  �<  �  >   G   �	  	N   �  B"i  o     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  ]  -      n�  �  �  ]  U    �  �    U   )  ]  -   -   U    �  �"5  ;  �   PJ�  2�  L8   �  M@   pos N@   �  P�  SF  Q�   �1 R  (=9 SE  0R�  U]  8y�  V8  @�� W8  H �  ��  �\ �-   m  �U    o  ��  �  �    @   8  )  @   8  @    >  �  2  R  X  c  )     :-   �  J�  x Lc   y Mc   )  Oo  	�  B   s�  M   uc   }  uc  V  vc  /  vc   t
  x�  �J  N   �;  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  N    ��  N   �  	G   B� 
8  L  <    >  s  >  v	  U     �  ;  	�  �  (N/  �  P)   Z�  Q)  �  S/  s  T�   [  U5  ?1  WG     �  )    Y�  �  =  N   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  �N  b   "�  �  �  %  <�  x >)   len ?<  *� @>   %  B�  	�    `    '  G   G   '  U    �  �  q:  @  G   Y  G   G   U    �  f  l  �  G   G   U    �  `�  �  �   �% �  ?1  �G   �&  ��  !  ��   I  �-  ()  �Y  0R   �U   8�  ��  @ �    �  ��  	  �   :  @  G   T  U   T   �  �  g  m  x  �   �  ?�  �  �  �  8  @    �  Y�  �  G   �  �  @   U    s  ��  �  G   �  �  �   (  W  0�\  �  ��   e� �-  �� �x  �� ��  �� ��   �� �Z  ( �'  ��  �!  l>  �  ��  �  -  �>  	�  �  �  ��   	�  �
  �)  �  �<  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   �0  D4   b   �o	  xx ��   xy ��  yx ��  yy ��   a  �,	  	o	  z'  ��	  m  ��   ss  ��   �  ��	    ��	  �	  �	  U    �  �
  �U  �U      ��	   %  ��	  �  $
  "
  �   [
  �� "
   �@ #
  �U  $U    �  7�
  �; 9
   ��  :
   L  <[
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=U  ��  ?c   �  @c  ~  Bc  �  Cc  �  Dc   5  Fc  (B  Gc  0�  Hc  8 �	  J�  
   s�  �  u�   ��  v�  �  xc  �
  zc  (  {c   �  }b  �  �#�  �  k  `	��  R�  	�]   (  	��  |  	��  �  	��  �  	��  �  	�c&  v  	��
  �  	�,  (�%  	��  07&  	�s&  8G   	��  X �  �"�  �  h  	�  �M 	J&   k  	�  R�  	]   �  �"�  �  %  8	;,  �� 	=P&   �M 	>�!    	?�
   r$  	@�  0 5  �$9  ?  %  �	�  �� 	P&   �M 	]&  �  	�   �  	=  (�� 	
�  h�� 	�  p�� 	�  x K  � �  �  �  �,�  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6  (A  7  0T  9�  8  :  @�  <�  H�  =  PE-  ?
  X�!  D�  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R�  ��� S;  �K1 W�  �R�  X]  �Jy  Y)  �%  [�
  ��	  ]
  �    ^U   ��8  `t  � L   �  �    X��  �  ��   E-  �
  N ��  �8  �%  P �  *%�  �  �  0t;  k  v�   �  w�  �@ x�  ݖ y�  E-  z
   N |U  0�  }�  pR  ~�  x�  �  �ߣ  ��  ��I ��  ��  ��  �h  ��  ��S  �;  �4  ��  �8  ��  �  �U    �  �-   �  �c  o  �c  �L �U    �8  �_  ( �
  L#H  N  W  H�  �  J�   = KZ    L�  d  M�   �  N   �Z  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  (0  ON  #   g)�  �  �   �	�  =  	�o	   L  	��   $  	��  0�  	�p"  8m  	�#�#  h�  	�u  pآ  	�C  tG   	��  x �  �  ;  �?  d�  �
  �)2  8  �   H	�q  �  	�U    "  	��  �!  	��   ~	  8f�  �
  h�   (  i�  �� k�  �� l�    nc  �  oc   �  pc  (�  qc  0 y  sq    �$
    �  0
'_  �N  
)�   ?1  
*�  }0  
+�  i/  
,�  � 
-o	   �  �)l  r     H	��  ��  	��   ?1  	��  (  	�i  4  	�o	  \  	��  0  	�U   @ +!     tag �   �U  	   �  �     `  N   
K  w%   }#  �&  h  �  &     
  E   9
�  � ;
K   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  X  �  N   ��  :   �   ^$  1  �!  �!   :  ��  � ���  ��  ��   �]  ��  @�  ��  j ��  L� ��  N� ��  P� ��  R�0 ��  Te ��  V� ��  X� ��  Z ��  [\ ��  \��  ��  ^��  ��  `�<  ��  b�X  ��  d� ��  f( ��  h�N  ��  j� ��  l ��  m� ��  n� ��  o� ��  p� ��  x ��  �� ��  � ��  �ݖ ��  �?1  ��  �� ��  �� ��  �� ��  �� ��  �M ��  � �  �  @   ; �    @    � �  � �)    �  �	  �#  �=  C  	  R  �   I$  �^  d  o  �   �&  �{  �  %  �  �  �   �   �!  H�  �  ��   S"  ��     �  �"  ��  �  ��   ;  �  (%  �1  0�   �R  8��  �o  @ �  R  ��  x  =�	  H  E#N  	=  �  @J�  �  L�   �  M�  �� O  .� PD  �  Q�   �  Ra  (�!  S�  08'  T�  8   W!�  �  -  (l  k  n�   �M o  ߣ  p�  �  q�   I  k  )*  0  	  D  �  �   w   .P  V  a  �   �  1m  s  �  �  �  H   |	  K  6�  �  �  �  �   �  �  :�  �  	  �  �  �   �  >*  "  Y�  �  	    ,  �  �  H   �  _$  *  	  H  ,  �  �  H   $  fT  Z  o  ,  �  �   �  l{  �  	  �  ,  �  	   #  x�  �� � $   �  � �  H  � �  P�  �   X9!  � H  `l� � o  h  �   p \    ��  �  H
2d  �S  
4;   �  
5/  (  
6/  04  
7�  88  
8�  @ �  
:  �  �
=�  R�  
?]   �  
@�  n  
A�  �  
B�  1$  
Ci  2�  
Ed  �� 
Fd  `�L 
HU   � �  
J�  p  P     
  	  -  )  �  �  �     �  &9  ?  J  �   �%  *V  \  	  k  �   �%  -w  }  �  �   {  1�  �  	  �  �   �  4�  �  �  �   l  8�  �  	  �  �  �   �  <�  �  	     �  �   �  @   $   	  B   �  �  �  C   �  GN   T   	  r   �  �  �  /   �'  N~   �   	  �   �  )   �  S�   �   	  �   �  �  �  C  �    �  &  ���!  �� �$   i'  ��  H   ��  P  ��  X�A ��  `Y �-  h�#  �J  p�  �k  x�  ��  �  ��  ���  �   �U�  �B   ��!  �r   ���  ��   ��  ��  �&  ��  �   ��   	�!  �&  ��!  �   �>  ��!  'O  ��   xC  �   s/  ��!  	�!  �  0tp"  �  v	   a   w	  �'  x	  !  y	  �#  z	   �  {	  ( �  }"  �  U'�"  �"  m  D   t�"  �  v�   A  w�  �  x�  &  y�   !  {�"  �  ��"  �"  	  #  }"  �  #   �	  �  �#  %#  5#  }"  #   �'  �A#  G#  	  e#  }"  �  i  e#   �"  �!  �#  ��  )�"   ��  )#  �  )5#   }  k#  	�#  O  ;�#  _� =%�#   ݰ  >%}"   �#  �  @�#  �#  cA  	�,$  $  /  	�4$  �� 	�g   �M 	�4$   ?<  	�,E$  	4$  �$  �5  P	��$  �  	��   �� 	��$  �Y 	�%  �H 	�/%  U@ 	�U%   �9 	�#�%  (�A  	�#�%  0�^  	�#�%  8�^  	�#&  @N7  	�#-&  H 	K$  ��  	�$  (Z  	��$  �$  	  %  �#  	   17  	�%  $%  /%  �#   �G  	�;%  A%  �  U%  �#  P   %G  	�a%  g%  �  {%  �#  {%   P  �@  	��%  �%  �  �%  �#  �#  P  P   �;  	��%  �%  i  �%  �#  P  P   �W  	��%  �%  {%  &  �#  ]   *;  	�&  &  {%  -&  �#  ]  P   �T  	�&  g�  	�K$  	9&  $  �  	�  	  �  s&  @    0  �&  @     �  	�%\  �(  N   9'  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  VD'  �\ X�   �  Y�  x  Z�   �7  \'  	D'  < #}'  �  %�   � '�   � )U'  � ,�'  �  .�   � 0�  � 1�   ' 3�'  1  63(  �  8�   � 9�  q :�  
v <�   >�  � @�  y A�   � D�'  �  G�(  F@ I�(    K�  ` L�  9 M�   �  �(  @    � P?(  < S�(  � U�   i V�  t W�   X�   Y�   Z�    \�(  M _-)  F@ a�   x  b�   � d)  E  g{)  � i�   �  j�  � k�  ݖ l�   N n9)  � ���)  x  ��   � �  2 ��)  �W ��  �d> �  � �  � ��)  �)  !] �3*  �� �   v�  ��)  �"� �;   "�� �g   � �?*  �)  
1  �.�!  N   ��,  �>  �B YS <S tX �X A: h; B dD 	�J 
�A %V 0L �F M �H �> �T �Z R �;  _9 !�E "�O #�P $p: %< &(N '�R (;U 0	X 1Q @W AQW Q�C R�D S�= TML U�B VG W�X X(P `FF abT b�E c�T pAM �O ��> �? ��L ��N ��: �ZP �XG �V= �bM ��M �H; �3O ��H �4H �3K ��S �HD ��U ��> ��Z �d[ ��T ��[ �{T ��Y ��< ��Q ��Z �gR �FA ��J �oV �/> ��V �=R ��P �xH ��? ��= ��G �?Y �3; ��? ��A ��R � D  �,  �,  	  �,  �  �,     V $�,  	�,  S $�,  � &�,    P'  �,  @    	�,  #0 + �,  	�H     P'  '-  @    	-  # 7 '-  	�H     P'  R-  @    	B-  #y D R-  	`H     P'  }-  @    	m-  # X }-  	@H     #� g }-  	 H     P'  �-  @    	�-  #� v �-  	 H     #6 � '-  	�~H     P'  �-  @   % 	�-  # � �-  	@~H        [S.  
H ]�$   N� ^P  .� _P    a`.  .  $� �"E&  	�}H     %* �@$  $� i&�,  	�}H     "  �.  @    	�.  $� s#�.  	�}H     &E*  �	�|H     '� |%  �C     
       �P/  (~ |)�  [a Wa (�1  })  �a �a )�C     0D  *U	�}H     *T�T  '� ]	  �C     �       ��/  +�  ],�  U+� ^,�,  T,v�  `�)  �a �a  '� �	  �C     i      ��1  ( �!�  b �a (�  �!�  xb tb (�^ �!�  �b �b (:1  �!C  c c ,�  �3*  �c �c ,v�  ��)  .d (d ,� �	  yd wd -p ��)  �d �d -len ��  ke ge ,�I ��1  �e �e ,x  ��  8f .f ,K �i  �f �f .�u  WC     /��  �1  ,R�  5]  g g ,�  6�  Tg Ng ,D 7�)  �g �g ,x� 8�)  �g �g 0�C     1       ]1  ,�� M�)   h �g  1�C     =D  *T~ ����*Q0*X0*Y�L  1C     ID  *Uv0  �  2� �	  2  3�  �&�  4req �&�  %�  �3*  %� �  %�� �  %� �	  %�  ��   '� �	  �C     L       ��2  (�  ��  )h #h (-U ��  yh uh ,�  �3*  �h �h ,� �  �h �h 1�C     VD  *T0  'k �	  @C     k      �4=  (Jy  �!)  i �h (� �!�  ni fi (� �!�  �i �i (G  �!�  �k �k (G  �!  �k �k ,�  �3*  l  l $� �	  ��,R�  �]  l gl ,�  ��  �m {m .�u  ��C     .�0  �kC     0C     �       �3  ,v�  ��)  Yn Wn 5-C     cD  �3  *U} *T�*Q�� 1hC     a@  *Tw   /��  �5  ,�� �  �n |n ,v�  �)  �n �n ,� �  Jo Do /��  �4  ,��   �o �o $�  �  \,  !�  �o �o 5�C     oD  �4  *T~ *QH 5�C     oD  �4  *T| *QH 1AC     oD  *TH*Q~   0�C     S       35  $�� Hg  ��1$C     |D  *U	�}H     *T0*Q��*R0  54C     =D  h5  *U} *T *Q0*R1*X0*Y��} 5jC     cD  �5  *U} *Tv*Q~  5�C     �D  �5  *Qv  5�C     �D  �5  *U|  1�C     =D  *U} *T1*Qv *X| *Y~   6�>  �C      p�  ��<  7�>  p �o 8�>  9p�  :�>  ��};�>  �q �q ;�>  �r �r :?  ��};?  �s �s <!?  �C     <*?  	C     <3?  ;C     =<?   �  <<  :=?  ��}=J?  ��  n8  ;O?  �t �t ;\?  �t �t ;i?  su iu ;v?  �u �u =�?  ��  27  ;�?  Gv =v ;�?  �v �v >�C     �D  5�C     �D  7  *U|  1C     �D  *U|   56C     �D  J7  *U|  5YC     �D  b7  *U|  5mC     �D  z7  *U|  5�C     �D  �7  *U|  5"C     �D  �7  *U|  5sC     cD  �7  *U} *T�*Q��} 5�C     �D  �7  *U| *T	~ <��}" 5�C     �D  8  *U| *T< 5�C     �D  )8  *U|  5�C     �D  A8  *U|  5C     �D  Y8  *U|  1C     a@  *T|   =�?  0�  �;  :�?  ��~:�?  ��:�?  ��~:�?  ��~:�?  ��~:�?  ��}:�?  ��}:�?  ��}:	@  ��;@  �v �v ;#@  yw qw ;0@  �w �w ;=@  Yx Ex ;H@  9y 3y ;S@  �y �y 5�C     �D  29  *U|  5C     �D  ^9  *U| *T	`H     *Q��~ 5�C     �D  �9  *U| *T	@H     *Q��} 5@C     �D  �9  *U|  5^C     �D  �9  *U| *T	 H     *Q��~ 5�C     �D  :  *U| *T��}�
��3$ $ &��}"# 5�C     �D  /:  *U| *T	 H     *Q��} 5%C     �D  O:  *U| *T��} 5FC     �D  {:  *U| *T	 H     *Q��~ 5�C     �D  �:  *U| *T} 
��3$ $ &��}"# 5�C     �D  �:  *U| *T	 H     *Q��} 5�C     �D  �:  *U| *Ts  5C     �D  ";  *U| *T	 H     *Q��~ 5TC     �D  O;  *U| *Tv 
��3$ $ &s " 5rC     �D  {;  *U| *T	 H     *Q��} 5�C     �D  �;  *U|  5�C     �D  �;  *U| *T	�~H     *Q�� 5IC     cD  �;  *U��}*T�*Q��} 1�C     a@  *T|   5�C     �D  <  *U|  1�C     �D  *U| *T	�H     *Q��}  5�C     �D  Y<  *U| *T0 5�C     �D  �<  *U| *T	�H     *Q��} 1�C     �@  *U    ?4=  kC      �  �7B=  �y �y 9�  ;O=  �y �y @\=  A4=  �  7B=  z z 9�  @O=  ;\=  Bz @z 5zC     �@  =  *U  1�C     �D  *Us       Bm �j=  3� ��  %�  �3*  %R�  �]   'g �P  �C     /       ��=  +
H �#S.  U+��  �#{%  T,n�  ��  mz ez ,E  �P  �z �z ,��  �P  P{ F{  '� v�  �C            �H>  +
H v#S.  U(��  w#P  �{ �{ ,n�  y�  | |  '7 e	  �C             ��>  +
H eS.  U+m  f	  T,�  h3*  *| (| ,v�  i�)  R| N|  2� 	  a@  3�  $3*  3� $�  %� 	  %Jy  )  %R�  ]  % }'  %�  �  C�u  VC�0  RCz �D%{ &�'  E�?  %� 3�  %� 5�  %\�  6�  %w�  7�  D%� T�  %.� T�    D%� �!3(  %� �!�(  %d �!�(  %� �+�(  % �5�(  %� �!-)  %& �--)  %1 �9-)  %� �!{)  %� ��  % �%�  %� �6�  Fi ��  Fj ��  Fk ��     G� �	  �@  Hv�  ��)  HJy  �)  I� �	  I� �  IK �i  I�  ��  .�u  	C      J� �PC     l       ��A  K�  �3*  �| �| LR�  �]  �| �| LJy  �)  } } Lv�  ��)  1} -} 5�C     �D  SA  *Tv� 5�C     �D  kA  *U|  1�C     �D  *U| *Tv   M�1  �C     �       �kB  7�1  n} h} 7�1  �} �} ;�1  ~ ~ ;�1  J~ F~ ;�1  �~ �~ N�1  ;2  �~ �~ O�1  @C            7�1  4 0 7�1  q m P@C            @�1  @�1  @�1  @�1  @2  )GC     2  *U�U*T0    Ma@  pC     �       ��C  7r@  � � 7~@  ~� n� ;�@  5� /� ;�@  �� ~� ;�@  T� P� ;�@  �� �� =a@  0�  ZC  7~@  � ܂ 7r@  4� .� 90�  ;�@  �� �� @�@  @�@  @�@  Q�@  5�C     �D  9C  *Uv  )C     E  *U�T*Q�U#�   5�C     �D  rC  *Uv  1�C     �D  *Uv *T	@~H     *Qs  M4=  �C     A       �0D  7B=  �� �� ;O=  � � @\=  A4=  @�  7B=  |� v� 9@�  @O=  ;\=  ʄ Ȅ 5�C     �@  D  *Us  1�C     �D  *Uv     R�*  �*  [S�6  �6  �R�D  �D  	�RP  P  	�S�K  �K  vRjO  jO  R�3  �3  	1T�D  �D   S�O  �O  2R�N  �N  �RF  F  mR9  9  cR�3  �3  �RxL  xL  �R�N  �N  �SF\  F\  �R�J  �J  �R�*  �*  � ]   ~@  �  F $"    C     U$      �� X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �	  	N   �  B"]  c     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  Q  -      n�  �  �  Q  U    �  ��  �  U     Q  -   -   U    �  �")  /  �   PJ�  2�  L,   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S9  0R�  UQ  8y�  V,  @�� W,  H �  ��  �\ �-   m  �U    o  ��  �  �    @   ,    @   ,  @    2  �  2  F  L  W     .|  Y/    :-   �  J�  x Ld   y Md   )  Op  	�  B   s�  M   ud   }  ud  V  vd  /  vd   t
  x�  �J  N   �<  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  N    ��  N   �  	G   B� 
,  L  0    2  s  2  v	  U     �  <  	�  �  (N0  �  P)   Z�  Q)  �  S0  s  T�   [  U6  ?1  WG     �  )    Y�  �  =  N   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  �O  b   "�  �  �  %  <�  x >)   len ?0  *� @2   %  B�  	�    `    (  G   G   (  U    �  �  q;  A  G   Z  G   G   U    �  g  m  �  G   G   U    �  `�  �  �   �% �  ?1  �G   �&  ��  !  ��   I  �.  ()  �Z  0R   �U   8�  ��  @ �    �  ��  	  �   ;  A  G   U  U   U   �  �  h  n  y  �   �  ?�  �  �  �  ,  @    �  Y�  �  G   �  �  @   U    s  ��  �  G   �  �  �   )  W  0�]  �  ��   e� �.  �� �y  �� ��  �� ��   �� �[  ( �'  ��  �!  	l2  �  	��  �  -  	�2  	�  �  �  	��   	�  �
  	�)  �  	�0  �  	�G   
  	�N   �  	�-   \#  	�@   �  	 -   �  	,G   \&  	7U   �0  	D4   b   	�p	  xx 	��   xy 	��  yx 	��  yy 	��   a  	�-	  	p	  z'  	��	  m  	��   ss  	��   �  	��	    	��	  �	  �	  U    �  	�
  �U  	�U      	��	   %  	��	  �  	$
  #
  �  	 \
  �� 	"
   �@ 	#
  �U  	$U    �  	7�
  �; 	9
   ��  	:
   L  	<\
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @
=V  ��  
?d   �  
@d  ~  
Bd  �  
Cd  �  
Dd   5  
Fd  (B  
Gd  0�  
Hd  8 �	  
J�  
   
s�  �  
u�   ��  
v�  �  
xd  �
  
zd  (  
{d   �  
}c  �  
�#�  �  k  `��  R�  �Q   (  ��  |  ��  �  ��  �  ��  �  �?$  v  ��
  �  �-  (�%  ��  07&  �O$  8G   ��  X �  
�"�  �  h  �  �M &$   k  �  R�  Q   �  
�"�  �  %  8;-  �� =,$   �M >�    ?�
   r$  @�  0 5  
�$:  @  %  ��  �� ,$   �M 9$  �  �   �    (�� 
�  h�� �  p�� �  x K  
� �  �  �  �
,�  �   
.�   �  
/�  O  
1�  C  
2�  �  
4�   d> 
6  (A  
7  0T  
9�  8  
:  @�  
<�  H�  
=  PE-  
?
  X�!  
D�  h:  
F�  �  
G�  ��  
H�  ��  
I�  ��  
K�  �  
L�  �U  
N�  ��  
O�  �)�  
Q�  ��  
R�  ��� 
S<  �K1 
W�  �R�  
XQ  �Jy  
Y  �%  
[�
  ��	  
]
  �    
^U   ��8  
`u  � L  
 �  �    X
��  �  
��   E-  
�
  N 
��  �8  
�&  P �  
*%�  �  �  0
t<  k  
v�   �  
w�  �@ 
x�  ݖ 
y�  E-  
z
   N 
|V  0�  
}�  pR  
~�  x�  
�  �ߣ  
��  ��I 
��  ��  
��  �h  
��  ��S  
�<  �4  
��  �8  
��  �  
�U    �  
�-   �  
�d  o  
�d  �L 
�U    �8  
�`  ( �
  
L#I  O  W  
H�  �  
J�   = 
K[    
L�  d  
M�   �  N   
�[  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  
�  (0  
OO  #   
g)�  �  �   ��  =  �p	   L  ��   $  ��  0�  �Q   8m  �#�!  h�  �v  pآ  �7  tG   ��  x �  �  <  �?  
d�  �
  
�)3  9  �   H�r  �  �U    "  ��  �!  ��   ~	  8
f�  �
  
h�   (  
i�  �� 
k�  �� 
l�    
nd  �  
od   �  
pd  (�  
qd  0 y  
sr    
�$    �  0'`  �N  )�   ?1  *�  }0  +�  i/  ,�  � -p	   �  
�)m  s     H��  ��  ��   ?1  ��  (  �j  4  �p	  \  ��  0  �U   @ +!  
  tag 
�   �U  
	   �  
�    `  N   

L  w%   }#  �&  h  �  &     

  E   
9
�  � 
;
L   ��  
<
�  �  
=
�  �  
>
�  �#  
?
�   �  
L
(�  Y  �  N   
��  :   �   ^$  1  �!  �!   :  
��  �  �	  �#  �  $  	  3  �   I$  �?  E  P  �   �&  �\  b    v  �  v   �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  �  (%  �  0�   �3  8��  �P  @ �  R  �|  x  =�	  H  E#/  	  �  @J�  �  L�   �  M�  �� O�  .� P%  �  Q�   �  RB  (�!  So  08'  T�  8   W!�  �  -  (l�  k  n�   �M o�  ߣ  p�  �  q�   *  k  )    	  %  �  �   w   .1  7  B  �   �  1N  T  i  �  i  I   }	  K  6{  �  �  �  �   �  �  :�  �  	  �  �  �   �  >  "  Y�  �  	  �  -  �  �  I   �  _    	  )  -  �  i  I   $  f5  ;  P  -  �  �   �  l\  b  	  {  -  �  	   #  x��  �� �    �  � �  H  � �  P�  � �  X9!  � )  `l� � P  h  � �  p ]    �{  �  H2E  �S  4<   �  50  (  60  04  7�  88  8�  @ �  :�  �  �=�  R�  ?Q   �  @�  n  A�  �  B�  1$  Cj  2�  EE  �� FE  `�L HU   � �  J�  Q  P   �  �  	      �  �  �     �  &     +  �   �%  *7  =  	  L  �   �%  -X  ^  i  �   {  1u  {  	  �  �   �  4�  �  �  �   l  8�  �  	  �  �  �   �  <�  �  	  �  �  �   �  @�    	  #  �  �  �  7   �  G/  5  	  S  �  �  �  0   �'  N_  e  	  y  �     �  S�  �  	  �  �  �  �  7  �   �  &  ���  �� �   i'  ��  H   ��  P  ��  X�A ��  `Y �  h�#  �+  p�  �L  x�  �i  �  ��  ���  ��  �U�  �#  ��!  �S  ���  �y  ��  ��  �&  ��  �   ��  	�  �&  ��  �  �>  ��  'O  �v   xC  �   s/  ��  	�  �  0tQ   �  v	   a   w	  �'  x	  !  y	  �#  z	   �  {	  ( �  }�  �  U'j   p   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {u   �  ��   �   	  �   ^   �  �    �	  �  � !  !  !  ^   �    �'  �"!  (!  	  F!  ^   �  j  F!   �   �!  �!  ��  )�    ��  )�   �  )!   }  L!  	�!  O  ;�!  _� =%�!   ݰ  >%^    �!  �  @�!  �!  cA  �,�!  �!  /  �"  �� �h   �M �"   ?<  �,!"  �"  �5  P��"  �  ��   �� ��"  �Y ��"  �H �#  U@ �1#   �9 �#]#  (�A  �#�#  0�^  �#�#  8�^  �#�#  @N7  �#	$  H 	'"  ��  ��!  (Z  ��"  �"  	  �"  �!  	   17  ��"   #  #  �!   �G  �#  #  �  1#  �!  D   %G  �=#  C#  �  W#  �!  W#   D  �@  �i#  o#  �  �#  �!  �!  D  D   �;  ��#  �#  j  �#  �!  D  D   �W  ��#  �#  W#  �#  �!  Q   *;  ��#  �#  W#  	$  �!  Q  D   �T  ��#  g�  �'"  	$    �  �  �  �  O$  @      _$  @     �  �%]  �(  N   9�$  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  V %  �\ X�   �  Y�  x  Z�   �7  \�$  	 %  $ N   J\%  D$  � n% �"  �# Q1%  � v�%  � x\%   u ~�%   !y�%  C0 zv  �  {7  �$ |D   �# �h%  �  '
&  � )�   ߣ  *�  �  +�  x  ,�     .�%  �& ."&  �%  � 1]&  ��  3�   .� 4�  _>  5&   � 7(&  � 7u&  (&  � :�&  F@ <�    =�  �\ >�   � @{&  � @�&  {&  !H�&  C0 J  "l K�  "ul L�   �& C.'  F@ E    F�  �\ N�&   ! P:'  �&  �# S�'  r$ U�   �" V�  5$ W�  �0 X�  �1 Y�   | [@'  " ^(  r$ `�   �" a�  5$ b�  �0 c�  �1 d�  % e�  
�� f�   ]( h�'  �' h(  �'  = �k�(  7( m�   ( n�  � o�  1 p�  � q�  � r�  H s�  � t�  � u�  �% v�  �! w(   = x(  8�! y(  P9 z(  h ' |"(  E% |�(  "(  & ,)  enc ��   )�  ��   o �8)  )  #� P�9*  �� �   �' �W  �$�% �  H$B! ��   P$( ��   X%toc �]&  `$�! ��(  x$D �G   �$2�  �.'   $�$ ��  $N �(  $� ��  $� �,)   $1 ��  ($'# ��  0$� �<  8$�� �h  @ � �E*  >)  
�%  (.�  N   ��,  �  � E' A(  5# �& K  [$ 	�! 
( x! �  � �! �$ � �% a' h W%   !� "x" #x $� %�& &�( '�' (k( 0?& 1� @� AM Q�" R� Sp Ti UG V W� Xq& `�  a� b�  c? p& �3 � �� � �U � �� �� ��% �% ��  �B �� �S! �+ �K �� �, ��# �� ��$ �� �# �l ��' ��" ��( �� �x' �� �� �B  �$  �� �� �Q  � �| �� �' �." �R# �l  �v# �Z" ��% � �$  �,  �,  	  �,  �  �,  �,   v  �  %�,  �,  	  �,  �  v  �,   �%  �( *-  	�,  ,& *5-  6' ,�,   z+ -�,   n)  A-  G-  	  e-  �  v    j   �)  $q-  w-  	  �-  �  v  U    nk  )�-  	�-  �;  )�-  �=  +5-   z+ ,e-   M" (B�-  �� D�"   � E�  � F,)     H
.  �-  &(( �!$  	 �H     '� �#-  	��H     'a �-  	��H     �  d.  @    	T.  '8% #d.  	��H     (K*  =	��H     ,%  �.  @    	�.  &i! C�.  	��H     ,%  �.  @    	�.  &� P�.  	��H     ,%  �.  @    	�.  ' �.  	��H     '[& �.  	`�H     ,%  </  @    	,/  '" /</  	@�H     ,%  h/  @    	X/  '� �h/  	 �H     '� �h/  	 �H     ,%  �/  @    	�/  '  '�/  	��H     '�& =�/  	��H     ) U0  *buf U!,  +? V!4   ,-c Z2    ) BB0  *buf B ,  +? C 4   ,-c G2    )! ,v0  *buf ,#,  +? -#4   ,-val 1N     .� 5	  0,C     �      ��B  /Jy  5  %� � /�  69*  �� p� /�  7�  �� o� 0�� 9�  �� �� 0� :	  �� �� 0R�  ;Q  �� �� 0� <j  � � 1�u  u�>C     2��  V6  0ZX t.'  #� � 2@�   3  0�� �  � ލ 0�$ ��  �� l� 0� �,�  �� s� 3�<C     �Y  �1  4U| 4T} 4Q	��H     5�H  s  3�<C     �Y  	2  4U| 4T} 4Q	Z�H     5�H  s  3'=C     �Y  <2  4U| 4T} 4Q	K�H     5�H  s  3o=C     �Y  o2  4U| 4T} 4Q	�H     5�H  s  3�=C     �Y  �2  4U| 4T} 4Q	$�H     5�H  s  3>C     �[  �2  4U 4QH 3J>C     �[  �2  4U  3�@C     �[  �2  4T�;$4QN  6UAC     �[  4U 0$0&4T24Q3  2P�  �3  0( c.'  f� `� 'B! c).'  P3l>C     �Y  �3  4U| 4T} 4Q	1�H     5�H  s  3�>C     �Y  �3  4U| 4T} 4Q	B�H     5�H  s  3�AC     �[  �3  4U 4Q~  6�AC     �[  4U 4Q~   7�B  �9C      ��  ~�5  8 C  �� �� 9��  :C  ��~;C  � �� ;'C  �� �� ;4C  � ۑ ;AC  E� ?� ;MC  �� �� :ZC  ��:gC  ��<tC  ��  5  ;uC  � � <�C   �  �4  ;�C  C� A� =�C  �>C     &       �4  ;�C  h� f�  6�;C     �[  4Qv   6O;C     �[  4U| 4Q��~  3�9C     �Y  55  4Uv 4T} 4Q	�H     5�H  s  3=:C     �Y  h5  4Uv 4T} 4Q	�H     5�H  s  3w:C     �Y  �5  4Uv 4T} 4Q	�H     5�H  s  3�:C     �Y  �5  4Uv 4T} 4Q	�H     5�H  s  >�:C     �[    3�;C     �Y  6  4Q	�H     5�H  s  3-<C     �[  96  4U��~4T 4Q04R14X04Y~  6@C     �[  4U��~4Q~   7�J  X,C      ��  ?�7  8�J  �� �� 8�J  ?� /� 9��  :�J  ��;�J  �� � ;�J  �� �� ;�J  R� B� ;�J  &� � ;�J  b� \� ?K  v-C     <
K  P�  &7  ;K  �� �� ;K  � � @!K  ��  ;"K  R� J�   3],C     �[  C7  4Uv 4T0 3�,C     �[  o7  4Uv 4T	��H     4Qs� 3	-C     �[  �7  4U��~4T 4Q04X04Y�� 3k-C     �[  �7  4Uv 4T	��H     4Q}  6�-C     �[  4U��~   7�G  �-C      ��  J\;  8�G  � ә 8�G  ,� � 9��  ;�G  �� {� ;�G  ڝ ʝ ;�G  �� �� ;�G  r� d� ;H  +� � :H  ��:H  ��:)H  ��~;6H  >� .� ;CH  �� � ;PH  �� �� ?]H  6/C     <fH  �  9  ;gH  �� �� =tH  6C     8       9  AuH  6>6C     �[  4U| 4Q��~  6�6C     �[  4U| 4Q��~  3�-C     I  J9  4Uv 4R14X��4Y�� 3.C     �[  h9  4Uv 4T  3>.C     �[  �9  4Uv 4T��~ 3�.C     �[  �9  4U| 4TH4Q} 4R~ 4X} 4Y��~ 3/C     �[  �9  4Uv  3A/C     �[  �9  4U| 4T  3L/C     �[  :  4U| 4T}  3�2C     	\  1:  4Uv 4T  3�4C     \  X:  4Uv 4T��~��~9 3 5C     	\  x:  4Uv 4T��~ 3�5C     �[  �:  4U| 4T14Q} 4R~4X} 4Y��~ 3�5C     #\  �:  4Uv 4T} 4Q~  3�5C     �[  
;  4U| 4TH4Q04R��~4X04Y��~ 3�?C     \  -;  4Uv 4T��~	� >V@C     �[  6�@C     \  4Uv 4T4��~3   7�H  j/C       `�  O�;  8I  ʣ ƣ 8�H  
� � 8�H  D� @� 9`�  ;I  ~� z�   7G  �/C      ��  Zj=  8'G  �� �� 8G  � � 9��  :4G  ��~;AG  �� }� :NG  ��:[G  ��;hG  ֥ ̥ ;uG  J� H� ;�G  w� m� A�G  ?�G  3C     3�/C     I  x<  4Uv 4R44X��4Y�� 30C     �[  �<  4Uv 4T~  3W0C     0\  �<  4Uv 4T��~ 3�0C     �[  �<  4U| 4TH4Q04R} 4X04Y��~ 31C     J  	=  4Uv 4Q~  3�2C     	\  '=  4Uv 4T~  33C     �[  ?=  4U|  >�4C     =\  6�4C     �[  4Uv 4T��~   7<F  x1C      ��  _i?  8[F  � � 8NF  l� N� 9��  :hF  ��~;uF  �� �� ;�F  � � A�F  :�F  ��:�F  ��;�F  ĩ �� ;�F  *�  � ;�F  �� �� ;�F  �� �� ?�F  b7C     3�1C     I  J>  4Uv 4R84X��4Y�� 3�1C     J\  g>  4Uv 4T8 3�1C     W\  >  4Uv  3�1C     d\  �>  4Uv  3�1C     q\  �>  4Uv  3B2C     �[  �>  4U| 4T84Q04R} 4X04Y��~ >}2C     	\  3�2C     �[  ?  4Uv 4T|  >�4C     W\  3�6C     	\  <?  4Uv 4T��~ 3m7C     �[  Z?  4U| 4T~  >v?C     �[    7VE  }7C      0�  d�B  8uE  � � 8hE  g� S� 90�  :�E  ��~;�E  =� 5� :�E  ��:�E  ��;�E  �� �� ;�E  $� � ;�E  u� m� ;�E  ߮ ծ ;�E  ^� T� ;�E  ׯ ѯ ;F  (�  � ;F  �� �� ;F  ΰ İ ;%F  O� ?� ?2F  R9C     3�7C     I  �@  4Uv 4R 4X��4Y�� 3�7C     J\  �@  4Uv 4T> 3�7C     W\  �@  4Uv  3�7C     ~\  �@  4Uv  3 8C     ~\  �@  4Uv  38C     ~\  A  4Uv  38C     ~\  A  4Uv  3&8C     ~\  3A  4Uv  358C     q\  KA  4Uv  3�8C     �[  �A  4U��~4T@4Q04R} 4X04Y��~ 3�8C     J\  �A  4Uv 4T} 1$ >9C     ~\  3P9C     �\  �A  4Uv  3a9C     �[  �A  4U��~4T��~ 3?C     q\  B  4Uv  3>?C     �[  >B  4U��~4T@4Q��~4R} 4X��~4Y��~ >�?C     �\  3�?C     �\  cB  4Uv  3�?C     �\  {B  4Uv  3�?C     �\  �B  4Uv  6�?C     �\  4Uv    3�/C     �C  �B  4Uv 4Ts 4Q2 6�>C     �C  4Uv 4Ts 4Q
   B�# �	  �C  Cpcf �"9*  D� �	  D�  ��  DR�  �Q  DZX �.'  Enn �4   Elen �4   DV` ��C  DϚ  ��C  ,Es �   ,Esrc �   ,Emm #4       �   �C  @    4   �C  @    .�! S	  `*C     �      �VE  /Jy  S  � �� /�  T9*  k� c� /� U�  в ʲ 'ߣ  W�  �P'�  W�  �X0� X	  � � 0�! Y�(  I� A� 1� ��+C     3�*C     I  �D  4Uv 4R�Q4X�P4Y�X 3�*C     �[  �D  4Uv 4T�L 3�*C     �[  �D  4Uv  3d+C     J  �D  4Uv 4Qs� 3�+C     J  E  4Uv 4Qs� 3�+C     J  :E  4Uv 4Qs� 6,C     J  4Uv 4Qs�  B�! �	  <F  FJy  �!  F�  �!9*  D� �	  DR�  �Q  Dߣ  ��  D�  ��  Ds �G   DO% �G   D�' �G   D�% �G   Dl# ��  D�& ��  Ei �G   Ej �G   Ek ��  D= �,)  G�   B�% (	  �F  FJy  (  F�  )9*  D� +	  DR�  ,Q  D�P  -�F  D�  .�F  Dߣ  /�  D�  /�  D�( 0�  D�( 0�  Ei 0)�  D� 0,�  G� � �  �  G  @    BW �	  �G  FJy  �  F�  �9*  D� �	  DR�  �Q  Dߣ  ��  D�  ��  DN �(  D�$ ��  D�$ ��  Ei �*�  G� " B.! �	  �H  FJy  �"  F�  �"9*  D�O ��&  D2�  �.'  DD ��  D? � �  Ei �-�  Dߣ  ��  D�  � �  D� �	  DR�  �Q  D� ��  DV` �  G� �,D r�  ,D�D ��     B� �.'  �H  F�  �(9*  FZX �(�  D2�  �.'  D;�  �j  Ei �G    B%% �j  I  F_>  �"&  F� �"�  F� �"�  Ei ��   .� u	  �&C     �       �J  /Jy  u&  �� �� /_>  v&&  ;� 3� /� w&�  �� �� /� x&�  #� � /
�  y&J  �� �� /�Y  z&J  S� C� 0� |	  � � Hi }�  �� �� 1�0  ��&C     6�&C     \  4U�U  �  B&$ ?	  �J  FJy  ?  Fߣ  @�  F.$ A(  D� C	  1�u  o*C     I|J  D�S H�J   ,D�( U!�'    ,%  J _	  1K  +Jy  _  +�  `9*  K� b	  -toc ci&  K_>  d&  KR�  fQ  -n g�  K�  i�  G�u  ,-i ��  K�# ��  ,-tmp �
&     L! 6�!C            �`K  M~ 6�  U .x &	  �!C            ��K  M~ &�  U .-   0'C     
       �L  /~ &�  �� �� /F@ &v  <� 8� N:'C     �\  4U	��H     4T�T  .�( �	  �!C            �TL  M~ �"�  UMn  �"v  TM�\ �"  Q .�( �	  �!C            ��L  M~ �"�  UMn  �"v  TM�\ �"  Q/�R  �"j  y� u�  .2' �	  �!C            �M  M�  �%9*  UMA! �%�,  TM' �%�,  Q .�' c	  p)C     U       ��M  /�  c+9*  �� �� /# d+v  �� � /�# e+�,  K� A� 0ZX g.'  Ĺ �� 6�)C     �Y  4Q�T5�H  �U  .�$ �	  @#C     =      �P  / �!�  � �� /�  �!�  �� v� /�^ �!�  � � /:1  �!7  �� s� 0�  �9*  S� I� 0Jy  �  ˼ ü 0� �	  3� '� 0�I �P  �� �� 0.$ �(  J� B� 0Ӏ ��  �� �� G�u  WO�/  %C       %C     A       R	�N  8�/  � � 8�/  P� J� @0   �  ;0  �� ��   OB0  �%C       �%C     d       CQO  8[0  Ŀ �� 8O0  � �� @g0  0�  ;h0  c� M�   O0  B&C       B&C     4       N	�O  8)0  �� �� 80  �� �� @50  `�  ;60  5� 3�   3v$C     �\  �O  4Us0 3�$C     �\  �O  4Us 4T|  3�$C     �[  �O  4U}  6�$C     #\  4U} 4Q|   �  .g �	  @"C     �       �*Q  /�  �&�  `� X� Preq �&�  �� �� 0�  �9*  � � 0�� �  �� �� Q� �	  0�  ��  v� n� R*Q  �"C      �"C     ;       �8IQ  �� �� 8<Q  �� �� S�"C     ;       ;VQ  !� � 6�"C     �\  4Us 4T0    B� �	  dQ  F�  ��  F-U ��  D�! ��(   .�! 	  BC     E      ��T  /Jy  !  S� G� /g !�  �� �� /�  !�  �� �� /G  !�  � �� /G  	!  >� :� 0�  9*  �� w� 0� 	  H� 8� 1�0  �DC     G�u  �2��  �R  0	*  	  �� �� 3WBC     �\  pR  4U~ 4T|  6CDC     �\  4U~ 4T|   T�CC            �R  0� /	  C� A� 6�CC     �\  4U~ 4T|   2��  �S  0( r  l� f� 0B! s  �� �� 0�T  tj  �� �� T�BC     �       AS  Hs y�   2� 0�  9�  '�� �h  �@6�CC     �\  4U	 �H     4T04Q�@4R0   7�T  4BC      p�  �S  8�T  W� U� 9p�  ;�T  �� z� AU  6LBC     X  4Us    7�T  �CC      @�  l-T  8�T  �� �� 9@�  ;�T  � � AU  6�CC     X  4Us    O�T  DC      DC            ��T  8�T  /� +� SDC            ;�T  l� h� AU  6DC     X  4Us    30BC     v0  �T  4U| 4Ts 4Qv  6�BC     v0  4U~ 4Ts 4Qv   )1 �+U  +g ��  K�  �9*  KR�  �Q  ,-i ��  ,KZX �.'     U�$ ��  � C     �       �&V  VV �"�!  �� �� W�" �#W#  TX
H ��-  �� �� X� �,)  !� � Ymin ��  J� D� Ymax ��  �� �� Ymid ��  � � X�j ��  �� �� XE  ��  1� '� Z�u  �<!C     9��  X� ��  �� ��   U� h�  @ C     y       ��V  VV h#�!  9� 5� W�j i#D  TX
H k�-  v� r� X� l,)  �� �� Ymin m�  �� �� Ymax m�  � � Ymid m�  }� s� XE  n�  �� �� 9p�  X� v�  G� =�   [e ]  C            �>W  WV ]�!  UX
H _�-  �� ��  UG L	    C            ��W  WV L�!  UW=R  M	  TX
H O�-  �� �� X�  P9*  � �  \*Q  �!C     N       �X  8<Q  Z� T� 8IQ  �� �� ;VQ  �� �� 6"C     �\  4Uv 4T�T  \�T  @'C     �      ��Y  8�T  � � A�T  ;U  �� �� =U  �'C            �X  ;U  �� �� =U  �'C     E       �X  ;U  /� +� 3�'C     �[  �X  4U}  6�'C     �[  4U}   6(C     �[  4U}   3c'C     �[  �X  4U}  3}'C     �[  �X  4U}  3"(C     �[  Y  4U}  39(C     �[  +Y  4U}  3M(C     �[  CY  4U}  3a(C     �[  [Y  4U}  3x(C     �[  sY  4U}  3�(C     �[  �Y  4U}  >�(C     �\   \�T  �(C            ��Y  8�T  k� e� ;�T  �� �� AU  N�(C     X  4U�U  \�H   )C     h       �WZ  8�H  � 	� ]�H  ]�H  ;�H  �� �� ;�H  � � ;�H  [� S� 6/)C     �\  4T|   \J  �)C     �       ��[  8$J  �� �� 81J  /� '� 8>J  �� �� ;KJ  +� %� T�)C            	[  ;nJ  z� v� 6�)C     �[  4U�U4T!`�H     ��H     �T4 $0.( 4Qs   @J  ��  81J  �� �� 8>J  � � 8$J  d� `� 9��  ;KJ  �� �� ^XJ  @|J  ��  :}J  �k6*C     �[  4U�U4T	@�H     4Q�k     _jO  jO  
_�?  �?  ^`�D  �D   a�K  �K  va�O  �O  2a�6  �6  �_9  9  c_�N  �N  �aF\  F\  �_�P  �P  �_�F  �F  �_ _   _  h_E1  E1  r_>Q  >Q  �_-4  -4  �_�3  �3  �_\  \  �_RH  RH  �_xL  xL  �_?  ?  �_�N  �N  �_�*  �*  [_�D  �D  �_T)  T)  �_P  P  �a�% �% [a^ ^ X_�3  �3  1_�U  �U  ^aBi  Bi   3q   (F  �  k0 $"  `DC     �B      B� :G  �9   X  ^� �L   �i L   int �i {S @�   g
  �       	@   v  #	@   �  &	@   |
  )	@    h  ,	@   (�  -	@   0�	  2X   8�  5X   < 	�   �  �   �
  8"h   
  K  	�   
�  L  
�  M  S  -  �  >   X   �	  	_   �  B"n  	t     ��  R   �f    �� ��  �N ��  �6  ��   �  Y�  	�  f   �  b  9      n�  	�  �  b  f    �  �
  	  f   .  b  9   9   f    �  �":  	@  �   PJ�  2�  L=   �  ML   pos NL   �  P  SF  Q   �1 R  (=9 SO  0R�  Ub  8y�  V=  @�� W=  H �  �  �\ �9   m  �f    o  ��  �  �  	  L   =  .  L   =  L    	C  �  C  2  \  	b  m  .     :9   �  J�  x Lm   y Mm   )  Oy  �  B   s�  M   um   }  um  V  vm  /  vm   t
  x�  �J  _   �E  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  _    ��  _   �  	X   B� 
=  L  A    C  s  C  v	  f     �  E  �  �  (N9  �  P:   Z�  Q:  �  S9  s  T�   [  U?  ?1  WX     	�  	:    Y�  	�  =  _   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  �X  b   "�  	�  �  %  <�  x >:   len ?A  *� @C   %  B�  �    `  	  1  X   X   1  f    	�  �  qD  	J  X   c  X   X   f    �  p  	v  �  X   X   f    �  `�  �  �   �% �  ?1  �X   �&  �  !  �   I  �7  ()  �c  0R   �f   8�  ��  @ 	�  	$  �  ��  %  �   D  	J  X   ^  f   ^   	�  �  q  	w  �  �   �  ?�  	�  �  �  =  L    �  Y�  	�  X   �  �  L   f    s  ��  	�  X   �  �  �   	2  W  0�f  �  ��   e� �7  �� ��  �� ��  �� ��   �� �d  ( �'  �  �!  lC  �  ��  �  -  �C  �  	�  �  ��   �  �
  �:  �  �A  �  �X   
  �_   �  �9   \#  �L   �   9   �  ,X   \&  7f   �0  D@   b   �y	  xx �	   xy �	  yx �	  yy �	   a  �6	  y	  z'  ��	  m  ��   ss  ��   �  ��	    ��	  	�	  �	  f    �  �
  �U  �f      ��	   %  ��	  �  $&
  	,
  �   e
  �� "
   �@ #
  �U  $f    �  7�
  �; 9
   ��  :
   L  <e
  _   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @	=_  ��  	?m   �  	@m  ~  	Bm  �  	Cm  �  	Dm   5  	Fm  (B  	Gm  0�  	Hm  8 �	  	J�  
   	s�  �  	u�   ��  	v�  �  	xm  �
  	zm  (  	{m   �  	}l  �  	�#�  	�  k  `
��  R�  
�b   (  
��  |  
��  �  
��  �  
��  �  
�H$  v  
��
  �  
�6  (�%  
��  07&  
�X$  8G   
��  X �  	�"�  	�  h  
�  �M 
/$   k  
�  R�  
b   �  	�"�  	�  %  8
;6  �� 
=5$   �M 
>�    
?�
   r$  
@�  0 5  	�$C  	I  %  �
�  �� 
5$   �M 
B$  �  
�   �  
'  (�� 

�  h�� 
�  p�� 
�  x K  	� �  	�  �  �	,�  �   	.�   �  	/�  O  	1�  C  	2�  �  	4�   d> 	6  (A  	7  0T  	9�  8  	:  @�  	<�  H�  	=  PE-  	?
  X�!  	D�  h:  	F�  �  	G�  ��  	H�  ��  	I�  ��  	K�  �  	L�  �U  	N�  ��  	O�  �)�  	Q�  ��  	R�  ��� 	SE  �K1 	W�  �R�  	Xb  �Jy  	Y.  �%  	[�
  ��	  	]
  �    	^f   ��8  	`~  � L  	 �  	�    X	��  �  	��   E-  	�
  N 	��  �8  	�/  P �  	*%�  	�  �  0	tE  k  	v�   �  	w�  �@ 	x�  ݖ 	y�  E-  	z
   N 	|_  0�  	}	  pR  	~	  x�  	�  �ߣ  	��  ��I 	��  ��  	��  �h  	��  ��S  	�E  �4  	��  �8  	�  �  	�f    �  	�9   �  	�m  o  	�m  �L 	�f    �8  	�i  ( �
  	L#R  	X  W  	H�  �  	J�   = 	Kd    	L�  d  	M�   �  _   	�d  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  	�  (0  	OX  #   	g)�  	�  �   �
�  =  
�y	   L  
��   $  
��  0�  
�Z   8m  
�#�!  h�  
�  pآ  
�H  tG   
��  x 	�  	�  	E  �?  	d�  �
  	�)<  	B  �   H
�{  �  
�f    "  
�  �!  
��   ~	  8	f�  �
  	h�   (  	i�  �� 	k	  �� 	l	    	nm  �  	om   �  	pm  (�  	qm  0 y  	s{    	�$  	  �  0'i  �N  )�   ?1  *�  }0  +�  i/  ,�  � -y	   �  	�)v  	|     H
��  ��  
��   ?1  
��  (  
�s  4  
�y	  \  
��  0  
�f   @ +!  	
  tag 	�   �U  		   �  	�  	
  `  _   	
U  w%   }#  �&  h  �  &     	
  E   	9
�  � 	;
U   ��  	<
�  �  	=
�  �  	>
�  �#  	?
�   �  	L
(�  	b  �  _   	�  :   �   ^$  1  �!  �!   :  	��  �  �	  �#  �'  	-  	  <  �   I$  �H  	N  Y  �   �&  �e  	k      �     	�   �!  H�  �  ��   S"  ��     �  �"  �	  �  �	   ;  �  (%  �  0�   �<  8��  �Y  @ 	�  R  ��  x  =�	  H  E#8  '  �  @J�  �  L�   �  M�  �� O  .� P.  �  Q�   �  RK  (�!  Sx  08'  T�  8   W!�  	�  -  (l  k  n�   �M o  ߣ  p�  �  q�   	3  k  )  	  	  .  �  �   w   .:  	@  K  �   �  1W  	]  r  �  r  R   	�	  K  6�  	�  �  �  �   	�  �  :�  	�  	  �  �  �   �  >  "  Y�  	�  	    6  �    R   �  _  	  	  2  6  �  r  R   $  f>  	D  Y  6  �  �   �  le  	k  	  �  6  �  	   #  x��  �� �    �  � �  H  � �  P�  �   X9!  � 2  `l� � Y  h  � �  p 	f    ��  �  H2N  �S  4E   �  59  (  69  04  7�  88  8  @ �  :�  �  �=�  R�  ?b   �  @�  n  A�  �  B�  1$  Cs  2�  EN  �� FN  `�L Hf   � �  J�  	Z  P   �  	�  	    .  �  �  �     �  &#  	)  4  �   �%  *@  	F  	  U  �   �%  -a  	g  r  �   {  1~  	�  	  �  �   �  4�  	�  �  �   l  8�  	�  	  �  �  �   �  <�  	�  	  �  �  �   �  @  	  	  ,  �  �  �  H   �  G8  	>  	  \  �  �  �  9   �'  Nh  	n  	  �  �  .   �  S�  	�  	  �  �  �  �  H  �   		  &  ���  �� �   i'  ��  H   ��  P  ��  X�A ��  `Y �  h�#  �4  p�  �U  x�  �r  �  ��  ���  ��  �U�  �,  ��!  �\  ���  ��  ��  ��  �&  ��  �   ��  �  �&  ��  	�  �>  ��  'O  �   xC  �   s/  ��  �  �  0tZ   �  v	   a   w	  �'  x	  !  y	  �#  z	   �  {	  ( �  }�  �  U's   	y   m  D   t�   �  v�   A  w�  �  x�  &  y�   !  {~   �  ��   	�   	  �   g   �  �    	�	  �  �	!  	!  !  g   �    �'  �+!  	1!  	  O!  g   �  s  O!   	�   �!  �!  ��  )�    ��  )�   �  )!   }  U!  �!  O  ;�!  _� =%�!   ݰ  >%g    	�!  �  @�!  	�!  cA  
�,�!  	�!  /  
�"  �� 
�q   �M 
�"   ?<  
�,*"  	�"  �5  P
��"  �  
��   �� 
��"  �Y 
��"  �H 
�#  U@ 
�:#   �9 
�#f#  (�A  
�#�#  0�^  
�#�#  8�^  
�#�#  @N7  
�#$  H 0"  ��  
��!  (Z  
��"  	�"  	  �"  �!  	   17  
�#  		#  #  �!   �G  
� #  	&#  �  :#  �!  U   %G  
�F#  	L#  �  `#  �!  `#   	U  �@  
�r#  	x#  �  �#  �!  �!  U  U   �;  
��#  	�#  s  �#  �!  U  U   �W  
��#  	�#  `#  �#  �!  b   *;  
��#  	�#  `#  $  �!  b  U   �T  
��#  g�  
�0"  $  	  �  
�  	�  �  X$  L      h$  L     �  
�%f  �3  5�$  !num 7�  !str 8   +P  :u$  �J  =�$  key ?�$   �U  @@    �7  D$�$  	�$  O  H�$  	�$  �  %  %   	�$  �Z  K%  	%  s  .%  %  %   �S  (O�%  �� Q�   �  R�  �6 S�  �B  U�$  3  V%  >) X�%    	�$  �6 Z.%  e-  \ �%  	.%  �) N�%  �- PX    z/ QX   i* RX   �7 SX    �5 U�%  �%  	�%  	�   "s8&  C0 u�   !l v9   !ul wL    0 nz&  F@ p�    ߣ  qX   �6 rX   �\ y&   :) {8&  z&  �* ��&  ��  �A   �  �A  �, �:  ��  �:  �0 �:  �1 �:  
 J6 ��&  �, 8�i'  F@ ��    = �9   6 �A  �7 �A  bbx ��&  �I �=   bpr �L   (Ӏ �A  0 1 ��&  �. @��'  pad �A   bpp �A  �S �9   end �9   �^ ��'  �* �L    �7 �L   (bbx ��&  0 	i'  -7 �u'  #X7 8� ��)  F@ ��    bbx ��&  � �L   �$ �L    � �L   (�, �X   0/ �A  4� �9   8�0 �9   @�1 �9   H�* �L   P�7 �L   X�^ ��'  `�7 �L   h�6 �L   p/ ��'  x�1 �L   ��+ �L   ��O ��)  �n* ��   �.0 �L   ���  ��'  ��8  �f   �v. ��)  �$�7 ��)  �@ $�  �A  �� %bpp �A  � $R�  �b  �� $k, ��)   � $j, �L   � $�1 ��%  �  	z&  L   �)  &L   �� o/ ��'  _   �,  O.  �/ �0 H0 �- �7 a1 6 �+ �2 	Q- 
-5 T6 �4 3 -6 �8 �+ G1 4 �3 i-  �4 !3* "?+ #z1 $5 %�3 &*1 '#3 ( , 0�/ 1�5 @W/ Ad3 Q7 RC, S�, T�+ UU4 VZ. W�0 X�) `�5 aQ* b�* cz5 p�4 �`5 ��3 ��2 ��* ��- ��8 ��6 �D5 ��, ��- �=7 �72 ��) �n) �+ ��+ �A3 ��1 ��1 �u6 ��6 ��, ��/ �1 �/ ��- �[+ �3 ��5 ��7 �4 �`8 �!+ ��/ �d7 �{4 �p2 �) �;/ �8 ��) �V2 ��/ ��* ��. �/ � '*. >�%  �&  8,  L   R (,  (2- P 8,  	 �H     ).- �S   S;8 �l,  	r,  	  �,  �   L   L   f   f    {.  ��,  �F �&   �  �L   �6 �L   R�  �b   �2 ��,  #u8 x@ ��-  ?1  �L    cnt  L   row L   �1 :  o8 :  u4 :  �* :  �- :   9 	:  "la �   (�7 9   0v�  �-  8�@ &  @(5 �)  H*�$ �,  H@ *R�  b  h@ *�  L   p@  	�)  �4 �,  �   .  L     �-  +�4 r.  	 �H     J  9.  L    ).  ,a2i �9.  	��H     J  e.  L    U.  +0 �e.  	`�H     +\3 �e.  	@�H     J  �.  L    �.  +, ��.  	0�H     $ _   J�.  D$  � n% �"  �# Q�.  � v!/  � x�.   u ~!/   "yO/  C0 z  �  {H  �$ |U   �# ��.  �$  g/  	m/  	  �/  �  �/  �/   	  �  %�/  	�/  	  �/  �    �/   	O/  �( *�/  �/  ,& *�/  6' ,[/   z+ -�/   �8 ,0  enc .�   )�  /�   - 1�/  -�/ 84�0  �� 6"   B! 8�   �.( 9�    .�8 ;�-  .$7 =�0  .� ?E  .�� @q   .�. B�  0 	0  64 D�0  	*0  
�  G.�  *2 (6 1  
H 8�"   � 9�  � :�0    �) <1  	�0  (�. �*$  	��H     +�. �#�/  	ЇH     �  O1  L    ?1  +�5 �#O1  	��H     /�0  �	��H     0I) �  KC     
       ��1  1~ �&�  �� �� 1F@ �&  � �� 2KC     &p  3U	��H     3T�T  0�0 �	  �GC            �?2  4�  �%�0  U4A! �%�/  T4' �%�/  Q 0�5 g	  �SC     �       �3  1�  g+�0  @� <� 1# h+  � y� 1�# i+�/  �� �� 5ZX k�)  �� �� 6�0  ��SC     7�I  �SC       ��  p8�I  �� �� 8�I  �� �� 9��  :�I  ;�SC     `k  3T�T    0�, 	   HC     �      �F4  1 !�  6� *� 1�  	!�  �� �� 1�^ 
!�  +� %� 1:1  !H  |� t� <bdf �0  �� �� 5�  �  � � =� 	   5�I F4  ^� R� 5)�  i'  � �� <bpp X   ]� Y� 6�u  [ HC     >�HC     3p  14  3Us  ;[IC     @p  3Us0  	�  ?. �	  �4  @�  �&�  Areq �&�  B�  ��  B�� �  B�8 ��-  B� �	  B�  ��   02 �	  �GC     G       �25  1�  ��  �� �� 1-U ��  � � 5�8 ��-  @� >� ;�GC     Mp  3T�T  0�2 Q	  `ZC     4      �E  1Jy  Q!.  s� c� 1m6 R!�  E� !� 1�  S!�  �� �� 1G  T!�  � � 1G  U!  I� E� 5� W	  �� �� B�  X�0  5R�  Yb  �� �� 5v�  [�-  �� �� +�� \�%  ��~6�u  ��gC     6�0  ��^C     C��  @  5ZX ��)  )� � C��  �9  5�� �  A� 3� 5�$ ��  �� �� 5� �,�  �� �� 5�\ �9   �� �� D�I  PcC       �  �7  8�I  �� �� 8�I  �� �� 9 �  :�I  ;ccC     `k  3Uv 3T	��H        E�I  �cC      �cC            ��7  8�I  � � 8�I  @� >� F�cC            :�I  ;�cC     `k  3Uv 3T	Z�H        E�I  �cC      �cC            	8  8�I  e� c� 8�I  �� �� F�cC            :�I  ;�cC     `k  3Uv 3T	K�H        E�I  dC      dC            �8  8�I  �� �� 8�I  �� �� FdC            :�I  ;3dC     `k  3Uv 3T	�H        E�I  rdC      rdC            /9  8�I  � 	� 8�I  9� 7� FrdC            :�I  ;�dC     `k  3Uv 3T	$�H        >LhC     Zp  9  3QH >xhC     Zp  D9  3T} 0$0&3Q~ 0$0& >iC     Zp  `9  3T23Q3 ;�iC     Zp  3T�;$3QN   G�dC     �       �9  <cur T�'  `� \� <n UL   �� �� ;�dC     gp  3Uw 3T@3Q03X03Y��~  C0�  �<  5( o�)  �� �� 5B! o-�)  9� 5� 5�T  ps  w� o� C�  |;  <s ~  �� �� C@�  �:  +�� �q  ��;:kC     sp  3U	��H     3T03Q��3R0  >AjC     �p  �:  3U~ 3Q��~ >fjC     �p  �:  3U~ 3Q��~ >�jC     �p  �:  3Uv 3T	S�H      >�jC     �p  ;  3Uv 3T	Y�H      >�jC     �p  ;;  3T	4hH      >�jC     �p  `;  3Uv 3T	^�H      ;kC     �p  3T	g�H       C��  �;  +�� �q  ��;�gC     sp  3U	��H     3T03Q��3R0  D�I  `gC      ��  t%<  8�I  � � 8�I  A� ?� 9��  :�I  ;wgC     `k  3Uv 3T	1�H        7�I  �gC      ��  v8�I  f� d� 8�I  �� �� 9��  :�I  ;�gC     `k  3Uv 3T	B�H         D�I  L`C      @�  ��<  8�I  �� �� 8�I  '� !� 9@�  :�I  ;p`C     `k  3Uv 3T	~�H        E�I  `C      `C            �`=  8�I  r� p� 8�I  �� �� F`C            :�I  ;�`C     `k  3Uv 3T	�H        DF  �`C      ��  �-@  8�F  �� �� 9��  H�F  ��~I�F  9� '� I�F  �� �� I�F  E� C� I�F  z� j� H�F  ��I�F  (� "� I�F  {� q� H�F  ��J�I  aC      aC     %       �o>  8�I  �� �� 8�I  � � FaC     %       :�I  ;AaC     `k  3U| 3T	�H        J�I  PaC      PaC            ��>  8�I  A� ?� K�I  FPaC            :�I  ;haC     `k  3U| 3T	�H        L�I  waC      ��  �9?  8�I  q� m� K�I  9��  :�I  ;�aC     `k  3U| 3T	�H        L�I  �aC       �  ��?  8�I  �� �� K�I  9 �  :�I  ;�aC     `k  3U| 3T	�H        MG  0�  @  IG  	� � MG  `�  @  IG  A� ?� N!G  [eC     <       �?  I"G  f� d�  ;�bC     �p  3Q~   ;:bC     �p  3U} 3Q��~  O�aC     �p    >�`C     �p  M@  3Uw 3Q��~ ;�bC     gp  3Uw 3T 3Q03R13X03Y��~  DZJ  �ZC      ��  l�D  8�J  �� �� 8�J  d� P� 8yJ  b� L� 8lJ  \� J� 9��  I�J  1� #� I�J  �� �� I�J  `� D� H�J  ��~P�J  �^C     P�J  �_C     Dif  v[C       ��  �SA  8�f  �� �� 8wf  �� ��  D�b  v[C      ��  ��C  8�b  �� �� 8�b  �� �� 8�b  P� @� 8�b   	  	 9��  H�b  ��I�b  � 	 � 	 I	c  8	 (	 Ic  	 �	 I#c  �	 �	 I0c  U	 Q	 I=c  �	 �	 IJc  �	 �	 IWc   	 �	 Idc  �	 �	 Iqc  �	 �	 I~c  �	 �	 I�c  	 		 H�c  ��P�c  m\C     M�c  ��  �B  I�c  �	 �	 ;L\C     gp  3U��~3T13Q} 3Rs 3X 3Y��~  >�[C     gp  �B  3U��~3T13Q03R
 3X03Y��~ >�[C     �p  C  3U��~3T } "3Q��}}  >z\C     �p  2C  3U��~ Q!_C     eC  3U��~3Tv 3Q��~3R��3X��~ Qe_C     �C  3Tv 3Q��~3R��3X��~ ;�eC     �p  3U 3Q}    EJ  �_C      �_C            3	D  8J  �	 �	 F�_C            :'J  :4J  :?J  :LJ  ;�_C     �g  3Uv    >�ZC     �p  CD  3Uv 3Tx@ 3Q��~ >�]C     gp  aD  3T13Y��~ >�_C     �p  zD  3Uw  >�_C     f  �D  3U��~ >�_C     �p  �D  3Uw  ;`C     �p  3Uw 3T    >�ZC     �p  �D  3U~ 3T0 >�^C     E  �D  3Us  ;�hC     E  3Us   R�3 6`OC     �       �F  1m6 6�   	 	 5�  8�0  �	 	 5R�  9b  �	 �	 EJ  �OC       �OC     
       A�E  8J  		 		 F�OC     
       :'J  :4J  :?J  :LJ  O�OC     �g    >�OC     �p  �E  3Uv  >�OC     �p  
F  3Uv  >�OC     �p  "F  3Uv  >�OC     �p  :F  3Uv  >�OC     �p  RF  3Uv  >PC     �p  jF  3Uv  ;#PC     �p  3Uv   S�2 �	  2G  Tbdf �"�0  '� �	  '�  ��  'R�  �b  'v�  ��-  'ZX ��)  'V` �2G  Unn �@   Ulen �@   'Ϛ  �BG  VWs �   VWsrc �   VWmm $@       �   BG  L    @   RG  L    X. ��  �FC     �       �MH  Y8 �#�!  4		 0		 Z�" �#`#  T[
H � 1  q		 m		 [� ��0  �		 �		 \min ��  �		 �		 \max ��  )
	 
	 \mid �!�  �
	 �
	 [E  ��  	 	 [�j ��  �	 �	 ]�u  �UGC     9��  [� ��  D	 :	   XL8 [�  `FC     y       �$I  Y8 [#�!  �	 �	 Z�j \#U  T[
H ^ 1  	 		 [� _�0  H	 F	 \min `�  o	 k	 \max `�  �	 �	 \mid `!�  	 
	 [E  a�  �	 �	 9p�  [� i�  �	 �	   ^�8 P@FC            �eI  Z8 P�!  U[
H R 1  �	 �	  X5, @	   FC             ��I  Z8 @�!  UZ=R  A	  T[
H C 1  �	 �	 [�  D�0  �	 �	  ?�8 �	�)  J  @v�  �	'�-  @F@ �	'  Bd0 �	J   	@   _�) >	ZJ  @v�  >	�-  BZX @	�)  Wi A	L   B�^ B	�'  BR�  C	b   ?%* �	  �J  @Jy  �".  @v, �"b  @�@ �"&  @v�  �"�J  B�2 �L   Wp ��J  BR�  �b  B� �	  `�u  %	`�0  2	 	�-  	�-  0�. j	  �pC     �      ��R  1+ j$�   	 	 12 k$L   k	 A	 1�2 l$L   $	  	 1B- m$f   w	 ]	 1w* n$f   �	 �	 +�[ pL   ��}5�@ q�R  	 �	 Wp r�J  5v�  s�-  2	 *	 <s t�   �	 �	 5R�  vb  ;	 )	 5� w	  	 �	 6�u  �NvC     C`�  �L  <i �@   �	 �	 5ZX ��)  �	 �	 >HrC     �p  `L  3U~ 3T  ;�rC     �p  3Tv 3Q~ 3R   G�xC     L       �L  <bpp LA  	 	 O�xC     �a   G=wC     �       �M  +�- i�R  ��}>iwC     q  M  3U��}3T	��H      >|wC     �k  4M  3T	e�H     3Q��}a+^  �Q >�wC     q  ZM  3U��}3T	��H      ;�wC     �k  3T	q�H     3Q��}a+^  �Q  E�b  !sC       !sC            �&�M  8�b  =	 ;	 F!sC            :�b  O8sC     �f    D�a  �sC       ��   N  8b  b	 `	 9��  :b  OtC     �f    E�a  tC      tC            yN  8b  �	 �	 FtC            :b  OtC     �f    D_  IuC       ��  -�O  8%_  �	 �	 82_  �	 �	 8_  /	 )	 9��  I?_  |	 x	 HL_  ��}HY_  ��}If_  �	 �	 Is_  �	 �	 P�_  �uC     b�_  Dif  �uC       �  �AO  8�f  �	 �	 8wf  �	 �	  >�uC     �p  YO  3Us  >�uC     �p  ~O  3U��}3Ts 3Q|  >�uC     �c  �O  3U��}3T	ۃH     3Q��}3R|  >�uC     f  �O  3U��} ;�yC     f  3U��}   D�b  �vC       p�  E"P  8�b  �	 �	 9p�  :�b  O�vC     �f    E�b  �vC      �vC            F{P  8�b  	 	 F�vC            :�b  O�vC     �f    E�b  �vC      �vC            G�P  8�b  @	 >	 F�vC            :�b  O�vC     �f    O�qC     �_  >rC     �p  	Q  3U 3T8� 3Q��} >sC     �c  >Q  3U}Ȁ3T	��H     3Q�U3R�T >�sC     �c  sQ  3U}Ȁ3T	��H     3Q�U3R�T O.tC     �a  O<tC     �a  >�tC     �c  �Q  3U| 3T	��H     3Q�U3R�T >�tC     �o  �Q  3U|  >�tC     yo  �Q  3Tt  >�tC     �p  R  3Uv  >uC     gp  6R  3Uv 3T13Q03X03Y��} >EuC     �p  NR  3T|  >tvC     �c  �R  3U}Ȁ3T	��H     3Q�U3R�T >,xC     gp  �R  3Uv 3TH3Q03X03Y��} >~xC     �p  �R  3U 3T(3Q��} ;�xC     �p  3T   	`,  �   S  L    0?4 	  �lC     d      �vW  1+ )�   g	 c	 12 )L   �	 �	 1�2 )L   	 	 1B- )f   _	 A	 1w* )f   �	 �	 +�+ L   ��~5�@ �R  �	 �	 <p 	�J  V 	 : 	 5F@ 
�   �!	 s!	 5�\ �   5"	 +"	 +�- �R  ��~5� 	  �"	 �"	 6�u  cPnC     E�I  �lC       �lC     %       �T  8�I  �#	 �#	 8�I  $	 $	 F�lC     %       :�I  ;mC     `k  3T	e�H        D�I  mC       p�  +�T  8�I  :$	 6$	 8�I  �$	 �$	 9p�  :�I  ;8mC     `k  3T	q�H        D�^  �nC       ��  NV  8�^  �$	 �$	 8�^  R%	 J%	 8�^  �%	 �%	 8�^  B&	 :&	 8�^  �&	 �&	 9��  I�^  `'	 V'	 I�^  �'	 �'	 I�^  )	 �(	 I�^  �)	 �)	 7�`  �nC      ��  %	8�`  *	 *	 8�`  �*	 {*	 9��  I�`  �*	 �*	 >oC     q  �U  3U| 3T��" ;?pC     q  3U| 3T��"     >�mC     �k  0V  3T| a+^  �Q >7nC     q  UV  3Uw 3T	��H      >HnC     �k  �V  3T	q�H     3Qw a+^  �Q >{nC     q  �V  3Uw 3T	��H      >�nC     �k  �V  3T	e�H     3Qw a+^  �Q >foC     �c  W  3U~ 3T	��H     3Q| 3Rv  >�oC     �o  W  3U~  >�oC     yo  7W  3Tw  >�oC     �k  RW  a+^  �Q ;pC     �k  3T| 3Qs a+^  �Q  0�* �	  �yC     I      ��]  1+ �%�   +	 +	 12 �%L   c+	 S+	 1�2 �%L   ,	 ,	 1B- �%f   y,	 u,	 1w* �%f   �,	 �,	 <c �X   !-	 -	 5�7 �X   �-	 �-	 <s ��   .	 .	 <bp �=  q.	 g.	 <i �L   �.	 �.	 +�[ �L   ��5&0 �!L   �/	 �/	 <p �J  �/	 �/	 5)�  �'  l0	 X0	 5v�  �-  J1	 :1	 5R�  b  �1	 �1	 +� 	  ��6�u  ��{C     6�. �2�C     C��  DY  <sw �A  52	 -2	 ;s�C     Zp  3T@   C��  �Y  5�7 �L   �2	 �2	 ;��C     gp  3U| 3T13Q03X03Y��  D�b  �zC       ��  -$�Y  8�b  �2	 �2	 9��  :�b  O�zC     �f    D�a  ӂC      ��  �Z  8b  �2	 �2	 9��  :b  O�C     �f    E�b  VC       VC            d'hZ  8�b  .3	 ,3	 FVC            :�b  OeC     �f    E�b  ��C       ��C            t'�Z  8�b  S3	 Q3	 F��C            :�b  O�C     �f    D�a  ��C       `�  �[  8b  z3	 v3	 9`�  :b  OǂC     �f    >szC     �c  5[  3UvȀ3T	��H     3Qs 3R~  >�{C     �_  M[  3U}  >#|C     �p  e[  3U|  >\}C     gp  �[  3U| 3T83Q03X03Y�� >~C     q  �[  3Q83R	 FC      >3~C     �p  �[  3U|  >N~C     �c  \  3U} 3T	��H     3Qs 3R~  >b~C     �o  \  3U}  >l~C     yo  2\  3Tt  >�~C     gp  `\  3U| 3T13Q03X03Y�� >�~C     �p  x\  3Ts  >:C     �c  �\  3UvȀ3T	��H     3Qs 3R~  >�C     �c  �\  3UvȀ3T	��H     3Qs 3R~  O�C     "b  >��C     �c  ]  3UvȀ3T	��H     3Qs 3R~  >��C     �c  Q]  3UvȀ3T	��H     3Qs 3R~  O��C     �a  O�C     �a  O�C     "b  >��C     gp  �]  3U| 3T83Y�� >��C     gp  �]  3U| 3T83Y�� >%�C     �p  �]  3U|  ;A�C     Zp  3T@   ?�2 N	  �^  @v�  N%�-  @F@ O%�   @�\ P%�   @�2 Q%L   Bd0 SJ  BZX T�)  Wfp T�)  BR�  Ub  B� V	  `�u  � ?;0 X   _  @+  �   @2  L   @F@  &  @�\  &  @v�   �-  B: X   Wsp �   Wep �   Wp �)   ?�, �	  �_  @v�  �-�-  @�@ �-&  @�2 �-L   Wlen �@   BF@ ��_  B�$ ��,  BR�  �b  B� �	  `�u  `�0   �   �_  L   � 0- �	  �JC     �       ��`  1v�  �$�-  �3	 �3	 1&- �$�   4	 4	 clen �$L   \4	 T4	 <cp ��   �4	 �4	 5R�  �b  �4	 �4	 +� �	  �L6�u  ��JC     >�JC     gp  l`  3T13Y�L ;�JC     �p  3T} 3Qv   ?v+ t�)  �`  @F@ t"�   @v�  u"�-  Bd0 wJ   ?�6 B	  4a  @F@ B%�   @ߣ  C%X   @v�  D%�-  Wn F@   Wp G�)  BR�  Hb  B� I	  `�u  n 0�3 .X    FC            ��a  da .  Udb /  T<c1 1�'  	5	 5	 <c2 1�'  .5	 ,5	  0�) :  @EC     �       ��a  cs �   [5	 Q5	 <v :  �5	 �5	 <neg :  U6	 K6	  ?<. �A  "b  As ��   Wv �A   0�) �9   `DC     �       ��b  cs ��   �6	 �6	 <v �9   P7	 D7	 <neg �9   �7	 �7	  ?�4 �L   �b  As ��   Wv �L    ?*) 		  �c  @Jy  	&.  @�  
&`,  @w* &f   Alno &�c  Wcb `,  B�2 L   B* L   B�	 X   B: X   B38 %X   BӀ -   B�S -   Wend %-   By�  *-   B�8 2-   Wbuf �   BR�  b  B� 	  `�u  �VB6^  R�    	L   ?%, �	  ud  @�$ �#ud  @_, �#�   @+ �#�   @2 �#L   B�4 �L   Bt� �X   Wsp ��   Wep ��   Wend ��   B�2 �{d  B� �	  6�u   �PC      	�,  �   �d  L    ?�6 v�   �d  @�$ v#ud  Ac w#X   @L- x#�c  Wi zL   Wj zL   Wdp {�   VWfp ��     _^) [0e  @�$ [#ud  An \#L   Wi ^L   Wu ^L    0�1 9	  �IC     �       �f  1�$ 9$ud  c8	 [8	 1��  :$L   �8	 �8	 +� <	  �\6�u  U�IC     9�  54. AL   9	 9	 5�8 BL   X9	 N9	 5G. CL   �9	 �9	 5R�  Db  #:	 :	 ;JC     gp  3T83Y�\   R�1 +PJC     )       �if  1�$ +!ud  w:	 o:	 5R�  -b  �:	 �:	 OhJC     �p   _9 "�f  @�$ "!ud  @R�  #!b   e�b   KC     y       ��f  8�b  ;	 ;	 I�b  i;	 a;	  e�a  �KC     g       ��f  8b  �;	 �;	 Ib   <	 <	  eL4  LC     �       ��g  8^4  �<	 ~<	 8k4  �<	 �<	 Ix4  &=	 "=	 I�4  `=	 \=	 I�4  �=	 �=	 f�4  I�4  �=	 �=	 gL4  �LC            8k4  B>	 >>	 8^4  >	 {>	 F�LC            :x4  :�4  :�4  :�4  :�4  2�LC     �4  3U�U3T0    eJ  �LC     �      �j  8J  �>	 �>	 I'J  ?	 
?	 I4J  S?	 /?	 I?J  �@	 �@	 ILJ  qA	 oA	 >�LC     �p  Wh  3Us  >�LC     *q  oh  3Ts  >�LC     �p  �h  3Us  >MC     �p  �h  3Us  >gMC     �p  �h  3Us  >�MC     �p  �h  3Us  >�MC     �p  �h  3Us  >�MC     �p  �h  3Us  >NC     �p  i  3Us  >NC     �p  /i  3Us  >8NC     �p  Gi  3Us  >LNC     �p  _i  3Us  >|NC     �p  wi  3Us  >�NC     �p  �i  3Us  >�NC     �p  �i  3Us 3T|  >�NC     *q  �i  3Uv��"3Ts  >OC     �p  �i  3Us  >*OC     �p  �i  3Us  ;JOC     �p  3Us 3T|   e�c  @PC     '      �`k  8�c  �A	 �A	 8�c  ,B	 (B	 8�c  oB	 eB	 8�c  �B	 �B	 :
d  :d  :$d  :0d  :<d  :Id  fVd   h�c  @�  8�c  >C	 6C	 8�c  �C	 �C	 8�c  ED	 =D	 8�c  �D	 �D	 9@�  I
d  E	 E	 Id  �E	 vE	 I$d  #F	 F	 I0d  lG	 TG	 I<d  fH	 `H	 HId  ��IVd  �H	 �H	 Pcd  �RC     >�QC     0e  Ik  3U|  ;�RC     0e  3U|     e�I  pSC     4       ��k  8�I  aI	 WI	 8�I  �I	 �I	 I�I  ,J	 (J	 ;�SC     q  3U�T  e�]  pTC     �      �yo  8^  rJ	 bJ	 8^  5K	 #K	 8^  �K	 �K	 8+^  �L	 �L	 I8^  �L	 �L	 IE^  �M	 �M	 IR^  �M	 �M	 I^^  N	 yN	 Hk^  ��Px^  RZC     E�b  `VC      `VC            u�l  8�b  �N	 �N	 F`VC            :�b  ;vVC     �f  3U|    E�b  @WC      @WC            �m  8�b  �N	 �N	 F@WC            :�b  ;VWC     �f  3U|    D�`  �XC      ��  �an  8�`  O	 O	 8�`  RO	 NO	 8�`  �O	 �O	 9��  I�`  �O	 �O	 Ia  P	 P	 Ia  YP	 UP	 Ha  ��P*a  �XC     >�XC     q  �m  3Uv 3T~  >\YC     gp  �m  3U 3TH3Y�� >�YC     �p  �m  3Uv  >�YC     gp  %n  3U 3T13Q03R��3X03Y�� >�YC     �p  En  3Tv 3Q�� ;ZC     �p  3Q~ 3R    >�TC     q  yn  3Uv  >UC     q  �n  3Uv 3T~  >,VC     �p  �n  3U}  >XVC     �p  �n  3U} 3T| 3Q�� >�VC     gp  �n  3U} 3TH >$WC     �p  o  3U} 3T| 3Q�� >uWC     �p  .o  3R}  >�WC     "b  Fo  3U|  >�XC     "b  ^o  3U|  ;�XC     q  3Uv 3T~   e�d  �kC     �       ��o  i�d  Ui�d  TI�d  �P	 �P	 I�d  �P	 �P	 I�d  3Q	 1Q	 j�d   g�d  �kC     E       I�d  XQ	 VQ	   e�d  0lC     I       �&p  ie  U:e  :$e  je   k�*  �*  [k�U  �U  
�k�D  �D  
�kP  P  
�kjO  jO  	l�6  �6  �k�3  �3  
1k�?  �?  ^lBi  Bi  m�D  �D   l�K  �K  vl�O  �O  2k�R  �R  �lF\  F\  �l�Z �Z k9  9  cl�-  �-  `l�,  �,  nl  gld\  d\  zl_T  _T  XlUP  UP  h   �L  �  9 $"   �C     ��      	� X  ^� �@   �i int G   �i S   {S @
�   g
  
�      
 	4   v  
#	4   �  
&	4   |
  
)	4    h  
,	4   (�  
-	4   0�	  
2G   8�  
5G   < 	�   �  �   �
  
8"a   
  
K  	�   
�  
L  
�  
M  S  �9  ?  -   O  @    .�  �[  -  �[  �n  �  n  >   G   �	  	S   �  �  B"�  	�     ��  R   �_    �� ��  �N �  �6  �5   �  Y�  	�  _     �  -      n  	%  5  �  _    �  �A  	G  _   e  �  -   -   _    �  �"q  	w  �   PJ  2�  Lt   �  M@   pos N@   �  P8  SF  Q8   �1 RD  (=9 S�  0R�  U�  8y�  Vt  @�� Wt  H �  �8  �\ �-   m  �_    o  �  �  �P  	V  @   t  e  @   t  @    	z  �  z  2  �  	�  �  e     :-   �  J�  x L�   y M�   )  O�  �  B   s'  M   u�   }  u�  V  v�  /  v�   t
  x�  �J  S   �|  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  S    ��  S   �  	G   B� 
t  L  n    z  s  z  v	  _     �  |  �  �  (Np  �  P[   Z�  Q[  �  Sp  s  T�   [  Uv  ?1  WG     	�  	[    Y  	�  =  S   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "�  	�  �  %  <)  x >[   len ?n  *� @z   %  B�  )    `H  	N  h  G   G   h  _    	6  �  q{  	�  G   �  G   G   _    �  �  	�  �  G   G   _    �  `�O  �  �O   �% �U  ?1  �G   �&  �;  !  �;   I  �n  ()  ��  0R   �_   8�  �'  @ 	  	[  �  ��  \  �   {  	�  G   �  _   �   	�  �  �  	�  �  �   �  ?�  	�  �  �  t  @    �  Y�  	�  G     �  @   _    s  �  	   G   4  �  4   	i  W  0��  �  ��   e� �n  �� ��  �� ��  �� �   �� ��  ( �'  �:  �!  lz  �  ��  �  -  �z  �  	�  �L  ��  �  ��   �  �
  �[  �  �n  �  �G   
  �S   !	  �  �-   \#  �@   �   -   �  ,G   W	  \&  7_   �0  D4   b   ��	  xx �J	   xy �J	  yx �J	  yy �J	   a  ��	  �	  z'  �
  m  ��   ss  �	   �  ��	    �
  	#
  .
  _    �  �Y
  �U  �_      �
   %  �.
  �  $s
  	y
  �   �
  �� "f
   �@ #f
  �U  $_    �  7�
  �; 9f
   ��  :f
   L  <�
  S    �-  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=�  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  J-  
   s  �  u�   ��  v�  �  x�  �
  z�  (  {�   �  }�  �  �#(  	.  k  `��  R�  ��   (  �	  |  �	  �  �	  �  �!	  �  ��$   v  ��
   �  ��  ( �%  ��  0 7&  ��$  8 G   �	  X �  �"�  	�  h  )  �M k$   k    R�  �   �  �"6  	<  %  8;�  �� =q$   �M >�    ?�
   r$  @"  0 5  �$�  	�  %  �  �� q$   �M ~$  �  �   �  y  (�� 
�  h��   p�� $  x K  �   	  �  �,�  �   .2	   �  /2	  O  12	  C  22	  �  42	   d> 6]  (A  7]  0T  9	  8  :c  @�  <	  H�  =i  PE-  ?Y
  X�!  D'  h:  F		  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q5  ��  R�  ��� S�  �K1 W)  �R�  X�  �Jy  Ye  �%  [�
  ��	  ]Y
  �    ^_   ��8  `�  � L   �  	�    X�5  �  �   E-  �Y
  N �G  �8  �|  P �  *%B  	H  �  0t�  k  v   �  w  �@ x5  ݖ y!	  E-  zY
   N |�  0�  }J	  pR  ~J	  x�  �  �ߣ  ��  ��I ��  ��  �	  �h  �	  ��S  �|  �4  �!	  �8  �T  �   �_     �  �-    �  ��   o  ��   �L �_     �8  ��  ( �
  L#�  	�  W  H�  �  J   = K�    L		  d  M		   �  S   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  (0  O�  #   g)�  	�  �   ��]  =  ��	   L  ��   $  �	  0�  ��   8m  �#"  h�  ��  pآ  �z  tG   �	  x 	�  	  	�  �?  d  �
  �)�  	�  �   H��  �  �_    "  �O  �!  �G   ~	  8fG  �
  h		   (  i		  �� kJ	  �� lJ	    n�  �  o�   �  p�  (�  q�  0 y  s�    �$a  	g  �  0'�  �N  )	   ?1  *		  }0  +	  i/  ,	  � -�	   �  �)�  	�     H�,  ��  �"   ?1  �!	  (  ��  4  ��	  \  ��  0  �_   @ +!  W  tag >	   �U  i	   �  ,  	W  `  S   
�  w%   }#  �&  h  �  &     
j  E   9
  � ;
�   ��  <
2	  �  =
2	  �  >
!	  �#  ?
!	   �  L
(  	�  �  S   �O  :   �   ^$  1  �!  �!   :  �  �  �i	  �#  �t  	z  W	  �  �   I$  ��  	�  �  �   �&  ��  	�  \  �  �  �   	�   �!  H�U  �  �>	   S"  �2	     �U  �"  �J	  �  �J	   ;  �U  (%  �h  0�   ��  8��  ��  @ 	�  R  ��  [  x  =
  H  E#�  y  �  @J   �  L2	   �  M�  �� OZ  .� P�  �  Q�   �  R�  (�!  S�  08'  T  8   W!  	  -  (lT  k  n   �M oT  ߣ  p�  �  q�   	�  k  )f  	l  W	  �     5   w   .�  	�  �      �  1�  	�  �     �  �   	�	  K  6�  	�  �     �   	'  �  :�  	  W	           �  >f  "  Y0  	6  W	  T  �  5  O  �   �  _`  	f  W	  �  �  5  �  �   $  f�  	�  �  �  5  �   �  l�  	�  W	  �  �  >	  i	   #  x�?  �� � [   �  � �  H  � $  P�  � T  X9!  � �  `l� � �  h  � ?  p 	�    ��  �  H2�  �S  4|   �  5p  (  6p  04  7!	  88  8T  @ �  :Q  �  �="  R�  ?�   �  @!	  n  A!	  �  B!	  1$  C�  2�  E�  �� F�  `�L H_   � �  J.  	�  P   @  	F  W	  i  e    	  	  d   �  &u  	{  �     �%  *�  	�  W	  �  �   �%  -�  	�  �  �   {  1�  	�  W	  �  5   �  4�  	�    5   l  8  	  W	  (  �     �  <4  	:  W	  N  �  >	   �  @Z  	`  W	  ~  5  �  !	  z   �  G�  	�  W	  �    !	  !	  p   �'  N�  	�  W	  �    e   �  S�  	�  W	  	    !	  !	  z  	   	J	  &  ���  �� �[   i'  �2	  H   �2	  P  �2	  X�A �4  `Y �i  h�#  ��  p�  ��  x�  ��  �  ��  ���  �N  �U�  �~  ��!  ��  ���  ��  ��  �  �&  �(  � �&  ��  	  �>  �'   'O  ��   xC  �U   s/  ��  '   �  0t�   �  vi	   a   wi	  �'  xi	  !  yi	  �#  zi	   �  {i	  ( �  }8   �  U'�   	�   m  D   t!  �  v2	   A  w2	  �  x2	  &  y2	   !  {�   �  �!  	!  W	  8!  �   !	  8!   	
  �  �J!  	P!  `!  �   8!   �'  �l!  	r!  W	  �!  �   !	  �  �!   	!  �!  �!  ��  )!   ��  )>!  �  )`!   }  �!  �!  O  ;"  _� =%"   ݰ  >%�    	�!  �  @�!  	"  cA  �,1"  	7"  /  �_"  �� ��   �M �_"   ?<  �,k"  	#  �5  P�#  �  �>	   �� �#  �Y �8#  �H �U#  U@ �{#   �9 �#�#  (�A  �#�#  0�^  �#$  8�^  �#($  @N7  �#S$  H q"  ��  �7"  (Z  �#  	$#  W	  8#  %"  i	   17  �D#  	J#  U#  %"   �G  �a#  	g#  !	  {#  %"  �   %G  ��#  	�#  !	  �#  %"  �#   	�  �@  ��#  	�#  !	  �#  %"  %"  �  �   �;  ��#  	�#  �  $  %"  �  �   �W  �$  	$  �#  ($  %"  �   *;  �4$  	:$  �#  S$  %"  �  �   �T  �4$  g�  �q"  	[  �  �  	E  �  �$  @    l  �$  @    	�$  �  �$     	�$  W	  �$    !	  i	  !	   	�$  !	  �$    ]   !�  �%�  �(  S   9�%  x,   �V  �K  *  	�Z  `Y  �,  /+  �N  �O   X  �[  �H  �I  �P  �U  �F  r9   �M  V�%  �\ X�   �  Y�  x  Z		   �7  \�%  �%  �6  `S�&  �<  UJ	   �Q  VJ	  a(  X2	  VA  Y2	  Q) [		   nX  \		  "�D  ^�&  (�5  _�&  8M   a�  H}  b�  JV  c�  L/  d�  N7K  f		  P>D  g		  R�:  i�  T�3  j�  V=]  k�  X 2	  �&  @    �5  m�%  �Q  8��'  �  �J	   �Z  ��  %?  ��  
L/  ��  �<  �		  �Y  ��  �7  ��  �)  ��  �O  ��  �H  ��  vH  ��  ^  ��'  �>  ��  $�7  �		  &0>  �_   (�+  �_   0 �  �'  @    �H  ��&  �?  8A�(  �  CJ	   �Z  D�  %?  E�  
L/  F�  S.  H		  �W  J�  �W  K�  C  L�  �O  M�  �H  N�  vH  O�  ^  Q�'  �>  S�  $�B  T		  &0>  Z_   (�+  [_   0 �]  ]�'  �B  �|�*  ��  ~		   �)  �  �)  �		  �.  �		  U  �		  �V  ��  
�0  ��  �6  ��  �C  ��  U?  ��  6P  ��  �C  ��  &L  ��  *J  ��  �L  ��  HP  ��  N*  ��*   [2  �>	  0k2  �>	  8.  �>	  @{2  �>	  HQ2  �+  P�0  �		  Tp4  �		  VmU  �		  X�Z  ��  Z ?  ��  \:  ��  ^�I  �		  `E8  �		  b�;  �>	  h�;  �>	  p�O  ��  xDF  ��  zfV  �		  |�9  �		  ~[9  �		  ��G  �		  �zQ  �		  � �  +  @   	 �  +  @    {D  ��(  �1  @��+  �I  �J	   6Y  �J	  �^  ��  S  ��  )  �>	  @3  �>	   �0  �>	  (4C  �>	  0�C  �>	  8 aM  �$+  �I  @��,  �  �J	   _7  �>	  )  �		  �O  �		  �n �		  �T  �		  EF  �		  I  �		  �K  ��,  N:  ��,  ,L  ��,  4�E  ��  :�Z  ��  ;�Z  ��  <^  ��  = �  �,  @    �  �,  @    �  �,  @    eU  ��+  �9  (7�-  ��  9J	   a@  :		  b<  ;		  
8  <		  .  =		  �H  >		  �Q  ?		  X  @		  �.  A		  �;  B		  ))  C		  eH  D		  I_  E		  �B  F		   !3  G		  " �)  I�,  �(  S   e.  �-   �D  �1  yA  �>  5  �L  }N   KK  q�-  	2	  �  IV.  F@ K]   I�  L2	  K�  M2	   ԃ  O!.  �b  hh�.  `h  j!	   m�  k!	  dh  l�.   V.  �.  @    ��  nb.  �j  0�/  F@ �]   I�  �J	  def �J	  K�  �J	  tag �>	   c  �!	  ( )�  ��.  �  �P/  �  �	   c  �!	  Cg  �!	   �~  �/  z�   ��/  `h  �!	   m�  �!	  L�  �!	  dh  ��/  e  ��/   	/  	P/  J�  �\/  �R   F0  tag H>	   ��  IJ	  .� J2	  �P  K0   	>	  DG  M�/  T cs0  �^  e>	   [>  f		  �Q g		  
�N h		  0R i		  x  k>	   �I m0  �L m�0  	0  f3   ��0  Tag �>	   Q  �>	  .*  �>	  �K  �>	   �J ��0  gW  ��0  	�0  zC X��1  ��  �>	   �O �>	  ss  �>	  [>  �		  ݖ �		  iA �>	   �y  �		  (�O �		  *rF �>	  0�; �>	  8�U �>	  @�? �>	  H�G �>	  P �F ��0  P 0�2  Tag �>	   .*  �>	  }W �>	  �U �>	  Q  �>	   qY �>	  ( �S �2  	�1  �^   �2  k@  		   aE  		  p0  		  �>  		  H  		  �/  >	  �� �2   	�  �2  �F  "2  9  �2  	"2  �<  0�2  H  2		   �/  3>	  �� 8�2   qS  :�2  2R  :3  	�2  A9  0U�3  ߣ  W		   �E  X!	  �^  Y!	  =Y Z�3  <  [!	  �=  \�3   Jy  ]e  ( 	�2  	�2  rY  _3  ;J _�3  	3  �1  ~�3  �.  �		   �L  �		   Z  ��3  	�3  �V  �+4  ��  �		   f>  �		  Y  ��3   �)  ��3  ��  ��4  �  �		   ��  �		  ~  ��  �  ��  �  �		  5  ��  
B  ��  �  �		   �w  �84  !T ��4  	84  �A  /�5    1�   �  2�  �N  3�  o=  4�  D4  5�  �^  6�  `*  7�  �0  8�  �G  9�  �D  :�  	I:  ;�5  
 �  �5  @    �@  =�4  			  �\  �6  +  ��5   Y�  ��5  �
  ��  (  ��  �F  ��  �C  ��   <)  �6  	�5  �,  `6  �  		   AK  		  z8  �5  V `6   	f6  	�  �R  6  �W �6  	6  	F  .�6  �  0		   �P  1f6   ">  3�6  �W 3�6  	�6  "I�6  #�K Kl6  #`B L�6   �[   E'7  �z  G�   =Y N�6   �6  P�6  �S PA7  	�6  O]  a!T7  	Z7  �(  7N  (��7  >) ��2   -N  ��2  V` ��2  TE  �>	  �/  �!	   �z  ��  $ G  �_7  7[ ��7  	_7  &8  � �7  	�7  eS  poI<  �� qo   ^  s0  � �^  u>	   [>  v		    �W  w�0  ( � y�&  0 �=  z�'  � �,  |�-  � ��  ~�  � �(  �(  � AK  �		  0 XL  ��3  8$os2 �+  h p�  ��+  � T  ��2  0 #9  �>	  8 !H �/>  @ �+  �`>  H @.  ��>  P �E  ��>  X �P  ��>  ` @  ��>  h $S  �_   p s  �_   x$mm �_   �$var �_   � Q  �_   � <B �+4  � 2Y ��,  � =  �>	  � =  �6  � UV  �'7  � �(  �>	   =  ��2    /:  �>	  ( �?  ��2  0 �]  �>	  8$cvt �?  @ �R  �I<  H 5$  �Y
  P ��  ��  ` HT  �>	  h �*  �>	  p �J  ��  x �+  ��  y �  �G7  � �C  ��  � �-  ��  � j7  �!	  � kN  �>	  � �F  �>	  � #7  �>	  � �(  ��2  � rE  ��2  � QZ  �>	  � 4  �!	  � �@  �>	  � :L  ��2  � �G  ��2  � �]  �>	  � �W  �?  � �/  �!	  � �B   ?    �I  �2   s-  >	   �*  !	   ,  �   ,  �   $bdf 	�7  ( �T  >	  P #F  >	  X �U  >	  ` �K  >	  h �=  �V<  	\<  W	  k<  _    �Q  �"x<  	~<  �\  xc/>  �  e�7   �  f�?  )�  g5  �V  h"  :1  j>	   �^ k!	  (Jy  me  0�  n	  8�  p�  <�!  q'  @R0  r	  `�  s	  duN t	  h6  u�  lpp1 v�  ppp2 w�  �2�  z�?  �Xc  {�?  � �6  }�?   )  ~�2   �8  >	    �L �_   ( C  �	  0 ��  �	  4$pp3 ��  8$pp4 ��  H y�  ��2  X �� ��2  ` U  ��
  h �I  �<>  	B>  W	  `>  �7  >	  e  0    1  m>  	s>  W	  �>  k<  !	  >	  !	   �M  +�>  	�>  W	  �>  k<   �<  :�>  	�>  �>  k<   y*  S   =?  4   �^  J  b8  �T   lK  H�>  	�  	!	  |T  @?�?  R�  A�   �  B		  n  C�  
Z�  D		  �  E�  org Gp  cur Hp  ��  Ip   s  K�2  ([  L�5  0c+  N		  8 R8  P?  RG  T'�?  	�?  [  O  _ �?  	�?  LL  Y�  E@  	@  W	  7@  e  �7  	  	  d   ��  k@  �y  �O@  	U@  `@  �7   �m  �l@  	r@  W	  �@  �7  >	  2	  �2  0   t�  "�@  	�@  W	  �@  �7  >	  !	  !	  e  �@  �@   	�  	�4  ن  @�@  	�@  W	  A  �7    0   �}  ZA  	 A  W	  9A  �7  >	  9A   	G  kp  sLA  	RA  W	  kA  �7  !	  kA   	]  T�  �~A  	�A  W	  �A  �7  e  �   �m  ��A  	�A  �A  �7  �  !	  ?  �5   1z  ��A  	�A  W	  �A  �7  		  kA   �a  �B  	B  �  ,B  �7  		  ,B  ,B   		  sz  �?B  	EB  W	  YB  �7  e   �w  O@  �m  !sB  	yB  	  �B  �7  !	  !	   3b  �2SD  !H 4"/>   �A 6"@  �M 7"7@  Y 8"C@  ��  9"�   K ;"`@  (�; ?"2B  0|G @"qA  8H A"2B  @"I B"2B  H�Y C"2B  P�Z D"2B  X�S F"2B  `�< G"YB  h�9 J"2B  p7B L"2B  x-Y M"2B  �(K Q"2B  �Z S"�@  ��i  V"?A  �s  W"YB  �U�  \"fB  ��@ b"2B  �x> c"qA  ��j  e"2B  ��w  f"YB  ��V h"�@  ��= i"A  ��D k"�A  �tW m"�A  ��9 n"�A  � ��  p�B  SD  ~c  trD  	SD  
�'  g  S    ��F  �>  �B XS ;S sX �X @: g; B cD 	�J 
�A $V /L �F M �H �> �T �Z R �;  ^9 !�E "�O #�P $o: %< &'N '�R (:U 0X 1Q @W APW Q�C R�D S�= TLL U�B VG W�X X'P `EF aaT b�E c�T p@M �O ��> �? ��L ��N ��: �YP �WG �U= �aM ��M �G; �2O ��H �3H �2K ��S �GD ��U ��> ��Z �c[ ��T ��[ �zT ��Y ��< ��Q ��Z �fR �EA ��J �nV �.> ��V �<R ��P �wH ��? ��= ��G �>Y �2; ��? ��A ��R � $ S   !J�F  D$  � n% �"  �# !Q�F  � !v$G  � !x�F   u !~$G   %!yRG  C0 !z�  �  !{z  �$ !|�   �# !��F  �$ " jG  	pG  W	  �G    �G  �G   	�  �  "%�G  	�G  W	  �G    �  �G   	RG  �( "*�G  �G  ,& "*�G  6' ",^G   z+ "-�G   �]  #*.H  	ZH  J>  X#XZH  �P  #Z3   2�  #\�  @�� #]�  H�D  #^�H  P� #_W	  T H  \4  S   #F�H  �C    ]  �]   RU  #L_H  AZ #aH  &I  $:�H  �8  $<>	   ߣ  $=2	   `K  $?�H  'B  $C�H  	�H  W	  �H  �  �H   	�H  �  $GI  �H  b:  $G(I  '�  $I�H    �: (%"]I  
H %$#   �U  %%�2  ?1  %&	    �? %((I  �: %(uI  	(I  �Z %*,�I  {I  {I  	�I  |= h%1�I  �M %3_$   ߣ  %4!	  P|Z %5�I  X'�  %6�H  ` �I  L %.�I  	�I  W	  J  �2  �G   > %8�I  J  %X `%�=J  �I %��H   �  %�!	  X �U %�J  =J  J %�ZJ  	J  
�R %�-J  f.  &&�$  <B  &,�$  %�  &0�J  �J  �3  &0�J  tW &2!lJ   i�  &3!xJ   FO  ')�$  ��  ',�J  �J  Y  ',�J  6 '.�J    �Q  ((K  	K  W	  *K    >	  2	  �2  0   �+  (26K  	<K  _   PK    .   �7  (:\K  	bK  W	  �K    !	  0  0  0   �W (A�K  �K  �Y  (A�K  $\  (C�J   �5  (D*K  �A (EPK   ��  )'�K  	�K  W	  �K    �K   	�.  jd  )+L  		L  W	  L    L   	#L  	�/  �g  )/5L  	;L  W	  TL    !	  .   �{  )6`L  	fL  W	  L    !	  	    l  )=5L  �n  )B`L  �x  )G�L  	�L  W	  �L    !	   1j  )K5L  �}  )P�L  	�L  W	  �L    ?  �L  �L  L   		  ��  )Wu  �b  P)Z�M  h  )\�K   �v  )])L  ��  )^L  ��  )_�L  .�  )`�K   �  )aTL  (V�  )b�L  0��  )c�L  88�  )f�L  @��  )gM  H M  h�  )Z�M  	�M  &�? ��K  	��H     &�X ��J  	��H     �  �M  @    �M  &F ��M  	��H     oJ �N  	!N  G   0N  G    �   @N  @    0N  '�P �@N  	��H     '*W ,�J  	x�H     '�V 6I  	p�H     'JN c�G  	`�H     3   �N  @    �N  '"C s�N  	 �H     '�9 �`D  	 �H     (xD  �	��H     ��  *#O  	O  �  O  �   d�  *)#O  	)O  �  8O  !	   0�  */#O  K�  *6lO  �> *8�   �^ *9!	   �  *;DO  Ѽ  *>$�O  	�O  ў  (*@�O  
H *B#   ��  *C!	  XT *D�O    	lO  ��  *N�O  	�O  �  �O  i	  !	   B�  *V�O  	�O  P  i	  �   ��  *ZP  	P  W	  GP  �  xO  !	  �O  �O  i	   ��  *bSP  	YP  !	  mP  xO  �   ��  *fyP  	P  �  �P  xO  �#   ��  @*j	Q  �\ *l �N   8` *n P  �\ *o GP  �_ *p mP  �T *r O   }�  *s 8O  (ʬ  *t  Q  0�  *u  Q  8 �P  ��  *jQ  		Q  	u  i  +'2Q  	8Q  W	  QQ    !	  ,B   4�  +,2Q  \�  +12Q  �l  +82Q  ~�  +=2Q  ŋ  +B2Q  �w  +G2Q  H�  +Nu  ȅ  @+QR  ��  +S&Q   ��  +TQQ  �n  +U]Q  Rs  +WiQ  ��  +XuQ   F}  +Y�Q  (�|  +Z�Q  0��  +\�Q  8 �Q  w�  +Q,R  	R  4< }>R  	DR  ]  XR  �2  �   )�; �J  	 �H     *D NJ  	��H     $@ P�S  
H �]I   VH ��  (Z: �!	  ,5�  �!	  0)c  �!	  4H �!	  8�E �!	  <u~  �	  @U ��2  H �> �S  	�R  *)G J  	 �H     *�9 �J  	��H     *�R �J  	 �H     *EP }J  	��H     �Y P��S  
H �]I   pw  ��  (VH �>	  0Z: �!	  8= �>	  @�@ �>	  H +? ��S  	�S  *MJ �	J  	 �H     
B P
qT  
H 
]I   pw  
�  (VH 
>	  0Z: 
!	  8= 
>	  @�@ 
>	  H @ !
~T  	T  *cH 'J  	��H     �W H~�T  
H �]I    Z �>	  (>V ��  0L[ ��#  8R�  ��  @ @ ��T  	�T  *b<  J  	 �H     +`J  �	��H     �I  =U  @   	 -U  '�V �=U  	@�H     �: X�V  �  ��7   Jy  �e  �I ��@  N ��4  ~I ��   )= ��  !�F ��  "�U  �>	  (�K  �>	  0�N �>	  86X �>	  @�C ��2  H.Z ��2  P UC �YU  T[ �8V  	YU  jB �KV  	QV  W	  yV  +V  �2  �2  	  	  !	   ,Z :W	  P%D     +      �R[  -�  :1�7  �Q	 {Q	 --U ;1>	  R	 �Q	 -�^ <1!	  �R	 �R	 -:1  =1!	  rS	 dS	 -Jy  >1e  $T	 T	 .map ?1�@  U	 �T	 /N @1�@  � 0� BW	  �U	 �U	 1x'D     !      jX  '�3 JR[  ��~2Ui  x'D      x'D            M5X  3�i  �V	 �V	 3�i  �V	 �V	 3ti  kW	 iW	 3gi  �W	 �W	 4x'D            5�i  �W	 �W	 5�i  #X	 X	 6�i  �(D     7�i  %(D     S       X  5�i  |X	 pX	  8�'D     � 9U|    8�(D     h\  9U��~9T} 9Q09R09X09Y~ F%1  : 	Y  '�D r�  ��~0k  s  Y	 Y	 ;�(D     � �X  9U��~ ;�(D     � �X  9U| 9T 9Q��~9R1 ;�(D     � �X  9U| 9T��~ <d)D     �  =b[  �%D      � ]3�[  RY	 PY	 3�[  wY	 uY	 3�[  �Y	 �Y	 3�[  Z	 �Y	 3�[  yZ	 sZ	 3�[  �Z	 �Z	 3t[  *[	 "[	 >� 5�[  �[	 �[	 5�[  �\	 �\	 5�[  �\	 �\	 ?�[  ?\  5\  ]	 ]	 5\  t]	 j]	 5*\  ^	  ^	 57\  _	 _	 6B\  �&D     ;&D     � 
Z  9U|  ;&D     
 'Z  9U| 9T8 ;+&D      ?Z  9U|  ;6&D      WZ  9U|  ;A&D     $ oZ  9U|  ;�&D     � �Z  9U|  ;�&D     
 �Z  9U| 9T ���� ;�&D     1 �Z  9U|  ;�&D     1 �Z  9U|  ;�&D      �Z  9U|  ;�&D     1 [  9U|  ;�&D     $ #[  9U|  ;s'D     $ ;[  9U|  8)D     $ 9U|     V  b[  @     @}F �W	  h\  A�  �1�7  A-U �1>	  A�^ �1!	  AJy  �1e  Bmap �1�@  AN �1�@  A��  �1�  CXR �!	  C��  �!	  C��  �+!	  CE> �	  CS> �	  C�@ ��  C=? �	  C� �W	  Dp ��2  E|N �FCS )�  CD�  *		    ,�P �W	  @�C     (      �na  -�3 �/+V  �_	 �_	 -�^ �/!	  �`	 �`	 -�s �/	  �a	 �a	 -��  �/	  Xb	 Jb	 -Q�  �/!	  �b	 �b	 -��  �/�  �c	 oc	 Gp ��2  ��03o  ��2  dd	 `d	 05�  �>	  �d	 �d	 0�S �!	  /e	 e	 Hend �!	  �e	 �e	 0�X �!	  �f	 �f	 0�? �)!	  rg	 Zg	 0�S �>	  di	 Pi	 0�S � >	  Oj	 7j	 0<G �/>	  Uk	 Mk	 E��  �I�K �C     I�9 ���C     :`�  ?^  '�C ->	  R8��C     &h  9Uu 9Tt 9Q 9Rr   :��  �^  Hmm K>	  l	 l	 '�  K>	  T>��  0n�  Z!	  jl	 ^l	   :P�  _  C�C o>	  Hmm o>	  ]m	 Wm	 0�  o#>	  �m	 �m	 :��  �^  0n�  �!	  �m	 �m	  88�C     &h  9Uu 9Tt 9Q 9Rr   =na  �C      0�  �3�a  o	 o	 3�a  po	 jo	 3�a  �o	 �o	 3�a  p	 p	 3�a  [p	 Wp	 J�a  J�a  3�a  �p	 �p	 >0�  5�a  q	 q	 5�a  �q	 �q	 Kb  ��5b  6r	 0r	 Kb  ��6'b  �C     60b  /�C     L9b  ��  �`  5:b  �r	 r	 LGb   �  /`  5Hb  �r	 �r	 5Ub  Cs	 As	 5bb  ps	 fs	 5ob  t	 t	  M�h  z�C      0�  ��`  3�h  >t	 :t	 3�h  xt	 tt	 >0�  5�h  �t	 �t	 5�h  +u	 u	 5i  v	 v	 5i  �v	 �v	 5"i  �v	 �v	 6/i  /�C     <��C     >   N��C     9Uv 9Qs 9R} 9X~ 9Y|   ;5�C     � a  9U  ;M�C     K ,a  9U 9Ts 9Q�� ;@�C     X Ka  9U 9T�� 8K�C     &h  9Uu 9Tt 9Qs     @�B QW	  b  A�3 Q0+V  A�  R0!	  A��  S0>	  A�  T0>	  A�s U0	  A��  V0	  AQ�  W0!	  A��  X0�  C� ZW	  CJy  [e  Dp \�2  C3o  ]�2  C�U  ^�2  E�u  �E�0  �FC��  � >V  FC��  �!	  C�  �!	  C�Q �!	  C�D �!	     ,�K �W	  p�C     K      �ed  -�3 �2+V  w	 	w	 .p �2�2  ~w	 pw	 -�� �2�2  x	 x	 -�s �2	  ^x	 Vx	 -��  �2	  �x	 �x	 -Q�  �2!	  ,y	 $y	 0� �W	  �y	 �y	 0:= �!	  �y	 �y	 Hnn �!	  1z	 -z	 0~  ��  kz	 iz	 0�  ��  �z	 �z	 0�  ��  �z	 �z	 05  ��  �z	 �z	 0B  ��  {	 {	 0�  ��  8{	 6{	 I�0  ��C     I�u  ��C     4�C     =       0n�  �!	  a{	 _{	 Gdx ��  QHdy ��  �{	 �{	 8R�C     h\  9Us 9Xv 9Y0   ,AQ QW	  ��C     �      �7f  -�3 Q5+V  �{	 �{	 .p R5�2  $|	 |	 -�� S5�2  �|	 �|	 -�s T5	  _}	 M}	 -��  U5	  %~	 ~	 -Q�  V5!	  �~	 �~	 O� XW	   0+ Y�2  �~	 �~	 0�  Z	  s	 i	 0��  Z	  �	 �	 0�  Z	  y�	 g�	 0�S Z'	  ��	 z�	 Hh Z2	  *�	 �	 0UO Z5	  Ƃ	 ��	 0�L [!	  ��	 ��	 0Q [!	  ă	 ��	 0�I \�@  �	 �	 0�P ]		  \�	 H�	 I�u  ��C     >@�  0�@ ��2  =�	 +�	 Hw �	  �	 ��	   ,�U �W	  ��C     -      �&h  -�3 �6+V  ��	 ��	 .p �6�2  +�	 !�	 -�� �6�2  ��	 ��	 -�s �6	  A�	 1�	 -��  �6	  �	 ��	 -Q�  �6!	  ��	 ��	 O� �W	   0+ ��2  ى	 ˉ	 0�  �	  t�	 p�	 0��  �	  ��	 ��	 0�  �	  �	 ��	 0�S �'	  g�	 c�	 Hh �2	  ��	 ��	 0�L �!	  \�	 X�	 0Q �!	  ��	 ��	 0�I ��@  �	 �	 I�u  &ߨC     :��  �g  0�@ ��2  8�	 2�	 Hw �	  ��	 ��	  >�  0�@ 	�2  ��	 ��	 Hw 
	  /�	 -�	 0�< !	  h�	 R�	   ,�M �W	  �C     �       ��h  /�3 �1+V  UPpp �1�h  T-�� �1�2  U�	 O�	 Pbig �1�  RHp ��2  ��	 ��	 0N ��4  #�	 !�	 E�0  � 	�2  @�I 1W	  9i  A�3 11+V  A��  21�  C� 4W	  C��  5!	  C�  5!	  Dmap 6�@  C�  7>	  E�u  z Q�B *Ui  A�3 *)+V   @2D �W	  �i  A�3 �.+V  A�  �.�7  A-U �.>	  AN �.�@  C� �W	  CJy  �e  E�u  $FDp �2    ,�=  W	  ��C     )      �ol  -�   2�7  O�	 G�	 --U !2>	  ��	 ��	 -N "29A  �	 �	 :��  �j  0�V :�2  ��	 ��	 0�; ;�  ��	 �	 03: <�  d�	 Z�	 ;��C     e �j  9T@B$ 8
�C     e 9T@B$  >��  0Jy  �e  ޒ	 Ԓ	 Cx  �!	  0EN �		  Q�	 O�	 0:� �		  x�	 t�	 C��  �%		  0+  �ol  ��	 ��	 0�J ��  ؓ	 ֓	 0� �W	  �	 �	 Hp ��2  ~�	 z�	 ;�C     � mk  9U}  ;-�C     
 �k  9U} 9T4 ;��C     1 �k  9U}  ;��C     1 �k  9U}  <��C     $ ; �C     e �k  9T} 9Q~  ;�C     e l  9T} 9Q~  ;B�C     e !l  9T} 9Q~  ;X�C     e ?l  9T} 9Q~  ;q�C     e Xl  9T@B$ 8��C     e 9T@B$   	�'  ,�V W	  ��C     
       � m  -�  -�7  ̔	 Ȕ	 .req -  	�	 �	 -,U -0  H�	 B�	 R��C     r 9U�U9T�T9Q09R�Q  S�U 
��C     /       �_m  -�  
�7  ��	 ��	 0Jy  e  �	 �	 8ǯC     X 9Ts�	  Tj= 2W	  ��C     �      �q  U�  2!�7  �	 �	 UJy  3!e  ~�	 t�	 V� 5W	  �	 �	 &x-  6>	  ��V�q  7>	  ��	 �	 W�u  �:@�  [n  Xp b�2  ؘ	 Θ	 V��  cJ	  ^�	 X�	 V�/  d>	  �	 �	 V.� e!	  ��	 ��	 8'�C     K 9Uv 9Q|   :�  �o  V��  �		  ��	 ��	 V?1  �		  �	 �	 V�/  �>	  Z�	 T�	 V.� �!	  ��	 ��	 ;��C     
 �n  9Uv 9T8 ;��C     1 �n  9Uv  ;��C     1 o  9Uv  ;��C      o  9Uv  ;��C     $ 1o  9Uv  ;1�C      Io  9Uv  ;=�C     � ao  9Uv  8c�C     K 9Uv 9T~ 2$#����9Qs�	  :p�  9p  &�K  �>	  ��Y0�C     �o  9Us 9TTDBC9Qv 9R�� YJ�C     �o  9Us 9TTDBE9Qv 9R�� Yd�C     $p  9Us 9Ttadb9Qv 9R�� 8��C      9Uv   Y�C     cp  9Us 9TCLBC9Qv 9R�� ;W�C     X �p  9Uv 9T|  ;��C      �p  9Uv  Y��C     �p  9Us 9TCLBE9Qv 9R�� Y��C     �p  9Us 9Tcolb9Qv 9R�� N��C     9Us 9Txibs9Qv 9R��  @�G 	�W	  �q  A�  	�%�7  Bidx 	�%!	  AD@ 	�%kA  C� 	�W	  C=Y 	�47  Cߣ  	�J	  Cs  	�Q  ZEnd 	3[�q  C>) 	y6  FCi�  			    FC>) 	#�6    S�C 	� �C           ��r  -�  	�#�7  �	 ݛ	 0R�  	��  F�	 D�	 0=Y 	�47  s�	 k�	 0ߣ  	�J	  �	 ޜ	 1p�C     �       �r  0>) 	�y6  /�	 -�	 Hn 	�		  ]�	 U�	 ;�C     � �r  9U}  ;��C     � �r  9U}  8��C     � 9U}   4 �C     (       0>) 	��6  ��	 ��	 8�C     � 9U}    ,�< 	~W	  �D     n      ��y  -�  	~�7  ��	 �	 0Jy  	�e  :�	 ,�	 0� 	�W	  �	 ϟ	 0ߣ  	�J	  ��	 ��	 'H< 	�>	  ��0y? 	�>	  ��	 �	 I�u  	�oD     M5z  �D      `�  	��w  3^z  ��	 ��	 3Rz  9�	 -�	 3Fz  ˢ	 ��	 >`�  5jz  ��	 ��	 Kvz  ��5�z  أ	 У	 5�z  c�	 U�	 5�z  �	 �	 5�z  ѥ	 ��	 6�z  �D     6�z  �	D     \�z  L�z  ��  �t  5�z  6�	 2�	 ;�D     � �t  9U~ 9T29Q09R 9X09Y�� ;�D     
 �t  9Uv 9T 1$ ;<D     1 �t  9Uv  ;aD     $ �t  9Uv  8G
D     $ 9Uv   L�z  ��  <u  5�z  r�	 n�	 ]�z  pD     %       5�z  ��	 ��	   L�z  0�  �v  5 {  
�	 ��	 L
{  ��  Cv  5{  ��	 ��	 L{  ��  �u  5{  ^�	 Z�	 8�D      9Uv   ;D      �u  9Uv  ;4D     � �u  9U~ 9T19Q09R}����9X09Y�� ;UD     � v  9Uv 9Q}  ;�D      'v  9Uv  8�D     � 9Uv 9T��  ;�D     � ~v  9U~ 9T89Q09R	���
��9X09Y�� ;`
D     � �v  9U~ 9T89Q09R09X09Y�� 8�
D     � 9U~ 9T19Q09R19X09Y��  78{   
D            w  59{  ��	 ��	 80
D     � 9U~   7%{  w
D     0       Cw  5*{  ��	 ��	  ;�D     � bw  9Uv 9T�� ;�	D     � �w  9U~ 9T�� 8�	D     � 9U~ 9T��   M�y  �D        	�)y  3�y  �	 �	 3�y  �	 �	 3�y  O�	 K�	 >  5�y  ��	 ��	 K�y  ��5�y  Ū	 ��	 5�y   �	 �	 6�y  	D     6�y  �	D     7z  s	D     G       ox  5
z  ��	 ��	 ^z  @  5z  �	 �	   7%z  �
D            �x  5&z  c�	 a�	  ;�D     � �x  9Uv 9T�� ;;	D     � �x  9U} 9T19Q09R��~9X09Y�� ;c	D     � y  9Uv 9T��~9Q�� 8�	D     � 9U}    YD     Sy  9Us 9Ttsop9Qv 9R�� ;0D      ky  9Uv  8LD     � 9Uv 9T   @[B 	;W	  5z  A�  	;�7  AJy  	<e  Ay? 	=>	  CR�  	?�  C� 	@W	  C�  	B	  C�X 	Cf6  E�u  	xE�0  	u[%z  Dn 	Z	  FDidx 	_2	    FC>) 	l�6    _�K 	�W	  F{  `�  	��7  `Jy  	�e  `y? 	�>	  aR�  	��  a� 	�W	  a�  	�	  aAK  	�		  az8  	��5  aTT 	�`6  E�u  	5E�0  	1E��  	([�z  bn 	�	   [�z  bn 	�	  Fbidx 	�	    [%{  bn 	�		  Fblen 	�!	  Fbd 	�	     [8{  C>) 	y6   FDn 	*		    c{D �0�C     �      ��}  U�  �$�7  ��	 ��	 U�(  �$�  ��	 �	 Un�  �$!	  5�	 -�	 US �$?  ��	 ��	 UD�  �$�5  �	 ��	 &� �W	  ��VJy  �e  ��	 ��	 V� �ol  ߮	 ݮ	 V�P �>	  �	 �	 Vx-  � >	  ԯ	 Я	 V-N  �,>	  �	 
�	 Xk �		  ��	 ��	 Xvar �# R  �	 �	 IB #��C     : �  �|  dv �_   P :P�  #}  Hf +  A�	 =�	 Ga ,	  ��Gb -	  ��Y��C     �|  9Us 9T 9Q�� Y�C     }  9Us 9T 9Q�� NV�C     9Us 9T 9Q��  ;��C     � E}  9U��9T�� ;ĶC     � f}  9U��9T�� ;!�C     � �}  9U�� ;C�C     � �}  9U��9T�� ;l�C     � �}  9U��9T�� ;��C     � �}  9Uw  8ǷC     � 9T��  TtG |W	  ��C     t       �  U�  |!�7  ��	 w�	 UJy  }!e  �	 ��	 U�(  ~!�  ��	 ��	 V� �W	  Ͳ	 ǲ	 V� �ol  �	 �	 &�U �"-  	 �H     e�0  ��C     :�  �~  Xv �_   T�	 P�	 N��C     9Us�|9Taehv9Qv 9R0  ;��C     � 	  9Uv 9T	 �H     9Qs  N'�C     9Taehh  �%  -  @      Tp> FW	  ��C     u       �5�  U�  F!�7  ��	 ��	 UJy  G!e  ��	 ��	 U�(  H!�  v�	 p�	 V� JW	  ȴ	 ´	 Xtag K>	  �	 �	 &x-  K>	  �HVIG L0  n�	 j�	 V�H M0  ��	 ��	 e�0  d�C     Y�C      �  9U�U9Qv 9R�H 8��C      9Uv   ,/B YW	  @�C     B      ��  -�  Y!�7  �	 ޵	 -Jy  Z!e  ��	 ��	 0� \W	  5�	 3�	 0R�  ]�  _�	 Y�	 Hj _!	  ��	 ��	 05�  _!	  з	 η	 0T `�3  ��	 ��	 I�u  �n�C     Yf�C     "�  9Uv 9Tpsag9Qs 9R0 ;��C     
 ?�  9Us 9T4 ;��C     1 W�  9Us  ;��C     1 o�  9Us  ;��C     $ ��  9Us  ;�C     � ��  9U| 9T49Q09R} 9X09Y�L ;%�C     
 ځ  9Us 9T} 2$ ;\�C     1 �  9Us  ;h�C     1 
�  9Us  8y�C     $ 9Us   ,%Y W	  ��C     J       ��  -�  !�7  V�	 J�	 -Jy  !e  �	 �	 '�O "#�  	@�H     0� 7W	  ��	 ��	 02Y 8(�  ��	 ��	 I�u  C��C     Y��C     �  9Us 9TTLCP9Qv 9R0 R�C     � 9U�T9T	@�H     9Q�U#�  �%  #�  @    �  	�,  ,�Z �W	  ��C     J       ��  -�  �!�7  ^�	 R�	 -Jy  �!e  ��	 �	 0� �W	  ��	 ��	 0�Z ��  û	 ��	 ' G �"'�  	��H     Y��C     �  9Us 9Ttsop9Qv 9R0 R��C     � 9U�T9T	��H     9Q�U#�  	�+  �%  '�  @   
 �  @�Y @W	  ��  A�  @ �7  AJy  A e  C� CW	  Dos2 D��  '�S F"��  	 �H     'JV {"�  	��H     '\V �" �  	��H     '�S �"�  	��H     I�u  �XD      	+  �%  ��  @   + �  �%  �  @    ��  �%   �  @    �  @�G W	  p�  A�  !�7  AJy  !e  C� W	  I�u  )�D      S�< �0�C     
      ���  -�  ��7  `�	 Z�	 0R�  ��  ��	 ��	 0>) ��3  ׼	 Ѽ	 1T�C     X       @�  0� ��2  2�	 ,�	 0�� ��2  �	 }�	 ;��C     � %�  9Uv  8��C     � 9Uv 9Ts   4��C     S       0� �3  ��	 ��	 0�� �3  ��	 �	 ;��C     � ��  9Uv  8 �C     � 9Uv 9Ts    ,�S $W	   �C     Z      �A�  -�  $!�7   �	 �	 -Jy  %!e  ��	 �	 '� 'W	  ��0R�  (�  ��	 ��	 0�P )>	  ;�	 5�	 '>k  )>	  ��0wA *>	  ��	 ��	 0�R *">	  �	 �	 0>) +�3  g�	 _�	 '�M -"Q�  	 �H     '1T 9" �  	�H     '%S H"f�  	�H     I�u  ���C     :��  8�  0� �3  ��	 ��	 0�� �3  ��	 ��	 8��C     � 9Us 9T	�H     9Q   :��  ��  0� ��2  :�	 2�	 0.� �!	  ��	 ��	 ;L�C     � ��  9Us 9T	�H     9Q  8��C     � 9U| 9T 9Y��  YR�C     �  9U~ 9Teman9Qs 9R�� ;x�C      ��  9Us  ;��C     � &�  9Us 9T	 �H     9Q~� ;��C     � U�  9U| 9T 9Q09X09Y�� ;�C     
 m�  9Us  ;��C     $ ��  9Us  ;�C     � ��  9Us 9T}  ;,�C     �   9Us 9T�� ;]�C     � ��  9U| 9TH9Q09R 9X09Y�� ;��C     
 �  9Us  ;�C     $ &�  9Us  8�C     � 9Us 9Tv  �%  Q�  @    A�  �%  f�  @    V�  ,I �W	  ��C     �       ���  -�  �!�7  K�	 C�	 -Jy  �!e  ��	 ��	 0� �W	  4�	 &�	 0�< ���  ��	 ��	 'rI �"�  	��H     '�O �"��  	`�H     I�u  ��C     Y��C     I�  9Us 9Tpxam9Q| 9R0 ;�C     � t�  9U| 9T	��H     9Q}  8l�C     � 9U| 9T	`�H     9Q}   	�-  �%  ��  @    ��  , K �W	  @D            �*�  -�  �!�7  @�	 <�	 -Jy  �!e  }�	 y�	 RGD     ��  9U�U9T�T9Qdehb  ,�; �W	  PD            ���  -�  �!�7  ��	 ��	 -Jy  �!e  ��	 ��	 RWD     ��  9U�U9T�T9Qdaeh  @�Q ^W	  �  A�  ^+�7  AJy  _+e  Btag `+>	  C� bW	  C� c�  '� e"/�  	��H     I�u  �D      	�&  �%  /�  @    �  ,�J W	  ��C     �       ���  -�   �7  8�	 0�	 .tag  >	  ��	 ��	 -x   2	  
�	 �	 -B�  �2  ]�	 S�	 -ss    0  ��	 ��	 '� "W	  P0Jy  #e  @�	 <�	 0>) $�0  z�	 x�	 0�  %>	  ��	 ��	 E�u  HM]�  ��C       `�  +z�  3n�  �	 �	 3n�  �	 �	 3z�  R�	 P�	 >`�  5��  y�	 u�	 5��  ��	 ��	   fW�C     � f��C     �  ,�@ OW	   D     �      �j�  -�  O%�7  ��	 ��	 -Jy  P%e  C�	 ;�	 '$S  Rs0  ��'� SW	  ��~0R�  T�  ��	 ��	 Hnn U		  �	 �	 07F U		  l�	 V�	 'N W"z�  	 �H     I�u  ��D     :@ �  0� ��0  l�	 V�	 Hi �		  ��	 ��	 0�B ��  ��	 ��	 ;bD      ȏ  9Us  ;mD      ��  9Us  ;yD      ��  9Us  8�D      9Us   M�  �D      � ~��  3��  �	 �	 3��  �	 �	 3��  G�	 A�	 3��  ��	 ��	 >� 5��  ��	 ��	 5��  �	 �	 5˒  ��	 {�	 5ג  ��	 ��	 5�  U�	 K�	 5�  ��	 ��	 5��  $�	 �	 \�  L&�  � v�  K'�  ��L3�   M�  ?4�  ;�D     � �  9Us  ;D     �  �  9Us 9T��~ 83D     � 9Us 9Tv 
��#4$ $ &w "  8�D     � 9Us 9T	 �H     9Q��  8D     � 9Us 9Tw    ;@D      ��  9Us  ;RD     � ʑ  9Us 9T��~ ;�D     � ��  9Us 9T	 �H     9Q�� ;�D     � %�  9U~ 9T 9Q09X09Y��~ ;�D     � =�  9Us  ;D     
 U�  9Us  8�D     $ 9Us   �%  z�  @    j�  _"D �W	  C�  `$S  �!0  `Jy  �!e  `pw  �!�5  a� �W	  bnn �		  a7F �		  a�; �!	  a[ �!	  a�T �,!	  ax  �>	  &�V �"z�  	 �H     E�u  3Fa>) ��0  Fa�  ��     TH ~W	  �C     V       �]�  U�  ~"�7  ��	 ��	 gtag ">	  ��	 ��	 UJy  �"e  -�	 '�	 Uss  �"0  �	 y�	 V>) ��0  ��	 ��	 a� �W	  e�u  ��C     h]�  �C        �  �G�  3n�  ��	 ��	 3n�  H�	 B�	 3z�  ��	 ��	 > �  5��  ��	 ��	 5��  �	 �	   R+�C     � 9U�Q  _�T 8�0  ��  `�  8#�7  itag 9#>	  a� ;�0  a�� <�0   TK? �	  ��C           �Ȗ  j�  �!�7  UU�U  �!!	  H�	 B�	 UB7  �!!	  ��	 ��	 VE  �	  ��	 ��	 V.� �!	  ��	 v�	 V� �!	  ��	 ��	 Xp ��2  b�	 D�	 V3o  ��2  ��	 ��	 I�C .�C     I�Y (��C     >@�  V2�  ��2  ��	 ��	 V�@ ��2  V�	 T�	 V��  �!	  ��	 y�	 Vss  �!	  k�	 [�	 V*� �!	  ��	 ��	 V�; �!	  ��	 ��	 V�\ �	  	�	 ��	 >��  a�M �>	  :p�  ��  Xmin �!	  ��	 ��	 Xmax �!	  ��	 ��	 >��  Xmid �!	  7�	 -�	 Xq ��2  ��	 ��	 Xkey �>	  I�	 A�	   >�  0+; 
!	  ��	 ��	 >@�  Hkey >	  �	 ��	      krU ��  `�  ��7  aJy  �e   T�9 ,W	  `�C     E      ��  U�  ,!�7  �	 ��	 UJy  -!e  Y�	 M�	 V� /W	  ��	 ��	 &x-  0>	  ��Xp 1�2  X�	 0�	 V3o  2�2   �	 ��	 Xnn 3!	  )�	 #�	 V[>  3!	  x�	 t�	 V�8 4�  ��	 ��	 V�L 4�  �	 �	 e�u  ���C     e�C �`�C     :��  Ә  V�; X!	  \�	 V�	 Vss  X!	  ��	 ��	 V*� X%!	  ��	 ��	 Vߣ  X/!	  -�	 +�	 V,H Y�2  \�	 T�	 V� Z�  ��	 ��	 4�C     [       V.� �>	  �	 �	 V+< �>	  _�	 Y�	 4*�C     /       VV ��  ��	 ��	    Y��C     ��  9Us 9Tnrek9Qv 9R�� 8��C     K 9Uv 9Qs�
  ,Q< NW	  ��C            ���  -�� N#�  =�	 7�	 -+�  O#�H  ��	 ��	 0
H Q%"  ��	 ��	 0�M R{I  1�	 -�	 l��C     9U�U9T�T  ,vQ �W	  ��C           �q�  -�  �!�7  s�	 i�	 0>) ��2  ��	 ��	 0�� ��2  t�	 j�	 '>[ �-	  ��~Gp ��2  ��~0k  �  ��	 ��	 >��  '�� �  ��0x  �  /�	 +�	 >��  '
H (�2  ��~'ߣ  (-	  ��~'�M (w�  ��~'�M (�I  ��~> �  'pw  'IJ  ��'� 'd	  ��~1��C     +       �  '_I )%"  ��~8��C     � 9Q��9R��~  ;!�C      C�  9U��9Qw 9R0 ;>�C      \�  9U�� N��C     9T��     	�I  q�  ,AB �  ��C            ��  -yW +xO  n�	 j�	 -��  �+�#  ��	 ��	 0�  ��7  ��	 ��	 0s  �Q  �	 
�	 l��C     9U�U9T�T  ,�I s!	  ��C            ���  -yW s,xO  8�	 4�	 -��  t,�  u�	 q�	 0�  v�7  ��	 ��	 0s  wQ  ��	 ��	 l��C     9U�U9T�T  S�K g0�C     (       ��  -yW g&xO  �	 ��	 0�  i  R�	 P�	 0R�  j�  x�	 v�	 <G�C     �  ,rK SW	  P�C     &       ���  -yW S&xO  ��	 ��	 -m  T&i	  ��	 ��	 0�  V�7  1�	 /�	 0R�  W�  V�	 T�	 0s  XQ  }�	 {�	 lv�C     9T�U9R	pD     9X0  ,�= F�  pD     (       ���  -�  F�7  ��	 ��	 .idx G!	  ��	 ��	 'D@ I]  �hmq  tD       tD            L3@q  "�	 �	 33q  s�	 o�	 3&q  ��	 ��	 4tD            ?Mq  ?Zq  ?gq  ?tq  \�q  8�D     � 9U�U9T�T9Q�h    ,�G ��#  @�C     P      ��  -
H �'iI  ��	 ��	 -R�  �'�  �	 ��	 -X6  �'�  ��	 ��	 Hp ��2  b�	 >�	 Hi �	   �	 ��	 0 P �>	  c�	 _�	 0P �>	  ��	 ��	 :��  �  0�W ��T  ��	 ��	 0f>  ��  s�	 o�	 0fI ��  ��	 ��	 0N ��  ��	 ��	 0�W ��  9�	 +�	 0QH ��  ��	 ��	 Hdp ��2  V�	 H�	 Hdi �!	  ��	 ��	 Hni �!	  !�	 �	 Hk �!	  ��	 ��	 Hret ��#  ��	 ��	 M"�  ��C      @�  ���  34�  ��	 ��	 >@�  5?�  &�	 "�	 5L�  ��	 ��	   ;��C     ��  ��  9U 9Q�T n/�C     С  Ӡ  9U�U9Q�T Rd�C     �  9U�U  8c�C     ��  9Uu 9Tt   ,�< {�#  ��C     �       �С  -
H {+iI  �	 ��	 .p |+�2  ��	 ��	 -R�  }+�  ��	 ~�	 0�W �T  ��	 ��	 CfI ��  Hi �!	  S�	 O�	 Hret ��#  ��	 ��	 8ƺC     ��  9U| 9Ts9Q�Q  ,�K V�#  йC     �       �"�  -
H V'iI  ��	 ��	 .p W'�2  ��	 n�	 -R�  X'�  N�	 F�	 0�W Z�T  ��	 ��	 0f>  [�  _ 
 Y 
 Hcnt \!	  '
 !
 Hq ]�#  �
 z
 10�C     6       ��  Huni h�  �
 �
  M"�  ׹C      ��  `��  34�  (
 
 >��  5?�  �
 �
 5L�  O
 I
   ;�C     ��  �  9U|  8��C     ��  9T1  @,A D!	  Z�  Bp D'�2  Cf>  F�  Dtot G!	   ,�P �#  ��C           ���  -
H 'iI  �
 �
 -R�  '�  
 
 -�@  '�  c
 S
 0�W "�T  
 
 0.� #�  y
 u
 Hp $�2  �
 �
 Hq %�#  }
 q
 :��  ��  0?C -�  
 
 0 P .>	  w
 q
 0P />	  �
 �
 ;�C     -�  r�  9Uu 9Tt  8w�C     c�  9Uu 9Tt   8��C     ��  9U| 9T}9Q�T  ,gC �#  ��C     �       ���  -
H "iI  )
 
 -R�  "�  �
 �
 0�W �T  	
 	
 0.� �  �	
 �	
 Hp 	�2  �	
 �	
 0E  
�#  �

 �

 Hi �  �

 �

 8��C     ��  9U| 9Tv9Q�T  ,|R �	  ФC     x       �y�  -
H �,iI  
 	
 -�j �,�  T
 F
 -X6  �,�  �
 �
 Hp ��2  s
 k
 0 P �>	  �
 �
 0P �>	  %
 
 ;�C     ��  @�  9Uu 9Tt  ;�C     c�  ^�  9Uu 9Tt  8=�C     -�  9Uu 9Tt   ,�9 �!	  @�C     �       ���  -
H �(iI  �
 �
 -�W  �(iI  �
 �
 -�j �(�  �
 �
 -X6  �(�  L
 B
 Hp ��2  �
 �
 0 P �>	  
 
 0P �>	  d
 ^
 ;^�C     ��  K�  9Uu 9Tt  ;��C     -�  i�  9Uu 9Tt  o��C     ~�  9U�T RȤC     c�  9Uu 9Tt   ,�W ��2  ��C     �       �c�  -2�  �'�2  �
 �
 /I= �'�  T0; ��  
 
 Hmax ��  Y
 K
 Hmin ��  
 
 >�  Hmid ��  X
 N
 Hp ��2  �
 �
 0?C �>	  x
 p
   ,�C �!	  �C     �       �-�  -2�  �1�2  �
 �
 /��  �1�  T0fI ��  5
 3
 Hmax ��  �
 }
 Hmin ��  
 
 >��  Hmid ��  `
 V
 Hp ��2  �
 �
 Huni ��  r
 j
   ,;I b!	  @�C     �       ��  -2�  b.�2  �
 �
 /��  c.�  T0f>  e�  
 
 Hmax f�  g
 Y
 Hmin f�  %
 !
 >��  Hmid q�  f
 \
 Hp r�2  �
 �
 0�S s>	  �
 �
 Hcnt t!	  O
 K
   ,TU TW	   �C            �N�  /
H T%iI  U/+�  U%�H  T ,�F H�  �C     	       ���  /
H H$iI  U/��  I$�#  T ,�= <!	   �C            �Ҫ  /
H <$iI  U/��  =$�  T ,�B �W	    D           �U�  ->) �%�2  �
 �
 -pw  �%�G  
 
 Hp ��2  �
 o
 0ss  �>	  ~
 z
 0 Z �>	  �
 �
 : �  �  Hn �>	  �
 �
 0~9 �>	  
 
 >P�  0?C �>	  �
 �
 0 P �>	  
 
 0P �>	  �
 u
 :��  ͬ  0�Y ��2  
 
 0f>  �>	  $ 
  
 Hi �>	  � 
 � 
 0S �>	  !
 � 
 :��  ��  02�  >	  i!
 e!
 Hcnt >	  �!
 �!
 ;D     $ |�  9Us 9T8 8,D     $ 9Us 9T8  ;�D     $ ��  9Us 9T8 8D     $ 9Us 9T8  :0�  �  Hndp �2  "
 �!
 0fI >	  �"
 �"
 Hi >	  9#
 -#
 0'Q >	  �#
 �#
 :��  ��  Huni #>	  +$
 %$
 Hgid $>	  z$
 v$
 ;1D     $ x�  9Us 9T8 ;QD     $ ��  9Us 9T8 8�D     $ 9Us 9T@  ;�D     $ ̭  9Us 9T8 8�D     $ 9Us 9T8  ;QD     $ �  9Us 9T8 8mD     $ 9Us 9T8   ;� D     $ ;�  9Us 9T8 8-D     $ 9Us 9T8  ,�> �W	  СC     !       ���  /
H ��T  U->) ��2  �$
 �$
  ,�O �W	  p�C     X       �K�  -
H � �T  %
 %
 -H[ � �  %
 u%
 -R�  � �  �%
 �%
 0�<  ��  t&
 p&
 '� �W	  �\8��C     � 9U�Q9T49Rv 9Y�\  S�Y ���C     1       ���  -
H ��T  �&
 �&
 0R�  ��  '
 '
 <�C     �  ,O W	  ��C            ���  /
H %iI  U/+�  %�H  THp �2  O'
 K'
  @^Z �
�  >�  A
H �
$iI  A��   $�#  C�W qT  Cn�  !	   ,nE �
!	  ��C            ���  -
H �
$iI  �'
 �'
 -��  �
$�  �'
 �'
 8��C     ��  9U�U9T�t9Q0  ,F �
!	  ��C     	      ��  -
H �
*iI  (
 (
 -��  �
*�#  �(
 �(
 -�@ �
*�  C)
 ;)
 0n�  �
!	  �)
 �)
 Hp �
�2  h*
 Z*
 0�@ �
�  +
 	+
 0��  �
�  �+
 �+
 0�S �
�  �+
 �+
 Hend �
�  �,
 �,
 Hmax �
�  �-
 �-
 Hmin �
�  B.
 <.
 Hmid �
�  �.
 �.
 >p�  0�  �
  �/
 �/
 0�W �
qT  �/
 �/
 8�C     �  9Uu    S�Z n
�C     �       ��  /
H n
qT  U0�  p
  T0
 R0
 Hp q
�2  �0
 x0
 0�S r
>	  1
 �0
 Hend r
>	  �1
 �1
 0�@ r
>	  U2
 O2
 0��  r
%>	  !3
 3
 Hn s
>	  F3
 D3
 0n�  t
!	  o3
 i3
 I�0  �
p�C      ,_F 4
W	  ��C     2      ���  ->) 4
%�2  14
 '4
 -pw  5
%�G  �4
 �4
 Hp 7
�2  /5
 5
 0ss  8
>	  �5
 �5
 0�@ 9
>	  d6
 ^6
 1P�C     �       L�  Hn M
>	  �6
 �6
 0�S M
>	  7
 7
 Hend M
>	  U7
 Q7
 0�@ M
 >	  �7
 �7
 0k� M
*>	  �7
 �7
 ;w�C     $ �  9U 9T8 ;��C     $ 2�  9U 9T8 8��C     $ 9U 9T@  ;P�C     $ i�  9U 9T8 8 D     $ 9U 9T8  ,[ %
W	  ПC            �˴  /
H %
qT  U->) &
�2  [8
 W8
  ,I �	W	  ��C            � �  /
H �	%iI  U/+�  �	%�H  THp �	�2  �8
 �8
  @�J �	�  g�  A
H �	$iI  A��  �	$�#  C�W �	�S  Cn�  �	!	   ,�L �	!	  ��C            �յ  -
H �	$iI  �8
 �8
 -��  �	$�  9
 9
 8��C     յ  9U�U9T�t9Q0  ,[O P	!	  `�C     !      �L�  -
H P	*iI  \9
 L9
 -��  Q	*�#  :
 :
 -�@ R	*�  �:
 �:
 0n�  T	!	  �:
 �:
 Hp U	�2  x;
 h;
 0�@ V	�  D<
 @<
 0��  W	�  �<
 �<
 0�S X	�  =
 =
 Hend X	�  b>
 T>
 0XM X	�  �?
 �?
 Hmax Y	�  u@
 k@
 Hmin Y	�  A
 	A
 Hmid Y	�  eA
 YA
 >@�  0�  �	  ZB
 VB
 0�W �	�S  �B
 �B
 8��C     L�  9Uu    S�@ 	P�C     	      �9�  /
H 	�S  U0�  	  #C
 C
 Hp 	�2  eC
 [C
 0�S 	>	  �C
 �C
 Hend 	>	  D
 D
 0XM 	>	  TD
 PD
 0��  	%>	  �D
 �D
 Hn 	>	  1E
 -E
 0n�  	!	  qE
 gE
 I�0  J	)�C     E��  '	 ,�: �W	  p�C     j      ��  ->) �%�2  �E
 �E
 -pw  �%�G  mF
 cF
 Hp ��2  �F
 �F
 0ss  �>	  �G
 �G
 0�@ �>	  $H
 H
 1��C     �       ��  Hn �>	  tH
 pH
 0�S �>	  �H
 �H
 Hend �>	  �H
 �H
 0XM � >	  @I
 >I
 0k� �*>	  �I
 �I
 1!�C     -       ��  Hd ��  �I
 �I
 8I�C     $ 9U~ 9T@  ;�C     $ ��  9U~ 9T8 8��C     $ 9U~ 9T8  ;��C     $ չ  9U~ 9T8 8��C     $ 9U~ 9T8  ,_@ �W	  0�C            �7�  /
H ��S  U->) ��2  RJ
 NJ
  ,v< pW	  �C            ���  /
H p%iI  U/+�  q%�H  THp s�2  �J
 �J
  ,K@ G�  `�C     �       �U�  -
H G$iI  �J
 �J
 /��  H$�#  T0>) J�2  K
 K
 0��  K�  aK
 ]K
 0n�  L!	  �K
 �K
 Hp M�2  �L
 �L
 C�S N�  C.� O�  Hidx P�  �M
 �M
  ,�H ,!	   �C     3       ��  /
H ,$iI  U-��  -$�  GP
 CP
 0>) /�2  �P
 �P
 0E  0!	  �P
 �P
 Hp 1�2  �P
 �P
 0�S 2�  OQ
 KQ
 0.� 3�  �Q
 �Q
 Hidx 4�  qR
 kR
  ,rZ W	  ��C     �       ��  ->) %�2  S
 S
 -pw  %�G  �S
 �S
 Hp �2  ?T
 /T
 0ss  	>	  �T
 �T
 0.� 	>	  xU
 pU
 :��  ۼ  0n�  !	  �U
 �U
 8-�C     $ 9U| 9T@  ;��C     $ ��  9U| 9T8 8e�C     $ 9U| 9T8  ,�Q �W	   �C            �g�  /
H �$iI  U/+�  �$�H  THp ��2  �V
 �V
  ,�; ��   �C     �       �x�  -
H �#iI  �V
 �V
 /��  �#�#  T0�  �   W
 W
 0E  ��  dW
 XW
 0��  ��  �W
 �W
 0n�  �!	  ~X
 hX
 0>) ��2  qY
 mY
 Hp ��2  �Y
 �Y
 0�@ ��  �Z
 �Z
 C�S ��  Dend ��  0XM ��  [
 [
 E��  � ,�N `!	  ��C     e       �@�  -
H `#iI  �[
 �[
 -��  a#�  �[
 �[
 0>) c�2  \
 \
 OE  d!	   Hp e�2  d\
 V\
 0�@ f�  ]
 ]
 C�S g�  Dend g�  0XM g�  []
 U]
  ,; �W	   �C     �      ���  ->) �$�2  !^
 ^
 -pw  �$�G  �^
 �^
 Hp ��2  j_
 N_
 0KW  �2  �`
 �`
 0ss  �  a
 a
 0�@ �  �a
 �a
 :�  k�  Hn �  :b
 .b
 0�S �  �b
 �b
 Dend �  0XM !�  hc
 dc
 0.� +�  �c
 �c
 0k� 2�  Xd
 Nd
 >`�  Hhi !	  �d
 �d
 Hlo !	  ^e
 Te
 :��  3�  Hd *�  �e
 �e
 ;�C     $ ��  9U} 9T@ ;p�C     $ ��  9U} 9T8 ;��C     $ ��  9U} 9T8 ;I�C     $ �  9U} 9T8 8a�C     $ 9U} 9T8  ;��C     $ P�  9U} 9T8 8��C     $ 9U} 9T8   ;��C     $ ��  9U} 9T8 ;}�C     $ ��  9U} 9T8 8��C     $ 9U} 9T8  ,�U �W	  `�C     $       ��  /
H �$iI  U/+�  �$�H  THp ��2  wf
 uf
  ,�J r�  ��C     �       ��  -
H r#iI  �f
 �f
 /��  s#�#  T0>) u�2  �f
 �f
 0E  v�  eg
 [g
 0��  w�  �g
 �g
 0n�  x!	  �h
 �h
 Hp z�2  �i
 �i
 0�S {!	  �j
 �j
 0.� |!	  l
 l
 Hidx }!	  Gm
 Am
  ,K \!	  @�C     I       ���  /
H \#iI  U-��  ]#�  �m
 �m
 0>) _�2  �m
 �m
 0E  `!	  
n
 n
 Hp a�2  6n
 .n
 0�S b!	  �n
 �n
 0.� c!	  [o
 Qo
 Hidx d!	  1p
 /p
  ,oP 6W	  �C     �       ���  ->) 6$�2  bp
 Tp
 -pw  7$�G  q
 �p
 Hp 9�2  �q
 �q
 0ss  :!	  )r
 %r
 0.� :!	  ir
 er
 1}�C     E       ��  0n�  L!	  �r
 �r
 8��C     $ 9Uv 9T@  ;��C     $ ��  9Uv 9T8 8��C     $ 9Uv 9T8  ,`K �W	  �C     $       � �  /
H �$iI  U/+�  �$�H  THp ��2  Ts
 Rs
  @"M ��  i�  A
H �#iI  A��  �#�#  Cn�  �!	  FCYI �S    ,#[ �!	  ИC     :       ���  -
H �#iI  �s
 ys
 -��  �#�  �s
 �s
 ;��C     O�  ��  9U�U9T�t9Q0 <�C     ��   ,�E �!	  ��C     P      �O�  -
H �)iI  @t
 4t
 -�N �)�#  �t
 �t
 -�@ �)�  ju
 bu
 0�  ��7  �u
 �u
 0�� ��2  �u
 �u
 0�R �!	  (v
 &v
 0�S �!	  |v
 Tv
 Hend �!!	  Fx
 x
 0x  �&!	  dz
 Dz
 0� �	  �{
 �{
 Hmax �!	  O}
 A}
 Hmin �!	  �}
 �}
 Hmid �!	  t~
 J~
 0�; �!	  �
 �
 0�j �!	  ��
 ��
 0n�  �!	  K�
 #�
 Hp ��2  ��
 @�
 : �  ��  Hi !	  ��
 k�
 :��  ��  0C !	  c�
 [�
 0�Y �2  ǉ
 ��
  > �  0�R >!	  /�
 '�
 0gU >"!	  ��
 ��
   >��  0YI �S  f�
 b�
 ;r�C     �  !�  9Uu  ;ВC     �  9�  9Uu  8�C     ��  9Us    ,cN 9!	  ��C     �      ���  -
H 9)iI  ��
 ��
 -�N :)�#  �
 ݋
 -�@ ;)�  %�
 �
 0�  =�7  ��
 ��
 0�� >�2  Ռ
 ӌ
 C�R A!	  0�S A!	  �
 �
 Hend A"!	  E�
 A�
 0x  A'!	  ��
 {�
 0� B	  ��
 ��
 Hi C!	  �
 ��
 0�; C!	  ��
 ��
 0�j D�  �
 �
 0n�  E!	  ��
 ��
 Hp F�2  $�
  �
 Hq G�2  `�
 ^�
 E��  i>��  Hr l�2  ��
 ��
   ,�D wW	   �C     	      ���  ->) w$�2  �
 ��
 -pw  x$�G  �
 ��
 Hp z�2  �
 �
 0ss  {!	   �
 �
 0��  }�2  ՗
 Ǘ
 0�D }�2  ��
 ��
 0�P  } �2  ��
 ژ
 0�o  }*�2  /�
 )�
 0	E }3�2  ��
 |�
 0�; ~!	  י
 ϙ
 0� W	  G�
 7�
 :p�  ^�  0�Q �!	  �
 ��
 0�N �!	  ��
 ��
 00R �!	  �
 �
 ;�C     $ D�  9U~ 9T8 8��C     $ 9U~ 9T8  :��  �  0�S �!	  ��
 ��
 Hend �!	  �
 �
 0x  �!	  ��
 �
 Hn �%!	  ��
 ��
 0>E �!	  ��
 ��
 0; �!!	  �
 
�
 0� �	  ��
 ��
 09Z ��2  &�
 �
 0��  ��2  �
 ٢
 0!= ��2  ��
 ��
 0�p  ��2  o�
 _�
 :��  ��  Hi !	  �
 �
 Hidx !	  F�
 >�
 8�C     $ 9Uv 9T@  ;-�C     $ ��  9U��9T8 ;��C     $ ��  9U��9T8 ;K�C     $ ��  9U��~9T8 8t�C     $ 9U��9T8  ;��C     $ -�  9U~ 9T8 ;��C     $ J�  9U~ 9T8 ;!�C     $ g�  9U~ 9T8 ;=�C     $ ��  9U~ 9T8 ;U�C     $ ��  9U~ 9T8 8��C     $ 9U~ 9T8  S%: @�C     W      ��  -
H S  �
 ӥ
 0�  �7  ��
 ��
 0�� �2  Φ
 ̦
 0�j !	  �
  �
 I�0  p�C     I�D g��C     >@�  0�D "�2  �
 ק
 Hend #!	  ��
 ��
 0� $	  #�
 �
 :0�  ��  Hp +�2  ��
 ��
 >p�  0n�  4!	  ��
 ��
   :��  ��  0n�  G!	  1�
 )�
  8��C     �  9Uu    ,nL �	  �C     '      ���  /
H �!S  U-�E �!!	  ��
 ��
 0>) ��2  ˪
 ɪ
 Hp ��2  �
 �
 05�  �!	  ͬ
 ˬ
 >��  0x  �!	  ��
 �
 4ČC     0       0�  ��7  ��
 ��
 0�� ��2  ��
 ��
    , P �W	  ��C     (       �2�  /
H �S  U/>) ��2  THp ��2  ޭ
 ܭ
  ,�< AW	  ��C     $       ���  /
H A$iI  U/+�  B$�H  THp D�2  �
 �
  ,�I ��  P�C     R      �g�  -
H �#iI  .�
 *�
 -�N �#�#  k�
 g�
 0>) ��2  ��
 ��
 0n�  �!	  Ю
 Ʈ
 0E  ��  H�
 B�
 0�j ��  ��
 ��
 0�X ��2  p�
 h�
 I�u  9��C     I�M 0̊C     :��  �  Hp ��2  ܰ
 ̰
 0�S  !	  ��
 ��
 0.� !	  "�
 �
 0� 	  ��
 ��
 0x  !	  J�
 >�
 0�: !	  �
 �
 Hpos !	  q�
 o�
 Hidx !	  ��
 ��
  ;q�C     ��  -�  9Uy 9Tx  ;ǊC     ��  K�  9Uy 9Tx  8�C     ��  9Uy 9T
   ,�G �!	  ��C     �       ���  -
H �#iI  �
  �
 -��  �#�  C�
 =�
 0>) ��2  ��
 ��
 0E  �!	  е
 ʵ
 0�X ��2  !�
 �
 1ƉC     z       ��  Hp ��2  v�
 j�
 Hidx �!	  
�
  �
 0�S �!	  ��
 ��
 0.� �!	  x�
 n�
 0� �	  L�
 F�
 0x  �!	  ڹ
 ֹ
  8��C     ��  9Tx   ,�X ��2  P�C     `       �t�  ->) �&�2  �
 �
 -��  �&�  k�
 e�
 OE  ��2   I�u  ���C     >P�  0�: �!	  ��
 ��
 0�Z �!	   �
 �
 Hp ��2  ��
 ��
 0��  ��2  �
 �
 Hsub ��2  <�
 8�
   ,�W (W	  ��C     v      ���  ->) ($�2  ��
 r�
 -pw  )$�G  W�
 K�
 Hp +�2  ��
 ܽ
 0ss  ,!	  &�
 �
 Hn .!	  ��
 ��
 0��  .!	  5�
 +�
 0&; /�2  ��
 ��
 0��  0�2  2�
 .�
 0	E 1�2  r�
 h�
 :��  ��  Hidx D!	  ��
 ��
 8)�C     $ 9U~ 9T8  : �  ��  0�H [!	  ��
 ��
 0U [!	  ��
 ��
 0x  [(!	  O�
 M�
 0� \	  ��
 ��
 :0�  j�  Hids r�2  �
 �
 :@�  P�  0�� |�2  D�
 B�
 Hidx }!	  q�
 g�
 8��C     $ 9U~ 9T@  8�C     $ 9U~ 9T9  8��C     $ 9U~ 9T8  ;8�C     $ ��  9U~ 9T8 ;��C     $ ��  9U~ 9T8 8��C     $ 9U~ 9T8  T\E �W	   �C     $       �)�  j
H �$iI  Uj+�  �$�H  TXp ��2  /�
 -�
  TMK ��  ��C     3       ���  j
H �#iI  Uj��  �#�#  TV>) ��2  X�
 T�
 V�j ��  ��
 ��
 VE  ��  ��
 ��
 Vn�  �!	  �
 
�
  TbQ �!	  ��C            ��  j
H �#iI  Uj��  �#�  TV>) ��2  r�
 p�
  _,E aW	  c�  `>) a$�2  `pw  b$�G  bp d�2  ass  e!	  Fbn t!	  bidx t!	    TQZ @W	  ��C            ���  j
H @iI  Uj>) A�2  T TIX �W	  @�C     �      ���  U�  �,�7  ��
 ��
 Un  �,�  3�
 '�
 U�C �,�G  ��
 ��
 Xbdf ��7  U�
 I�
 V�  ��  ��
 ��
 V� �W	  Q�
 ;�
 Xp ��2  K�
 =�
 V.� �!	  ��
 ��
 V�V ��2  ,�
 &�
 VE �v	  ��
 ��
 e�u  �N�C     W�C �:0�  ��  V9� �!	  ��
 ��
 V-� �!	  ��
 ��
  :`�  S�  V� �!	  ��
 ��
 >��  V ��  q�
 o�
 V�\ ��  ��
 ��
 ;ñC     0 6�  9Uv  8�C     < 9U��9T0   h��  U�C       ��  ���  3��  	�
 �
 3��  \�
 V�
 >��  5��  ��
 ��
 K�  ��5�  ��
 ��
 \�  6$�  p�C     7,�  ��C     �       L�  5-�  S�
 E�
 57�  ��
 ��
 5C�  .�
 *�
 5O�  l�
 j�
 5[�  ��
 ��
 5g�  ��
 ��
 ]s�  8�C             5t�  ��
 ��
   ;Z�C     C�  |�  9U} 9T FDB9Q��9R�� ;~�C     K ��  9U��9Q~  8}�C     X 9U��9T~    8��C     H 9Uv   _uO >W	  ��  `�  >&�7  `Jy  ?&e  bbdf A�7  ass  B>	  a� CW	  W�u  �WL �Fbp T�2  a��  U!	  a�/  V!	  aV` W>	  a.� X!	  a�V Y�2  Fa��  o!	     k�Y )��  `�  )$�7  bbdf +�7  FaJy  0e    SY �@�C     q      �O�  -�  ��7  ��
 ��
 0R�  ��  �
 �
 0$S  �eD  A�
 =�
 : �  I�  0Jy  �e  y�
 w�
 8�C     X 9Ts�  M��  ��C      ��  ���  3��  ��
 ��
 >��  5��  ��
 ��
 ]��   �C     H       5��  3�
 1�
 86�C     X 9Ts�
    MȖ  ��C      ��  ��  3Ֆ  Z�
 X�
 >��  5�  �
 }�
 8��C     X 9Ts�
   Yr�C     "�  9Us  Y��C     6�  9Us  ;��C     � N�  9Uv  ;��C     � f�  9Uv  ;\�C     � ~�  9Uv  Y}�C     ��  9Us  ;��C     � ��  9Uv  ;��C     � ��  9Uv  ;��C     � ��  9Uv  ;��C     � ��  9Uv  ;��C     � 
�  9Uv  ;�C     � "�  9Uv  ;w�C     � :�  9Uv  8��C     � 9Uv   ,�M nW	  ��C     �      ���  -Jy  n"e  ��
 ��
 -�  o"�7  ��
 ��
 -� p"	  ��
 ��
 -G  q"	  �
 ��
 -G  r"d  m�
 e�
 '� tW	  ��~0�A vW	  ��
 ��
 0�N x�  ��
 ��
 0aJ y�  �
 �
 0~J z�  ��
 ��
 0_? {�  ��
 ��
 0J |�  a�
 [�
 0$S  ~eD  ��
 ��
 I�u  ���C     :P�  ��  Hi �	  ��
 ��
  :��  ��  0�� c  .�
 "�
 0?1  d2	  ��
 ��
 :P�  ��  Hm �	  ��
 ��
 0�G ��  1�
 +�
 :��  ��  0�� ��  �
 {�
 =<�  '�C       ��  �3[�  ��
 ��
 3N�  ��
 ��
 >��  5��  �
 ��
 5��  F�
 B�
    4��C     C       '��  ��  ��8��C     � 9U	��H     9T09Q 9R0   : �  d�  0.� �!	  ��
 ��
 >0�  0R�  �  ��
 ��
 0	Y  		  ;�
 /�
 0�H �  ��
 ��
 'N G  ��0�B  ?  9�
 -�
 0�: 	!	  ��
 ��
 0�M 	!!	  �
 �
 :`�  ��  0�� c  i�
 g�
 N��C     9U} 9T~ 9Q   ;��C     � ��  9Uw 9T 9Q09R 9X09Y��~ ;�C     � )�  9Uw 9T49Q09R 9X09Y��~ 87�C     � 9Uw 9T49Q��~9R��~9X��~9Y��~   M]�  P�C       ��  ���  3n�  ��
 ��
 3n�  ��
 ��
 3z�  ��
 ��
 >��  5��  M�
 I�
 5��  ��
 ��
   p]�  ��C            ��  Jn�  Jn�  Jz�  4��C            5��  ��
 ��
 ?��    M]�  ��C       �  �{�  3n�  ��
 ��
 3n�  ��
 ��
 3z�  �
 �
 > �  5��  J�
 F�
 5��  ��
 ��
   8��C     ��  9U}   M]�  ��C       ��  ���  3n�  ��
 ��
 3n�  ��
 ��
 3z�  �
 	�
 >��  5��  k�
 g�
 5��  ��
 ��
   p]�  ��C             �D�  Jn�  Jn�  Jz�  4��C             5��  >�
 :�
 ?��    p]�  ��C     *       ���  Jn�  Jn�  Jz�  4��C     *       5��  v�
 t�
 ?��    Yc�C     ��  9U} 9Txibs9Qv 9R0 Y��C     ��  9U} 9Tv  Y��C     ��  9U} 9Tv  Y��C     �  9U} 9Tv  Y��C     %�  9U} 9Tv  Y��C     ?�  9U} 9Tv  Y�C     Y�  9U} 9Tv  Y'�C     s�  9U} 9Tv  Y4�C     ��  9U} 9Tv  YE�C     ��  9U} 9T�U ;��C      �  ��  9U} 9T19Qv  Y#�C     ��  9U} 9Tv 9Q0 Y=�C     	�  9U} 9Tv 9Q0 Y[�C     (�  9U} 9Tv 9Q1 Yx�C     G�  9U} 9Tv 9Q1 Y��C     a�  9U} 9Tv  ;��C      �  ��  9U} 9TE9Qv  ;�C      �  ��  9U} 9TF9Qv  ;;�C      �  ��  9U} 9T2 Yb�C     ��  9U} 9Tv  ;�C      �  �  9U} 9T@9Qv  ;e�C      �  $�  9U} 9TA9Qv  ;��C      �  G�  9U} 9T19Qv  ;��C      �  j�  9U} 9TA9Q}0 ;��C      �  ��  9U} 9T@9Qv  Nj�C     9U} 9Txibs9Qv 9R0  ,�A VW	  `D     (      �[�  -Jy  V"e  ��
 ��
 -�  W"�7  +�
 �
 -� X"	  �
 �
 -G  Y"	  u�
 m�
 -G  Z"d  ��
 ��
 0� \W	  E�
 A�
 0k  ]  ��
 }�
 0$S  ^eD  �
 ��
 0�  _	  _�
 S�
 :� ��  0~ u�  ��
 ��
 0�O  ui	  �
 �
 8�D     T 9T	�BH     9Q1  1 D     @       V�  0�I {�  T�
 R�
 ;-D     a 5�  9Us 9T	�.H      8<D     T 9T	�1H     9Q0  1�D     (       ��  0�I ��  y�
 w�
 ;D     a ��  9Us 9T	�.H      8D     T 9T	�1H     9Q0  :  ��  0R�  ��  ��
 ��
 '|Y �>	  ��~0��  �>	  �
 �
 0x  �>	  B�
 <�
 0�m  �		  ��
 ��
 0$~  �		  ��
 ��
 0�|  �		  ?�
 +�
 0J �		  �
 �
 0� �	  t�
 d�
 0FC ��2  8�
 "�
 0�D ��2  5�
 !�
 :p ��  0?W �>	  �
 	�
 0�D �>	  Q�
 K�
 0�: �)>	  ��
 ��
 Hp ��2  ��
 ��
 Hi  !	  l�
 d�
 ;�D      8�  9Us  ;kD     � a�  9Us 9T| 9Q} 9R4 ;D     � ��  9Us 9T| 9Q~ 9Rv  8D     n 9U 9T~ 9Qv   YD     ��  9U} 9Travf9Qs 9R��~ ;DD     � ��  9U| 9T  ;OD     � �  9U| 9T~  YcD     :�  9U} 9Tfylg9Qs 9R0 Y{D     b�  9U} 9T2FFC9Qs 9R0 Y�D     ��  9U} 9T FFC9Qs 9R0 ;�D     y ��  9U| 9T��~9Q��~ ;�D     y ��  9U| 9T��~9Q��~ ;=D     � ��  9Us 9T��~ ;[D     � �  9Us 9T��~ ;~D     � 7�  9Us 9T2 ;�D     � W�  9Us 9T��~ ;�D     � w�  9Us 9T��~ ;�D     � ��  9Us 9T��~ 8!D     � 9Us 9T��~  M[�  �D        ��  3z�  ��
 ��
 3m�  ��
 ��
 >  5��  ��
 ��
 K��  ��~5��  ��
 ��
 5��  ��
 ��
 6��   D     M��  KD      � ��  3�  p�
 d�
 3�  p�
 d�
 3��  �
 ��
 >� 5�  ��
 ��
 K"�  ��~K/�  ��~5<�  X�
 D�
 5I�  D�
 .�
 5V�  A�
 /�
 5c�  -�
 �
 5p�  b�
 N�
 5}�  c�
 3�
 5��  q  c  5��    
 5��    6��  TD     L.�  0 ��  5/�  � � L<�  � _�  K=�  ��~8�#D     � 9Us 9Q��~  ;-#D     � w�  9U  ;F#D     
 ��  9U  ;�#D     $ ��  9U  <T$D     �  L��  � ��  ?��  5��  9 / 5��  � � 5��  � �  L�  @ ��  5�  y o ;�D      !�  9U  ;�D      9�  9U  ;�D      Q�  9U  ;�D      i�  9U  ;	D      ��  9U  8.D     $ 9U   L�  � ��  5 �  � �  ;iD     � ��  9U 9T	 �H     9Q��~ ;7D     y ��  9Us 9Q��~ ;_D     � �  9Us  ;kD     � 3�  9Us 9Tw  ;BD     y X�  9Us 9TP9Q��~ ;�D     � ��  9Us 9T09Q09X09Y��~ ;6D     � ��  9Us 9T89Qw 9Xw 9Y��~ ;bD     
 ��  9U  ;KD     � ��  9Us 9Tv  ;SD     � �  9U~  ;^D     � %�  9Us 9T~  ;1 D     $ =�  9U  ;I D     � h�  9Uw 9Q89R	��C      ;%"D     � ��  9Us 9T19Q��~4$#9R��~9Xv 9Y��~ ;	$D     � ��  9U~ 9Tv  <0$D     �   L��  � ��  5��  9 5 ;�D     � �  9U 9T	@�H     9Q}� ;jD     � I�  9U��~9T89Q09X09Y��~ ;�D     
 a�  9U  ;�D      y�  9U  8�D     $ 9U   ;D      ��  9U  ;D     � ��  9U 9T��~ ;?D     � ��  9U 9Ts  85D     y 9U��~9T89Q��~   ;�D     � ,�  9Us 9T	�1H      ;�D     � D�  9Us  N�D     9U} 9Ts   @,I �W	  ��  AJy  �e  A�  ��7  CR�  ��  C� �W	  Dtag �>	  Cx  �>	  '/Q �"�  	@�H     E|N �FDn "	    @�L �W	  M�  AJy  �e  A�  ��7  CR�  ��  C� �W	  CHJ ��1  C_>  �2  C�8  �M�  C: �>	  C$S  ��2  C�S  �e  C: ��2  C�F �>	  Dnn �	  C[N �>	  '? �"��  	 �H     E�u  �[�  C�N �!	  C> �!	  C^A �,!	  Dx �8!	   [�  C>) 2   [.�  C>) 12   FC>) �2  FCW �>	     	2  ,DT vG   ��C            ���  Pa v!U  UPb w!U  T0�9 y2  r p 0: z2  � � 0�E |>	  � � 0�E }>	  � �  SA h��C     )       �<�  -Jy  h!e    0R�  j�  b ` <��C     �  @= "�   �  A  "G   Ad  #G   �A %��    'G    d  (G   = )�   �F +h�  ��  ��  ��  @   
 ��  '�J .��  	`�H     Dcur @��  	��  C�� @��   TlW �W	  ��C     �      ��  U�  �"�7  � � U7Y �"		  @ 2 UF@ �"kA  � � VR�  ��  I E &� �W	  ��VE  �]  �  Xn �		  	 	 Xrec ��2  �	 �	 V�Q �	  �
 �
 V�E �	  � � V�K �	  
 � V�B �	  � � V�> �	  X H V5M ��    V�I �2R  � | I�u  ��C     1��C     �       ��  0Jy  
e  x v ;��C     � ��  9U| 9T 9Q09X09Y�� ;��C     � ��  9U~  ;��C     � ��  9U|  8�C     � 9U~   N��C     9Us 9T|   T�L \]  �C     �       � �  U� \(�2  � � UR�  ](�  � � V�� _]  0 * Xlen `!	  � z V� `!	  � � Xn `!	    V�1 a�2  � � &� bW	  �\8�C     � 9U�T9T19Q09Rs����9X09Y�\  T�@ 9]  ��C     �       ���  U� 9(�2  � � UR�  :(�     V�� <]  r l Xlen =!	  � � V� =!	    Xn =!	  O E V�1 >�2  � � &� ?W	  �\8ƸC     � 9U�T9T19Q09R|����9X09Y�\  ,|M �\  P�C     
       �b�  -~ �$�  #  -;  �$�  ` \ RZ�C     � 9U	 �H     9T�T  ,_X @W	  0�C     t       �L�  -�  @&�7  � � -A! A&�G  9 - -' B&�G  � � '= DRG  �@'d�  D RG  �P0� EW	  ] U ;P�C     ��  $�  9Us 9T	1�H     9Q�P 8p�C     ��  9Us 9T	B�H     9Qw   @�K ��  ��  A�  ��7  C;�  	  Dwin 	  C�Q 	  CE  �   @�? �  <  A�  "�7  C� W	  CR�  �  Dmm �M  C�u  !	  C�  		  C2�  
#L  C;�  	  Dwin 	  C�Q 	  Di !	  Dj !	  CE  �   Dp �   EuS �EYY �[��  Dlen !	   [��  C$S  deD  CϽ  f2	  CCg  g!	  C�  i�   FCc  {!	  Ca> }�   Ds ~�     [  Cdh  ��/  FDt ��     FCߢ  ��  Cx�  �<  Dh ��#  FDv ��     �  L  @    @ E ��   �  A�  �	  Bbuf ��   Dp ��   Dq ��   Dtmp ��  C�Y �	  C�Q �	  Di �	   �   �  @    ,�9 P�  ��C     �       �j -�  P �7  � � Pid Q 		  T.win R ,B  � � /�Q S ,B  RHn U	  O I >�  0F@ ]�2  � �   q�L �   ��C     J      �� -R�  %�     -Jy  %e  � � -� %�2   � -e: %N  k c -�@ %�  � � '� W	  ��0E  �   ? 1 Hr ]  � � Hp  f6  _ [ Hlen !!	  � � ;��C     y v 9Us 9Q�� ;��C     � � 9U}  ;��C     
 � 9U}  ;^�C     $ � 9U}  ;��C     � � 9Us 9T�� 8��C     � 9Us   q0C ��   `�C     -      �t -R�  �#�  � � -Jy  �#e  s k -� �#�2  � � -e: �#N  A 9 -�@ �#�  � � '� �W	  ��0E  ��   � � Hr �]  � � Hp �f6    � Hlen �!	  : 6 ;��C     y � 9Us 9Q�� ;��C     �  9Uv  ;��C     
 / 9Uv  ;9�C     $ G 9Uv  ;^�C     � _ 9Us  8y�C     � 9Us   Q�N %� Bkey %*U  Blen &*Z   Aߢ  '*�  Bout (*_   C�U  *�  C�F +N   Dh1 -�  Dh2 .�  Dh3 /�  Dh4 0�  Dc1 2�  Dc2 3�  Dc3 4�  Dc4 5�  C 7� Di 9
G   [~ Dk1 >�  Dk2 ?�  Dk3 @�  Dk4 A�   FC��  j�  Dk1 l�  Dk2 m�  Dk3 n�  Dk4 o�    	�  @�Y �  � Bh �   ,n@ G   ��C            � .c G   t p  T1@ �G   ��C     "       �[ rc �G   UXcc �S   � �  TU �!	  �D     �       �� U�  �$  � � Ula �$]  @  8  Ve5  ��7  �  �  Xi �!	  
! ! V5? �!	  G! A! 4D     /       &��  �]  �HV� �W	  �! �! sq  D      D            �� 3@q  �! �! 33q  " " 3&q  3" 1" 4D            ?Mq  ?Zq  ?gq  ?tq  \�q  8*D     � 9Uv 9Ts 9Q�H   8;D     � 9U}    _�O �W	   `�  �$  `�^ �$!	  `B� �$i	  `(5  �$!	  a��  �]  a� �W	   _�A yW	  j `�  y�7  iidx z!	  itag {0  `x  |0  `ss  }0   TA L_    �C     �       �� j�  L �7  Ugtag M .  Z" V" V>) O_   �" �"  t @D     V       �_	 u- U39 �" �" uE QuQ Ru] X] dD     ,       3] K# I# 3Q p# n# 3E �# �# 39 �# �# 3- �# �#   t �  �D     U       �u
 32�  ($ $ 3?�  �$ �$ KL�  P1�D            �	 5Z�  |% r% R�D     ��  9U�U9T�T9Q1  7 �  �D            a
 3?�  �% �% 32�  2& .& 4�D            5L�  m& k& ]�	 �D            ?Z�  8�D     ��  9Us     R�D     O�  9Q1  t �   D     ?       �& 32�  �& �& 3?�  �& �& 5L�  g' a' KY�  PL �  ��   3?�  �' �' 32�  �' �' >��  ?L�  5Y�  ( ( 8*D     L�  9Uu    RD     յ  9Q1  t��  @D     ?       �� 3	�  @( :( 3�  �( �( 5#�  ) ) K0�  PL��   �  � 3�  a) ]) 3	�  �) �) > �  ?#�  50�  �) �) 8jD     �  9Uu    RXD     ��  9Q1  t%�  �D     \       �� 37�  �) �) 3D�  o* c* 5Q�  �* �* L%�  0�  t 3D�  J+ F+ 37�  �+ �+ >0�  5Q�  �+ �+ \^�  8�D     K 9Uv 9Qs�   N�D     9Us 9Tpamc9Qv 9Rs�  vq  PD     Q      �� 3&q  �+ �+ 33q  �, �, 3@q  �- �- 5Mq  �. �. 5Zq  �. �. 5gq  �/ �/ 5tq  k0 _0 \�q  L�q  p  l 5�q  �0 �0 7�q  �D     /       W 5�q  11 /1  8hD     �r  9Us   L�q  �  � 5�q  X1 T1 8�D     �r  9Us   YzD     � 9U0 N	D     9U}   tq  �D     &       �9 3&q  �1 �1 33q  �1 �1 3@q  >2 82 ?Mq  ?Zq  ?gq  ?tq  R�D     � 9U�U9T�T9Q�Q  t� �D     r       �� 3� �2 �2 3� �2 �2 3� :3 .3 3� �3 �3 ? ? hq  �D      �  �� 3@q  X4 V4 33q  �4 �4 3&q  �4 �4 >�  ?Mq  ?Zq  ?gq  ?tq  \�q    ^�  3� *5 $5 3� y5 s5 3� �5 �5 3� 6 6 > K �X5 r6 l6 wq  �D            �� J@q  J3q  J&q  4�D            ?Mq  ?Zq  ?gq  ?tq  \�q  8�D     � 9U�U9T�T9Q�X   8�D     � 9Uv 9Qs ����    t��  �D     B       �� 3��  �6 �6 3��  F7 :7 3Ɍ  �7 �7 5֌  "8  8 ?�  L��  @ � 3Ɍ  G8 E8 3��  s8 m8 3��  �8 �8 >@ K֌  P5�  9 9 \�  R2D     � 9U�T9T	��H     9Q�U#�   N
D     9Us 9T�Q9Qv 9R0  t,�  `D     �       �C 3>�  x9 l9 3K�  :  : 5X�  �: �: ?e�  L,�  �  3K�  *; "; 3>�  �; �; >� 5X�  < < 5e�  �< �< \΄  ;�D     � � 9U| 9T	 �H     9Q}  ;D     � � 9U| 9T	��H     9Q}  ;(D     � � 9U| 9T	��H     9Q}  RTD     � 9U�T9T	��H     9Q�U#�   N�D     9Us 9T2/SO9Q| 9R0  t�  �$D     �       �j 3�  �< �< 3(�  �= �= 54�  2> (> 5>�  �> �> 7�  �$D     :       3 3(�  �> �> 3�  ? ? 4�$D     :       54�  Y? W? ?>�  ]J�  �$D     :       5K�  �? |? 5U�  �? �? 8%D     $ 9Uv 9T@    ;-%D     $ P 9Uv 9T8 8<%D     $ 9Uv 9T8  tL�  �)D     
      �� 3^�  B@ 2@ ?k�  ?x�  ?��  x��   LL�  @ c 3^�  �@ �@ >@ 5k�  >A <A Kx�  ��K��  ��5��  jA fA ;�)D     �   9Uv 9Tt 9Q��9Rr  ;"*D     � A 9R	��C     9X1 8�+D     j 9R	��C     9X1   =��  8*D      p 3��  �A �A >p K��  ��5��  B B 5��  YB SB K��  ��K��  ��K��  ��5�  �B �B K�  ��K&�  ��53�  $C C 5>�  �C �C 5I�  �C �C 5V�  E �D 6a�  .D     6j�  �+D     L��  � @ 5��  VG PG ?��  5��  �G �G K��  ��L��  �  5��  �G �G K��  ��5��  H H Y�*D     � 9Uv 9Q�� <�*D     H ;+D     y � 9U~ 9Q�� ;6+D      � 9U|  8�+D     � 9U~   Y�/D     + 9Uv 9Q�� 8�/D     H 9U   L��    $ 5��  BH :H L��  P � 5��  �H �H =L  K,D       � �3k  4I ,I 3^  �I �I >� 5x  �I �I 5�  tK bK K�  ��5�  9L /L 5�  �L �L 5�  �M �M    ;�+D     y  9U~ 9Q�� <,D       L  	 � 5  fN `N K  ��5"  �N �N Mt ".D      P	 �� 3� /O 'O 3� �O �O 3� ,P $P 3� �P �P >P	 5� �P �P 5� GQ ;Q 5� R R 5� "S S 5� T T 5� �T �T 5  �U �U 5 "V V 5 �V zV 5$ �V �V 50 >W 6W 5= �W �W 7H �.D     �       � 5M �W �W 5Y �X �X 5e EY AY 5q �Y }Y  L~ �	 � 5 DZ >Z 5� �Z �Z 5� a[ Q[ 5� $\ \ 5� �\ �\  M� �0D      
 �

 3� �] �]  M� �0D      �
 �
3 3� 	^ ^  M� �0D      � �
\ 3� A^ ?^  =� 1D      � �
3� h^ d^    ]-  x1D     '       5.  �^ �^   Ls�  0 � 5x�  	_ _ ;g2D     �  � 9Uv 9Tt 9Q��9Rr  ;�2D     �  9R	��C     9X0 ;�2D     H ( 9U|  ;3D     �  S 9Uv 9Tt 9Q��9Rr  ;63D     �  ~ 9Uv 9Tt 9Q��9Rr  8\3D     j 9R	��C     9X0  Nk*D     9Uv 9T��9Q��9R09X��    y9  9  cz�A �A ,FzR R ,�z�9 �9 ,�y�U  �U  �y�3  �3  �yRH  RH  �yxL  xL  �y?  ?  �yT)  T)  �y�*  �*  �y�J  �J  �yjO  jO  yL  L  �yF  F  mzF\  F\  -�z�6  �6  -�yE1  E1  ry?U  ?U  �y>Q  >Q  �y _   _  hy�N  �N  �y`I  `I  xy�F  �F  �y�3  �3  1zU  U  #kz�X �X 'z%[  %[  #zz��  ��  .z�[ �[ ."z�O  �O  .2yKM  KM  Yy�R  �R  {�  �  0 z�K  �K  -vzIE IE /�{�D  �D  0 y�U  �U  ^z_T  _T  1Xy�X  �X  Xy�:  �:  Sy!,  !,  Uy�*  �*  [zBi  Bi  .yq]  q]  -zz;�  ;�  . #  �S  l�  �o $"  �3D     *�      X� L�i :G  �@   LX  ^� �S   L�i mint n,{S @�   
g
  �    
   	G   
v  #	G   
�  &	G   
|
  )	G    
h  ,	G   (
�  -	G   0
�	  2Z   8
�  5Z   < �   L�  %�   �
  8"c   	  K  �   	�  L  	�  M  LS  L-  L�  >   Z   �	  	-   �  B"i  o  ,   ��  
R   �a    
�� ��  
�N ��  
�6  ��   �  Y�  �  &a   �  ]  @      n�  �  0�  ]  a    �  �    &a   )  ]  @   @   a    �  �"5  ;  �   PJ�  2�  L8   �  MS   ?pos NS   �  P�  SF  Q�   �1 R  (=9 SE  0R�  U]  8y�  V8  @�� W8  H o�  ��  d�\ �@   dm  �a    o  ��  �  �    &S   8  )  S   8  S    >  L�  2  R  X  0c  )     :@   ,�  J�  1x Lc   1y Mc   )  Oo  %�  ,B   s�  
M   uc   
}  uc  
V  vc  
/  vc   t
  x�  k	  (q  �  -    ��  -   �  	Z   B� 
8  L  <    >  s  >  v	  a     �  �  %q  �  (N�  �  P5   Z�  Q5  �  S�  s  T�   [  U�  ?1  WZ     �  5    Y�  �  K=  -   �C  �   /M
  pmoc/5  stib/	  ltuo/|  tolp 	  �  b   "]  c  ]�  %  <�  ?x >5   ?len ?<  *� @>   %  Bh  %�    `�  �  0�  Z   Z   �  a    �  �  q�  �  &Z     Z   Z   a    �    #  08  Z   Z   a    �  `��  �  ��   �% ��  ?1  �Z   �&  ��  !  ��   I  ��  ()  �  0R   �a   8�  ��  @ ~  �  p�  �8  %�  �   �  �  &Z     a      P  �    $  0/  P   �  ?<  B  0W  P  8  S    �  Yd  j  &Z   �  P  S   a    s  ��  �  &Z   �  P  �   �  W  0�  �  �C   e� ��  �� �/  �� �W  �� ��   �� �  ( �'  ��  �!  l>  �  �8  L�  -  �>  %?  K  �  ��   %V  �
  �5  �  �<  �  �Z   
  �-   �  �@   \#  �S   �   @   �  ,Z   \&  7a   �0  DG   �H  Q4   b   �3	  ?xx ��   ?xy ��  ?yx ��  ?yy ��   a  ��  %3	  z'  �p	  m  �P   ss  �   �  �E	    ��	  �	  0�	  a    �  ��	  �U  �a      �}	   %  ��	  �  $�	  �	  �   
  �� "�	   �@ #�	  �U  $a    �  7J
  �; 9�	   ��  :�	   L  <
  e-   (��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=  ��  ?c   �  @c  ~  Bc  �  Cc  �  Dc   5  Fc  (B  Gc  0�  Hc  8 �	  J�  
   s{  �  ug   ��  vg  �  xc  �
  zc  (  {c   �  }&  �  �#�  �  Yk  `�J  R�  �]   (  �  |  �  �  �  �  ��  �  ��"  6v  �J
  6�  ��  (6�%  �J  067&  ��"  86G   �  X �  �"W  ]  h  �  �M �"   k  �  R�  ]   �  �"�  �  %  8;�  �� =�"   �M >r    ?J
   r$  @�  0 5  �$�    %  �t  �� �"   �M �"  �  C   �  �  (�� 
P  h�� �  p�� �  x K  � �  �  �  �,H  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9  8  :�  @�  <  H�  =�  PE-  ?�	  X�!  D�  h:  Fs  �  Gg  ��  Hg  ��  Ig  ��  Kg  �  Lg  �U  Ng  ��  Og  �)�  Q�  ��  RH  ��� S�  �K1 W�  �R�  X]  �Jy  Y)  �%  [J
  ��	  ]�	  �    ^a   ��8  `+  � L   U  [    X��  �  �t   E-  ��	  N ��  �8  ��  P �  *%�  �  Y�  0t�  k  v�   �  wt  �@ x�  ݖ y�  E-  z�	   N |  0�  }�  pR  ~�  x�  �  �ߣ  �C  ��I �q  ��  �  �h  �  ��S  ��  �4  ��  �8  ��  �6  �a    6�  �@   6�  �c  6o  �c  6�L �a    6�8  �	  ( �
  L#    W  HY  �  Jt   = K    Ls  d  Ms   K�  -   �  �   /�  bmys/=  cinu/�  sijs/w    bg/O  5gib/p  snaw/M  ahoj/�    bg/�  sijs/�    bg/q  5gib/�  snaw/�	  ahoj/  BODA/4   EBDA/�	  CBDA/  1tal/�  2tal/   nmra �	  Y  #   g)8  >  �   ���  =  �3	   L  ��   $  �  0�  �;!  8m  �#�"  h�  �,  pآ  �C  tG   �  x V  {  �  �
  �)�  �  �   H�  �  �a    "  ��  �!  ��   ~	  8f�  �
  hs   (  is  �� k�  �� l�    nc  �  oc   �  pc  (�  qc  0 y  s    �$�  �  ,�  0'	  
�N  )   
?1  *s  
}0  +  
i/  ,  
� -3	   �  �)       H�  ��  ��   ?1  ��  (  �   4  �3	  \  ��  0  �a   @ +!  �  ?tag �   �U  �   �    �  K`  -   
�  w%   }#  �&  h  �  &     
�  E   9
W  � ;
�   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(d    K�  -   ��  :   �   ^$  1  �!  �!   :  �j  K�F  -   �  �D   ;?  �O   S  �9   �  ��  �#  ��  �  &�    J   I$  �     0+  J   �&  �7  =  &�  Q  J  Q   �   ,�!  H��  
�  ��   
S"  ��  
   ��  
�"  ��  
�  ��   
;  ��  (
%  ��  0
�   �  8
��  �+  @ b  R  �W  %�  x  =�	  H  E#  %�  ,�  @J�  
�  L�   
�  MC  
�� O�  
.� P  
�  Qw   
�  R"  (
�!  SO  0
8'  T�  8   W!�  �  ,-  (l�  
k  n�   
�M o�  
ߣ  pC  
�  q�   
  k  )�  �  &�    �  �   w   .    0"  �   �  1.  4  0I  �  I  �   @	  K  6[  a  0q  �  q   �  �  :�  �  &�  �  �  �   �  >�  "  Y�  �  &�  �  �  �  �  �   �  _�  �  &�  	  �  �  I  �   $  f    00  �  �  q   �  l<  B  &�  [  �  �  �   ,#  x��  
�� � �   
�  � C  H
  � �  P
�  � �  X
9!  � 	  `
l� � 0  h
  � �  p     �[  ,�  H2%  
�S  4�   
�  5�  (
  6�  0
4  7�  8
8  8�  @ �  :�  ,�  �=�  
R�  ?]   
�  @�  
n  A�  
�  B�  
1$  C   
2�  E%  
�� F%  `
�L Ha   � �  J�  1  P   �  �  &�  �  )  t      �   �  &�     0  t   �%  *    &�  ,  H   �%  -8  >  0I  H   {  1U  [  &�  j  �   �  4v  |  0�  �   l  8�  �  &�  �  H  W   �  <�  �  &�  �  H  �   �  @�  �  &�    �  H  �  C   �  G    &�  3  t  �  �  �   �'  N?  E  &�  Y  t  )   �  Se  k  &�  �  t  �  �  C  �   �  ,&  ��r  
�� ��   
i'  ��  H
   ��  P
  ��  X
�A ��  `
Y ��  h
�#  �  p
�  �,  x
�  �I  �
  �j  �
��  ��  �
U�  �  �
�!  �3  �
��  �Y  �
�  ��  �
&  ��  � �&  �~  �  }\  P&�  �  ]pR  qB  i�  �  0�  �  t  �  �   a   @   A  �  �  0�  �  a    4H  �      0   �  t   �U  �#   )   &�  L   �  �  H  �  C   ,�*   ��   
n*  �$�   
�5  �$�  
XO  �$�  
��  �$    ^~ �L   %�   ,�>  ��   
'O  �Q   
xC  ��   s/  ��   %�   �  0t;!  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�   �  U'T!  Z!  ]m  ,D   t�!  
�  v�   
A  w�  
�  x�  
&  y�   !  {_!  �  ��!  �!  &�  �!  H!  �  �!   p	  �  ��!  �!  0 "  H!  �!   �'  �"  "  &�  0"  H!  �     0"   �!  �!  o"  ��  )�!   ��  )�!  �  ) "   }  6"  %o"  O  ;�"  _� =%�"   ݰ  >%H!   |"  �  @�"  �"  �  �  ]  �  (J  �"  -S    (�  �"  -S    �  �%  ^,� -   N=(  �  â � (fa A�` i� {G� ��� �[� ��m ��� �U� �v l� R .�� 8� X�~ xE{ ��} �� ��� �#} �ݦ ��� � 4� T:� tφ �� �
� ��w �T� �� 4"� M@� �� ��� �wp �� ��� �i >9� ^�k ~�� � �� ��� �H� �  ȧ )�� Bxv [z� trh ��� �Ug �̮ �^ �{x ;j 5N� U�] uw� �Xs ��u ��� �� �� 5�f U�� uT� �w� ��_ ��� ��  � 1Ӱ FԬ Xϯ jOz ��s ��a �cw �0� 	� -	�` A	�t a	^} �	�� �	�l �	k� �	B� �	� �	׏ 
?n :
�h Z
d� r
�| �
�v �
;w �
+y �
�� �
 � �
�� Ǔ 1h� �Db ��` ��^ �� ��� �Qr �ܐ %� �� ,� :�u JA� Zv� d�b x?� �Wt ��[ ��� �i �ҙ �r .x� G@� R� rMp �o �7\ �� �>} ` :�� Z�� rAl ��� �� �Uc ��� �}� ��� ��j M� &� N$� v�� �� ��� �:� ��� )� "1z ,W� E�d O�� r�s ��` �z� �i� ��z � %�k -x\ A�� Me^ m� �� ��| �M� �� �;� c� �� !�� )ɥ 5Ǥ Ut uA� ��� �<� _�� (� (�z (�\ ) � #  (�   U(  Q %J(  �n U(  K� -   ?�)  ��  ̲ (d 	� (� �z nf t{  �� $h� +*� .8o 5�� :�� ?^� E[� K�g P`� S)� Xn _թ d4� g�o nD� tn� zr ~� �1� ��~ � � �L� �� �c� �� ��� �Ñ �1� �sc �}d �� ��� �� ��r �o� �� �ob �#� �z� ��� �] ��c ��� �� ��� �l� �z� �� �� � A� �g(  <� �*  �� �=(   2�  �s   �� ��)  %*  (*  ,*  Q %!*  �e �,*  ,�� Ms*  1org Oc   1cur Pc  1fit Qc   �� S>*  s S�*  >*  � �&�*  �*  Y�� x2 N�+  R�   P]   ��  R�  ͩ  Sc  ��  U�  =�   Vc   �   X  (2]   Y  ,�   Z�<  0n   \  8[   ]  <[   ^�@  @dh   `�@  H6�x  bP  6;�  cP  6N  e<,   6˴  gc  (6ʩ  hc  06B�  po@  8 ,D� 0�,  
�  �t   
�� ��  
�� ��  
ͩ �c  
=�  �c   
Q,  ��  (
?1  �P  , �y ��+  � �6,  �+  s� �(H,  N,  ȱ H��,  Nh ��3   �m �,  J� �   89� ��3  @ h� ��,  �,  &�  �,  <,  t   �� ��,  �,  0�,  <,  *,   w ��,  �,  0�,  <,   �� �-  -  0!-  <,  !-  !-   c  �� �3-  9-  &�  M-  �*  <,    � �Y-  _-  &�  }-  �  �*  }-  <,   �  Kgk -   �-  aj  �a շ �g �  � �-  �^ @A.  � �-   $\ (�  D� (�,  �d (�,  �j (�,   "� (�,  (� ('-  0j� (M-  8  � !�-  %A.  0� #,e.  %S.  N.  Kܱ -   <�/  Ԍ  N� �� � �� f x� �j on �t 	!� 
O� �� 
� �� Ō �f �� Ȑ �{ \� 1� \� �h � �^ �� 	� yj 	t >� �� M�  w� !�t "�{ #n� $İ %� &k� '�� (nd )4_ *}� +�� ,� ->� .�� /�| 0� 1r� 2�v 3Yx 4ƫ 5�n 6�� 7v� 8%~ 9 �� Ck.  `� F0  N� HP   k� IP   � K�/  %0  s O)20   0  l (R�0  Ƭ T�/   �z W%0  �e X%0  � Z   ж \Q    E� ^80  %�0  �\ `%�0  %�0  �0  K�� -   �1  <a  �c \ ?d 0� �h \� �u �� ݅ 	�n 
 �� ��0  Kș -   �,3  ��  8� � ʋ 4� ȸ ǣ �p �� z} 	�h 
� ч y �� �� ִ 4i } [f +| � �� �� K� d � �n 0� �� nr �� Ƃ  ہ !y~ "�� #�{ $� %۸ &�� '�v (�r )� *� +� ,n� -:� .1� /�^ 0f� 1a� 2y� 3�i 4�} 5g 6� 7�� 8�� 9[] :�� ;� <3~ =~� >�l ?� @� A[d B�� C� D~n E�� F\� G)a H�u I�� Jhx KH� L� M�_ NH� OH� PXy Q�y R�� Sjp T �n �1  [� ��3  ��  �,3   � ��-  Ƭ ��/  Is ��)  *� �1   j �93  %�3  b� �$�3  %�3  �3  %� �'�3  �3  Ud� �!i}4  
�  !kt   
� !l�  
� !mc<  
�} !u�  
N !wi<   2'� !{s  �2� !~c  �2�� !�c  �2o� !�c  �2x� !�c  �2h� !��  �2~ !�5  � .f �N,  RZ(  "	@�H     _1*  "�	��H     ,�k H##	5  
�� #%�"   
�� #'�  
B� #(�  
�{ #*    
�  #,   !
X;  #-	5  $ (  5  -S    Zh #/%5  �4  	�  #2�  (`.  B5  Q %75  	�� !!B5  	ٽ $!�0  	g� $'�0  	� $-�0  	�� $3�0  	� $9�0  	�� $@�0  	Rm $F�0  	�� $L�0  	m $R�0  	]� $X�0  	�� $^�0  	� $d�0  	)� $j�0  	 j $p�0  	M� $v�0  	Hq $|�0  	� $��0  	�� $��0  	-� $��0  	0� $��0  	�a $��0  	�� $��0  	�� $��0  	� $��0  	w $��0  	�� $��0  	$� $��0  	ۜ $��0  	� $��0  	�\ $��0  	,h $��0  	�� $��0  	�v $��0  	wt $��0  	n� $��0  	�� $��0  	�_ $��0  F] $�0  9� $�0  ;k $�0  �q $�0  3� $�0  � $ �0  "� $&�0  �� $,�0  t| $3�0  g� $:�0  �y $@�0  i� $G�0  W� $M�0  � $S�0  �x $Y�0  _ $a�0   $g�0  X� $m�0  b� $s�0  �� $}�0  (�0  8  Q %8  	Ѡ !+8  	�� %V�3  	� %]�3  	�n %d�3  	�b %k�3  	�p %r�3  	�� %y�3  	}� %��3  	�� %��3  	f %��3  	1� %��3  	� %��3  	� %��3  	�� %��3  	�� %��3  	 %��3  	U� %��3  	�e %��3  	�� %��3  	m� %��3  	�� %��3  	Fv %��3  	<� %��3  	Q� %��3  	ne %��3  	[| %��3  	Ș %��3  	�� %��3  	݋ %��3  	̍ %��3  	!� %��3  	]� %��3  	Ah %��3  	K� %��3  	C� %��3  	�m %��3  	)� %��3  	@� %��3  	n] %��3  	�� %��3  	9x %��3  	_ %��3  	�� %��3  	�� %��3  	r� %��3  ա %�3  �� %	�3  �� %�3  �� %�3  �\ %�3  ϊ %�3  �� %�3  r� %�3  �x %�3  �x %�3  �q %�3  !e %�3  �[ %�3  �� %�3  �� % �3  >� %'�3  >t %7�3  :� %>�3  _v %E�3  a %L�3  n %S�3  ի %Z�3  (l %a�3  L^ %h�3  �z %o�3  �� %v�3  �� %}�3  ֳ %��3  �b %��3  
� %��3  '� %��3  �[ %��3  �f %��3  � %��3  l� %��3  z� %��3  ޹ %��3  �� %��3  �� %��3  u %��3  (�3  R<  Q %G<  	nm !5R<  s  (<,  y<  -S   S ^-g -    !�<  |�  �z �  �  *y<  ^�w Z    /�<  @� e� f�� � f�l ~ ��  7�<  �|  �#�<  �<  ,�� P ��=  
?1   �s   
�  �,  
L�  �,  1ox  �c  1oy  �c  1fx  �g  1fy  �g  1x  �c   1y  �c  (1u  �c  01v  �c  8
�@  ��<  @
��  ��<  H Η  �#�=  �=  Ʒ P �>  ?1   ?   ?dir  ,  ?pos  g  �  g  �a  g  Li  	g  �   
g  
c�  �>  ^�  �=  ʊ  �=   	s  �=  (F�  c  0?len  c  8N�  �<  @k�  �<  H ��  �#�>  �>  A� X `?  dh  g   ��  c  ?pos  c  ?1    ?  ?dir  !,  ��  "�   �  $*  (ʊ  %�>  0	s  &�>  8F�  '  @N�  )�=  Hk�  *�=  P ��  ��<  6�  �=  ޖ  ,�>  g�	 A�?  �k  C�?   6�y  D�?  � (l?  �?  -S    (y?  �?  -S    Y�\ �	 1O@  �j  3   2n  4  �k  5�=  ��  :  (�  ;  �y  <�>  ��  >�<   B�  E�?  ( u  H�?  �a  Hi@  �?  g@ l�@  [   n�@   �   o�@  @ (�<  �@  -S    (`?  �@  -S   _ �<  (O@  �@  -S    1�  r�*  	� &N.  ,8s H&M5A  1ref &Os*   
#� &Ps*  
  &Qc  0
�  &Rc  8
?1  &S�  @ �p &U�@  Ѩ &UMA  �@  U x �G&X�A  
�� &Z�   
� &[c  
�� &]�  
�q &^�A  2k &_c  �2��  &`c  �2�p &a   �2v� &d�  �2�  &eB  �2�{ &g�  �G2v &hc  �G (s*  B  -S    (5A  B  -S   � �i &jSA  Dr &j0B  SA  U�l ��&mlB  
�� &o}4   
U�  &p�  H
dh  &qlB  P (B  |B  -S    -m &s6B  b� &s�B  6B  	�] 'N.  ,nu 8'@�B  1ref 'Bs*   
#� 'Cs*  
?1  'D�  0 � 'F�B  }� 'F�B  �B  U�f 88'I�C  
�� 'K�   
� 'Lc  
�� 'N�  
�q 'O�A  2k 'Pc  �2��  'Qc  �2�p 'R   �2� 'U   �2v� 'V�  �2�  'W�C  �2�{ 'Y�  (82v 'Zc  08 (�B  �C  -S   � �� '\�B  �x '\�C  �B  UY� �p'_D  
�� 'a}4   
U�  'b�  H
dh  'cD  P (�C   D  -S    �k 'e�C  ]\ 'e8D  �C  e-   (��F  B^  �� 4` � Oo � k� � &j � 	� 
� q ٗ �c B� έ �p h � ި ��  � !�g "�~ #�c $4� %k� &+� 'V� (0q 0rl 1G� @W� A�� Qe� R� S�y T�� U�n V�h W4u X�] `.] a�d bO` c� p7� �ʚ �X� �\� �ʻ ��w �C_ �|� �:� ��� ��g ��� �� �}u �r� � �C� �� �;� � � �m� �w� ��� �� ��� �� �tg ��� �� ��� �]� ��w �G� �� �8� �ț �fo �tz ��_ �,� ��l �Ҫ ��� ��e ��o ��^ �� � +s ) C  %�F  ,�� p)"^G  1x1 )$c   1x2 )$c  1t1 )%c  1t2 )%c  
�� )&c   
�g )&c  (
x )'c  0
yk )'c  81w0 )(c  @
6� )(c  H
�� )(c  P
p )*�  X
9� )+c  `
Pk ),�F  h
g )-�F  l H� )/�F  �b )/vG  �F  _�B  %		@�H     	M� *N.  R�G  :	 �H     ( 0  �G  Q %�G  	� $!�G  	�{ $'�G  	L~ $-�G  	�j $3�G  	 c $9�G  	�� $@�G  	{ $F�G  	�� $L�G  	�� $R�G  	n_ $X�G  	�q $^�G  	�� $d�G  	� $j�G  	�� $p�G  	u� $v�G  	\_ $|�G  	�c $��G  	� $��G  	\e $��G  	@m $��G  	�� $��G  	�� $��G  	b $��G  	,� $��G  	�y $��G  	�^ $��G  	� $��G  	�� $��G  	]n $��G  	� $��G  	� $��G  	�� $��G  	�� $��G  	� $��G  	U� $��G  	h $��G  	K� $��G  f� $�G  �� $�G  �� $�G  6� $�G  � $�G  k� $ �G  �f $&�G  �w $,�G  �w $3�G  �� $:�G  � $@�G  5� $G�G  �� $M�G  �_ $S�G  � $Y�G  I| $a�G  7� $g�G  ӟ $m�G  �� $s�G  �� $}�G  	�� $!�G  	U� $'�G  	�� $-�G  	Be $3�G  	յ $9�G  	�e $@�G  	z $F�G  	� $L�G  	�t $R�G  	!k $X�G  	�~ $^�G  	� $d�G  	� $j�G  	!� $p�G  	�s $v�G  	�� $|�G  	Ԓ $��G  	3p $��G  	�r $��G  	� $��G  	O� $��G  	w� $��G  	� $��G  	*b $��G  	m� $��G  	(� $��G  	w� $��G  	�� $��G  	ܝ $��G  	�� $��G  	I� $��G  	x $��G  	מ $��G  	#� $��G  	�� $��G  	޺ $��G  	�� $��G  +{ $�G  � $�G  ;g $�G  Af $�G  
� $�G  �i $ �G  �� $&�G  �� $,�G  c� $3�G  S� $:�G  �� $@�G  z� $G�G  m $M�G  k� $S�G  �p $Y�G  �k $a�G  �� $g�G  � $m�G  �y $s�G  Tu $}�G  	| +N.  S5  	��H     _5  	��H     k5  	@�H     w5  	 �H     �5  	��H     �5  	��H     �5  	@�H     �5  	 �H     �5  	��H     �5  	��H     �5  	@�H     �5  	 �H     �5  	��H     �5  	��H     �5  	@�H     6  	 �H     6  	��H     6  	��H     +6  	@�H     76  	 �H     C6  	��H     O6  	��H     [6  	@�H     g6  	 �H     s6  	��H     6  	��H     �6  	@�H     �6  	 �H     �6  	��H     �6  	��H     �6  	@�H     �6  	 �H     �6  	��H     �6  	��H     �6  	@�H     �6  	 �H     7  	��H     7  	��H     7  	@�H     )7  	 �H     67  	��H     C7  	��H     P7  	@�H     ]7  	 �H     j7  	��H     w7  	��H     �7  	@�H     �7  	 �H     �7  	��H     �7  	��H     �7  	@�H     �7  	 �H     �7  	��H     �7  	��H     �7  	@�H     �7  	 �H     8  	��H     /8  	��H     ;8  	p�H     G8  	P�H     S8  	0�H     _8  	�H     k8  	��H     w8  	��H     �8  	��H     �8  	��H     �8  	p�H     �8  	P�H     �8  	0�H     �8  	�H     �8  	��H     �8  	��H     �8  	��H     �8  	��H     �8  	p�H     9  	P�H     9  	0�H     9  	�H     +9  	�H     79  	пH     C9  	��H     O9  	��H     [9  	p�H     g9  	P�H     s9  	0�H     9  	�H     �9  	�H     �9  	оH     �9  	��H     �9  	��H     �9  	p�H     �9  	P�H     �9  	0�H     �9  	�H     �9  	�H     �9  	нH     :  	��H     :  	��H     :  	p�H     ':  	P�H     3:  	0�H     ?:  	�H     L:  	�H     Y:  	мH     f:  	��H     s:  	��H     �:  	p�H     �:  	P�H     �:  	0�H     �:  	�H     �:  	�H     �:  	лH     �:  	��H     �:  	��H     �:  	p�H     �:  	P�H     ;  	0�H     ;  	�H     ;  	�H     );  	кH     6;  	��H     C;  	��H     P;  	p�H     ];  	P�H     j;  	0�H     w;  	�H     �;  	�H     �;  	йH     �;  	��H     �;  	��H     �;  	p�H     �;  	P�H     �;  	0�H     �;  	�H     �;  	�H     �;  	иH     <  	��H     <  	��H      <  	p�H     -<  	P�H     :<  	0�H     RG5  
M	 �H     R#8  
[	 �H     RW<  
i	`�H     R;M  u	 �H     _�@  �	�H     ,̀ x,%cV  
�  ,(t   
9� ,)�3  
  ,,�*  
N ,-<,  
#(  ,.    
[� ,/3	  (
[k ,0�  H1pp1 ,1�  X1pp2 ,2�  h r ,5�U  }� ,5{V  �U  �q -��V  �  -�t   ?map -�c<   �d -��V  R� -��V  �  -�t   �� -��   �s -��V  n)  .�V  W  &�  !W  J  Q  �      �)  .$-W  3W  &�  LW  J  Q  a    nk  .)]W  %LW  ,�;  .)�W  
�=  .+�V   
z+ .,!W   9�� �XW  	��H     (�   �W  -S    %�W  9�� ��W  	��H     q� =�   	��H     +5  F	 �H     )�G  /; 	�H     ){J  /A 	 �H     )�G  /H 	��H     )�J  /S 	 �H     )�G  /l 	�H     )�J  /s 	�H     )�G  /z 	аH     )�J  /� 	��H     )�G  /� 	��H     )�J  /� 	��H     )�G  /� 	��H     )�J  /� 	`�H     )H  /� 	@�H     )�J  /� 	0�H     )H  /� 	 �H     )�J  /� 	 �H     )H  /� 	�H     )�J  /� 	ЯH     )'H  /� 	��H     )�J  /� 	��H     )3H  /� 	��H     )�J  /� 	��H     )?H  /� 	��H     )�J  /� 	p�H     )KH  /� 	`�H     )K  /� 	P�H     WH  / 	 �H     K  / 	�H     cH  / 	��H     #K  /* 	`�H     oH  /7 	P�H     /K  /= 	H�H     {H  /C 	 �H     ;K  /L 	�H     �H  /S 	 �H     GK  /] 	��H     �H  /c 	�H     SK  /k 	حH     �H  /q 	��H     _K  /x 	��H     �H  / 	��H     kK  /� 	��H     �H  /� 	��H     wK  /� 	@�H     �H  /� 	0�H     �K  /� 	 �H     �H  /� 	�H     �K  /� 	��H     �H  /� 	��H     �K  /� 	`�H     �H  /� 	@�H     �K  /� 	0�H     I  /� 	 �H     �K  /� 	�H     �H  /� 	ЫH     �K  /� 	��H     �H  / 	��H     �K  / 	p�H     I  / 	`�H     �K  / 	@�H     #I  / 	 �H     �K  /B 	��H     /I  /X 	`�H     �K  /` 	P�H     ;I  /f 	�H     �K  /x 	ШH     GI  /~ 	��H     L  /� 	��H     SI  /� 	��H     L  /� 	��H     _I  /� 	`�H     L  /� 	�H     kI  /� 	ЧH     +L  /� 	��H     wI  /� 	��H     7L  /� 	��H     �I  /� 	��H     DL  /� 	��H     �I  /� 	��H     QL  /� 	p�H     �I  /� 	`�H     ^L  /� 	P�H     �I  /� 	@�H     kL  /� 	0�H     �I  /� 	 �H     xL  / 	 �H     �I  /	 	�H     �L  / 	�H     �I  / 	ЦH     �L  / 	��H     �I  /# 	��H     �L  /* 	p�H     �I  /2 	`�H     �L  /8 	@�H     �I  /A 	0�H     �L  /G 	 �H     J  /R 	�H     �L  /X 	��H      J  /b 	��H     �L  /h 	��H     J  /q 	`�H     �L  /w 	P�H     -J  /} 	@�H     �L  /� 	0�H     :J  /� 	 �H     �L  /� 	 �H     GJ  /� 	�H     M  /� 	��H     TJ  /� 	��H     M  /� 	`�H     aJ  /� 	P�H     !M  /� 	 �H     nJ  /� 	 �H     .M  /� 	�H     (�F  ^`  -S   ? %N`  Ah� 	-^`  	�H     Z�[ 	��a  !k 	�%jG  !  	�%�*  `dim 	�%�<  !�� 	�%�  !� 	�%!-  dh  	�\@  �  	��<  �{ 	��  v 	�c  *nn 	�  2]  	�  �j 	�#  *X1 	�  *X2 	�  *w 	�  �� 	��F  �k 	��=  #]a  *X 	�   #pa  �� 	Z    #�a  ,� 	.�  4� 	/c  xx1 	0c  xx2 	0c   p 	`�  9� 	ac    VVi 	H�;D     �      �d  Nk 	H.jG  UN�� 	I.�  T+� 	J.c  Z_ T_ axx1 	K.c  �_ �_ axx2 	L.c  �_ �_ +�� 	M.�F  &`  ` N�k 	N.�=  � N�j 	O.  �1x 	Q  z` r` k 	Q  $a "a � 	Q%  Sa Ga :nn 	R  b b A�� 	Sd  ��}   c  �� 	]c  bb Xb �g 	^c  Dc 8c :w 	_c  6d 0d  3�<D     h       �c  :len 	yc  �d �d :y0 	zc  
e �d :y 	{c  *f  f :idx 	|  }g wg r��  �<D      ` 	z��  �g �g ��  �g �g ` ��   h h  �  ch _h    � :idx 	�  �h �h � F� 	��F  i i �� 	��F  �i �i    (�F  d  -S   @ b�v ��  �d  N �(<,  א �(a   4idx �(-   �  �(�d  ��  �(�d  �  �t  �^ ��   �  sM� iQ  @�D     �      ��e  Gp i+Q  �i �i N j+<,  *k $k א k+a   �k vk .� l+�e  l 
l �  nt  �l �l ch o�  m m ��  o�  n �m buf p�e  `o To   6 ze  ȳ  v�  �o �o   @6 �e  ȳ  {�  dp Xp  W��D       -   �  tǅ ^�e  �  ^#t  4buf _#a   R�  a]   b?� Pa   0f  �  P"t  � R�  R�  S]  buf T�e   bl� A�  wf  9� A+�3  Nh B+�3  �� C+c<  B� D+    @�~ ��  �|D     �      ��q  ~ �+5  q �p  �+�  �q �q �  �+H   r r �^ �+�  mr Yr :1  �+C  Vs Ls � �  �s �s R�  ]  <t 4t 9  (�q  ���9��  )�q  ���,y  @}D      `# 1�p  my  �t �t ay  �u �u Uy  qv gv Iy  �v �v =y  �w �w `# yy  
x �w �y  
y y �y  ]y Wy �y  �y �y �y  �y �y �y  �z �z �y  { { "�y  ����y  P{ B{ h�y  @�y  �{ �{ �y  *| "| B	z  ��D     Bz  D     |  �}D      �# 0�h  8|  �| �| ,|  �| �|  |  } } �# D|  M} E} :�D     _�  Uv T�șQ���   ��  �}D      �# @�i   �  �} �} -�  ~ ~ �  e~ _~ �  �~ �~ �# :�   �~ G�  � � T�  K� C� a�  i� a� "n�  ��B{�  ��D     .��  0$ ��  )� #� Y�D      �i  U���Q�� X��D     �i  U��� X؁D     �i  U��� �D     ) U���    '�z  p$ �k  "�z  ��"�z  �����  !D      �$ pj  ��  z� x� ��  �� �� �$ ��  ҂ ΂  �  � �   ��  BD       % �j  ��  R� P� ��   % ��  z� v�  �  �� ��   ��  '�D      0% 2k  ��  �� �� ��  "� � 0% ��  ^� Z�  �  �� ��   ��  W�D      `% A#jk  ��  ބ ܄ ��  � � `% ��  -� )�  �  p� l�   �D     5 �k  Uv  ��D     A �k  Uv Q0 ��D     N �k  Uv T}  ��D     [ U���T}   �z  2�D      �% ��n  {  �� �� {  � � {  #� � �% *{  e� a� 6{  �� �� B{  �� � N{  I� G� Z{  �� �� "f{  �ؘ"r{  ���~{  � � �{  a� [� �{  �� �� "�{  ��B�{  �~D     '�{  �% lm  �{  � � �{  6� 4� C��  \�D      & �0m  ��  [� Y� ��  �� �� & ��  Ɖ   �  	� �   \�D     ��  Tm  8�w  ���8�w  v  ��D     h T���  5�{  ӃD     �       Wn  �{  F� D� �{  s� q� C��  �D      @& ��m  ��  �� �� ��  ي ׊ @& ��   � ��  �  C� ?�   �D     ��  n  8�w  ���8�w  v  -�D     h 3n  T��� w�D     h U�Șv T�Ș  ��D     h zn  U�B$T�Ș X�D     �n  U T���Q�ؘ ��D     u �n  Uv  ӄD     N Uv T���   'z  �& 'o  " z  ��&�D     � o  U���  �D     [ U���T���  ��  ��D      �& �}o  ��  �� ~� ��  �� �� �& ��  ы ͋  �  � �   '.z   ' #p  3z  Q� O� @z  v� t� Mz  �� �� Zz  �� �� gz  � � tz  � � �z  N� J� �z  �� �� H�z  0�D     @       �z  H� F� �z  m� k�   5�z  ��D     P       Wp  �z  �� �� �z  �� ��  Xs~D     sp  U T��� X�~D     �p  U| T  �~D     � �p  Uv Tw � y�D     A �p  Us� u�D     Uw �T| Qv R    ]�  }D      0' ."q  x�  � �� k�  � �  Q|  2}D      �' /Xq  j|  ,� *� ^|  S� O�  �{  ��D      �' 4�q  |  �� ��  ƀD     S�  U|   (�@  �q  -S     (cV  �q  -S     =+� ��;D            ��q  D~ �"J  U @�s ��  @;D     H       �-r  D~ �"J  U~ �5  �� ��  @�� ��  pbD     
       ��r  ~ �"J  ߏ ۏ ;  �"Q  � � OzbD     � U	��H     T�T  @�q K�  �D     �      �'u  ~ K!J  e� U� n  L!Q  � � �\ M!a   _� ;� � O�  ڒ Β ~ P5  p� `� �� Q�  3� !� B� R�  	� �� �{ T   ߕ ͕ 3 �D     !       �s  ZX Z"'u  �� �� 99� ["�3  �h0�D     �v  T�hQ�U  3 �D            �s  val f-u  �� �� Nh h�3  1� /�  3T�D            )t  val q-u  m� i�  3p�D     (       t  ZX z!3u  �� �� 99� {!�3  �h��D     �v  T�hQ�U  3e�D            �t  val �9u  � ��  3��D     @       �t  X;  �?u  � � val �?u  0� ,�  $�D            �  �   h� f� val �9u  �� ��   �V  �  �V       Pق y�  �v  !~ y!J  !n  z!Q  !�\ {!�  !�R  |!   � ~�  ~ 5  #�u  �� �-u  *ss ��  Nh ��3    #�u  B� �-u   #�u  ZX �!3u  9� �!�3   #v  *s �Q  *w �@    #%v  �{ �9u   #�v  X;  �?u  *x1 �  *y1 �  *x2 �  *y2 �  *x3 �   *y3 �$  *x4 �(  *y4 �,  *dp �	5  *s �Q  *ep ��   *i �Z     #�v  s /Q  nsd 0@    �  ;9u    S$� J�  ��D     f       �w  +�  J2t  �� �� +p� K2w  8� ,� +~ L25  Ǚ �� � N�  D� <� A9� O�3  �XڈD     _�  T�X  �3  E�� WC  ,y  ��  W+oV  �  X+t  ��  Y+c  ~ [5  :  ]s  :� ^�  ?� ^�  � _�  �} _�  �� _1�  �� _>�  Ŷ `  x1 a  y1 a  x2 a  y2 a  x3 a   y3 a$  x4 a(  y4 a,  I�r �I�r �I�� �#�x  G� �  �� �  x �   #y  G� �  �� �  x �   G� �  �� �  x �    P�t ��  �z  !��  �$oV  !~ �$5  !�  �$t  !�^ �$�  !:1  �$C  � ��  �  �H  =� ��   ��  �� �	  �V  ��    ��*  �m �,  �d �<,  � ��  Nh ��3  | �S.  I�u  JI�� #.z  :e �3	   #�z  �i �c  w� �c  �� �#c  �] �c  �� �c  dh  �\@  ~ ��>  ~ ��>  x� �c  ]� �c    #�z  x� �c  ]� �c   �!  �  o� �    P\� Z�  �{  !��  Z6oV  !�  [6t  !�d \6<,  � ^�   `�  9� a�3  | bS.  4  d�{  { fc  �m gc  -� i   	Y  l�  ?� m�  �j o3	  [�u  �#�{  yi ��  o� �)�   F� ��  x� �)�    �  Z�� I|  !��  IoV   P�� ,�  Q|  !��  ,oV  !~ -5  !�  .t  � 0�   Ze  w|  !��   "oV  !  !"�*   E�� ��  }  �^ �*�    �*�*  �S  �*}-  N �*�B  � ��  dim �Z   dh  �$B  J�u  �D     k �^G  �� ��  � �c    7`{ p�    p'�*  4dim q'�<  dh  s\@  �y t�>  M� u�>  � v�  c� w�>  YK  x�>  N� y  Nh �3  � ��0  � �   #~  �� �*  ~ ��>  ~ ��>  � �?  �t �?    #  ~ ��>  #�~  �b c  �� c  $� &c  �} c  �;  c  	*  #c  � +c  �� 2c   (� Vc  �b Vc  �� V#c  $� V/c  �} Wc  �} Wc  ؊  W%c  �k  W-c  � nc  �� nc     #z  ~ ��>  ~ ��>  F~ ��>  *� �c  �� �c  �� �c  � �$c   � c  AT  :�>  ;  :�>     7"� X�    X-�*  2�  Y-�>  	s Z-�>   =ڀ 9jD     I       ���    9.�*  �� �� Gdim :.�<  � �� ڣ ;.�>  6� 2� .� <.�>  u� o� ��  >c  Ǜ �� �� >c  � � ^� ?c  \� Z� NjD     `�  Q�T8��  �U  EI� t
c  ��    t
/�*  4dim u
/�<  ��  v
/c  �� w
/c  �� x
/�  >| y
/�  N {
�B  dh  |
$B  ��  }
c  �b ~
  �(  
  Ik� .#��  � �
c  �� �
c  :� �
�     |�  �
c  � c     vDy C
c  ,�  �q C
"*  .� D
"�  ��  E
"c  n G
�  mi H
c  �m I
c  ��  J
c  w O
c  ��  P
c    @Ԏ �	�  p:D     �       ��  D  �	)�*  UDN �	)�B  T�� �	�  �� � �x �	P  ՜ Ϝ ;� �	#P  &�  � �  �	t  w� u� ;*�  x:D      � �	8�  �� �� 8�  �� �� E�  �� ��   7�{ x	�    x	7�*  N y	7�B  dh  {	\@  c� |	�>  M� }	�>  Nu ~	$B  �� 	�  bb �	�  �| �	*  � �	   S� �	c  �� �	AA  � �	   �� �	$   �� �	5   ��  �	c  �� �	        E� a	�  H�    a	2�*  �� b	2�  �q c	2H�  4dim d	2�<  � f	�   s*  @2� ��  �VD     5      ���    �0�*  � � Gdim �0�<  � u� dh  �\@  �� � �  �  v� n� R�  ]  � ՟ � $B  �� � Nh �3  � 	�0  � � �    E� =� �k �=  �� �� �� �=  �� �� seg �=  Y� C� �� �  >� :� k c  �� u� �� c  � � H� c  m� g� J�u  Y	�XD      � �  ;�  S�>  �� �� ee T  �� �� 3`XD     )       <�  c� g�>  !� � ��  hc  s� m�    9c� x�>  ��F��  YD      YD            ���  ��  ��  ѥ ͥ $YD            ��  � �  �  u� q�   �XD     ֹ  U��R���X��Y��   3iYD     i       W�  ;�  ��>  �� �� ee �  � � P c� ��>  -� '� ��  �c  � y�    � W�  �y ��>  ۧ ٧ M� ��>  � � c� ��>  R� J� � ih �  ƨ �� �� �  � � � s �   f� `� @ ~ 	�>  �� �� ,� 	�=  � � $�ZD     :       t� 	c  �� �� Kc 	c  �� ��      ��  �WD      p I��  ��  ۪ ٪ ��   � �� p ��  <� 8�  �  � {�   `WD     h ň  U@ uWD     h �  U Ts  �WD     h Ts   =G� r�8D     �      ���    r0�*  �� �� �� s0�  �� �� �q t0H�  8� 4� Gdim u0�<  u� q� dh  w\@  �� �� �k x�=  5� 3� �� y�=  Z� X� � zc  �� }� B� z"c  � �� w�d z-c  ��N  z9c  Q� O� �� {�=  z� t� ,� {�=  Ǯ î   �} �c  � �� �} �c  O� G� ` min �c  ί ʯ max �c  /� +� len �c  �� �� � ��  �c  �� �� � �c  � � F� �#c  4� 2� � � �c  [� W�      @q� ��  �ED     �	      �s�    �3�*  �� �� Gdim �3�<  � � N ��B  {� y� dh  �\@  �� �� R�  �]  �� x� � ��  �� � zx  ��=  � �� 9� �l?  ��~� ��@  n� ^� �� ��@  &�  � �� ��<  {� s� �e �!�<  �� ۷ �� �c  %� � J�u  iLD     3�FD     "       y�  oI ��<  x� r� �� ��<  ȹ Ĺ  3tOD     ,       ��  oI ��<  '� � �� ��<  �� ��   0 ��  oI ��<  Ϻ �� k� ��<  �� �� �� �Z   ;� � ,` c  �� �� �s c  ʾ �� �a c  ۿ Ϳ Li c  �� v� � s  �� �� 0� s  Z� B� �l 	c  t� ^� E 
c  y� a� Џ    �� y� 1t �=  ~� n� '` c  2� (� �s c  �� �� �a c  \� @� Gi c  �� �� � s  �� �� +� s  J� ,� �l c  �� �� @ c  �� �� � u 2c  =� 1� v 2c  �� �� ;E�  0ID       n�  c� W� b�  � � V�  �� ��  "z�  ��~��  �� �� B��  OD     .��  � ��  �� �� ��  � � ��  �� �� {JD     � c�  U��~TPY��~ �ND     � U��~TPQ0X0      $�MD     �       �k <�=  E� C� ^� =�=  j� h� @ N� B�<  �� �� k� C�<  � � �x Dc  R� F� q� Ec  �� �� 3 ND     &       K�  p J�<  :� 6�  $LND     &       p Y�<  {� w�     =�� ��8D            ���  DN �2�B  UD�m �2!-  TD{ �2!-  Q =� ��`D     <       �N�  N �,�B  �� �� �m �,*,  '� � �`D     N�  ,�  Us Tv Q0 O�`D     N�  U�UT�TQ1  =-� \ \D     U      �ӕ  N \0�B  �� �� �m ]0*,  M� E� Gdim ^0�<  �� �� �� `�  w� m� � ac  �� �� dh  b$B  6�  � nn c�  �� ��  � ��  �x ~$B  �� �� �� AA  ?� 9� � ��  �c  �� �� A�  �c  �� �� � �c  � � �� ��  P� L� :� ��  �� �� 3�_D     �       _�  � �c  �� �� ��  �c  T� P� ,� ��  �� �� ��  !`D      ` �J�  ��  �� �� ��  � � ` ��  8� 2�  �  �� ��   �_D     � U   ;��  �]D     	  ���  �� �� ��  �� ��  ��  !� �  �  d� `�      � 4�  ��  �*  �� �� M��  ]D      ]D            ���  ��  �� �� $]D            ��  �� ��  �  1� -�       =�  �� AA  ��  c   @ v�  �k  +c  n� l�  ��  �^D       � Ĕ  ��  ��  �� �� � ��  �� ��  �  (� $�   ��  %_D      � %��  ��  ��  � ��   �    ;��  _D      P  ��  ��  P ��  g� c�  �  �� ��    3u_D     K       ��  �� gAA  i h�  $�_D     '       b rAA    ;��  1]D      � ��  ��  �� �� � ��  � �  �  J� F�    @ȹ D�  @�D     M      ��  N D+�B  �� �� �  E+t  �� �� gm G�  [� S� �  ��D      �@ P��  8�  �� �� +�  �� �� �@ E�  � � R�  �� �� "_�  ��l�  �� �� y�  T� P� "��  ����  �� �� �e  ��D      �@ .�  �e  �� �� �@ "f  ��f   � �� "f  %� #� ��D      T8Q��   '��  @A 0�  ��  L� H� "��  ��Fd  #�D      #�D            $�  ed  �� �� Xd  �� �� Kd  �� �� >d  �� �� 1d  $� "� $#�D            rd  I� G� d  q� o� @�D     � T~ Q
R��   �D     �d  U Tv Q| R��  M�e  k�D      k�D            ;�e  �� �� �e  �� �� $k�D            �e  �� �� z�D     ) T|      w�D     � Ę  Us Tcinu ��D     � �  Us T�� ��D     ��  �  Uv Ts  ��D     Й  Uv Ts   7޻ 	��  N 	3�B  �  
3t  "�    V�    �  �  ρ �  R\ a   ]� ˙  p Q  �^ �  � -     (�   ˙  -S    %��  =R� 7p�D     �      ��  N 71�B  	� � �  81t  E� A� 9�� :�  ��y9E� ;�  ��|�� =�  �� }� A� >�  B� 2� �� @AA  � �� � A�  �� �� dh  B$B  �� �� �S  C�  =� )� sc E�3  )� '� bss G�)  U� M� bs H�  �� �� �� Jc  (� $� R\ La   h� `�  �< k�  p ZQ  �� �� �� [!-  �� �� � \!-  �� ��   ]c  a� M� �  ^c  H� 4�  @= g�  �^ ��  � � ��  ��  N� @� ]� �  � �� T� �!  � � p �5  �� �� �  ��  >� �c  �� �� �i �   Z� L� i �-   � �� 9� �-   ��x �= B�  y� �c  �� �� �o  �   �� ��   > �  nn �  �� �� N� �  �� �� k� �  _  Y  P> Y� �  �  �  pp �  �  �     �> ��  �q +c  � � �� ,  � � �@ ,  � � ,� -   � �� -)  � � �� .   � �r .*  � x ��  /c  )
 �	 ? �� �c  � � P? �\ �c  N� �  � � k� �  d R hit �   1  � �  � � '] �  c Y �� �   � � �? l2r �    � d �c  m _     Fd  ��D      ��D            �(�  ed  t r Xd  � � Kd  � � >d  � � 1d    $��D            rd  6 4 d  a _   йD     � U~ Q1  S�D     �d  T��wQw R��x  3��D     :       ��  ref �c  � � #� �c  � � U� �   � �  i��  ǿD     r       ��  ��  ��  $ǿD     r       ��  $  ��  ��  r p   j��  9�D     s       ���  ��  $9�D     s       ��  � � ��  ��  � �     �? "�  i ��  9�x ��  ��x �@ ��  a �!-  < 6 b �!-  � �  x�  @ �2�  %�  @ ?�  � � J�  * ( U�  .b�  @@ c�  Q M n�  � �     �e  ϸD      �< V~�  �e  �< "f  ��|f  "f  � � ԸD      T8Q��|   M�e  λD      λD            ��e  � � �e    $λD            �e  5 3 �D     ) Tw     (c  �  -S   2 *  (AA  �  -S   	 7�} {�  .� &�  >) &{�  i �  j �  �8  AA  a c  b c    AA  V�� =�D     Z      �~�  +N =2�B  f ^ +�  >2t  � � A  A�q  ���|[�u  � �: 4�  � P�  J D �^ Q�  � � :dim RZ   	 � A��  S~�  ���}�m T*,  � � Nh Z�3  � � � [�0     R\ ^a   � � :p _Q  � � 3��D     B       {�  A� r-   ���}kd  ̵D      ̵D            �R�  ed  8 6 Xd  8 6 Kd  8 6 >d  ^ \ 1d  � � $̵D            rd  � � d  � �   ��D     �d  Us Tv Q| R���}    < z�  dh  �$B  � � �\ �\@  S O :seg ��=  � � �� ��=  � � ʊ �#�=   u A� ��  ���| 0< �  ��  �c  � �  ��D     ��  5�  U} Ts  ��D     ��  ]�  U} T0Q0Rs  ?�D     ��  U���|Tt    p< ��  dh  �$B       3� �c  �  �   C�e  y�D      P; f�  �e  #! !! P; "f  ���}f  H! F! "f  m! k! ~�D      T8Q���}   C�e  յD      �; ���  �e  �! �! �e  �! �! �; �e  " " �D     ) w�  T|  h�D     ) T|    C*�  a�D      �; �Ϧ  8�  F" B" 8�  F" B" E�  ~" |"  ��D     � �  U~ T Q1 %�D     � �  U���}T0Q
�� y�D     ��  U} Ts�  C]�  5�D       �: Ji�  x�  �" �" k�  �" �"  �D     S�  U}   (|B  ��  -S     ywq `��  !N `0,D  !�m a0!-  !{ b0!-   S�� R�  ��D            �\�  +�^ R(�  # # +  S(�*  E# A# +�S  T(}-  �# ~# +N U(,D  �# �# O��D     K�  U�UT�TQ�QR�R  S� I�  �8D            ���  N  I'�*  U+N J',D  �# �# O�8D     ��  Uu T�T  VX� @�VD            ��  +N @*,D  9$ 5$ +�m A**,  v$ r$ O�VD     �  U�UT�T  S�� $�  ��D     l       ���  +N $),D  �$ �$ +�  %)t  % % gm (�  �% }% ȴD     � ��  Us Tcinu �D     � ��  Us T|  ��D     ��  ک  Uv Ts  
�D     ' Uv Ts�8%�  s   7� ch�    c,�*  4dim d,�<  �� e,�  � f,c  �  h�<  �a i�<  oI j�<   =Õ ��sD     P      ��    �4�*  �% �% Gdim �4�<  @& 6& �  ��<  �& �& (� ��<  ' ' � ��@  p' f' �� ��@  �' �'  | ��  '( ( oI ��<  �( �( �k  ��<  "+ + c+  ��<  w+ k+ J� LtD     J�� <IuD     `" 4w  	�<  b 	 �<  , �+ �  �uD      �" 8	,�  ?�  x, t, 2�  �, �, &�  �, �, �  �" L�  W�  b�  n�  z�  ��  ��  ��  vD     ��  Rv    F�  RuD      RuD     ;       Dܬ  ?�  *- (- 2�  Q- M- &�  �- �- �  $RuD     ;       L�  W�  b�  n�  z�  ��  ��  ��  yuD     ��  T| Q��Rs    F�  �uD       �uD     5       H��  ?�  �- �- 2�  �- �- &�  �- �- �  7. 5. $�uD     5       L�  W�  b�  n�  z�  ��  ��  ��  �uD     ��  U~ Ts�Rs    M��  HvD      HvD     T       ?	�  ^. Z. Ԯ  �. �. Ȯ  �. �. $HvD     T       �  �. �. ��  y/ u/     7N� ���  4p1 ��<  4p2 ��<  1v  ��<  zf  ��<  p ��<  u �c  v1 �c  v2 �c  u1 �c  u2 �c  d1 �"c  d2 �&c  �� ��    7k\ ��  4p1 ��<  4p2 ��<  4ref ��<  p ��<  � �c   =p� ��QD     �      �h�    �6�*  �/ �/ Gdim �6�<  �/ �/ �  ��<  [0 Y0 (� ��<  �0 0 dh  �\@  �0 �0 �y ��>  e1 a1 M� ��>  �1 �1  | ��  �1 �1 Jd� k5SD     � oI ��<  (2 $2 c� ��>  p2 ^2   u  c  O3 ;3 ou  c  '4 4 fu  c  �4 �4 � c  �4 �4 0 min -�  �5 �5 max -�  6 �5 mid -!�  �6 �6 dh .c  ,7 $7  p ٰ  nn 9�  �7 �7  � AT  ]�>  �7 �7 ;  ^�>  ��  SD      � fV�  ��  68 48 ��  [8 Y8 � ��  �8 �8  �  �8 �8   WXTD     h      7_� �5�    �4�*  4dim �4�<  dh  �\@  �k ��=  �� ��=  seg ��=  #��  c� ��>  oI ��<  N� ��<  k� �!�<   c� ��>  oI ��<  N� ��<  k� �!�<    7�� z��    z'�*  �S  {'}-  oI }�<  �� ~�<  vec �  tag ��    @* ��  p=D     m      �*�    �)�*  9 9 �S  �)}-  �9 �9 9� ��  ���  ��<  �: �: �<  ��  0; "; �:  ��  �; �; �� ��  ?= 7= �� ��  �= �= ͩ �c  > > =�  �c  �> �> R�  �]  _? Y? J�u  r�@D     J�a H�DD        Ʒ  oI D�<  �? �? (� E�<  �@ �@ U�  H�  zA tA �x I  �A �A  ` W�  vec N�  tB nB tag O�   �B �B �� Pg  C C end Q�<  �C �C �� R�<  AD /D ^� S  E 
E � bX  Xc  rE pE hX  Xc  �E �E ��  �?D        `"�  ��  ��    ��  �E �E  �  7F 3F   ;��  �?D      ` a"��  ��  ` ��  vF rF  �  �F �F      � ��  � ��@  �F �F �� ��@  hG ZG end ��  H �G idx �5  kH cH  $�AD     �      �t �  �H �H � ��@  I I �� ��@  mI gI  � ��  N� ��<  �I �I �@ ��<   J J �� ��<  uJ iJ �o �!�<  K �J bX  �c  �K ]K hX  �c  �M �M   L� ��<  ;��  �BD      � ���  P P ��  �P wP � ��  Q Q ��  IQ EQ ȹ  �Q �Q      � ��  oT   c  �Q �Q n/   c  ZR VR bX  !c  �R �R hX  !c  bS ^S ,p #�<  �S �S Rx $�<  �S �S    ,p U�<  T T Rx V�<  ?T =T WAED     �    1>D       ޷  U~  `@D     � �  Uv T8R Y�� �@D     � Uv TPY��  7�m �S�    �,�*  N �,<,   =�f ��`D     "      �]�    �'�*  hT bT R�  �]  dim �Z   �T �T 3�`D     �       0�  dh  �\@  U U �`D     ) �  Uv  aD     ) �  Uv  HaD     ) �  Uv  yaD     ) Uv   �aD     ) H�  Uv  �aD     ) Uv   7�| ���    �'�*  R�  �']   E�� e�<  ֹ  4dx e!c  4dy f!c  ll hc  ss hc  dir i�<   S�� c�  �OD     8      �?�  +dh  c)\@  nU ^U +dh d)  !V V adir e)�<  �V �V +� f)   KW ;W +R�  g)]  
X �W +:� h)?�  �X �X A� j�  ��c� k�>  �Y �Y �y l�>  IZ GZ z�u  �vPD     p �<  y  wZ mZ �:  z  �Z �Z -� {  �[ �[ QD     � �  TXY�� |QD     � TXQ0X0Y��   �>  Pm` &�  ��  !dh  &,\@  !R�  ',]  !} (,��  � *�  zx  +�=  [�u  Y�<  8  �:  9  -� :    �=  E�o 
�   ��  9� 
�-�3  n�  
�-�   Eޤ 
��  ��  9� 
�2�3  n�  
�2�  �� 
�2�  K� 
�2��  N 
�<,  ��  
�,3  | 
�S.  Nh 
��3  � 
��  I�u  
�R�  
�]    <,  {z 
��aD     }       �_�  9� 
�)�3  �[ �[ � R�  
�]  W\ S\ nn 
��  3bD     :       H�  Nh 
�"�3  �\ �\ | 
�"S.  �\ �\ GbD     ) U|   OlbD     ) T�U   @�] 
P�  �yD     ?      �s�  �  
P)t  ] ] p� 
Q)w  s] k] ~ 
R)5  �] �] |� 
T�   R�  
U]  T^ R^ 9� 
V�3  �^ y^ J�u  
|�yD     s�  ezD      0# 
s]�  ��  �^ �^ 0# ��  _ _ ��  X_ T_ ��  �_ �_ ��  �_ �_ ��  %` ` ��  x` r` ��  �` �` B��  w|D     5��  �zD     4      ��  ��  �` �` ��  a a �  Ra Ja 5�  {D     k       J�  �  �a �a "$�  �� {D      .�  Uv T�� p{D      Uv Q��  H1�  �{D     }       2�  Lb @b ">�  ���{D      ��  Uv T~  |D      Uv T~ Q��   5^�  P|D     !       ��  c�  �b �b [|D      Uv T|   5q�  �|D     :       �  r�  �b �b  �zD     � ?�  Uv Tcinu �|D     � Uv T��   �yD      Q��  P� 
��  ��  !9� 
�;�3  � 
��  �  
�t  �� 
��  �� 
�c<  *ss 
��  *i 
��  |� 
��  I�u  
#L�  Nh 
��3  � 
��0  �a  
�%0  #1�  �j 
��  n�  
��   �j 
��  n�  
��    #^�  Nh 
��3   #q�  n�  
�   nn 
�    P�� )�  ��  !�^ )(�  !  *(�*  !�S  +(}-  � -�   S�� �  @8D     3       �K�  N  )�*  UNN )<,  T}*�  @8D      @8D            8�  c c 8�  c c E�  @c >c   E}� ��  ��  �^ �&�    �&�*  �S  �&}-  N �&,D  � ��  dim �Z   J�u  	z�D     k 	^G  �� 	�  � 	c    7� v��    v,�*  4dim w,�<  dh  y\@  �y z�>  M� {�>  c� |�>  �� }   seg ��=  #p�  oI ��<   � �c  oI ��<      7L� ���    �%�*  4dim �%�<  dh  �\@  �y ��>  M�  �>  � �  c� �>  YK  �>  � c  �}   �]    ^� c  I�u  i#p�  �� *  ~ �>  ~ �>   #��  ~ O�>   #��  ~ ��>  ~ ��>  F~ ��>  *�  c  ��  c  ��  c   AT  F�>  ;  F�>    @^l {c  @dD     \      ���    {'�*  kc cc c� |'�>  �c �c ~ }'�>  �d vd YK  ~'c  e 
e Gdim '�<  �e �e �b �c  'f f $� �c  �f �f �� �c  g �f �} �c  �g �g �} �c  �h �h ri �c  2j j � �c  Lk :k ͬ �c  Sl Kl � �%c  �l �l � �-c  am Qm x  �c  n n A�  �c  on en J�u  ��eD     �dD     �  Q�XR| v 8Z�  �U  7�� `��    `+�*  2�  a+�>  	s b+�>   7O� FH�    F,�*  4dim G,�<  ڣ H,�>  .� I,�>  ��  Kc  ^� Mc   E�� �c  ��    �-�*  4dim �-�<  ��  �-c  �� �-�  >| �-�  N �,D  dh  ��C  ��  �c  �b �  �(  �   Ik� ;� �c    @<� �c  �7D     w       ���  �q � *  �n �n .� � �  To Lo D��  � c  Qn ��  �o �o mi �c  �o �o �m �c  Mp Ep ��  �c  �p �p $�7D     "       w �c  q q ��  �c  <q 6q   @c M�  7D     �       ���  D  M%�*  UN N%,D  �q �q �� P�  �q �q �x QP  br Xr ;� Q#P  �r �r ;*�  7D      � T8�  Xs Vs 8�  Xs Vs E�  }s {s   =�� �p5D     �      �
�    �3�*  �s �s N �3,D  �s �s Gdim �3�<  t t dh  �\@  ]t Wt c� ��>  �t �t M� ��>  u u cjk ��C  Au =u �� ��  �u �u { �c  �u �u 3�5D           ��  bb �  Lv Jv �| *  tv pv S� c  �v �v � �� �B   w �v 0^    <w 8w �� (   �w �w $d6D     ~       ��  ,c  �w �w 3  -*  (x &x M��  �6D      �6D            ;��  ��  Mx Kx $�6D            ��  tx px  �  �x �x      ;��  �5D      ` ��  �x �x ��  ,y *y ` ��  ay ]y  �  �y �y    E�` ��  D�    �0�*  4dim �0�<  � ��   Eky ��  �    �.�*  4dim �.�<  dh  �\@  � ��  R�  �]  � ��C  �k ��=  �� ��=  seg ��=  �� ��  k �c  I�u  �#��  ;�  �>  mi c  ee   #s�  c� �>  ��  c  ʊ �=  ��  �=  �� !c  �� &�=      c� =�>    �y r�>  M� s�>  c� t�>  ih �  �� �  s �   ~ ��>  ,� ��=  t� �c  Kc �c        7�b 8�    8.�*  4dim 9.�<  dh  ;\@  �k <�=  �� =�=  �� >�<  �� ?�=  ,� ?�=  � @c  �| Ac  #��  ��  Sc  min Zc  max [c  len \c    �� ��=  � ��=  seg ��=  ʊ ��=      E�k �  ��    1�*  4dim 1�<  dh  \@  �k �=  �� �=  � �  seg �=  pt �<  k� �<  f0  �  f1 !�    =)r �P5D            ��  DN �.,D  UD�m �.!-  TD{ �.!-  Q =�� ��VD     C       ���  N �(,D  �y �y �m �(*,  Nz Fz �VD     ��  q�  Us Tv Q0 O�VD     ��  U�UT�TQ1  =2c ��TD     �      �	�  N �,,D  �z �z �m �,*,  { { Gdim �,�<  �{ �{ �� ��  �{ �{ � �c  �{ �{ dh  ��C  <| 2| nn ��  } }   �� ��B  ^} V} ��  �c  >~ :~    �  ؊  �c  �~ �~ �k  �c   �~ ��  �UD      0 ���  ��  5� 1� ��  o� k� 0 ��  �� ��  �  (�  �   �UD     h T   ��  8UD       0 �g�  ��  �� �� ��  �� �� 0 ��  ܁ ؁  �  � �   ��  wUD      p ���  ��  \� Z� ��  �� � p ��  �� ��  �  � �   ;��  �UD      � ���  (� &� ��  � ��  O� K�  �  �� ��     @ڔ m�  0�D     g       �
�  N m',D  Ճ ̓ �  n't  <� 4� gm p�  �� �� X�D     � ��  Us Tcinu g�D     � ��  Us T|  {�D     ��  ��  Uv Ts  ��D     ��  ��  Uv Ts  ��D     ' Uv Ts�8%�  s   7H� 2��  N 2/,D  �  3/t  "� 5   V� 5   �  6�  ρ 6�  R\ 8a   ]� ;˙  p <Q  �^ D�  � E-     =]q P�D     �      ���  N -,D  ݄ Մ �  -t  @� <� 96� �  ��y9�� �  ��|2� �  �� x� �� �  � � �	    �� �� �� !�B  v� n� � "�  ,� *� dh  #�C  U� O� �S  $�  �� �� sc &�3  �� �� bss (�)  Ȋ Ċ bs )�  � �� R\ +a   b� \�  �8 ��  p :Q  �� �� �� ;!-  A� 9� � <!-  �� ��   9 ��  �^ ^�  �� �� �� _c  ލ ֍ ]� `  L� <� �  a�  9� c-   ��x p9 �  nn �  �� �� N� �  <� 4� k� �  �� �� �9 pp �  � �   Fd  (�D      (�D            ���  ed  �� �� Xd  �� �� Kd  �� �� >d  �� �� 1d  � ߐ $(�D            rd  � � d  .� ,�   �D     �d  ��  Us T~ Q R��x ?�D     � U��xQ1  3B�D     ?       7�  ref c  S� Q� #� c  �� �� ��    �� ��  i��  �D     g       ���  ��  ��  $�D     g       ��  � � ��  ��  =� ;�   j��  ��D     k       ���  ��  $��D     k       ��  {� u� ��  ��  ɒ ǒ    �e  ��D      �8 6A�  �e  �8 "f  ��|f  "f  � � ��D      T8Q}    M�e  z�D      z�D            '�e  (� &� �e  M� K� $z�D            �e  t� r� ��D     ) T     V�� F�D     Z      ���  +N F.,D  �� �� +�  G.t  � � A  J�q  ���}[�u  � �6 f�  � Y�  �� �� �^ Z�  ڔ Ҕ :dim [Z   H� 8� A��  \��  ���~�m ]*,  �� �� Nh c�3  $�  � � d�0  _� [� R\ ga   Ȗ  :p hQ  � � 3s�D     B       ��  A� v-   ���~kd  ��D      ��D            ���  ed  w� u� Xd  w� u� Kd  w� u� >d  �� �� 1d   �� $��D            rd  � � d  � �   ��D     �d  Us Tv Q| R���~    8 ��  dh  ��C  6� 2� �\ �\@  �� �� :seg ��=  � � �� ��=  0� (� ʊ �#�=  �� �� A� ��  ���} 08 I�  ��  �c  2� 0�  |�D     ��  g�  U} Ts  ��D     ��  ��  U} T0Q0Rs  �D     ��  U���}Tt    p8 ��  dh  ��C  _� U� 3� �c  � �  C�e  Y�D      P7 oK�  �e  a� _� P7 "f  ���~f  �� �� "f  �� �� ^�D      T8Q���~   C�e  ��D      �7 ���  �e  қ Λ �e  � � �7 �e  F� B� īD     ) ��  T|  H�D     ) T|    C*�  A�D      �7 ��  8�  �� �� 8�  �� �� E�  �� ��  ԫD     � $�  U~ T Q1 �D     � J�  U���~T0Q
�p Y�D     ��  U} Ts�  C]�  �D       �6 S��  x�  � ߜ k�  � �  �D     S�  U}   ( D  ��  -S     V�� ��3D     �      ���  +.� �*-u  H� B� N>) �**  T+A�  �*c  �� �� :i ��  � � :j ��  �� �� n� ��  מ Ǟ ֺ �c  �� �� :sum �c   �� �8  �s*  � �  Zڑ ���  !.� ��  !>) �!-  *i ��  *j ��  �8  �c   P�6  �C  �  `a �C  `b �C  *ret �.  *tmp �.   <H�  �bD     �      ���  g�  �� s� t�  r� d� ��  � � ��  ?� =� Z�  Z�  ��  u� g� ��  $� � ��  � Ȥ ��  d� V� ��  � �� B��  �bD     '��    ��  ��  D� >�  .cD     ��  ��  Qq  PcD     ��  Qq   <5�  �fD     Q       �`�  P�  P�  C�  C�  ]�  �� �� j�  �� �� w�  ۩ ٩ ��   � ��  <��   gD           ���  ̀  7� #� ـ  2� � �  ͬ �� �  �� � \ �  � ��  ��  �  �� �� �  T� <� '�  C� � 4�  � ܲ A�  l� X� BN�  �gD     'W�  0 X�  \�  Ǵ �� .i�  ` j�  � � .w�  � x�  �� ��    .��  � ��  5��  �hD     8       ��  ��  L� F�  hD     ��  ��  Qq  �hD     ��  Qq    <��  `jD     K       ���  ��  �� �� ��  � ܷ ��  e� [� ��  ޸ ڸ 5��  �jD            ��  ��  � � ��  A� =� ��  ~� z� $�jD            ��  �jD     ��  8C�  s 8P�  v    wjD     ��  Us Tv   <
�  �jD     �      ���  �  �� �� )�  &� � 6�  �� �� �  �jD         ���  6�  ź �� )�  �� ��   C�  E� 5� P�  {� y� ]�  �� �� j�  � � w�  � � 5��   kD     L       ��  ��  >� 8� ��  �� �� ��  �� �� ��  �� �  �jD     ��  U T|    .
�  @ )�  <� 2� �  �� �� @ 6�  �  UkD      p �U�  +�  � � �  W� O� p 8�  �� �� E�  �� �� R�  �� �� _�  y� u� l�  �� �� y�  R� H� ��  �� �� ��  %� � 5��  �kD     �       ��  ��  �� �� .��  � ��  �� �� ��  F� B� ��  �� ��   '��  � ?�  ��  �� �� ��  G� A� .��  0 ��  �� �� .�  ` �  �� ��    �kD     h U�   ;D�  3nD      � �c�  !� � V�  �� �� � p�  �� �� }�  -� %� ��  �� �� ��  � � ��  �� �� ��  �� �� ��  C� 1� ��  � �� ��  J� 8� c��  '��  � ��  ��  �� �� ��  �� �� ��  �� �� .��    ��  Y� S� ��  �� �� .��  P  ��  �� �� .��  �  ��  5� /� ��  �� ~� .��  �  ��  �� �� ��  	� �      ��  �nD        ! ��  ��  .� ,� ��  S� Q�  ! ��  z� v�  �  �� ��   '��  P! ��  ��  �� ��  �  N� H� �  �� �� '�  �! ��  �  �� �� +�  �� �� .8�  �! 9�  8� 4� HF�  xoD     ^       G�  r� n� T�  �� �� .a�  �! b�  �� ��     Hs�  `qD     �       "t�  ��F��  �qD      �qD            OQ�  ��  ��  M� I� $�qD            ��  �� ��  �  �� ��   ~qD     ֹ  U��Q} 8$8&R0X��Y��   2rD     h U@      <�  prD           ���  �  6� ,� &�  �� �� 2�  +� '� ?�  i� a� L�  �� �� W�  i� Y� b�  � � n�  =� 9� z�  y� u� ��  �� �� ��  � �� ��  ?� 9� H��  sD     t       ��  �� �� ��  hsD       " ���  ��  ��  �� ��  " ��  �� ��  �  5� 1�   +sD     h T} v    <�w  �vD     �      �C�  �w  z� p� �w  �w  �w  �w  �� �� �w  �w  W� S� �w  �� �� �w  ,� (� �w  }� w� x  �� �� x  4� *� &x  �� �� 3x  � �� ?x  �� r� Kx   � � Wx  �� �� cx  �� �� ox  X� P� {x  �� �� �x  9� 1� B�x  xxD     B�x  �wD     B�x  yD     ��  /wD       # �j�  ��  �� �� ��  �� ��  # ��   � �  �  x� r�   5y  �wD     F       �  y  �� �� y  y  �� �� �wD     h ��  Ts  xD     � ��  U|  $ &Tv  $ &Q  $ & xD     h U~ ����Ts   5�x  xxD     h       ��  �x  � � �x  �x  X� V� �xD     h a�  Ts  �xD     � ��  U|  $ &T~  $ &Q��� $ & �xD     h U ����Ts   F��  �xD      �xD            �)�  ��  �� �� ��  �� �� $�xD            ��  �� ��  �  � �   5�x   yD     �       ��  �x  P� L� �x  �x  �� �� DyD     h y�  Ts  yD     � ��  U|  $ &T  $ &Q��� $ & �yD     h U���@$����Ts   	wD     h ��  U�B$ 7xD     h 
�  Ts  BxD     h "�  T}  yD     h Uv ����Ts   <Eu  ��D     4      �|�  Vu  �� �� bu  H� F� nu  {� k� zu  0� ,� h�u   �u  u� i� 3 �D     @       ��  �u  �u  � �� �' �u  =� 9�    ( ��  �u  w� s�  .Eu  @( zu  �� �� nu  F� >� bu  �� �� Vu  �� �� @( �u  .� *� �u  '%v  �( L�  *v  h� d� 6v  �� �� Av  �� �� Lv  �  � Wv  )� %� bv  d� `� mv  �� �� xv  �� �� �v  � � "�v  ��H�v  q�D     n       �v  9� 7� "�v  ���v  ��D      *�  U| T��Q: ��D      U| T��Q:   5v  ՋD            s�  v  ^� \�  5�u   �D     @       ��  �u  �� �� "�u  ���D     �v  T��Qv   5�v  ��D            ��  �v  �� ��  '�u  �( +�  �u  �� �� v  	� � ԍD      U| T0Q:  H�v  	�D            �v  A� ?� �v  f� d� �D      U| T0Q:     <y`  0�D     �      �2�  �`  �� �� �`  $� � �`  �� �� �`  7� /� �`  �� �� �`  0� *� �`  � {� �`  �� �� �`  �� �� �`  �  � 	a  W� Q� a  �� ��  a  +� � +a  �� �� 5a  �  � Aa  _� S� ~�`   5Ma  ��D            ��  Ra  �� ��  C��  ώD      �( 	���  ��  /� -� ��  T� R� �( ��  �� w�  �  /� '�   C��   �D      @) 	�.�  ��  �� �� ��  �� �� @) ��   �    ']a  �) I�  ba  �� ��  'pa   * Y�  ua  Y� W� �a  �� |� �a  x� j� �a  /� %� ��  ��D      @* 	X��  ��  �� �� ��  �� �� @* ��  �� ��  �  3� /�   u�D     h ��  T�� ��D     �a  Uu Tt Q'v t  $ &��t  $ &��?&"#��@&Rv X} Y	~ 2$~ "1$  H�a   �D     g       �a  p� n� �a  �� �� ��  �D      �* 	d��  ��  �� �� ��  � � �* ��  7� 3�  �  z� v�   ;��  ?�D      �* 	f��  �� �� ��  �� �� �* ��  � �  �  H� D�     <K�  �D     �      �Q�  ]�  �� �� j�  �� �� w�  p� l� ��  �� �� ��  �� �� ��  'K�  + ��  ]�  g� a� ��  �� �� w�  � � j�  m� c� + ��  �� �� ��  [� I� c��  ��  ��D      p+ 		%�  ��  (� � ��  �� �� p+ ��  � � ��  �� �� ��  �  k  ��  y w ��  � � ��  � � �  � � �  � �  �  � � -�  � � B:�  #�D     'C�   , ��  H�  T N U�  � � b�  	 	 ;��  4�D      `, ?�  �	 �	 �  �	 �	  �  �	 �	  �  �	 �	 �  �	 �	 ��  
 
 `, -�  +
 '
 :�  j
 h
 T�D     �  Q��~�8Z�  ~     'p�  �, g�  u�  �
 �
 ��   �D      - t	^�  �  �
 �
 �  �
 �
  �     �    �  = ; ��  d b - -�  � � :�  � � C�D     �  Q��~�8Z�      ��  x�D      P- �	�  �  � � �  � �  �     �    �  9 7 ��  ` ^ P- -�  � � :�  � � ��D     �  Q��~�8Z�      ٔD     ��  5�  U Ts Q} R0X0 p�D     ��  U Ts Q} R��~X��~�  '��  �- ��  ��  � � ��  B : ��  � � ��  � � ��  h d ��  � �  ��  r�D      �- ;	 �  ��  & $ ��  K I ��  K I ��  p n ��  p n  .��  0. ��  � � ��    F��  ��D      ��D            [��  ��  r p ��  � � ��  � � ��  � � ��  � �  F��  )�D      )�D            Y�  ��  � � ��    ��    ��  + ) ��  + )  W �D     �    ��  #�D      �. 		�  �  X N ��  � � �. �  H @ �  � � (�  v l 5�  G C B�   } .O�  �. P�  � � 5p�  ��D     L        �  q�  � � H~�  ��D     >       �      .]�  / b�  * &     5��  ��D     �       N�  "��  ��~"��  ��~"��  ��~��  ӗD       @/ 	"�  �  b ` �  � � �  � � 3�  � � &�  � � @/ @�  � � M�  4 2 Z�  ] W ;��  �D      p/ p��  ��  � � p/ ��  � �  �  > :     ��D     |�  U��~T��~Q��~R��~  ��D     
�  k�  U T1 ��D     ��  ��  U T��}Q1 �D     �  ��  U��~T|  �D     h�  ��  U��~T|  F�D     ��  8C�  { 8P�  ��}   �D     ��  �  U T��} r�D     
�  /�  U T0 ϓD     ��  U T��}Q0  <w|  ��D     =      �- �|   y �|  � � �|  +  �|   � �|  � � �|  �|  'w|  �/ �
 �|  { s �|  � � �|  e K �|  x l �/ �|    �|  �  �|  � � c�|  �  +�D      �/ �	N �      �  U  Q  �/ )�  �  �  6�  �  �  C�  ! ! P�  \! X! ]�  �! �! .j�  00 k�  �! �! w�  " 	" ��  c" Y" ��  �" �" '��  p0  ��  ?# 7# ��  �# �# ��  �# �# ƃ  �# �# .Ӄ  �0 ԃ  :$ &$ '�  �0 � �  �% �% M��  ��D      ��D            �	��  ��  �% �% $��D            ��  j& f&  �  �& �&    M��  0�D      0�D            �	��  ��  �& �& $0�D            ��  d' `'  �  �' �'     ;��  ��D       1 �	��  ��   1 ��   �       }  i�D       @1 �	 :}  �' �' -}  �( v( @1 G}  �) �) T}  |* v* a}  �* �* n}  �+ �+ {}  �, �, �}  �. t. �}  �0 l0 �}  �1 �1 �}  �1 �1 �}  2 2 '~  �1 � ~  {2 o2 '�~  P2 � �~  3 �2 �~  Q3 K3 �~  �3 �3 �~  �~  4 	4 �~  �4 �4 �~  �4 �4 �~  �5 |5 H�~  {�D     �       �~  :6 66 	  �6 ~6   '$~  �2 Y )~  �6 �6 6~  +7 )7 C~  P~  T7 N7 ]~  �7 �7 j~  �7 �7 w~  @8 :8 �~  �8 �8 M�D     �  U} T��}�Qs Rv   R�D     �  U} T��}�Qv Rs   '�}  �2 � �}  �8 �8 �}  �9 o9 �}  J: @: '�}  03 � �}  �: �: ~  7; /;  ��D     �  U T1Rv   '  p3 h   �; �; +  �; �; 8  6< 0< E  �< < R  �< �< _  9= 1= l  �= �=  .z  �3 {  > > F�  n�D      n�D            )� �  e> c> �  �> �> �  �> �> �  �> �> �  �> �>  .�  4 �  �> �> �  %? !? W��D     �     h�  �D      `4 �	# ��  f? ^? v�  �? �? `4 ��  5@ -@ ��  �@ �@ ��  <A 4A ��  �A �A 5��  �D     9       � ��  �A �A �  %B #B �  LB HB &�  �B �B  Hı  �D     9       ɱ  �B �B ֱ  �B �B �  #C C �  ]C [C    �  ��D       �4 �: -�  �C �C  �  �C �C �  D D �  BD <D �4 :�  �D �D '�  �4  -�  �D �D  �  E  E �  -E +E �  RE PE �4 :�  wE uE �D     ��   U Tv Q��}#hR0 �D     N�  U T0   ��D     ��  U T0   �  �D       5 �O	 -�  �E �E  �  �E �E �  �E �E �  F F 5 :�  PF LF '�  `5 4	 -�  �F �F  �  �F �F �  �F �F �   G �F `5 :�  %G #G �D     ��  	 U Tv Q~��R1 �D     N�  U T1   �D     ��  U T1   5�|  0�D     q       �
 "�|  ��~"}  ��~"}  ��~��  T�D       �5 �	W
 �  JG HG �  pG nG �  pG nG 3�  �G �G &�  �G �G �5 @�  �G �G M�  H H Z�  EH ?H ;��  p�D      �5 p��  ��  �H �H �5 ��  �H �H  �  &I "I     G�D     |�  U��~T Q��~R��~  `�D     �  �
 U Ts  j�D     h�  �
 U Ts  ��D     ��  8C�   8P�  ��~   �D     ��  �
 U T��~ �D     `�  Q��}�R��~X0Y| �  <0f   �D            �k \Bf  U\Of  T\\f  Qif  eI aI  <�e  �D            �� �e  �I �I "f  �lf  �I �I "f  J J *�D      T8Q�l  <�e  0�D            �' �e  EJ AJ �e  �J ~J �e  �J �J O<�D     ) T�T  <
�  @�D     �       �w �  �J �J %�  2�  hK ^K ?�  �K �K "L�  ��Y�  yL oL f�  �L �L "s�  ����  @M 8M �e  ��D       : @ �e   : "f  ��f  �M �M "f  �M �M ��D      T8Q��   '��  @:  ��  �M �M "��  ��Fd  ³D      ³D            M� ed  "N  N Xd  LN FN Kd  "N  N >d  �N �N 1d  �N �N $³D            rd  �N �N d  O O ߳D     � T Q
R��   ��D     �d  Us Tv Q| R��  M�e  �D      �D            d�e  4O 2O �e  $�D            �e  YO WO �D     ) T|     <d  ��D     :       � 1d  �O O >d  �O �O Kd  �O �O Xd  :P 6P ed  yP sP rd  �P �P d  �P �P ��D     � Tv Q
R�R  >)=  )=  gT�K  �K  0vTF\  F\  0�T�,  �,  �>cL  cL  >�-  �-  B>�:  �:  �>5<  5<  ?>;  ;  �>�1  �1  W>7  7  �
>�*  �*  [T�6  �6  0�>jO  jO  TtV  tV  1z>�=  �=  >B2  B2  /i0  _0  3 >-  -  M>uJ  uJ  7>�W  �W  �T�\  �\  2. ��   ][  �  �� $"  ��D     �<      �
 X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �	  	N   �  	B"]  c     	��  R   	�U    �� 	��  �N 	��  �6  	��   �  	Y�  �  U   �  Q  -      	n�  �  �  Q  U    �  	��  �  U     Q  -   -   U    �  	�")  /  �   P	J�  2�  	L,   �  	M@   pos 	N@   �  	P�  SF  	Q�   �1 	R�  (=9 	S9  0R�  	UQ  8y�  	V,  @�� 	W,  H �  	��  �\ 	�-   m  	�U    o  	��  �  	�    @   ,    @   ,  @    2  �  2  	F  L  W       
:-   �  
J�  x 
LW   y 
MW   )  
Oc  	�  B   
s�  M   
uW   }  
uW  V  
vW  /  
vW   t
  
x�  k	  (
e  �  
N    ��  
N   �  
	G   B� 

,  L  
0    
2  s  
2  v	  
U     �  
�  	e  �  (
N�  �  
P)   Z�  
Q)  �  
S�  s  
T�   [  
U�  ?1  
WG     �  )    
Yw  �  =  N   
�7  �   M
  pmoc5  stib	  ltuo|  tolp 	  
��  b  
 "Q  W  �  %  
<�  x 
>)   len 
?0  *� 
@2   %  
B\  	�    
`�  �  �  G   G   �  U    �  �  
q�  �  G     G   G   U    �  
    ,  G   G   U    �  `
��  �  
��   �% 
��  ?1  
�G   �&  
��  !  
��   I  
��  ()  
�  0R   
�U   8�  
��  @ r  �  �  
�,  	�  �   
�  �  G   �  U   �   D  �  
    #  D   �  
?0  6  K  D  ,  @    �  
YX  ^  G   w  D  @   U    s  
��  �  G   �  D  �   �  W  0
�  �  
�7   e� 
��  �� 
�#  �� 
�K  �� 
�w   �� 
�  ( �'  
��  �!  l2  �  �,  �  -  �2  	3  ?  �  ��   	J  �
  �)  	[  �  �0  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   �0  D4   b   �	  xx ��   xy ��  yx ��  yy ��   a  ��  		  z'  �\	  m  �D   ss  �x   �  �1	    �v	  |	  �	  U    �  ��	  �U  �U      �i	   %  ��	  �  $�	  �	  �   
  �� "�	   �@ #�	  �U  $U    �  76
  �; 9�	   ��  :�	   L  <
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=  ��  ?W   �  @W  ~  BW  �  CW  �  DW   5  FW  (B  GW  0�  HW  8 �	  J�  
   sg  �  u[   ��  v[  �  xW  �
  zW  (  {W   �  }  �  �#�  �  k  `�6  R�  �Q   (  �x  |  �x  �  �x  �  ��  �  �D!  v  �6
  �  ��  (�%  �6  07&  �T!  8G   �x  X �  �"C  I  h  �  �M +!   k  t  R�  Q   �  �"�  �  %  8;�  �� =1!   �M >,    ?6
   r$  @a  0 5  �$�  �  %  �`  �� 1!   �M >!  �  7   �  �  (�� 
D  h�� w  p�� c  x K  � m  s  �  �,4  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9x  8  :�  @�  <x  H�  =�  PE-  ?�	  X�!  D�  h:  Fl  �  G[  ��  H[  ��  I[  ��  K[  �  L[  �U  N[  ��  O[  �)�  Q�  ��  R4  ��� S�  �K1 W�  �R�  XQ  �Jy  Y  �%  [6
  ��	  ]�	  �    ^U   ��8  `  � L   A  G    X��  �  �`   E-  ��	  N ��  �8  ��  P �  *%�  �  �  0t�  k  vt   �  w`  �@ x�  ݖ y�  E-  z�	   N |  0�  }�  pR  ~�  x�  �  �ߣ  �7  ��I �e  ��  �x  �h  �x  ��S  ��  �4  ��  �8  ��  �  �U    �  �-   �  �W  o  �W  �L �U    �8  ��  ( �
  L#�  �  W  HE  �  J`   = K
    Ll  d  Ml   �  N   �
  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  E  #   g)$  *  �   ���  =  �	   L  ��   $  �x  0�  ��  8m  �#%!  h�  �   pآ  �7  tG   �x  x J  g  �  �
  �)�  �  �   H�  �  �U    "  ��  �!  ��   ~	  8f�  �
  hl   (  il  �� k�  �� l�    nW  �  oW   �  pW  (�  qW  0 y  s    �$�  �  �  0'�  �N  )x   ?1  *l  }0  +x  i/  ,x  � -	   �  �)       H�k  ��  �a   ?1  ��  (  �  4  �	  \  ��  0  �U   @ +!  �  tag �   �U  �   �  k  �  `  N   
�  w%   }#  �&  h  �  &     
�  E   9
C  � ;
�   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(P  �  �  N   ��  :   �   ^$  1  �!  �!   :  �V  �  ��  �#  ��  �  �  �  6   I$  ��  �  �  6   �&  ��  �  �    6     �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  ��  @ V  R  �  	�  x  =v	  H  E#�  	�  �  @J?  �  L�   �  M7  �� O�  .� P�  �  Q1   �  R�  (�!  S	  08'  TW  8   W!K  Q  -  (l�  k  nt   �M o�  ߣ  p7  �  q�   �  k  )�  �  �  �  ?  �   w   .�  �  �  ?   �  1�  �    ?    �   ,	  K  6    +  ?  +   �  �  :=  C  �  W  ?  ?   �  >�  "  Yo  u  �  �  �  �  �  �   �  _�  �  �  �  �  �    �   $  f�  �  �  �  �  +   �  l�  �  �    �  �  �   #  x�~  �� � �   �  � 7  H  � c  P�  � �  X9!  � �  `l� � �  h  � ~  p     �  �  H2�  �S  4�   �  5�  (  6�  04  7�  88  8�  @ �  :�  �  �=a  R�  ?Q   �  @�  n  A�  �  B�  1$  C  2�  E�  �� F�  `�L HU   � �  Jm  �  P     �  �  �    `  x  x  �   �  &�  �  �  `   �%  *�  �  �  �  4   �%  -�  �    4   {  1    �  $  �   �  40  6  A  �   l  8M  S  �  g  4  C   �  <s  y  �  �  4  �   �  @�  �  �  �  �  4  �  7   �  G�  �  �  �  `  �  �  �   �'  N�  �  �    `     �  S  %  �  H  `  �  �  7  H   �  &  ��,  �� ��   i'  ��  H   ��  P  ��  X�A �s  `Y ��  h�#  ��  p�  ��  x�  �  �  �$  ���  ��  �U�  ��  ��!  ��  ���  �  ��  �A  �&  �g  � �&  �8  N  �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }>  �  U'�  �  m  D   t   �  v�   A  w�  �  x�  &  y�   !  {�  �  �   %   �  >   �  �  >    \	  �  �P   V   f   �  >    �'  �r   x   �  �   �  �    �       �!  �   ��  )    ��  )D   �  )f    }  �   	�   O  ;!  _� =%!   ݰ  >%�   �   �  @�   !  �  �  I  �  6  T!  @    �  d!  @    �  �%  ��  ���"  ֤  �x   Ğ  �x  ��  �3  �  �3  	��  �3  
�  �3  ��  ��"  �  ��"  (��  ��"  <�  ��"  X��  ��  p��  �x  x��  �x  |��  ��"  ��  ��"  �R�  �3  ���  �3  ���  �  �F�  �  �V�  ��"  ���  ��"  ���  ��  �"�  ��  ��  ��  �@�  �#  � [  �"  @    [  �"  @   	 l  �"  @     [  #  @    [  #  @    ��  �q!  �  �#  �  ��  )$>#  D#   H�  p�{#  R�  �Q   ^� ��*  !�  �v*  8 ��  ,�#  �#  �  �#  Q  �#  �#    #  2#  ��  1�#  �#  �#  2#  �  �  �  �   ��  8�#  �#   $  2#   �  ;5$  M� ={#   �� >�#  Յ ?�#   y� A $  ��  AM$   $  �  h!_$  e$  ��  ��  u-v$  �$  ��  8V�$    XS$   j�  Y�$  =9 Zd%  �� [%  Q� \6%   �� ]B%  (�� ^�%  0 	|$  ��  ��$  %  %  S$   ��  �%  !%  6%  S$  �  H   K�  �%  å  �N%  T%  d%  S$  �   ��  
q%  w%  �  �%  S$  �   ?�  1�%  �%  �  �%  S$  �%  2#  �   �  r� `|$  1�  �!�%  �%  $�  ��  �-�%  k&  .�  8�k&    ��%   j�  �p&  =9 �'  �� ��&  +�  ��&   �� ��&  (�� �7'  0 	�%  ǡ  �}&  �&  �&  �%   ��  ��&  �&  �&  �%  �  x  H   ��  ��&  �&  �&  �%  �  �  D   !�  &�&  �&  '  �%  �  D   K�  D'  #'  �  7'  �%  �   	�  kD'  J'  �  h'  �%  �%  2#  �   7� ��%  ��  ��'  ��  ��'   X� ��'  l� ��'   A$  �'  6   �'  j$  �'  6   �'  �%  �'  6   �'  $�  �u'  	�'  �� @4(  org Bx   cur CW  fit DW   �� F�'  
� FL(  �'   G� �J{(  .� L�   �q M{(   4(  �(  @    `� OR(  �� O�(  R(   �� �R�(  3� T�(   !n� U�  �!I� V�  � ^� X�(  �� X�(  �(  �� 0\u)  �� ^x   v _x  n� `x  q� ax  x� cW  u~  dW  �� eW   ʿ fW  ( �� h�(  �� h�)  �(   �� k�)  .� m�   O� n�)   u)  �)  @    Z� p�)  @� p�)  �)   ]� 8tv*  �� v�)   !�� w�)  !�� x�)  !�� y�)  	!��  {�   !��  |x  (!l� }x  ,!��  ~x  0!��   4 � ��)  �� ��*  �)  �(  �*  @    �� ��*  ~� �G    �� �W  N� �W   �� ��*  )� ��*  �*  �� 4 +  	+  N� E>+  pos Gx   len Hx  ?1  I�   "$� N   7]+  � H�  � <>+  p� T�+  ��  V�   � W�    X�*   V� Zi+  R� Z�+  i+  �� ^�+  �� `�   �� a�  Ӏ b�+  �k  c�   3  9� e�+  :� e,  �+  �� iW,  �� k�   r� l�  �� m,   %� o",  �� oo,  ",  B� 0s�,    u�+   �� vW,  >� wW,    � yu,  J� y�,  u,  �� x-  R�  �Q   � ��  �  �D  �� �]+  ^� �-   �,  '-  @    �� ��,  � �?-  �,  �� !Q-  W-  <� 03�-  (� 5x   �b 6x  �� 7W  $� 8W  ?1  9�  S� :E-   Z ;x  ( ��  C.  �� E�   � F�  min GW  max HW   �� J�-  �� J.  �-  ҿ HM�.  � O�   ��  P�    QE-  `T  R�.  o� S�.  � T�   O� U�.  (Xc  V.  0I� Wc,  8"� Xc,  @ E-  .  h� Z .  � Z�.   .  �� ]$�.  �.  2� H��/  �� ��.   �@ ��.  � ��/  ?1  ��  B� ��  �� �    �� �   !�� �E-  (�� �W  00� �W  8�� �W  @ 4� ^$�/  �/  �� ��/  �S ��.   .� ��   G   a�/  �� #�� ^� #�� ~��  �� ���0  2]  ��   [  ��  �  ��.  [  ��/  R�  �Q  �S  ��%   9� �2#  (T� ��0  0�(  �  ��� �x  �� �x  ��� �  ��� �  �{� �  ��� �  ��� �  � �.  �0  @    $� ��/  �� ��0  �/  N   �?3  ��  I� �� �� V� o� �� �� �� }� 	l� 
W� �� � �� {� -� |� �� z� � X�  � !� "^� #f� $z� %�� &�� '~� (�� 0U� 1�� @#� A�� Q�� R� S�� TO� UU� V�� WN� X7� `S� a�� b�� c� p�� �� ��� �þ ��� �e� ��� �1� ��� �,� ��� �T� ��� ��� �� ��� ��� �E� �*� ��� ��� �� ��� �;� �� ��� ��� �q� �1� �k� ��� �پ �0� �|� ��� ��� �� ��� ��� �	� �W� ��� ��� �J� �,� ��� ��� �  �� �3  �� 1!   �� '-  ��   5$  �\� !�%  �p� "h'  � �� $�3  ?3  $d� `�'  	��H     %!  i�  	��H     &�� ��3  '_� �,�3   h'  (�� �`�D     �       �a5  )  ��%  -Q 'Q )^� ��  }Q yQ ).� �x  �Q �Q )�  �H  
R R *�� �a5  ��}+y �W  \R VR ,y
 �x  �R �R +n �x  �R �R -�:   �D       �D            �L5  .�:  OS IS .�:  �S �S .�:  �S �S .�:  �S �S / �D            0�:  1�D     }  2Uw 2T��}�2Q~ 2R��}   1��D     �  2U   W  q5  @    (�� ���D     9       �D6  3  ��%  U4;  ��D      ��D     8       �.8;  T T .+;  8T 6T -MC  ��D      ��D            B6  .[C  ]T [T  4MC  ��D      ��D            C.[C  �T �T    & � u`6  '_� u,`6   �%  (@� f �D     V       ��7  )  fS$  �T �T )^� g�  U �T )�  hH  TU NU *�� j�7  �P-�:  3�D      3�D            pl7  .�:  �U �U .�:  �U �U .�:  �U �U .�:  V V /3�D            0�:  1M�D     }  2Uv 2T| 2Q12Rw    5�D     �  5*�D     �   W  �7  @    (�� `@�D     9       �j8  3  `S$  U4;  @�D      @�D     8       b.8;  7V 5V .+;  ]V [V -MC  N�D      N�D            B78  .[C  �V �V  4MC  c�D      c�D            C.[C  �V �V    69� ;�  �8  '  ;3-  '�k  <�  7� >�  87R�  DQ  9dim E�,    &�� B9  '  '3-  '�� '�  'Ӏ 'D  7� �  :�0  489dim �,  7R�  Q  7�� �  7+; �    & � ��9  '  �$3-  '�k  �$�  '�� �$�  'Ӏ �$D  7� ��  :�0  89dim ��,  7R�  �Q  7�� ��  7+; ��    &�� �:  '  �3-  '�k  ��  7� ��  :�0  �87R�  �Q    &F� y�:  '  y 3-  '^� z �  '�� { H  7� }�  :�0  �89dim ��,  7R�  �Q  7.� �x  9idx ��:    x  �:  @    &�� I;  '  I3-  '^� J�  '.� Kx  '�� L,#  9dim N�,  87� b�  7R�  cQ    &�� <F;  '  < 3-  '�� = ]+   &`� 2o;  '  23-  'R�  3Q   &�� $�;  '  $3-  7R�  &Q   6�� �  �;  ;dim #�,  '�k  #�  'R�  #Q   6�� ��  V<  ;dim �+�,  '6� �+x  '�� �+x  '<� �+x  'R�  �+Q  7� ��  7.� ��  7�� �,  :�u   <�� ��  ��D     �      �Z?  =dim �*�,  �V �V =pos �*x  �W �W =len �*x  SX EX )R�  �*Q  �X �X )�� �*Z?  �Y �Y ,� ��  �Z �Z ,?1  ��  5[ ![ >�u  �p�D     ?�H ,� �,  \ 
\ +idx ��  L\ D\ +max ��  �\ �\ ,�� ��*  t] h] @�H  E�D      0I �>  .�H  ^ 	^ .�H  S^ M^ .�H  �^ �^ ?0I A�H  �^ �^ AI  1_ -_ BI  ��C%I  ��D     1��D     5I  2U}2T��2Q��   @MM  ��D      pI �D?  .vM  k_ g_ .jM  �_ �_ .^M  ` ` ?pI A�M  |` x` A�M  �` �` A�M  	a a D�M  E�M   �D       �D     `       `.�M  Xa Ta .�M  Xa Ta .�M  �a �a .�M  �a �a / �D     `       A�M  �a �a A�M  b b BN  ��12�D     '�  2U��2T<2R	�����2Y��     1d�D     �K  2Ts    x  <�� r�  pE     4      ��B  =dim r/�,  yb eb )�% s/D  dc Vc )D� t/�  d d )�� u/�  �d �d )�k  v/�  ^e Ze )R�  w/Q  �e �e ,� y�  Gf Cf >�u  ��E     @�B  wE       @] }+A  .�B  �f }f .�B  �f �f .�B  �f �f ?@] B�B  ��-C  �E       �E            iA  .C  Bg .g .C  3h h .#C  i i /�E            A0C  9i 5i F=C  �E            A>C  ti pi    1�E     5I  2U 2T~ 2Q��   GH  �E      p] �.QH  �i �i .DH  @j 6j .7H  �j �j .*H  &k k .H  �k �k ?p] A^H  �k �k AkH  Ll Fl DxH  @�H  �E      �] @AB  .�H  �l �l .�H  �l �l .�H  m m ?�] A�H  Um Om AI  �m �m BI  ��C%I  �E     1�E     5I  2U 2T~ 2Q��   H�H  �] �B  A�H  n n A�H  1n +n A�H  ~n |n A�H  �n �n A�H  Ao 7o  1�E     �|  2Uv2Tv2Qs 2R~ I�L  v     6� a�  C  ;dim a*�,  '�k  b*�  'R�  c*Q  7� e,   &n� NMC  ;dim N(�,  '�k  O(�  7.� Q�  87� V,    &`� +iC  '^� +$�,   &�  �C  '^�  $�,  'R�  !$Q   <�� ��  ��D     �      ��F  )>) �+c,  �o �o )R�  �+Q  Np Hp ,��  �x  �p �p ,��  �x  rq jq J� ��   >�u  u�D     @xG   �D      �I  �D  .�G  �q �q .�G  $r  r .�G  ^r Zr ?�I A�G  �r �r A�G  �r �r A�G  s s A�G  us qs A�G  �s �s A�G  �s �s A�G  5t -t   G�F  ��D       J .�F  �t �t .�F  �t �t .�F  �t �t .�F  u u .�F  ^u Zu ? J A�F  �u �u C�F  u�D     K�F  pJ A�F  �u �u AG  v v AG  jv hv A G  �v �v A-G  �v �v H:G  �J ;F  A?G  0w $w ALG  �w �w AYG  Dx >x @sL  ��D      K �F  L�L  L�L  .�L  �x �x ?K A�L  �x �x   1��D     �|  2U��#2T��#2Q���2R��  FgG  $�D     [       AhG  �x �x 1O�D     3�  2Q ����1$ ����"3$      6�� ��  xG  '>) �'c,  '��  �'�  '��  �'�  'R�  �'Q  7� ��  :�u  �M�F  7/� ��   87H� �,  7�� �,  7�� ��  7+; ��  7� �x  MgG  9pos ��  7�1 ��+  7x� ��+   87��  �,     6|� sx  H  '>) s0c,  '��  t0�  '��  u0�  7H� w,  7�� x,  9p1 y�+  9p2 z�+  7�� {�  7+; |�  7.� }�   6�� 6�  �H  '>) 6+c,  '�% 7+D  '%� 8+�  '�� 9+�  'R�  :+Q  7� <�  7� =,  :�u  l87�1 L�+  7�� Mx  7x� N�+  7�� Ox  9val Px    6�� �  /I  '>) &c,  'R�  &Q  'w� &/I  7� �  7.�  �  7� !,  :�u  . ,  N�� ��  ��D     �       ��J  O>) �'c,  by Zy OR�  �'Q  �y �y Ow� �'/I  Hz @z P.� ��  �z �z ,�  �  �z �z ,� ,  M{ G{ >�u  ��D     G�J  �D      �G 	.�J  �{ �{ .�J  �{ �{ .�J  �{ �{ .�J  �{ �{ ?�G A�J  !| | A�J  H| D| B�J  �L15�D     '�  2U�T2TH2R| ����2Y�L    QI� ��  �J  R>) �(c,  R.� �(�  RR�  �(Q  S�<  ��  S�:  ��  S� ��   T�� � �D     �       ��K  O>) �&c,  �| ~| OR�  �&Q  �| �| P.� ��  &} "} P� �,  c} ]} U'M  P�D      PE ��K  .@M  �} �} .4M  �} �} 1`�D     ?�  2Uv   1��D     ?�  2Uv 2Ts   N�� ��  ��D     Q       �sL  O� �,  ~ ~ Vidx ��  �~ �~ OR�  �Q  �~ �~ P� ��  w q Wp ��+  � � X�u  ���D     1��D     �|  2Uv2Tv2Q| 2R�QI�L  v   Y"� ��L  R� �,  Zidx ��  [p ��+   Q� �x  �L  R� �,  Zidx �x   Q�� ��  'M  R� �,  R.� ��  RR�  �Q  S�<  ��  S�:  ��  S� ��   YP� |MM  R� |,  RR�  }Q   Q%� R�  �M  R>) R'�+  RR�  S'Q  R�� T'�M  S� V�  S.� W�  S�� X�*  \�u  l �*  Q=� =�  N  R>) =(�+  R.� >(�  RR�  ?(Q  S�<  A�  S�:  B�  S� C�   Y�� 25N  R>) 2&�+  RR�  3&Q   Nc� Z�%  0�D            �fN  ]~ Z%6  U NO� Rj$   �D            ��N  ]~ R%6  U N�� JA$  �D            ��N  ]~ J*6  U N�� 4�  ��D     �       ��O  O~ 4%�3  � � PR�  6Q  #� !� Wph 7U   H� F� UF;  ��D       E :ZO  .a;  m� k� .T;  �� ��  ^�Q  ��D      ��D     !       <�O  .�Q  �� ��  ^D6  �D      �D     B       >�O  .R6  ߀ ݀  E�3  f�D      f�D     B       A.�3  � �   To� )� E     �       ��Q  O~ )%�3  3� -� _o;  � E      `\ .L};  ?`\ A�;  �� � @iC  � E      �\ )�P  .�C  �� �� LwC  @N  � E      �\ %�P  .(N  ˁ Ɂ LN  1E     ?�  2Uv   `� E     �J  �P  2Us� 2Tv  1� E     �J  2Us� 2Tv   GiC  E      ] *.�C  �� � .wC  � � -N  /E      /E            %�Q  .(N  =� ;� .N  b� `� 1;E     ?�  2Uv   `#E     �J  �Q  2Us�2Tv  1/E     �J  2Us� 2Tv      &�� �Q  '_� 2�Q   5$  (�� �@�D     �      ��U  )9� �'2#  �� �� )�� �'�  Ȃ  )�� �'�   � � )ͩ �'�  �� �� )=�  �'�  ܃ ҃ +dim ��(  W� Q� @�Z  ��D       pB �U  .'[  �� �� .[  �� �� .[  S� K� ?pB A4[  �� �� AA[  �� �� AN[  �� �� a[[  ��D     i       gS  A`[  �� � Gt  ��D       �B � .9t  p� l� ./t  �� �� ?�B ACt  � �� AOt  W� M�    Hn[  �B �T  As[  ݈ Ո @t  ��D      C ��S  .9t  =� ;� ./t  d� `� ?C ACt  �� �� AOt  � ߉   @t  ��D      @C �%T  .9t   � � L/t  ?@C ACt  G� C� AOt  �� ��   @t  ��D      pC �sT  .9t  Ǌ Ŋ L/t  ?pC ACt  � � AOt  1� -�   Gt  ��D      �C �.9t  n� l� L/t  ?�C ACt  �� �� AOt  ؋ ԋ    K�[   D A�[  � � A�[  }� y� A�[  �� �� A�[  � � A�[  � � A�[  Y� U� K�[  PD A�[  �� �� Gt   �D      �D �.9t  f� b� ./t  �� �� ?�D ACt  $� � AOt  �� ��       `}�D     _  �U  2U{ 2T0 1��D     _  2U{ 2T1  <�� ��  ��D     �      ��Y  )R�  �"Q  �  � )��  �"�#  n� h� )p� �"�#  �� �� ,9� �2#  � � *� ��  ��b�D     A      �Y  ,.� ��  w� s� ,�1 ��Y  �� �� c�L �V  +dim ��(  A� ?� ,x� �@(  o� g�  c�L �V  +dim ��(  Ғ В ,x� �@(  �� ��  b#�D     �       �Y  ,�� ��  a� _� ,� �[  �� �� -�Z  (�D       (�D     4       ��W  .�Z  � �� .�Z  =� 9� .�Z  w� u� /(�D     4       A�Z  �� �� F�Z  @�D            A�Z  ۔ Ք    -�Z  a�D       a�D     +       �HX  .�Z  \� Z� .�Z  �� � .�Z  �� �� /a�D     +       A�Z  ͕ ɕ F�Z  p�D            A�Z  
� �    -�Z  ��D       ��D     +       ��X  .�Z  �� �� .�Z  �� �� .�Z  ϖ ͖ /��D     +       A�Z  �� � F�Z  ��D            A�Z  3� -�    -�Z  ��D       ��D     ,       �jY  .�Z  �� �� .�Z  ӗ ї .�Z  �� �� /��D     ,       A�Z  � � F�Z  ��D            A�Z  \� V�    1��D     K�  2U
�  `��D     �[  �Y  2U��2Q��2X  1#�D     �[  2U��2Q~ 2X}   1�D     X�  2U} 2T
p2Q��  [  &4� kZ  '9� k%2#  87R�  oQ    &� $�Z  '�  $'�*  '�� %'x  '.� &'x  'P� ''�*  7>) )�)  7.� *�  7� +W  7Xc  ,�)  7�� -x   6v� [  �Z  ;num )�  '�D )�Z  '�� )[  7.� �  87I� [    g  &?� n�[  '�  n%�*  '�� o%�  '� p%W  7.� r�  9num s�  7>) t�)  Mn[  7A�  �x   M�[  7Xc  ��)   87&� ��)  79� ��)  7�� ��  7+; ��  7W� ��)  7r? ��)  87a�  �W     T�� � �D     �      �;^  O�  �#�*  ݘ ՘ O.� �#�  [� ?� O�  �#�Y  �� �� O�� �#�  �� � O�  �#�Y  p� f� O��  �#x  � � Or? �#x  O� I� P�� ��)  �� �� P�� � �)  ٜ ל P$� ��  � �� P?� � �  (� $� bk�D     J       -]  ,Xc  �)  f� ^� /p�D     @       ,� x  ̝ ȝ   cL s]  ,Xc  )�)  
� � /��D     :       ,� .x  n� l�   c@L �]  +dim ?x  �� �� +top ?x  � � +bot ? x  U� M� ,� ?%x  �� �� ,Xc  @�)  � �  `G�D     ��  ^  2U02Rr 2Xv IH^  �U 1W�D     ��  2U12T} 2Q~ IH^  �U  Y�� �_  R�  �*�*  R�� �*  R)� �*�  R�1 �*�Y  R�� �*�)  R�� �*�)  S$� ��  S?� ��  SN� �  \*_  �8S�m �x  S� �!x  S.� ��  SO� ��)  SXc  ��)  [top �  8S�� �x     Tx� )p�D     �       ��`  O9� )*2#  �� �� On� **�  � � Wdim ,�(  .� (� P3� -�(  �� �� P.� .�  6� 2� P��  /@(  v� n� P�� 0@(  � � P�� 1�  G� E� cB L`  Ww >W  �� |� P��  >W  ӣ ͣ _t  ��D      @B AL9t  ./t  #� !� ?@B ACt  K� G� AOt  �� ��    Et  ��D      ��D     !       6L9t  ./t  ˤ ɤ /��D     !       ACt  � � AOt  6� 2�    d� �  �a  '�� #3-  '�S  #�%  '9� #2#  '&  #�  7w� �0  7)�  �0  7� �  7^� !x  :�u  �87� A�(  7� B�(  7�� D�  7�� E�  7�� G�  7�� H�  7��  J�  7� K�  7�m M    &�� ��b  ')�  �2�0  '^� �2x  9dim ��(  7�� ��  7� ��  7� ��/  7[  ��  :�� 87�S ��.  7N� ��.  7�@ ��.  7oI ��.  7T� ��  87k� �W  76� �W  7� �$W  7�� �+W  7�� �W  7� �W  76� �$W  7@� ��     &� ��c  ')�  �3�0  '^� �3x  9dim ��(  7�� ��  7R�  �Q  7�� ��c  7Z� ��c  7�� ��  7�  ��.  7�� ��.  7oI ��.  Myc  7� �   M�c  7\+  �c   87AT  ?�.  7;  ?�.  9nn @�  89u aW     �.  �.  �c  @    &�� �Sd  ')�  �3�0  '^� �3x  9dim ��(  7�� ��  7.� ��  7oI ��.  87�� �E-  87� �W     &�� l�d  '�  l*�*  ')�  m*�0  7>) o�)  7Xc  p�)  7� q�  7v� r�  7oI s�.  89y xW  M�d  7� �W   87� �W     &�� �e  ')�  ,�0  '^� ,x  7>) #�.  7� $,  7�� %�  7N� &�  7�� 'x  9dim )�(  7�� *�  7A�  +x  M�e  7�@ <�  87.� A�  7oI B�.    M�e  7.� Q�  7oI R�.   87.� ^�  7oI _�.    &�� �9g  '>) �6�.  'oI �6�.  '.� �6�  'A�  �6x  '�� �6x  7`T  ��.  7��  ��  87I� �x  7�� �W  M�f  9nn ��  87�� �E-  9d �W    M�f  9nn ��  87�� �E-  9d �W    89nn ��  7i� ��  7�� � �  M	g  7�� �E-  9d �W   M'g  7�� �E-  9d �W   87�� E-      &�� 	�g  ')�  	)�0  9n �  :*_  y:�� L:�� =M�g  7N� �.  7oI �.  7AT  �.  7;  !�.   87oI T�.  7AT  T�.  7;  T!�.    6�� ��  -i  ')�  � �0  '�S  � �%  '�� � 3-  '9� � 2#  7� ��  7R�  �Q  :�u  M�h  7N� ��  7�@ ��  9n �%�  7�  ��.  7� ��/  87.� ��  7oI ��.    87�  ��.  7oI ��.  9vec ��  9n ��  87�� �x  7�� �x  9dxi �W  9dyi �W  9dxo �W  9dyo � W     &4� [�i  ')�  [%�0  '^� \%x  9n ^�  7oI _�.  9vec `�  7s  a�    &�� 9�i  ')�  9%�0  '^� :%x  9vec <�  7oI =�.  7.� >�   6S� G   (j  ;dx W  ;dy W  9ax !W  9ay !W  7E  "G    &*� Qj  ')�  �0  7R�  Q   &�� �k  ')�  �-�0  9n ��  :*_  87N� ��.  7�S ��.  9end � �.  7AT  �%�.  7;  �-�.  7oT  �W  7n/  �W  7bX  �W  7hX  �%W  7.� �x  7� �x  7�� �x    &� N|k  '>) N/�.  '9� O/2#  '^� P/x  ')�  Q/�0  7�� SE-  7.� T�   (u� �p�D     "      ��o  )�� � E-  �� q� )9� � 2#  ?� /� )^� � x  	� � ))�  � �0  A� 1� +dim ��(  � � ,�� ��  �� � ,� ��  Q� M� ?PM +pos �W  ˬ �� +len �W  P� 0� ,�� �x  �� �� ,y� �W  d� X� ,~� ��*  � � cPN �n  ,S� �E-  Գ γ c�N �m  ,�� �W  � � ,�� �%W  [� S� ,��  W  ˴ ɴ ,u~   %W   � �� @t  F�D      �N em  L9t  ./t  6� 4� ?�N ACt  s� o� AOt  �� ��   1.�D     |k  2U 2T| 2R}   b2�D     @       �m  ,� @W  �� � ,�� AW  =� 9� ,�� BW  �� � ,#� CW  Ķ ��  @=p  ��D       O WJn  .ip  � � .\p  b� N� .Op  ;� 7� Kvp  0O Awp  �� ��   G�o  �D      `O ]!.p  � � .p  >� <� ?`O A"p  i� c� A/p  Ĺ ��    @t  ��D       �M ��n  .9t  � � ./t  �� �� ?�M ACt  �� �� AOt  � ��   -t  ��D       ��D            �ao  .9t  >� <� ./t  t� p� /��D            ACt  �� �� AOt  � �   GZ  1�D        N �	.TZ  4� .� .GZ  �� �� .:Z  � ۼ .-Z  r� l� ? N AaZ  ν Ľ AnZ  T� L� A{Z  ¾ �� A�Z  ɿ �� A�Z  @� 8�     6� ��  =p  ;pos �,�  ;len �,�  7؊  ��  7�k  ��   6�� XW  �p  ;dim X.�(  ;len Y.W  '�� Z.  87� `W    Y�� �Wq  R>) �1�.  RF� �1,  S� �x  [val �x  Sy�  ��+  [idx ��  S�� ��  S.� ��  Mq  7�� E-  87+; �    89i1 5x  9i2 5x  76� 6E-  7�� 6E-  7`T  7�.    Q� ��  r  R>) �(�.  R  �(�+  RI� �(c,  R"� �(c,  RR�  �(Q  S.� ��  S� ��  \�u  �M�q  Sx� �E-  S�1 ��*   M�q  S� �,   8[idx ��    Y;� �er  R>) �/�.  RF� �/,  S� �x  [val �x  Sy�  ��+  [idx ��  S�� ��   T�� `��D     �       �7s  ]>) `*�.  UVidx a*�  �� �� P�� cE-  �� �� ?�A P�x u�.  \� V� P.� v�  �� �� P�� wE-  �� �� _�s  &�D       �A Lt  Lt  .t  � � .t  � �    Y,� Pis  R>) P.�.  S.� R�  S�� SE-   T�� ?��D     m       ��s  O>) ?(�.  D� >� OR�  @(Q  �� �� `��D     ?�  �s  2Uv  `��D     ?�  �s  2Uv  1��D     ?�  2Uv   Qg� 5x  t  R6� 5E-  R�� 6E-   Q�6  �7  \t  Za �7  Zb �7  [ret �"  [tmp �"   e�p  ��D     C      ��u  .�p  �� �� L�p  L�p  A�p  @� 4� A�p  �� �� A�p  <� 4� A�p  �� �� A�p  �� �� A�p  � � ^7s  ��D       ��D     -       �Iu  .Ds  �� �� .Ds  �� �� /��D     -       APs  L� J� A\s  w� o�   a�p  �D     .       �u  A�p  �� �� Fq  +�D            Aq  �� ��   Kq  �E Aq  (�  � A"q  �� �� A.q  �� �� A;q  �� �� AHq  �� ��   e�e   �D     �      ��w  .f  V� N� .f  �� �� ff  Xf*f  YL�e  L�e  A7f  �� �� ADf  � � KQf  �E ARf  M� 9� A_f  S� E� H�f  F w  A�f  �� �� A�f  E� =� A�f  �� �� H�f  PF �v  A�f  � � A�f  M� G�  a'g  m�D     #       �v  A(g  �� ��  K	g  �F Ag  �� �� Ag  � �   Hlf  �F Pw  Aqf  e� c� K}f  �F A~f  �� �� A�f  �� ��   F�f  ��D     X       A�f  � � F�f  �D     ;       A�f  A� =� A�f  }� w�     eWq  ��D     #      ��y  .hq  �� �� .�q  k� _� .�q  �� �� .�q  �� �� Ltq  Ltq  A�q  �� �� B�q  ��C�q  d�D     H�q  G Ix  A�q  �� �� A�q  �� ��  H�q  PG y  A�q  R� L� _r  ��D       �G �	.r  �� �� .r  �� �� .r  �� �� ?�G A(r  � � A4r  �� �� A@r  � �� ALr  W� M� AXr  �� �� 1.�D     er  2Uu 2T|    H�q  �G 8y  A�q  �� �� 1_�D     er  2Uu 2T|  `��D     '�  ly  2U| 2T82Q02R} 2X02Y�� `�D     '�  �y  2U| 2T02Q02Rw 2X02Y�� 1/�D     '�  2U| 2T 2Q02R}����2X02Y��  e�9  P�D     �       ��|  .�9  v� j� .�9  � �� g�9   K�9  0H .�9  �� �� .�9  E� ;� ?0H A�9  �� �� C:  u�D     K:  pH A:  � 	� @�B  ��D      �H �o{  .�B  G� E� .�B  o� k� .�B  �� �� ?�H B�B  �X-C  ��D      ��D            iM{  .C  �� �� .C  +� %� .#C  �� ~� /��D            A0C  �� �� F=C  ��D            A>C  �� ��    1��D     5I  2Us(2T| 2Q�X   4�B  ��D      ��D     '       �L�B  .�B  <� :� .�B  a� _� /��D     '       B�B  �X-C  ��D       ��D            i[|  .C  �� �� .C  �� �� .#C  � � /��D            A0C  4� 0� F=C  ��D            A>C  p� l�    1��D     5I  2Us� 2T| 2Q�X       e�L   �D     t       �}  .�L  �� �� .�L  )� � L�L  L�L  AM  �� �� AM  �� �� BM  �\1Y�D     '�  2U�R2T12Rs ����2Y�\  e�:  ��D     �       ��}  .�:  �� �� .�:  � � .�:  �� �� .�:  �� �� A�:  � � K ;  �I A;  �� �� A;  �� �� 1��D     V<  2U} 2X0   e�Y  @�D     Q       �.~  .Z  �� �� F�Y  H�D     H       .Z  a� [� FZ  H�D     H       AZ  �� �� h��D     ?�  2T�U    ej8  0�D     u       ���  .|8  �� �� .�8  s� i� A�8  �� �� Kj8  @K .�8  � � .|8  �� �� ?@K A�8  '� #� K�8  @K A�8  c� ]� A�8  �� �� @�;  J�D      �K H�  .�;  O� M� .�;  v� r� .�;  �� �� -C  J�D      J�D            �  .C  �� �� .C  �� �� .#C  \� Z� /J�D            A0C  �� � F=C  N�D            A>C  �� ��    1n�D     �C  2Us82T|   G�;  r�D      �K K.�;  � � .�;  T� P� .�;  �� �� -C  u�D       u�D            ��  .C  �� �� .C  E� ?� .#C  �� �� /u�D            A0C  �� �� F=C  y�D            A>C  �� ��    h��D     �C  2U�U#h      e;^  ��D     O      ���  .T^  `� X� .`^  �� �� .l^  � � fx^  Rf�^  XA�^  Q� M� A�^  �� �� A�^  � � C�^  ��D     .H^  U� S� K�^  �K A�^  �� }� A�^  � 	� A�^  Q� C� A�^  �� �� A�^  ;� 7� A�^  {� q� F_  ��D            A_  �� ��    e�`  ��D     �      �Ҕ  .�`  2� � .�`  �� �� .�`  _� [� .�`  �� �� B�`  ��}0a  Aa  � � Aa  �� �� C(a  �D     @�g  ��D      �O 9�  .h  �� ~� .
h  "� � .�g  �� �� .�g  e� W� ?�O B$h  ��|A1h  � � C>h  ��D     HGh  @P �  ALh  �� �� AYh  ;� 5� Afh  �� �� Aqh  �� �� A~h  @� <� K�h  �P A�h  �� v� A�h  �� ��   H�h  �P ��  A�h  _� U� A�h  �� �� A�h  +� !� A�h  �� �� K�h  �P A�h  � � A�h  �� �� A�h  �� �� Ai  � � Ai  �� z� Ai  �� �� @�i  ��D      0Q �"�  .�i  F� B� .�i  �� |� ?0Q Aj  �� �� Aj  :� 6� Aj  t� p�   @�i  %�D      `Q �#z�  .�i  �� �� .�i  /  %  ?`Q Aj  �  �  Aj  ` V Aj  � �   5�D     d�    @�i  ��D      �Q ��  .�i    .�i   s ?�Q A�i    A�i   w A�i  � �   iQj   R �"�  L_j  L_j  ? R Alj  %  Cwj  �D     K�j  0R A�j  � � A�j  � � A�j  � � A�j  } w A�j  � � A�j  ` T A�j  � � A�j  ^ L A�j  '	 	 A�j  �	 �	 Ak  
 
 Ak  f
 ^
 `��D     q�  ��  2U��{2T~ 2Q} 2R  1R�D     q�  2U} 2T��|2Q 2Rs     ` �D     '�  Q�  2Us 2TH2Q02X02Y��| `��D     '�  �  2Us 2T@2Q02X02Y��| `��D     �w  ̆  2U��~2Q��|# 2R��|#(2X��|Itq  ��|#I�q  ��|#8 1��D     �w  2U��~2Q��|#P2R��|#X2X��|Itq  ��|#HI�q  ��|#h   -(j  �D      �D     T       �Շ  .6j  �
 �
 /�D     T       ACj  �
 �
 `,�D     is  ��  2U��~2Ts  `<�D     is  ��  2U��~2Ts  `L�D     ?�  ��  2Us  1h�D     ?�  2Us    K1a  pR A2a    A?a  k e ALa  � � AYa  [ K Afa    Asa   � A�a  � � A�a  � � A�a  � m @t  #�D      �R P��  .9t  a _ ./t  � � ?�R ACt  � � AOt  � �   iSd   S {b�  Lnd  Lnd  Lad  ? S 0{d  A�d  5 1 0�d  A�d  u k A�d  � � K�d  `S A�d    a�d  ��D     |       <�  A�d  6 2  F�d  H�D            A�d  p l     -�i  ��D      ��D     �       m	݉  .�i  � � .�i  | l /��D     �       A�i  E 9 A�i  � � A�i  x t   i9g  �S p	��  LGg  ?�S ATg  � � C_g  ��D     Chg  ��D     Dqg  Hzg   T f�  Ag  n h A�g  � � A�g    A�g  F B  K�g  0T A�g  � | A�g  � � A�g  N D    -k  ��D       ��D     C       s	X�  .-k  � � .-k  � � .Tk  r l .Gk  � � .:k  � � /��D     C       Aak    Ank  y u 1
�D     |k  2UvP2Ts 2Q��|�2R��}   @�d  �D      �T y	u�  .e  � � .�d    ?�T Ae  c ] A!e  � � A.e    A;e  G ; AHe  � � AUe  3 / Abe  � � Aoe  � � H|e  �T ��  A�e  �  F�e  ��D     O       A�e  � � A�e  � � `��D     \t  c�  2U I�p  v  1�D     �u  2Uu 2Tt 2Qs 2R~ 2X��|�2Yy I�e      a�e  ��D     @       ֌  A�e      A�e  C  ?   a�e  �D     K       _�  A�e  }  {  A�e  �  �  `�D     \t  !�  2U  17�D     �u  2Uu 2Tt 2Qs 2R~ 2X��|�2Yy I�e     1N�D     K�  2U    i�c   U |	��  L�c  L�c  ? U 0 d  0d  0d  A'd  �  �  K4d  @U A5d  "! ! KBd  �U ACd  �! �! @t  ��D      �U �+�  L9t  ./t  j" f" ?�U ACt  �" �" AOt  �" �"   -t  p�D      p�D            �,��  L9t  ./t  )# '# /p�D            ACt  P# L# AOt  �# �#   5Q�D     ~�      @�b   �D       V }	Ő  .�b  �# �# .�b  B$ :$ ? V A�b  �$ �$ A�b  ?% 7% Ac  �% �% Ac  & 	& B%c  ��|A2c  �& �& A?c  l' h' ALc  �' �' AYc  ( ( Hyc  pV h�  A~c   ) �(  H�c  �V ]�  A�c  )) #) A�c  �) �) A�c  �) �) H�c   W ď  A�c  �* �* 5M�D     ~�   @t  ��D      @W L�  L9t  ./t  �* �* ?@W ACt  3+ /+ AOt  v+ r+   Gt  ��D      pW \L9t  ./t  �+ �+ ?pW ACt  �+ �+ AOt  7, 3,    afc  ��D     )       ��  Bkc  ��|1��D     '�  2U 2T82Q02X02Yv   1�D     ?�  2U 2Tv    @�a  .�D      �W ~	ޓ  .�a  x, r, .�a  �, �, ?�W A�a  !- - A�a  \- Z- A�a  �- �- A�a  �- �- Ab  5. 3. Cb  ��D     Kb  �W Ab  ^. X. A)b  �. �. A6b  0/ "/ ACb  �/ �/ APb  D0 >0 H]b   X +�  A^b  �0 �0 Akb  1 �0 Axb  �1 �1 A�b  �1 �1 A�b  n2 h2 A�b  �2 �2 A�b  ^3 Z3 A�b  �3 �3 @t  ��D      pX �(Z�  L9t  ./t  4 4 ?pX ACt  D4 @4 AOt  �4 �4   @t  p�D      �X ���  L9t  ./t  �4 �4 ?�X ACt  �4 �4 AOt  .5 *5   -t  1�D      1�D            ��  L9t  ./t  m5 i5 /1�D            ACt  �5 �5 AOt  �5 �5   1��D     K�  2U��|2T~   @t  ��D      �X �"y�  L9t  ./t  �5 �5 ?�X ACt  #6 6 AOt  f6 b6   4t  ��D      ��D            �L9t  ./t  �6 �6 /��D            ACt  �6 �6 AOt  7 
7      --i  ��D      ��D     �       �	f�  .Hi  M7 I7 .;i  �7 �7 /��D     �       AUi  �7 �7 A`i  �7 �7 Ami  8 8 Azi  48 28   `V�D     ~�  ��  2U��|2T| 2Qv  `z�D     �Q  ��  2R02X0 1��D     �Q  2T��|2Q��|2R02X0   e�`  ��D            �C�  .�`  [8 W8 .�`  �8 �8 .�`  �8 �8 .�`  9 9 0�`  0a  0a  0a  j��D     ��   e:  ��D           ���  .-:  U9 K9 .::  �9 �9 .G:  j: ^: gT:   K:   Y .G:  �: �: .::  P; D; .-:  U< M< ? Y AT:  �< �< Ca:  U E     Kj:  `Y Ak:  = = Ax:  �> �> 0�:  B�:  ��@�;  L�D       �Y �D�  L<  .<  �> �> .�;  G? A? .�;  �? �? .�;  �? �? ?�Y A%<  �@ �@ A2<  yA uA B?<  ��CL<  � E     @�L  ��D       �Y ���  .�L  �A �A .�L  �A �A .�L  �A �A K�L  PZ L�L  L�L  .�L  B B   @�L  ��D       �Z �\�  .�L  AB ?B .�L  AB ?B .�L  hB fB K�L  @[ L�L  L�L  .�L  �B �B   @�L  ��D       �[ ���  .�L  �B �B .�L  �B �B .�L  �B �B K�L  \ L�L  L�L  .�L  �B �B   `! E     5I  �  2U	s ��"#82T} 2Q�� `8 E     �K  
�  2Tv 2Q}  `� E     �K  (�  2T~ 2Q}  1� E     �K  2T| 2Q}    5��D     �  5�D     �  1�D     V<  2U~ 2Q| @&2R} 2Xv      e�8  �E     �       �Ǚ  .�8  +C !C .�8  �C �C .�8  D 
D 0�8  K�8   ^ .�8  �D �D .�8  E E .�8  |E rE ? ^ A�8  �E �E C9  (E     K9  @^ A9  5F +F A9  �F �F A&9  �F �F A39  G G `E     `?  ��  2Us2Tv 2Q02R| 2X02Y~  1$E     `?  2Us� 2Tv 2Q| 2R} 2X02Y~      eB9  @E     �       ��  .P9  XG NG .]9  �G �G .j9  TH LH .w9  �H �H 0�9  KB9  �^ .w9  ?I 5I .j9  �I �I .]9  (J J .P9  �J �J ?�^ A�9   K K C�9  �E     K�9  �^ A�9  `K VK A�9  �K �K A�9  	L L A�9  CL ?L `�E     `?  �  2Us2T} 2Q| 2Xv 2Y~  1�E     `?  2Us� 2T} 2Q02R| 2Xv 2Y~      k\  \  Vl�6  �6  �l�Z �Z lF\  F\  �k5<  5<  ?l�K  �K  vk-  -  MkV  V  AkjO  jO   �S   �a  �  !� $"  �E     S*      #F X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �	  	N     :-   �  J�  x LQ   y MQ   )  O]  	�  B   s�  M   uQ   }  uQ  V  vQ  /  vQ   t
  x�  k	  (_  �  N    ��  N   �  	G   B� 
_  L  0    e  s  e  v	  U     e  �  �  �  	l  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     �  )    Y~  	�  �  =  N   �C  �   M
  pmoc5  stib	  ltuo|  tolp 	  �  b   "]  c  �  %  <�  x >)   len ?0  *� @e   %  Bh  	�    `�  �  �  G   G   �  U    �  �  q�  �  G     G   G   U    �    #  8  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  �  0R   �U   8�  ��  @ y  �  �  �8  	�  �   �  �  G     U      P  �    $  /  P   �  ?<  B  W  P  _  @    �  Yd  j  G   �  P  @   U    s  ��  �  G   �  P  �   �  W  0�  �  �C   e� ��  �� �/  �� �W  �� ��   �� �  ( �'  ��  	  
�� &+   �  B"=  C     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  1  -      n�  �  �  1  U    �  ��  �  U   �  1  -   -   U    �  �"	    �   PJ�  2�  L_   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S  0R�  U1  8y�  V_  @�� W_  H �  ��  �\ �-   m  �U    o  ��  �  ��  �  @     �  @   _  @    2      *  �   �!  	le  �  	�B  �  -  	�e  	I  U  �  	��   	`  �
  	�)  �  	�0  �  	�G   
  	�N   �  	�-   \#  	�@   )H  	-   �  	 -   �  	,G   \&  	7U   �0  	D4   b   	�=	  xx 	��   xy 	��  yx 	��  yy 	��   a  	��  	=	  z'  	�z	  m  	�Z   ss  	��   �  	�O	    	��	  �	  �	  U    �  	��	  �U  	�U      	��	   %  	��	  �  	$�	  �	  �  	 )
  �� 	"�	   �@ 	#�	  �U  	$U    �  	7T
  �; 	9�	   ��  	:�	   L  	<)
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @
=#  ��  
?Q   �  
@Q  ~  
BQ  �  
CQ  �  
DQ   5  
FQ  (B  
GQ  0�  
HQ  8 �	  
J�  
   
s�  �  
uq   ��  
vq  �  
xQ  �
  
zQ  (  
{Q   �  
}0  �  
�#�  �  k  `�T  R�  �1   (  ��  |  ��  �  ��  �  ��  �  �h!  v  �T
  �  ��  (�%  �T  07&  �x!  8G   ��  X �  
�"a  g  h  �  �M O!   k  �  R�  1   �  
�"�  �  %  8;�  �� =U!   �M >J    ?T
   r$  @  0 5  
�$    %  �~  �� U!   �M b!  �  C   �  �  (�� 
P  h�� �  p�� |  x K  
� �  �  �  �
,R  �   
.�   �  
/�  O  
1�  C  
2�  �  
4�   d> 
6�  (A  
7�  0T  
9�  8  
:�  @�  
<�  H�  
=�  PE-  
?�	  X�!  
D�  h:  
F}  �  
Gq  ��  
Hq  ��  
Iq  ��  
Kq  �  
Lq  �U  
Nq  ��  
Oq  �)�  
Q�  ��  
RR  ��� 
S	  �K1 
W�  �R�  
X1  �Jy  
Y�  �%  
[T
  ��	  
]�	  �    
^U   ��8  
`5  � L  
 _  e    X
��  �  
�~   E-  
��	  N 
��  �8  
��  P �  
*%�  �  �  0
t	  k  
v�   �  
w~  �@ 
x�  ݖ 
y�  E-  
z�	   N 
|#  0�  
}�  pR  
~�  x�  
�  �ߣ  
�C  ��I 
�l  ��  
��  �h  
��  ��S  
��  �4  
��  �8  
��  �  
�U    �  
�-   �  
�Q  o  
�Q  �L 
�U    �8  
�  ( �
  
L#    W  
Hc  �  
J~   = 
K(    
L}  d  
M}   �  N   
�(  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  
c  #   
g)B  H  �   ���  =  �=	   L  ��   $  ��  0�  ��  8m  �#I!  h�  �6  pآ  �7  tG   ��  x `  �  	  �
  
�)�  �  �   H�%  �  �U    "  ��  �!  ��   ~	  8
f�  �
  
h}   (  
i}  �� 
k�  �� 
l�    
nQ  �  
oQ   �  
pQ  (�  
qQ  0 y  
s%    
�$�  �  �  0'  �N  )�   ?1  *}  }0  +�  i/  ,�  � -=	   �  
�)   &     H��  ��  �   ?1  ��  (  �*  4  �=	  \  ��  0  �U   @ +!  
�  tag 
�   �U  
�   �  
�  �  `  N   

�  w%   }#  �&  h  �  &     

�  E   
9
a  � 
;
�   ��  
<
�  �  
=
�  �  
>
�  �#  
?
�   �  
L
(n    �  N   
��  :   �   ^$  1  �!  �!   :  
�t  �  ��  �#  ��  �  �  �  T   I$  ��  �    T   �&  �    �  )  T  )   �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  �  @ l  R  �/  x  =�	  H  E#�  	�  �  @JX  �  L�   �  MC  �� O�  .� P�  �  QJ   �  R�  (�!  S"  08'  Tp  8   W!d  j  -  (l�  k  n�   �M o�  ߣ  pC  �  q�   �  k  )�  �  �  �  X  �   w   .�  �  �  X   �  1      X    �   J	  K  6.  4  D  X  D   �  �  :V  \  �  p  X  X   �  >�  "  Y�  �  �  �  �  �  �  �   �  _�  �  �  �  �  �    �   $  f�  �    �  �  D   �  l    �  .  �  �  �   #  x��  �� � �   �  � C  H  � |  P�  � �  X9!  � �  `l� �   h  � �  p     �.  	�  �  H2�  �S  4�   �  5�  (  6�  04  7�  88  8�  @ �  :�  �  �=  R�  ?1   �  @�  n  A�  �  B�  1$  C*  2�  E�  �� F�  `�L HU   � �  J�  	  P   �  �  �  �  �  ~  �  �  �   �  &�  �  �  ~   �%  *�  �  �    R   �%  -    !  R   {  1-  3  �  B  �   �  4N  T  _  �   l  8k  q  �  �  R  a   �  <�  �  �  �  R  �   �  @�  �  �  �  �  R  �  7   �  G�  �  �    ~  �  �  �   �'  N    �  1  ~  �   �  S=  C  �  f  ~  �  �  7  f   �  &  ��J  �� ��   i'  ��  H   ��  P  ��  X�A ��  `Y ��  h�#  ��  p�  �  x�  �!  �  �B  ���  ��  �U�  ��  ��!  �  ���  �1  ��  �_  �&  ��  � �&  �V  l  -   �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }b  �  U'�  �  m  D   t+   �  v�   A  w�  �  x�  &  y�   !  {�  �  �C   I   �  b   �  �  b    z	  �  �t   z   �   �  b    �'  ��   �   �  �   �  �  *  �    +   �!  �   ��  )7    ��  )h   �  )�    }  �   	�   O  ;6!  _� =%6!   ݰ  >%�   !  �  @!  <!  �  �  g  �  T  x!  @    �  �!  @    �  �%  N   ��#  :�  )� w� 9� 0� Q� �� �� u� �� 	t� 
�� |� �� �� �� �� z� �� R� �� �  x� !� "�� #�� $� %l� &�� 'K� (:� 00� 1}� @�� Ap� Q� R�� S)� T�� Uj� V�� W%� X�� `� aQ� b>� c@� pb� ��� �s� �6� ��� ��� ��� �R� �[� �[� ��� ��� ��� �� ��� ��� �^� ��� �3� ��� �i� �q� ��� �h� �� ��� ��� ��� �;� ��� �� ��� ��� ��� �� �� �� ��� ��� �<� ��� ��� ��� ��� ��� ��� �� �  Int 5G   
  6N   �  7)  �  80  �� 9-   �� 9"\  _#  :@   d� <e  c� <"_  �!  =�   �� I�$  x K$   y L$   �� NZ$  5� N   X�$  ��  g� �� _�  {� _�$  I� b�$  S� @eQ%  X g�   ʊ hQ%  x  i$  ?1  j�#  �  n$   �S o$  (�� q�#  0�@ tQ%  8 ]� c^%  �$  �� xQ%  3� y~%  Q%  �� ~�%  :� ��#   q�  ��#   O� ��%  [� �"�%  �� ��1(  �� ��#   H� ��#  �� ��#  � ��#  � ��#  �� ��#  �� ��#  �� �$   �� �$  (�� �$  0top �$  8� ��  @_� ��#  Darc ��(  H�� ��#  P�� �@$  XK� �@$  `C� �$  h�� �$  ph� �$  xF� �$  ��� ��#  ��� �M$  �
� �M$  �@� �Q%  �=�  Q%  �V� Q%  ��l  �$  ��  l  ��S  �  ��� 	$   �� 
$  �� �#  �� �(  �� �(   O� �(  (�� �(  0~� 3$  8W� M$  9�� �(  @/� �(  PI� �#  � T� �2>(  �%  �� �Q(  f(  1(  f(  f(   �#  �� �y(  �(  1(  �#  �  �  Q%  Q%   �� ��(  �(  1(   �$  D(  l(  �(  �$  �(  @   ` �%  �(  @    H� $
)  R�  &U     �� ()  �(  �� �*)  0)  ;)  �(   !%  �	��H     
|  �  "N)  �	 �H     #�� _�  �+E     $      �K+  $�� _(�  �L yL $ `(�  YM OM $�� a(�  �M �M $�\  b(�  qN eN %� d�  ��~&�S  eK+  O �N &�I fQ+  ZO PO &R�  g1  �O �O &�B  hQ  P P &M  iQ  �P �P %G  k�  ��~'�u  ��,E     (N,E     'S  �*  )Us )T2)Q��~ (m,E     4S  �*  )U )Q0)X0)Y��~ *�,E     �*  )T��~ (,-E     @S  �*  )U~ )T| )Q}  (K-E     @S  +  )U~ )T| )Q}  (l-E     MS  6+  )U  +�-E     MS  )U   �  l  ,�� Rp+E     /       ��+  $�� R&�  Q Q $ S&�  OQ IQ $C!  T&D  �Q �Q -�+E     YS  )U�T#�)T�Q  .�� 7�  /,  /�� 7+�  / 8+�  /:  9+  /� :+�  0� <�  '�u  K�-E      #a� *�  pE            ��,  $�� *%�  �Q �Q $�� +%�  1R -R $�U  ,%�  nR jR 1�E     )T�T)Q�Q  #��  �  @E     !       ��,  $��  !�  �R �R 2ZE     )T0)Q0  3#� GG   �'E     2      �q.  4�� G-P  S �R 4G  H-�  kS cS 5�S  Jq.  �S �S 5x� K�  0T $T 6Հ  Mw.  ���~6B� O�.  ���~7�(E     k       �-  8vec v�  �T �T 5�� w�  �T �T  9I0  })E      �d �:[0  0U *U ;�d <h0  �U }U =�Q  })E       e �8.  :R  �U �U :R  V �U  (V*E     v0  U.  )Uw )T0 +�*E     v0  )Uw )T1    �  �%  �.  @     $  �.  >@   � 3�� :G   0E            ��.  ?�� :!P  U?�� ;!&$  T?��  <!U   Q @� / E            �6/  ?�� /P  U?j� 0@$  T?��  1&$  Q @�� "�E            ��/  4�� "!
)  =V 7V 5R�  $1  �V �V -�E     MS  )T�U  3�� G   0+E     9       �'0  4R�  !1  �V �V 4� !'0  W W 6� �  �\5�� 
)  lW hW +R+E     eS  )Uv )T8)Q�\  
)  A[� �I0  B�� �!
)   C�O  ��  v0  BՀ  �1(  D� ��   3�� ZG   �E     \      �l:  4Հ  Z1(  �W �W 4� Z&M$  �X �X 8i \�#  $Y Y Ej \�#  X8k \�#  uY mY =�B  #E       ` hf5  :�B  �Y �Y :�B  �Z �Z ; ` <�B  �[ �[ <�B  p\ h\ F�B  �` �4  <�B  �\ �\ <�B  ] ] =�B  �E      0a ��4  :4C  O] E] :'C  �] �] GC  :C  h^ N^ ;�a <AC  ~_ r_ <NC  8` ` <[C  �a �a <hC  [c Uc <uC  �c �c <�C  Wd Kd <�C  �d �d <�C  +f f H�C  pE     I�C  I�C  I�C  J�C  �E            `2  K�C   J�C  �E            2  K�C   J�C  �E     B       �2  <�C  �g �g <D  �g �g JD  �E            �2  KD   +�E     �H  )U~   FiD  @b �3  <jD  �g �g <vD  ^h Zh <�D  �h �h <�D  i i <�D  wi qi <�D  �i �i J�D  OE            `3  K�D   J�D  XE            3  K�D   J�D  �E            �3  K�D   (�E     �D  �3  )U~  +�'E     �D  )U~ )Yv   JD  E            �3  K#D   F1D  pb n4  K6D  <CD  �i �i <ND  fj ^j JYD  �E            ;4  KZD   ([E     %G  S4  )U~  +�E     %G  )U~ )Rs   (�E     �H  �4  )U~ )Tv )Q|  +�E     %G  )U~ )Ts )Rv )X|    +\ E     6Q  )Uu   9\P  � E      �b �
:nP  �j �j ;�b <{P  �k �k <�P  Xl Ll L�P  �b <�P  �l �l <�P  8m *m (� E     �P  M5  )Uu  +� E     �P  )T}      9l:  ~!E       c �:~:  �m �m ; c <�:  \n Fn <�:  Ko Eo <�:  �o �o <�:  Bp p <�:  $r r <�:  Bs >s <�:  |s xs M�:  ��M�:  ��<�:  �s �s <;  �s �s <;  Zt Pt <!;  �t �t <-;  2u .u K9;  <E;  nu hu <Q;  �u �u M];  ��Mj;  ��Mw;  ��H�;  �$E     H�;  &E     H�;  �$E     =|B  ~!E     	 @c l
�6  :�B  �v �v  N|B  �!E      �!E     	       n
�6  :�B  �v �v  =|B  �!E      pc o
%7  :�B  �v �v  =.B  �!E      �c �
�7  :IB  w w :<B  Gw Aw ;�c <VB  �w �w <cB  5x -x <pB  �x �x   =�A  w%E      �c !�7  :B  �x �x :�A  y y ;�c <B  my ay < B  z �y   =�A  F#E      d �
48  :B  �z �z :�A  �z �z ;d <B  U{ G{ < B  | �{   =.B  �#E      Pd �
�8  :IB  �| �| :<B  �| �| ;Pd <VB  8} ,} <cB  �} �} <pB  ~ �}   =.B  �%E      �d �
�8  :IB  ;~ 7~ :<B  w~ q~ ;�d <VB  �~ �~ <cB  a ] <pB  � �   =�A  %E      �d P9  :B  � � :�A  � � ;�d <B  n� b� < B  	� ��   J�;  p&E     0       w9  <�;  �� ��  *�"E     �9  )U~ )T��)Q�� (�#E     wA  �9  )Uu  (�#E     wA  �9  )Uu  *�$E     �9  )U~ )T )Xs )Y}  *�$E     :  )U~  (&E     wA  :  )Uu  (&E     wA  3:  )Uu  *X&E     Y:  )U~ )T )Xs )Y}  2�&E     )U~     Cm� \
M$  �;  BՀ  \
1(  Oy ^
�#  D�� ^
�#  DG|  ^
 �#  OP `
Q%  OQ `
Q%  Di� `
Q%  D�� `
!Q%  D3� b
�#  Dw� b
�#  Otop b
!�#  Du� b
&�#  D�� b
.�#  Ox1 d
$  Ox2 d
$  Oxs d
$  Oe1 d
$  Oe2 d
#$  DI� f
d%  D� g
d%  Df� g
d%  P�� �
	P�� /P�� QD~� �
�#    @� N
E            ��;  ?Հ  N
1(  U @l� �	�E           �=  ?Հ  �	1(  URy �	/�#  �� �� Rx1 �	/�  � � Rx2 �	/�  ǂ �� 4�  �	/Q%  u� e� 4�� �	/Q%  9� )� 8e1 �	$  �� � 8e2 �	$  �� �� 8pxl �	$  �� �� 5�� �	@$  "� � 8f1 �	3$  Ň �� S�u  H
pE     T�E     �      5~� �	�#  6� (�   @'� �	`E     �       � >  ?Հ  �	1(  URy �	/�#  � � Rx1 �	/�  W� S� Rx2 �	/�  �� �� 4�  �	/Q%  �� �� 4�� �	/Q%  ;� 7� ;�_ 8e1 �	$  z� t� 8e2 �	$  � � T�E     :       8f1 �	3$  �� �� 5�� �	@$  �� �� 8p �	@$  � ��    @�� �	PE            �m>  ?Հ  �	1(  UUmin �	+f(  TUmax �	+f(  Q @� |	@E            ��>  ?Հ  |	1(  U @�� ��E     �      ��?  ?Հ  �1(  URy �-�#  4� $� Rx1 �-�  �� � Rx2 �-�  �� �� 4�  �-Q%  P� @� ?�� �-Q%  Y8e1 �$  � � 8e2 �$  �� � 8pxl �$  א ː 8c1 ��#  e� Y� 8f1 ��#  � �� S�u  v	�E     T�E     O      5~� 	�#  d� V�   @&� �PE     !      �	A  4Հ  �1(  J� D� Ry �-�#  �� �� Rx1 �-�  ד ӓ Rx2 �-�  � � 4�  �-Q%  N� J� 4�� �-Q%  �� �� 8e1 �$  Д Ĕ 8e2 �$  �� � 5�  �	A  \� V� 5~� �
�#  �� �� ;�_ 8c1 ��#  9� 5� 8c2 ��#  q� o� 8f1 �3$  �� �� 8f2 �3$  җ Η   3$  @�� � E     B       �wA  ?Հ  �1(  UUmin �)f(  TRmax �)f(  � � 5�  �$  K� E�  @R� EPE     �       ��A  4�$ Eq%  �� �� 8old G~%  �� � 5�� GQ%  X� R� 5�@ GQ%  �� ��  AA� ".B  B�$ "q%  B�,  #Q%  Oold %~%  D�� %Q%   A� |B  B�$ q%  B�,  Q%  Oold ~%  D�� Q%  Ox $   A�� ��B  Vl ��B   d%  C�� �M$  �B  BՀ  �1(  B� � �#  Oi ��#  D�S ��#  QD� �Q%  Oo �M$    C�� �M$  �D  BՀ  �1(  BN� �%�#  Bk� �%�#  B� �%�#  D/_  ��  D�C  ��  Dy>  ��  D�  ��  DoI ��  D�� ��  Ds  ��   Otag ��#  P��  �P�0  �P�S  )P�U  �W�C  D�8  �$   W�C  D�8  �$   WD  Ox $  Oy $  QD�8  $    W1D  D�8  '$   WiD  Dp>  ,�  Ox -$  Oy -$  QD�8  8$    QOx1 Y$  Oy1 Y$  Ox2 Y$  Oy2 Y$  Ox3 Y!$  Oy3 Y%$  W�D  D�8  j$   W�D  D�8  k$   QD�8  t$     3� 5M$  0E           �%G  4Հ  51(  � ۙ Rcx1 5$  �� �� Rcy1 6$  ˚ ǚ Rcx2 7$  � � Rcy2 8$  E� A� Rx 9$  �� ~� Uy :$  � 8y1 <$  Û �� 8y2 <$  ;� 3� 8y3 <$  �� �� 8y4 <$  +� #� 8x4 <$  �� �� 5q� <"$  � � 5�� <)$  `� Z� 5X� <0$  �� �� 5�� <7$  �� �� 5i� =�$  K� G� P�0  �X�_ �F  8o |M$  �� �� (E     6Q  �F  )Uu )Ty  +5E     �Q  )Uu )Tt )Qq   (dE     �J  �F  )Us )T3)Q	�E      Y�E     �O  +-E     �K  )Us )T3)Q	�E       3�� �M$  @
E     �      ��H  4Հ  �1(  ˟ �� Rcx �$  p� l� Rcy �$  �� �� Rx �$  � � Ry �$  '� #� 8y1 �$  h� `� 8y2 �$  � ء 8y3 �$  X� P� 8x3 �$  Т Ȣ 5�� �$  >� 8� 5�� �$$  �� �� 5i� ��$  �� �� P�0  X`_ �H  8o �M$  4� 0� (%E     6Q  }H  )Uu )Ty  +;E     �Q  )Uu )Tt )Qq   (jE     �J  �H  )Us )T2)Q	PE      Y�E     P  +E     �K  )Us )T2)Q	PE       3`� ZM$  `E     +      ��J  4Հ  Z1(  v� j� Rx Z$  � �� Ry [$  '� � N�L  �E      �E     Q       �*J  :SM  � � :FM  g� c� ::M  �� �� :.M  ɧ ǧ :"M  � � :M  � � :	M  S� O� T�E     Q       <`M  �� �� <mM  �� �� +�E     {M  )Us )R| )Xv    (0E     6Q  BJ  )Us  (�E     �Q  fJ  )Uu )Tt )Qq  (�E     {M  �J  )Us )R| )Xv  (�E     6Q  �J  )Us  +AE     �Q  )Uu )Tt )Qq   3#� +M$  �	E     a       ��K  4Հ  +1(  ٨ Ө 4�9  +$�#  )� %� 4�� ,$)  f� b� 4�� -$$  �� �� 4�� .$$  � 	� 8arc 0�(  `� ^� 5E  1M$  �� �� 5�� 1M$  �� �� +
E     �K  )Uv )R�X)X�R  ZW� �M$  �E            ��L  4Հ  �1(  ٪ ͪ 4�9  �"�#  e� a� 4�� �")  �� �� 4�� �"$  >� 2� 4�� �"$  ά Ƭ 8y1 �$  :� 0� 8y2 �$  �� �� 8e �$  p� f� 8e2 �$  � ߮ 8e0 �$  8� .� Of1 ��#  8arc ��(  �� �� D�� ��(  8top �$  �� v� [Fin �E      C�� wM$  {M  BՀ  w1(  Vx1 w$  Vy1 x$  Vx2 y$  Vy2 z$  B�� {$  B�� |$  DE  ~M$  D�� ~M$   34� �M$  �E     �      ��O  4Հ  �1(  �� u� Rx1 �$  C� 3� Ry1 �$  �� � Rx2 �$  ϳ ó Ry2 �$  e� Y� 4�� �$  �� � ?�� �$  � 8Dx �$  �� l� 8Dy �$  �� �� 8e1 ��#  � 	� 8e2 ��#  �� �� 8f1 ��#  � � 8f2 ��#  j� d� 5�  ��#  �� �� 8Ix �$  O� G� 8Rx �$  �� �� 8Ax �$  � � 8top �$  R� N� (fE     qS  &O  )U��)Q  (�E     ~S  FO  )T��)Q  (�E     qS  oO  )U��)T} s )Q  ++E     ~S  )T��)Q   @�� ��E     �       �P  ?2�  ��(  U8a �$  �� �� 8b �$  4� .� 8c �$  �� � 8d �$  � ��  @H� �PE     �       �\P  ?2�  ��(  U8a �$  l� `� 8b �$  �� �  C�� QM$  �P  BՀ  Q1(  On S�#  Op TQ%  QDu� ^�#  Otop ^�#    33� M$  pE     �       �6Q  ?Հ  1(  URy  �#  �� �� 5�� $  �� �� 8n  �#  4�  � ;0_ 8y2 .�#  � 
�   3�� �M$  �E     �       ��Q  ?Հ  �1(  U4� �M$  K� E� 8h �$  �� �� ; _ 5� �Q%  � �   3l� �M$  �E     �       ��Q  ?Հ  �1(  U?w� �"�$  T?� �"M$  Q A�� L&R  BՀ  L1(  Br� L%�#   \�+  �-E     S       �'S  :�+  <� 8� :�+  {� u� :�+  �� �� :,  
� � ],   J�+  .E            
S  :�+  X� V� :�+  �� ~� :,  �� �� :�+  �� �� T.E            <,  �� �� H,  .E     +.E     @S  )Us�   +�-E     �S  )Us�)T�Q  ^ZJ  ZJ  �_�6  �6  �^cL  cL  _F\  F\  �_�,  �,  �_�K  �K  v^jO  jO  
^�=  �=  ^�-  �-  B ]B   3g  �  �� $"  0.E     S      Gl d� �i :G  �G   X  ^� �4   int Z   �i {S @�   g
  �       	N   v  #	N   �  &	N   |
  )	N    h  ,	N   (�  -	N   0�	  2Z   8�  5Z   < 	�   �  
�   �
  8"o     K  	  �  L  �  M  S  �9  M  G   ]  4    -  �  >   Z   �	  	f     :G   �  J�  x L�   y M�   )  O�  
�  B   s  M   u�   }  u�  V  v�  /  v�   t
  x�  �J  f   �]  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  f    ��  f   �  	Z   B� 
�  L  d    �  s  �  v	  m     	�  �  �  ]  
�  �  (N^  �  P]   Z�  Q]  �  S^  s  T�   [  Ud  ?1  WZ     	�  	]    Y�  
j  l<  ��  	�  Z   �  �  m    	�  G  �  �:  '�  	�  Z   �  �  �  m    /\  G�  	�  Z     �  �  �  m    oF  0tv  ��  v|   ��  w�  F� x�  �� y�  �� {Z    � |�  ( V  ~  
v  =  f   ��  �   M
  pmoc5  stib	  ltuo|  tolp 	  ��  b   "�  	�  �  %  <"  x >]   len ?d  *� @�   %  B�  
"    `A  	G  a  Z   Z   a  m    	/  �  qt  	z  Z   �  Z   Z   m    �  �  	�  �  Z   Z   m    �  `�H  �  �H   �% �N  ?1  �Z   �&  �4  !  �4   I  �g  ()  ��  0R   �m   8�  �  @ 	�  	T  �  ��  
U  �   t  	z  Z   �  m   �   	�  �  �  	�  �  �   �  ?�  	�  �  �  �  4    �  Y�  	�  Z     �  4   m    s  �  	  Z   -  �  -   	b  W  0��  �  ��   e� �g  �� ��  �� ��  �� �   �� ��  ( �'  �3  
�  �� 0+�  �  	B"�  	�     	�  R   	�m    �� 	�  �N 	�.  �6  	�P   �  	Y  	  m   .  �  G      	n:  	@  P  �  m    �  	�\  	b  m   �  �  G   G   m    �  	�"�  	�  �   P	J-	  2�  	L�   �  	M4   pos 	N4   �  	PS	  SF  	QS	   �1 	R_	  (=9 	S�	  0R�  	U�  8y�  	V�  @�� 	W�  H �  	�S	  �\ 	�G   m  	�m    o  	�-	  �  	�k	  	q	  4   �	  �  4   �  4    2  	�	  	�	  �	  �   �!  
l�  �  
��	  �  -  
��  
�	  	�	  �  
��   
�	  �
  
�]  �  
�d  �  
�Z   
  
�f   �  
�G   \#  
�4   �  
 G   �  
,Z   \&  
7m   �0  
DN   �H  
Q;   b   
��
  xx 
�<
   xy 
�<
  yx 
�<
  yy 
�<
   a  
�}
  
�
  z'  
��
  m  
��	   ss  
�
   �  
��
    
�  	  (  m    �  
�S  �U  
�m      
�
   %  
�(  �  
$m  	s  �  
 �  �� 
"`   �@ 
#`  �U  
$m    �  
7�  �; 
9`   ��  
:`   L  
<�  f   �'  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=�  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  J'  
   s  �  u�	   ��  v�	  �  x�  �
  z�  (  {�   �  }�  �  �#"  	(  k  `��  R�  ��   (  �
  |  �
  �  �
  �  �
  �  ��"   v  ��   �  �}  ( �%  ��  0 7&  ��"  8 G   �
  X �  �"�  	�  h  #  �M �"   k    R�  �   �  �"0  	6  %  8;}  �� =�"   �M >�     ?�   r$  @  0 5  �$�  	�  %  �  �� �"   �M �"  �  �   �  T  (�� 
�  h��   p�� �  x K  �   	  �  �,�  �   .$
   �  /$
  O  1$
  C  2$
  �  4$
   d> 6J  (A  7J  0T  9
  8  :P  @�  <
  H�  =V  PE-  ?S  X�!  D  h:  F 
  �  G�	  ��  H�	  ��  I�	  ��  K�	  �  L�	  �U  N�	  ��  O�	  �)�  Q/  ��  R�  ��� S�  �K1 W#  �R�  X�  �Jy  Y�  �%  [�  ��	  ]S  �    ^m   ��8  `�  � L   �  	�    X�/  �  �   E-  �S  N �'  �8  �\  P �  *%<  	B  �  0t�  k  v   �  w  �@ x/  ݖ y
  E-  zS   N |�  0�  }<
  pR  ~<
  x�  �  �ߣ  ��  ��I ��  ��  �
  �h  �
  ��S  �j  �4  �
  �8  �4  �   �m     �  �G    �  ��   o  ��   �L �m     �8  ��  ( �
  L#�  	�  W  H�  �  J   = K�    L 
  d  M 
   �  f   ��  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  �  #   g)�  	�  �   ��J  =  ��
   L  ��   $  �
  0�  �B!  8m  �#�"  h�  ��	  pآ  �k  tG   �
  x 	�	  	  	�  �
  �)i  	o  �   H��  �  �m    "  �/  �!  �'   ~	  8f'  �
  h 
   (  i 
  �� k<
  �� l<
    n�  �  o�   �  p�  (�  q�  0 y  s�    �$A  	G  �  0'�  �N  )
   ?1  * 
  }0  +
  i/  ,
  � -�
   �  �)�  	�     H�  ��  �   ?1  �
  (  ��	  4  ��
  \  ��  0  �m   @ +!  7  tag 0
   �U  V
   �    	7  `  f   
�  w%   }#  �&  h  �  &     
J  E   9
�  � ;
�   ��  <
$
  �  =
$
  �  >

  �#  ?

   �  L
(�  	�  �  f   �/  :   �   ^$  1  �!  �!   :  ��  �  �V
  �#  �T  	Z  I
  i  �   I$  �u  	{  �  �   �&  ��  	�  <  �  �  �   	�   �!  H�5  �  �0
   S"  �$
     �5  �"  �<
  �  �<
   ;  �N  (%  �H  0�   �i  8��  ��  @ 	�	  R  ��  x  =  H  E#e  
T  �  @J�  �  L$
   �  M�  �� O5  .� P[  �  Q�   �  Rx  (�!  S�  08'  T�  8   W!�  	�  -  (l/  k  n   �M o/  ߣ  p�  �  q�   	`  k  )A  	G  I
  [  �  /   w   .g  	m  x  �   �  1�  	�  �  �  �  �   	�
  K  6�  	�  �  �  �   	  �  :�  	�  I
  �  �  �   �  >A  "  Y  	  I
  /  }  /  /  �   �  _;  	A  I
  _  }  /  �  �   $  fk  	q  �  }  /  �   �  l�  	�  I
  �  }  0
  V
   #  x�  �� � ;   �  � �  H  � �  P�  � /  X9!  � _  `l� � �  h  �   p 	�    ��  
   �  H2�  �S  4j   �  5^  (  6^  04  7
  88  84  @ �  :1  �  �=  R�  ?�   �  @
  n  A
  �  B
  1$  C�	  2�  E�  �� F�  `�L Hm   � �  J  	�  P      	&  I
  I  �    
  
  D   �  &U  	[  f     �%  *r  	x  I
  �  �   �%  -�  	�  �  �   {  1�  	�  I
  �  /   �  4�  	�  �  /   l  8�  	�  I
    �  �   �  <  	  I
  .  �  0
   �  @:  	@  I
  ^  /  �  
  k   �  Gj  	p  I
  �    
  
  ^   �'  N�  	�  I
  �    �   �  S�  	�  I
  �    
  
  k  �   	<
  &  ���   �� �;   i'  �$
  H   �$
  P  �$
  X�A �  `Y �I  h�#  �f  p�  ��  x�  ��  �  ��  ���  �.  �U�  �^  ��!  ��  ���  ��  ��  ��  �&  �  � �&  ��   	�  �  0tB!  �  vV
   a   wV
  �'  xV
  !  yV
  �#  zV
   �  {V
  ( �  }�   �  U'[!  	a!  m  D   t�!  �  v$
   A  w$
  �  x$
  &  y$
   !  {f!  �  ��!  	�!  I
  �!  O!  
  �!   	�
  �  ��!  	�!  "  O!  �!   �'  �"  	"  I
  7"  O!  
  �	  7"   	�!  �!  v"  ��  )�!   ��  )�!  �  )"   }  ="  
v"  O  ;�"  _� =%�"   ݰ  >%O!   	�"  �  @�"  	�"  	;  �  �  	   �  �"  4    G  #  4    !�  �%�  f   �U%  U�  h� �� j� �� K� �� u� p� �� 	E� 
;� � "� a� 8� q� ~� �� �� �� ��  B� !� "� #�� $�� %L� &�� '� (�� 0�� 1�� @F� A�� Q�� RF� S�� T�� U�� V'� W�� Xe� `�� a�� b�� c
� p^� �A� �N� �,� �� ��� ��� ��� �k� �x� ��� �c� �� � � ��� �Q� �X� �f� �H� ��� �3� ��� � � �� ��� � � ��� ��� ��� �� ��� ��� ��� ��� ��� ��� ��� �� ��� �/� ��� �#� �]� ��� ��� ��� ��� � � �G   z� �Z   
b%  �� �Z   x� ��%  	�%  �� ��%  x �b%   E� �b%  OD �t%  �@ ��%   � ��%  �� �&  �\  ��   �  �Z    �� ��%  8� ��?'  �P  �A   ex �b%  @ey �b%  D�� �b%  H%� �b%  L�� �b%  P,� �b%  TOD �t%  XE� �b%  \MV  �Z   `�� �?'  hz� ��%  pn� �p
  xv� �p
  �x �U%  �y �U%  ��S  �j  ��  �&  ��� �4  ��� �m   � 	�%  ;� �&  �� �_'  	&  O� ��'  R�  �m     �� ��'  	e'  "�R  ��  	��H     #�  �	��H     �  ,  !    ,  *  ",  $�'  	 �H     $�'  �	��H     $�'  �	 �H     %� uI
  0BE            ��(  &�� u-}  � � & v-/  W� S� &�� w-/  �� �� &�\  x-�  �� �� ';BE     *  (U�U(T�T(Q�Q(R�R(X4  %7� iI
   BE            �g)  &�� i+}  � 
� & j+/  K� G� &�� k+/  �� �� &�\  l+�  �� �� '+BE     *  (U�U(T�T(Q�Q(R�R(X3  %� ZI
   BE            �*  &�� Z'}  � �� & ['/  ?� ;� &�� \'/  ~� x� &�\  ]'�  �� �� 'BE     *  (U�U(T�T(Q�Q0�Q $@L$.( (R�R(X0  )�� ^I
   <E     �      �V.  *�� ^/}  +� � * _//  � � *�� `//  B� $� *�\  a/�  �� �� *�� b//  �� �� +� dI
  ��~,�S  eV.  x� `� ,�I f\.  �� �� ,R�  g�  �� �� ,�B  h�  U� 7� ,M  i�  �� �� ,3� j
  � �� ,�� k
  � �� +G  mU  ��~-�u  E�=E     .0f �,  ,+ �b.  � � ,/� �b.  5� )� /i �
  �� �� /j �
  &� "� ,�  �f   g� ]� ,��  �f   �� �� ,�  �Z   �� �� 0�>E     ,  (T��~ 1�>E     �A  *,  (U} (T	�(Q0 0?E     ?,  (T��~ 1@E     �A  b,  (U} (T*(Q0 0G@E     w,  (T��~ 1t@E     �A  �,  (Uw (T��~(Q��~ 1FAE     �A  �,  (T~ (Q��~ 2wAE     �A  (Uw (T~   .pf z-  3�  Z   �� �� 0�?E     -  (T��~ 1�?E     �A  0-  (U} (T0(QE 0�?E     E-  (T��~ 1�AE     �A  h-  (U} (T0(Q	� 4�AE     (T��~  1�<E     �A  �-  (Uw  1�<E     �A  �-  (U} (Tv (Q|  1�<E     �A  �-  (Us (T~ (Q  1=E      B  .  (Uw (Q0(X0(Y��~ 0�=E     .  (T��~ 1->E     �A  5.  (Uw  2�>E     �A  (U} (Tv (Q|   	j  	�  	�	  5�� Q�/E     /       ��.  *�� Q%}  /� +� * R%/  n� h� *C!  S%�  �� �� '�/E     B  (U�T#�(T�Q  6�� 6I
  @/  7�� 6*}  7 7*/  7:  8*�  7� 9*�  8� ;I
  9�u  J_HE      )E� *I
  �.E            ��/  *�� *$}   � �� *�� +$0
  P� L� *�U  ,$V
  �� �� :�.E     (T�T(Q�Q  )��  I
  P.E     !       �0  *��   }  �� �� 4j.E     (T0(Q0  %�� �Z   @.E            �S0  ;�� �(�  U;�� �(4   T;��  �(m   Q <�� �0.E            ��0  ;�� �&�  U;j� �&�  T;��  �&4   Q <�� ��.E            ��0  &�� � �  � � 3R�  ��  n� j� '�.E     �A  (T�U  %`� �Z   �;E     9       ��1  &R�  � �  �� �� &� � �  �� �� "� �I
  �\3�� ��'  M� I� 2�;E     �A  (Uv (T8(Q�\  %�� !Z   �3E     �      �m2  &�� !0�  �� �� &G  "0-   � �� 3�S  $m2  �� �� 3x� %H  �� |� "C!  &  ��}3�� &  �� �� "Հ  )s2  ��~1P4E     B  W2  (Tw  25E     �2  (U��~  	w  E'  �2  4     %%� �Z    1E     {      ��4  &Հ  �R'  � � 3}  �o%  b� ^� =/  �o%  3M   �o%  �� �� 3V  �o%  �� �� "B� ��4  ���~3�  �N   /� -� >n �N   \� R� >y �b%  � 
� "�� ��4  ���~3�� ��4  g� _� ?�e 3��  �b%  �� �� 3� �Z   d� ^� @�5  |2E      |2E     �       �4  A�5  �� �� B|2E     �       C�5  �� �� D�5  �e C�5  �� �� C�5  7� 1� C�5  �� �� C�5  �� �� 1�2E     �5  ]4  (U (Q| (R~  13E     �5  �4  (U (Q| (R~  2;3E     �5  (U (Q| (X1    1U2E     B  �4  (T0(Qw  2x2E     �4  (U    �%  �4  E4   � b%  �4  4    	b%  %�� �Z   �0E     h       ��5  &Հ  �R'  ,� (� "� �a   �l1�0E     #B  _5  (U�X 1�0E     /B  �5  (Us�(T	��H     (Qs  2�0E     �=  (U�X  F�� �5  GՀ  R'  Hy 
Z   I=�� �%  Hx b%  =E� t%  =OD t%    < � ��.E           �
7  &Հ  �R'  k� c� Jx � b%  �� �� Jy � b%  C� 7� &*� � t%  �� �� &A�  � b%  �� �� K�.E     &       �6  "�� �"  �j4/E     (U�Q(T1(Q�j  ?Pe >q ��  � �� >c ��  �� �� 2�/E     ;B  (Q	�X $ &   %�� �Z   �EE     *       ��7  &*�  �$�  9� 5� &3�  �$�  v� r� Jto �$�  �� �� &Հ  �$R'  �� �� 2�EE     P>  (U�RLN9  �UL[9  �TLh9  �Q  %A� �Z    HE     $       �:8  &�i  �$�  B� >� Jto �$�  � {� &Հ  �$R'  �� �� 2HE     �?  (U�QL�:  �UL�:  �T  %�� �Z   @;E     )       ��8  Jto �#�  � 
� &Հ  �#R'  M� G� 2b;E     <;  (U�T  %�� �Z   p;E     G       �39  Jto �#�  �� �� &Հ  �#R'  �� �� >x �U%  C� =� >y �U%  �� �� 2�;E     P=  (U| (Tv 8&(Qs 8&  F�� C!:  GՀ  CR'  G*�  C1�  G3�  D1�  Mto E1�  =�� G!:  Harc H^  Hdx IU%  Hdy IU%  Hdx_ IU%  Hdy_ IU%  Hdx1 JU%  Hdy1 JU%  Hdx2 JU%  Hdy2 J U%  HL KU%  Hs KU%  =�a KU%  N�� � �  1:  4   0 F�� 'y:  G2�  '!^  Ha )U%  Hb )U%  Hc )U%  Hd )U%   FX� ��:  GՀ  �R'  G�i  �1�  Mto �1�  =�� ��:  Harc �^  Hdx �U%  Hdy �U%  =�� �Z   =/, �Z    �  
;  4     F0� �<;  G2�  �!^  Ha �U%  Hb �U%   <� M�6E     �      �P=  &Հ  MR'  �� �� &� M$U%  �� �� &� N$U%  � 
� >dx PU%  T� F� >dy PU%  � �� >fx1 PU%  �� �� >fy1 PU%  &� �� >fx2 PU%  �� �� >fy2 P$U%  s� c� >ex1 Qb%  J� *� >ex2 Qb%  �� �� >ey1 Qb%  _� ;� >ey2 Qb%  �� �� OEnd �9E     . f �<  3�� �U%  �� �� 3�� �G   O� K� 3�� �G   �� �� 2Q8E     P=  (Us (T| (Q}   1�9E     P=  =  (U} (T| (Qv  1�:E     P=  /=  (U} (T���(Q|  2;E     P=  (U} (T (Qs   <� 96E            ��=  &Հ  9R'  �� �� Jex 9#b%  c� [� Jey :#b%  �� �� P�6E     �=   <��  0E     �       �P>  &Հ  R'  ,� (� 3�� ?'  m� e� 3�� �%  �� �� >x b%   � � -�Y -p0E     2�0E     GB  (T1  Q39  @BE     p      ��?  AA9  s� k� Rh9  Rh9  R[9  R[9  RN9  RN9  St9  ��yC�9  �� �� C�9  �� �� C�9  �� �� C�9  i� ]� C�9  3� '� C�9  �� �� T�9  C�9  K� E� C�9  �� �� C�9  �� �� C�9  � �� C
:  �� �� U:  PDE     V1:  PDE      �f ��?  A?:  �� �� ?�f CL:  A  1  CW:  �  �  Cb:  l f Cm:  � �   2DE     <;  (U��y(T| (Qv   Qy:  �EE           ��@  A�:   
 R�:  R�:  R�:  R�:  S�:  ��{C�:  � � C�:  ^ X C�:  � � C�:  � � C�:  � � V
;  GE      �f 	�@  A;    ?�f C%;  < 6 C0;  � �   1�GE     <;  �@  (Uv  2�GE     <;  (Uv   Q�.  0HE     S       ��A  A�.  � � A�.  / ) A/   { A/  � � W#/   X�.  gHE            �A  A�.   
 A/  4 2 A/  \ Z A�.  �  BgHE            C#/  � � U//  {HE     2{HE     �A  (Us�   2_HE     SB  (Us�(T�Q  YcL  cL  Z�K  �K  v[�D  �D   ZF\  F\  �YZJ  ZJ  �Z�6  �6  �Z�,  �,  �[i0  _0   Z�X �X 'ZN  N  {Zi0  i0  0Z+A  +A  #Y�-  �-  B <;   ]l  �  �� $"  �HE     �0      �� X  ^� 	�@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  �	  
	N   �  B"P  V     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  D  -      n�  �  �  D  U    �  ��  �  U     D  -   -   U    �  �"  "  �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S,  0R�  UD  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��    @       @     @    %  �  2  9  ?  J       :-   B   s�  M   uJ   }  uJ  V  vJ  /  vJ   t
  xV  k	  (#  �  N    ��  N   �  	G   B� 
  L  0    %  s  %  v	  U     �  �  	#  =  N   �s  �   M
  pmoc5  stib	  ltuo|  tolp 	  �5  b   "�  �  �  %  <�  x >)   len ?0  *� @%   %  B�  	�    `�  �    G   G     U    �  �  q!  '  G   @  G   G   U    �  M  S  h  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  �  ()  �@  0R   �U   8�  ��  @ 0    �  �h  	  �   !  '  G   ;  U   ;   �  �  N  T  _  �   �  ?l  r  �  �    @    �  Y�  �  G   �  �  @   U    s  ��  �  G   �  �  �     W  0�C  �  �s   e� �  �� �_  �� ��  �� ��   �� �A  ( �'  ��  �  -  �%  	W  c  �  �0  
  �N   �  �-   \#  �@   �  ,G   \&  7U   �0  D4   N   �
  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �   �  �%C  N   �^  ��  � Z P  &  ?� s� s� y� 	� 
2 C� �� e | �  � j� � " �  k !� "�  #�� $�� %� &�� '� (�� 0� 1�� @D  A Q�� R_ S� T0� U� V�� W� X  `>� a]  b�� cW p�� �� �+� �&� �w ��� ��� �Z� �M� �) � �]� �� �� ��� �� �< �� �+ �\� �E� �� �p ��� � � ��  �n� ��� �]� �� ��� �� ��� �7� �'� �m �� ��� �6� �� �� �o� ��� �� �� �� ��� � d� �%  � �N   	j  =� �@   �� �^  	�  �  �j  	�  X� �{  � �U   
�  ��  �   
{  ��   
�  �G   
�  �G   
   �G   �� ?    �  .  �  j  j   �� @:  @  P  �  �   �� pD   E   � Fj  �� G{  �� I  �� Jj   �� K{  (msg M�   0�l  N i  8� P  @� Q.  H�  R�  P� TG   X{� U{  `ݖ V{  h �  J (i  �� !�   sub +,  >� .G   � /j   1Z      �� WP  _� Y�  o  
�� 	G   
�� �   
! �   �� ��  �  {  �  {  �  j   �  (� #�  	�  p�   �  ?   2�  j   ?  K ^   �� ^   a  �   pad 
j   �� )m  �� p  �� �   sub /U  k� 0j  (�� 3j  ,i� 4	{  0� 52  8�� 6
  @end 7
  H�1 8
  Px� 9
  X�� :�  `��  ;	{  h � (#  �� 0�  �� !�   len $j  sub /@  �� 2^  �� 3^  � 42   5� 52  ( N   �  �D   ` ^ �� �� �� �� DRY � BAD 	 �� �   $,  >) %j   �N  &j  e ',  bb (j  tb )2   �  �  +O   � -O       "�  �  #
j  �� *�  8� .8    v  �  !@    	�  "R +�  	�I     "� /�  	 I      v  �  !@    	�  "� 2�  	�I     "�� 6�  	 I     #-� 
v  	#� v   �  0  $@   � 	  "3 0  	 �H      �  [  !@    	K  "* �[  	 �H      v  �  !@    	v  "�� �  	��H     N   �  >  LEN � Y R� �� LIT �� END Y� 	  �  &  G� '2   � (j   +@  get ,j   ��  -j   %n  � )�  lit *
j  �  .    v  ~  !@    	n  "Y ~  	@�H     N   �  ?  c  �� �� �� �� � �� d� ]� 	V� 
�� � N  � �  &,  was '{   � ({   $Z  �� %
j  ��  )  �� *
j   a  %�� � ��  �% �   Jy  �  R�  �D  �� �o  �S ��  �� ��  �&B� ��  �'pos ��  � &y�  �  � &�� �  �   W    $@   � W  �� �  `  (IE ��  `xE     �       �7  )R�  �'D  � � )U� �'  T J )W �'7  � � )� �'h  �	 �	 )� �'�  (
  
 *Jy  �o  ��~+err �G   �
 �
 ,�xE     7  �  -Uw -T? ,�xE     0#  
  -Uw -T4 ,�xE     >-  "  -Uw  .8yE     >-  -Uw   �  (�% o�  PuE           ��  )Jy  o"  a W )�% p"  � � /� r�  . * /R�  sD  j f +zip t  � � 0�u  ��vE     1�n �  /> ��  { q 1`o /  /� �  � � 1po   /.� ��  � | 2-  �wE      �o ��  3;  � � 4�o 5H    .�wE     >-  -U|   ,xwE     �  �  -U| -T0-Qv -R  ,�wE     �  �  -U| -T0-Q0-R0 ,�wE     �:  �  -U} -Tv  .xE     �:  -U} -T|   .#wE     �:  -U} -T -Q��  6�  ~vE       o �3  d X 4 o 7  ��5  � � 5,  � t ,�vE     �:  �  -Uv  ,�vE     �:  �  -Uv -T�� ,wE     �:  �  -Uv -T~  8UwE     �:     2V  �uE      �n ��  3�    3u  \ T 3h  � � 4�n 5�  (  5�  � � 9�  8wE     ,vE     �  f  -Uv  ,vE     �:  ~  -Uv  .^vE     7  -U|-T	�   ,�uE     �  �  -Uv  ,�uE     �:  �  -U} -T
� -Q�� .GwE     �:  -U} -T|   :�� W�  :  ;Jy  W-  <� Y�  <# Z�  <E  [�   =� J@   @uE     	       ��  )Jy  J&  4 0 )x  K&@   q m )B� L&  � � ).� M&@   � � +zip O  ( $ >IuE     �  -T�T-Q�Q-R�R  ?�  4 RE     �       ��  )Jy  4$  i _ +zip 6  � � /R�  7D    2-  RE       g =�  3;  U S 4 g 5H  ~ x .RE     >-  -Us   ,uRE     �:  �  -U| -Ts  .�RE     �:  -U|   : ��  L  @zip �!  @pos �!�  ;B� �!  ;.� �!�  <E  ��  <� ��  0�u  &�sE     A<� �    :�� ��  �  @zip �*  ;.� �*�  <� ��  <� ��   =C� ��  �qE     �      ��  Bzip �*  � � /�� ��  � � /� ��  J @ 4�l +err �G   � � 2�  drE      pm ��  3�   � 4pm 5�  } s 5�    � 5�   o C%rE     -Uv -Q| -R
    .ErE     0#  -U} -T0   :G |�  �  @zip |)  <�� ~�  <Jy    <�  ��   :�� `�  -  @zip `$  <Jy  b  <� c�  A<�� h�    D;� IV  @zip I#  <�� K�   :v  �  �  @zip #  ;Jy  #  ;�% #  <��  �  <� !�  E�u  C F ��  SE     .      �u   GJy  �$  P H H� ��  � � "�; �u   �\0�u  dSE     I�SE     =       y  Jlen �z  � � ,�SE     �:  d  -Us -Tv  .TE     ;  -Us   I�SE            �  Jc �z   � .�SE     ;  -Us -Tv   I�SE     "       �  +c z  G C .�SE     ;  -Us -Tv   , SE     �:     -Us -T0 ,BSE     ;  >   -Us -T�\-Q4 ,xSE     ;  [   -Us -T6 .9TE     ;  -Us -T2   W  �   !@    K�� ��RE            �%!  G�  ��  � � Lptr ��  � � M"  �RE      �RE            �35"    3)"  B > >�RE     �:  -U�U-T�T   Fk� ��  �RE            �"  G�  ��   { G��  �N   � � G�  �N   � � NB"  �RE      Pg �3k"  6 2 3_"  s o 3S"  � � 4Pg 5w"  � � 7�"  �l5�"  ` \ .SE     �:  -U�U-T�Q�����T����-Q�l    O> �B"  PR�  �D  P ��   Q� ��  �"  PR�  �D  P��  �j  P�  �j  Rsz ��  S� ��  Rp ��   FF {  �OE     2      �0#  G{� {  � � Lbuf �  � � Llen 
j  �  y  Js1 @   H!  ! Js2 @   �" �" Jk 	G   p$ h$  T�� �G   pWE     b      � -  Lz �{  % �$ Lf �G   t' l' Jr �G   �' �' Jb �j  �) �) U[.  "[E       �g ��,  3�.  �* 4* 3v.  	0 �/ 3l.  1 1 4�g 5�.  �1 U1 5�.  +4 �3 5�.  �6 e6 5�.  �; e; 5�.  �> �> 5�.  �@ S@ 5�.  �B �B 2�0  �aE      �h TT&  3�0  D �C 3�0  �G �G 3�0  �G �G 4�h 5�0  H H 5�0  UI EI 5�0  J �I 5�0  �K sK 5�0  cM 'M 5�0  �O �O 5�0  R �Q 51  �S yS 51  �V �V 51  X �W 5#1  Y �X ,�[E     �1  5%  -U| -Ts -Q	� ,dE     �1  W%  -U��~-T��~ ,fE     �1  y%  -U��~-T��~ ,�fE     �1  �%  -U| -Ts -Q1 ,�fE     �1  �%  -U| -Ts  ,�jE     �1  �%  -U| -Ts  ,[lE     �1  �%  -U| -Ts -Q	� ,nE     �1  &  -U| -Ts  ,�nE     �1  8&  -U| -Ts  .xqE     �1  -U| -Ts    Vn0  �[E      �[E            W�&  3�0  �[ }[ 3�0  �[ }[ 3{0  �[ �[  W/  �i �&  5/  �[ �[ 5/  �\ �\ 5/  o] k] 5(/  �] �]  Uh3  _E       @j ��'  3�3  E^ ?^ 3�3  �^ �^ 3�3  _ �^ 3�3  �_ �_ 3z3  n` f` 4@j 5�3  �` �` 7�3  ��5�3  la da X_E     �'  -TC-Q4 ,p_E     �3  �'  -U��~-TC-QC-R0-X0 X�_E     �'  -T��~ X�mE     �'  -T��~ C�nE     -T��~   W4/  �j q*  75/  ��7A/  ��7M/  ��7Y/  ��5e/  �a �a 2�2  �iE      k ;�)  343  b 	b 3(3  `b Xb 33  �b �b 33  Sc Ic 33  �c �c 3�2  ]d Sd 3�2  �d �d 3�2  3e -e 3�2  �e �e 4k 5?3  �e �e 7J3  ��5V3  �f �f ,o`E     �3  =)  -U��~�����2$��"-T���#-Q0-R	�I     -X	 I     -Y�� X�`E     S)  -T��~ X�iE     m)  -T
 -Q4 ,�iE     �3  �)  -U��-T��~�-Q
-R	�I     -X	 I     -Y�� X<jE     �)  -T��~ C�pE     -T��~   6.1  �`E       �k I3k1  Og Mg 3k1  Og Mg 3`1  tg rg 3U1  �g �g 3J1  �g �g 3?1  h h 4�k 5u1  Oh Mh C�`E     -T1-Q0    W�.  0l �+  5�.  vh rh 5�.  �h �h 5�.  �h �h 5�.  :i 6i U.1  �lE      �l �#C+  3k1  �i �i 3k1  �i �i 3`1  �i �i 3U1  j j 3J1  Xj Tj 3?1  �j �j 4�l 5u1  �j �j C�lE     -T1-Q0   Yi2  �lE      �lE             ��+  3�2  
k k 3�2  Bk @k 3�2  lk jk 3�2  �k �k 3{2  �k �k  .�oE     �1  -Ts -Q	�  ,;]E     �1  �+  -Ts -Q	� ,`E     �1  ,  -Ts -Q1 XIbE     *,  -T O 
�?5%O"#�-Q4 ,�bE     �1  H,  -U| -Ts  ,$cE     *;  h,  -Tv -Q��~ ,ucE     �1  �,  -Uw -Ts  ,�hE     �1  �,  -Ts  ,�hE     �1  �,  -Ts -Q	� ,�jE     �1  �,  -Ts  .)oE     �1  -Ts    .�gE     �/  -Ts   Q�� RG   >-  Zz S{  Zw TG   P��  U
  P� VG    T�� DG   @OE     ~       ��-  Lz E{  �k �k M2.  iOE      iOE     5       J3O.  Sl Ol 3D.  �l �l ,vOE     �/  �-  -Uv -Ts -Q0 C�OE     -Tv    F�� 6G   �NE     R       �2.  Lz 7{  �l �l .%OE     �/  -T�U-Q0  :�� wG   [.  @s xZ  @z y{   Q� wG   r/  Zs xZ  Zz y{  Zr zG   Rt |j  Rb }	{  Rk ~j  Rp 
  Rn �j  Rq �
  Rm �j  [/  Rbl �j  Rbd �j  Rtl �2  Rtd � 2   [4/  \h 2  \i j  \j j  \c j   A\bl 4j  \bd 4j  \tl 52  \td 52  \c 6O    Q� XZ  �/  Zz Y{  Zc Z�  Zw [j  Rs ]Z   ]#� C`NE     �       �h0  Ls DZ  m m Lz E{  mm gm Lc F	h0  �m �m Yn0  �NE      �NE            MN0  3�0  �m �m 3�0  �m �m 3{0  n n  C�NE     -U0-T0-Q0  �  Ox� ��0  Zc �O  Zz �{   Q�� PG   .1  Zs QZ  Zz R{  Zr SG   Rj Uj  Rt V2  Re Wj  Rb X	{  Rk Yj  Rp Z
  Rn [j  Rq \
  Rm ]j  Rf ^
  Rc _O   Qa� :O  �1  Zbl ;j  Zbd ;j  Ztl <2  Ztd =2  Zz >{  Rc @O   Fa� G   @TE     A      �i2  Ls Z  In An Lz {  �n �n Lr G   .o $o Jn j  �o �o Jp 
  p p Jq 
  vp fp X�TE     (2  -T -Q~  ,�TE     *;  F2  -T -Q~  X@UE     [2  -Tw  8bUE     *;   :�� �G   �2  @bl �,  @bd �,  @tl ��2  @td ��2  @z �{   �2  �  : GG   b3  @nl Hj  @nd Ij  @c J,  @bl K,  @bd L,  @tl Mb3  @td Nb3  @hp O2  @z P{  \r SG   \hn Tj  \v U
,   2  :� +G   �3  @c ,,  @bb -,  @tb .b3  @hp /2  @z 0{  \r 3G   \hn 4j  \v 5
,   FG _G   �HE     �      ��5  Lb `,  -q #q Ln aj  �q �q Ls bj  Ir Er Ld c�5  �r �r Le d�5  �r �r Lt eb3  �r �r ^m f,  � ^hp g2  �^hn h�5  �Lv i,  ;s 5s Ja qj  �s �s _c r�5  ��}Jf sj  ?t 1t Jg tG   u  u Jh uG   �u �u Ji vj  �v {v Jj wj  &x �w Jk xG   �y �y Jl yG   Pz Bz H� zj  �z �z Jp {
,  r{ .{ Jq |2  �~ �~ Jr }�  " �~ _u ~
6  ��~Jw G   )� � _x ��5  ��~Jxp �
,  �� � Jy �G   ;� '� Jz �j  V� B�  �  j   j  
6  !@     2  6  !@    `"  �RE            �l6  3)"  }� y� 35"  �� �� >�RE     �:  -U�U-T�T  `B"  �RE            �7  3S"  �� � 3_"  4� 0� 3k"  q� m� 5w"  �� �� 7�"  �l5�"  !� � .�RE     �:  -U�U-T�Q�����T����-Q�l  a -  �UE     �      ��8  3-  d� X� 3-  �� � b1-  pc%-  ��  Ur/  =VE       �g }28  3�/  �� �� 3�/  � ۈ 3�/  0� *� 4�g 5�/  �� y� X@VE     �7  -T1-Qp X]VE     �7  -T8-Q
� XyVE     �7  -T1-Q}  ,�VE     �/  8  -Uv -Ts -Q0 XWE      8  -Tv  C5WE     -Tv    X�UE     K8  -T1-Q( ,�VE     �-  c8  -Us  ,WE     >-  {8  -Us  .HWE     >-  -Us   `�  �sE     �      ��:  3�  � ݉ 3�  �� �� 3�  �� t� 3  +� � d   d   W�  �m �9  e�  3  Ό ƌ e�  e�  4�m 5  7� +� 5  �� �� f+  g<   n 5=  � ލ ,�sE     *;  l9  -U} -Q|  ,tE     *;  �9  -Qv  .*tE     �  -Us     2�  @tE      `n �,:  3�  1� -� 4`n 5  i� g� 5  �� �� h  �tE     O       :  5  ͎ ǎ .�tE     �-  -Us  8OtE     �:    iL  stE       stE     m       3k  $� � 3^  �� �� jstE     m       5x   �� 5�  �� �� .�tE     �  -Us     kF\  F\  �k�K  �K  vl9  9  cl�P  �P  �lF  F  mkkA  kA  {l-4  -4  �l _   _  hl?U  ?U  �lE1  E1  rm�D  �D   n�1.1.4  �   �r  �  h $"  `yE     �      � X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  �
  8"W   	  K�   �   	�  L�   	�  M�   S  -  �  
>   G   �  B"K  Q     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  ?  -      n�  �  �  ?  U    �  ��  �  U     ?  -   -   U    �  �"    �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S'  0R�  U?  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��  �  @       @     @       �  
2  4  :  E       :-   B   s�  M   uE   }  uE  V  vE  /  vE   t
  xQ  k	  (  �  N    ��  N   �  	G   B� 
  L  +       s     v	  U     
�  �    =  N   �n  �   M
  pmoc5  stib	  ltuo|  tolp 
	  �0  
b   "�  �  �  %  <�  x >$   len ?+  *� @    
%  B�  �  
  `�  �  	  G   G   	  U    �  
�  q  "  G   ;  G   G   U    
�  H  N  c  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  �  ()  �;  0R   �U   8�  ��  @ +  �  
�  �c  �  
�     "  G   6  U   6   {  
�  I  O  Z  {   
�  ?g  m  �  {    @    
�  Y�  �  G   �  {  @   U    
s  ��  �  G   �  {  �   
  W  0�>  �  �n   e� �  �� �Z  �� ��  �� ��   �� �<  ( 
�'  ��  �!  l   �  -  �   �  �+  �  �G   
  �N   �  �-   \#  �@   
�  ,G   
�0  D4   N   
�
  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �  	�%>  N   
�S    � � " & � �
 �  � 	]
 
x	 � � � n �
  �	 � �   i !Z "$ # $� %Q &� '
 (C 0� 14 @ A� Qg R� S� T�	 U� V� W� XB ` a* b� c� pT �� �� �
 �� �� �� �c	 �� �O	 �� �� �t � �
 ��	 �k �Y �> �� ��
 � �� �� �2	 �J �/
 �> �� �	 �� �> �p �� �� �� �4 � �8 �> �� �g �� �� �  �v ��	 � O N   2~  �
   � '  \ 9S  � �q�   t  s~   m tv  x v�  Y w�  * x�  � yK   u
 z�  (�� |�  0�� }v  4t ~�  8�� ��  <d ��  @& ��  D� ��  H�	 ��  L} ��  P��  ��  X  ��  `Q
 ��  h4� ��  p� ��  x~0 ��  �� ��  ��% �  �R�  �?  � ^  �  @    j  ^  ^  	  @   ?  
 ��  � �!  �  � F�  �% H   Jy  I  R�  J?  lzw K	  B� M�  � pos N�  �!y�  O�  �!�� P�    ^  �  "@   � � R�  '  #�  �   E     �      �A  $�l      P� H� $B�  �  �� �� $0  �  5� +� %E  �  �� �� %�	 �  �� �� %� �  � �� %} �  :� � &�u  �dE     'Eof ��E     &� A�E     (`q   )�� ^  ��*c 2  +A�E     (  �  ,T2 +_�E     5    ,T��,Q1 -ǀE     T  ,Us   ( q �  .c =2  l� `� %� >�  � � +�E     T  e  ,Us  +́E     �  }  ,Us  +��E     �  �  ,Us  -�E     �  ,Us   /e  �E     �q �0v  � � 1�q 2�  U� O� 2�  �� �� 2�  �� � 3�  ��+!�E     B  (  ,T3,Q��,Y�� -N�E     N  ,Q��    4V �0~E     �       ��  5�l  �"  1� +� 6R�  �?  � }� 7K  O~E     �p ��  0X  �� ��  +�~E     Z  �  ,Uv  -�~E     Z  ,Uv   42 �`|E     �       �K  5�l  �"  ˙ Ǚ 8�% �"  T9K  �|E     �|E     )       �0X  � �   :\ �e  ;�l  �#   <^ �G   �  ;�l  �)  = ��  =6^  ��  =R�  �?  =� ��   >� wG   `{E     �       �T  5�l  w(  0� &� 1 p 6R�  {?  �� �� ?� |�  �\6 }�  � ߚ 66^  ~�  ;� /� -�{E     B  ,T1,Y�\   >� <2  �yE     �      �#  5�l  <&  ћ ɛ 6�� >�  >� 0� 6x  ?�  � ֜ @p @�  �� }� 6E  Av  Н Ν A#  3zE     �o Z04  �� � 1�o 2@  1� -� -QzE     5  ,Ts    <�	 G   M  ;�l  $  =.� �   #^ [�   }E     $      ��  $Jy  [!  q� g� $�% \!  � � B� ^�   %R�  _?  c� _� .zip `�  �� �� &�u  ��}E     C�  �}E     `p {|  0"  C� ?� 0  }� y� 0
  �� �� 1`p 2.  � � 2:  -� '� DF  +�}E     O  `  ,Uv  -~E     �  ,U~ ,Tt    +0}E     O  �  ,Uv  +e}E     f  �  ,U| ,T
,Q�L -�}E     Z  ,U| ,T}   E�	 N@    �E     ,      ��  $Jy  N%  |� x� $x  O%@   �� �� $B� P%  <� 4� $.� Q%@   �� �� .zip S�  3� /� /�  ;�E     �q V0�  s� i� 0�  � � 0�  T� J� 0�  ͤ ɤ 1�q 2�  � � 2�  �� �� F�  ��E     G�  �q �  2�  ե ϥ Cg  �E     0r (f  0x   � � 10r 2�  I� C� 2�  �� �� 2�  �� �� -�E     �  ,Us,T~ ,Q
    +��E     r  ~  ,Q|  -��E     r  ,Qv   C�  ��E     `r   0�  � � 1`r 2�  � � 2�  .� ,� 7K  �E     �r �   0X  S� Q�  -�E     (  ,T0   /  b�E      �r 0"  �� x� 0  (� $� 1�r 2.  b� ^� G:   s r  2?  �� ��  HL  0s 2M  Ǩ �� 2Y  /� )� +��E     �  �  ,U ,T0,Q
  -�E     �  ,U ,T0,Q~        I@ ;�~E     L       ��  $Jy  ;#  ~� x� .zip =�  Ω ʩ %R�  >?  	� � C�  �~E     �p Dx  0�  B� @� -�~E     A  ,Us  -E     Z  ,U| ,Ts   <� ��    Jzip ��  Jpos ��  ;B� ��  ;.� ��  =E  ��  =� ��  K�u  -LM� �    <� ��  g  Jzip �(�  ;.� �(�  =� ��  NL  =� ��   L=� ��  =_ ��    <9 ��  �  Jzip �(�  Olzw �  =.� ��  =� ��   <		 ��  �  Jzip �"�  =Jy  �  =� ��   P� ��  Jzip �!�   <� l�  O  Jzip l!�  ;Jy  m!  ;�% n!  Olzw p  =� q�  Q�u  � >�
 W�  `yE     c       ��  5Jy  W#  s� e� 6� Y�  � � ?�; Z�  �nR�u  fsyE     +oyE     (  �  ,Us ,T0 -�yE     }  ,Us ,T�n,Q2  ^    @    SK  0|E     *       �(  TX  U U9  9  cU�R  �R  �V�6  �6  �V�Z �Z VF\  F\  �V�K  �K  vW�D  �D   UE1  E1  r �  'x  s�  �A $"  P�E     *�      (� :G  �9   SX  ^� �L   S�i tint S�i u{S @�   g
  �       	@   v  #	@   �  &	@   |
  )	@    h  ,	@   (�  -	@   0�	  2S   8�  5S   < �   S�  "�   �
  8"c   A  K  �   A�  L  A�  M  SS  S-  S�  "<  >   S   �	  	Z   � S   e- Z   �  B"�  �     ��  R   �a    �� ��  �N ��  �6  �   �  Y�  �  a   �  |  9      n    $  |  a    �  �$  *  a   H  |  9   9   a    �  �"T  Z  �   PJ�  2�  LW   �  ML   Epos NL   �  P  SF  Q   �1 R'  (=9 Sd  0R�  U|  8y�  VW  @�� WW  H j�  �  k�\ �9   km  �a    o  ��  �  �3  9  L   W  H  L   W  L    ]  S�  2  q  w  $�  H     :9   �  J�  +x L�   +y M�   )  O�  "�  B   s  M   u�   }  u�  V  v�  /  v�   t
  x�  k	  (�  �  Z    ��  Z   �  	S   B� 
W  L  <    ]  s  ]  v	  a     �    "�  �  (N  �  P5   Z�  Q5  �  S  s  T�   [  U  ?1  WS     �  5    Y�  �  Z=  Z   �b  �   4M
  pmoc45  stib4	  ltuo4|  tolp 	  �$  b   "|  �  U�  %  <�  Ex >5   Elen ?<  *� @]   %  B�  "�    `�  �  $�  S   S   �  a    �  �  q    S   /  S   S   a    �  <  B  $W  S   S   a    �  `��  �  ��   �% ��  ?1  �S   �&  ��  !  ��   I  �  ()  �/  0R   �a   8�  �  @ �  �  v�  �W  "�  �       S   *  a   *   o  �  =  C  $N  o   �  ?[  a  $v  o  W  L    �  Y�  �  S   �  o  L   a    s  ��  �  S   �  o  �   �  W  0�2  �  �b   e� �  �� �N  �� �v  �� ��   �� �0  ( �'  ��  �!  l]  "?  �  �a  "P  S�  -  �]  "h  t  �  ��   "  �
  �5  �  �<  "�  �  �S   "�  
  �Z   �  �9   \#  �L   �   9   �  ,S   \&  7a   �0  D@   �H  Q-   b   �f	  Exx ��   Exy ��  Eyx ��  Eyy ��   a  �#	  "f	  z'  ��	  m  �y   ss  ��   �  �x	    ��	  �	  $�	  a    �  ��	  �U  �a      ��	   %  ��	  �  $
  
  �   R
  �� "
   �@ #
  �U  $a    �  7}
  �; 9
   ��  :
   L  <R
  OZ   ,��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=L  ��  ?�   �  @�  ~  B�  �  C�  �  D�   5  F�  (B  G�  0�  H�  8 �	  J�  
   s�  �  u�   ��  v�  �  x�  �
  z�  (  {�   �  }Y  �  �#�  �  Pk  `�}  R�  �|   (  ��  |  ��  �  ��  �  ��  �  �"$  
v  �}
  
�  �#  (
�%  �}  0
7&  �2$  8
G   ��  X �  �"�  �  h  �  �M �#   k  �  R�  |   �  �"�  �  %  8;#  �� =$   �M >�    ?}
   r$  @�  0 5  �$0  6  %  ��  �� $   �M $  �  b   �  8  (�� 
o  h�� �  p�� �  x K  � �  �  �  �,{  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9�  8  :  @�  <�  H�  =	  PE-  ?�	  X�!  D  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  R{  ��� S2  �K1 W�  �R�  X|  �Jy  YH  �%  [}
  ��	  ]�	  �    ^a   ��8  `k  � L   �  �    X��  �  ��   E-  ��	  N ��  �8  �  P �  *%�  �  P�  0t2  k  v�   �  w�  �@ x�  ݖ y�  E-  z�	   N |L  0�  }�  pR  ~�  x�  �  �ߣ  �b  ��I ��  ��  ��  �h  ��  ��S  �  �4  ��  �8  �  �
  �a    
�  �9   
�  ��  
o  ��  
�L �a    
�8  �c  ( �
  L#?  E  W  H�  �  J�   = KQ    L�  d  M�   Z�  Z   �Q  �   4�  bmys4=  cinu4�  sijs4w    bg4O  5gib4p  snaw4M  ahoj4�    bg4�  sijs4�    bg4q  5gib4�  snaw4�	  ahoj4  BODA44   EBDA4�	  CBDA4  1tal4�  2tal4   nmra �	  �  (0  OE  #   g)x  ~  �   ���  =  �f	   L  ��   $  ��  0�  �'   8m  �#�!  h�  �P  pآ  �H  tG   ��  x   �  2  �?  d�  �
  �))  /  �   H�h  �  �a    "  �	  �!  ��   ~	  8f�  �
  h�   (  i�  �� k�  �� l�    n�  �  o�   �  p�  (�  q�  0 y  sh  �a  ��    �$    �  0'c  �N  )�   ?1  *�  }0  +�  i/  ,�  � -f	   �  �)p  v     H��  ��  ��   ?1  ��  (  �?  4  �f	  \  ��  0  �a   @ ��  ��  +!    Etag �   �U  �   �  �    Z`  Z   
\  w%   }#  �&  h  �  &     
$  E   9
�  � ;
\   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  i  Z�  Z   �	  :   �   ^$  1  �!  �!   :  ��  �  ��  �#  �.  4  �  C  }   I$  �O  U  $`  }   �&  �l  r    �  }  �   �   "�  �!  H�  �  ��   S"  ��     �  �"  ��  �  ��   ;  ��  (%  �"  0�   �C  8��  �`  @ �  R  ��  "  x  =�	  H  E#I  "8  �  @J�  �  L�   �  Mb  �� O  .� P?  �  Q�   �  R\  (�!  S�  08'  T�  8   W!�  �  -  (l  k  n�   �M o  ߣ  pb  �  q�   D  k  )%  +  �  ?  �  �   w   .K  Q  $\  �   �  1h  n  $�  �  �     s	  K  6�  �  $�  �  �     �  :�  �  �  �  �  �   �  >%  "  Y�  �  �    #  �  	     �  _  %  �  C  #  �  �     $  fO  U  $j  #  �  �   �  lv  |  �  �  #  �  �   #  x��  �� �    �  � b  H  � �  P�  �   X9!  � C  `l� � j  h  � �  p 2    ��  �  H2_  �S  4   �  5  (  6  04  7�  88  8  @ �  :  �  �=�  R�  ?|   �  @�  n  A�  �  B�  1$  C?  2�  E_  �� F_  `�L Ha   � �  J�  k  P   �    �  (  H  �  �  �     �  &4  :  $E  �   �%  *Q  W  �  f  {   �%  -r  x  $�  {   {  1�  �  �  �  �   �  4�  �  $�  �   l  8�  �  �  �  {  �   �  <�  �  �    {  �   �  @    �  =  �  {  �  H   �  GI  O  �  m  �  �  �     �'  Ny    �  �  �  H   �  S�  �  �  �  �  �  �  H  �   �  &  ���  �� �   i'  ��  H   ��  P  ��  X�A ��  `Y �(  h�#  �E  p�  �f  x�  ��  �  ��  ���  �  �U�  �=  ��!  �m  ���  ��  ��  ��  �&  ��  � �&  ��  �  a   �  0t'   �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�  �  U'@   F   Um  D   t�   �  v�   A  w�  �  x�  &  y�   !  {K   �  ��   �   �  �   4   �  �    �	  �  ��   �   $�   4   �    �'  ��   �   �  !  4   �  ?  !   �   �!  [!  ��  )�    ��  )�   �  )�    }  "!  "[!  O  ;�!  _� =%�!   ݰ  >%4    h!  �  @m!  �!  cA  �,�!  �!  /  ��!  �� �^   �M ��!   ?<  �,�!  �"  �5  P��"  �  ��   �� ��"  �Y ��"  �H ��"  U@ �#   �9 �#3#  (�A  �#c#  0�^  �#�#  8�^  �#�#  @N7  �#�#  H "�!  ��  ��!  (Z  ��"  �"  �  �"  �!  �   17  ��"  �"  $�"  �!   �G  ��"  �"  �  #  �!  U   %G  �#  #  �  -#  �!  -#   U  �@  �?#  E#  �  c#  �!  �!  U  U   �;  �o#  u#  ?  �#  �!  U  U   �W  ��#  �#  -#  �#  �!  |   *;  ��#  �#  -#  �#  �!  |  U   �T  ��#  g�  ��!  "�#    �  �    -1  B�  }  2$   L    +  B$   L    w�  �%2  �  8 Y�$  ��   [�   Ǧ   \�  ��   ]�  d>  ^�  ��   _�   I�   `�  (�   a?  0U   b�  2�   c�  4 ��   eO$  ��   p$�$  O$  ��  � �C&  ֤   ��   Ğ   ��  ��   �h  �   �h  	��   �h  
�   �h  ��   �C&  �   �S&  (��   �C&  <�   �S&  X��   ��  p��   ��  x��   ��  |��   �c&  ��   �c&  �R�   �h  ���   �h  ���   �?  �F�   �?  �V�   �s&  ���   �s&  ���   ��  �"�   ��  ��   ��  �@�   ��&  � �  S&   L    �  c&   L   	 �  s&   L     �  �&   L    �  �&   L    ��   ��$  o�   �#�&  �$  �   ��&  ��   �&  2]    h   U�   !�&  5�   "�   �  �   $�&  P��    *�'  m�   ,�   `h   -�  �   /�'  #�   0�'  (��   1�'  �
�   3�  
z�   4�  
��   6(  
��   7(  �
�   9�  (
Ԯ   ;'(  0
��   C7(  �
��   D�  � �  �'   L    �  �'   L    �&  (   L    �$  (   L    �&  '(   L    �  7(   L    �  G(   L    ��   FT(  	'  Z�  Z    0�(  ��   r�  �  E�  Ϊ   H�   8Z(  ��  !)$�(  �(  UH�  ��  !,�(  �(  �  �(  |  �(  �(   �&  �(  ��  !1�(  �(  $)  �(  �  �  �  �   ��  !8$)  *)  $5)  �(   �  !;j)  M� !=�(   �� !>�(  Յ !?)   ��  !Av)  5)  �  !h!�)  �)  U��  ��  !u-�)  *  ��  8!V*    !X|)   j�  !Y*  =9 !Z�*  �� ![8*  Q� !\_*   �� !]k*  (�� !^�*  0 "�)  ��  !�'*  -*  $8*  |)   ��  !�D*  J*  $_*  |)  �  �   K�  !�D*  å  !�w*  }*  $�*  |)  �   ��  !
�*  �*  �  �*  |)  �   ?�  !1�*  �*  �  �*  |)  �*  �(  	     1�  !�!�*  �*  U$�  ��  !�-+  �+  .�  8!��+    !��*   j�  !��+  =9 !�,,  �� !��+  +�  !��+   �� !�,  (�� !�S,  0 "+  ǡ  !��+  �+  $�+  �*   ��  !��+  �+  $�+  �*  �  �  �   ��  !��+  �+  $,  �*  �  �  y   !�  !&,  ,  $,,  �*  �  y   K�  !D9,  ?,  �  S,  �*  �   	�  !k`,  f,  �  �,  �*  �*  �(  	   ��  !��,  ��  !��,   X� !��,  l� !��,   j)  �,  }   �,  �)  �,  }   �,  +  �,  }   �,  $�  !��,  �  !� -  �,  j�3  "5B-  Qnum "7�  Qstr "8�   +P  ":-  �J  "=v-  +key "?B-   �U  "@@    �7  "D$�-  N-  O  "H�-  �-  �  �-  �-   B-  �Z  "K�-  �-  ?  �-  �-  �-   �S  ("O1.  �� "Q�   �  "R�  �6 "S�  �B  "U�-  3  "V�-  >) "X1.    v-  e-  "\ C.  �-  ��  ##U.  [.  U  j.  �   d�  #)v.  |.  �  �.  �   0�  #/v.  K�  #6�.  �> #8U   �^ #9�   �  #;�.  Ѽ  #>$�.  �.  ў  (#@/  
H #B�"   ��  #C�  XT #D/    �.  ��  #N$/  */  �  >/  �  �   B�  #VJ/  P/  $`/  �  �   ��  #Zl/  r/  �  �/  |  �.  �  /  >/  �   ��  #b�/  �/  �  �/  �.  U   ��  #f�/  �/  U  �/  �.  -#   ��  @#j\0  �\ #l I.   8` #n `/  �\ #o �/  �_ #p �/  �T #r j.   }�  #s �.  (ʬ  #t s0  0�  #u s0  8 "�/  ��  #jm0  \0  C  7�   $F�0  ~�  $H�   ̰  $I�  V�  $J�  �H $L�0  �  $M�0   �  �  b�  $Oy0  �  $O�0  y0  ��  $W1  ��  $Y�    ��  $[�0  L�  $^u2  �  $`�$   8�  $a1  8-�  $b�&  @�  $c�   E�  $e�(  (= $f�0  0�  $hu2  P
�  $iu2  X��  $ju2  `��  $l�  h��  $m{2  ph�  $n�2  x��  $o7.  ��  $q�  �V $r�0  �� $s{2  �'�  $t�2  ���  $vh  ��  $wh  ���  $xf	  �w�  $y�  �;�  $z  �* ${�   ܲ  $}�   h  u2  �  �  $1  �  $�2  1  ��  ($��2  �9  $��   ��  $��  ɲ  $��  �  $��  �  $��    T�  $� 3  �2  ��  $�D3  ��  $��   ��  $��  +x $��  +y $��   �  $�P3  3  z�  X$��3  ��  $�?   ��  $�  �Z  $��  (%?  $��  0L�  $��2  8)�  $��  @W�  $�D3  HѺ  $��  P b�  $��3  V3  �  $�!�3  �3  L6�  x$��4  �� $�   �6  $��2  �s  $��  Q  $��  Y�  $��  B�  $��4   �  $��4  @�  $�G(  P�  $��  X�  $��  \�  $��  `�  $��&  h2�  $��  p ^  �4   L    2  �4   L    �6  `%S�5  �<  %U�   �Q  %V�  a(  %X�  VA  %Y�  Q) %[�   nX  %\�  "�D  %^�5  (�5  %_�5  8M   %a�  H}  %b�  JV  %c�  L/  %d�  N7K  %f�  P>D  %g�  R�:  %i�  T�3  %j�  V=]  %k�  X �  �5   L    �5  %m�4  �Q  8%��6  �  %��   �Z  %��  %?  %��  
L/  %��  �<  %��  �Y  %��  �7  %��  �)  %��  �O  %��  �H  %��  vH  %��  ^  %��6  �>  %��  $�7  %��  &0>  %�a   (�+  %�a   0 �  �6   L    �H  %��5  �?  8%A�7  �  %C�   �Z  %D�  %?  %E�  
L/  %F�  S.  %H�  �W  %J�  �W  %K�  C  %L�  �O  %M�  �H  %N�  vH  %O�  ^  %Q�6  �>  %S�  $�B  %T�  &0>  %Za   (�+  %[a   0 �]  %]�6  �B  �%|:  ��  %~�   �)  %�  �)  %��  �.  %��  U  %��  �V  %��  
�0  %��  �6  %��  �C  %��  U?  %��  6P  %��  �C  %��  &L  %��  *J  %��  �L  %��  HP  %��  N*  %�:   [2  %��  0k2  %��  8.  %��  @{2  %��  HQ2  %�:  P�0  %��  Tp4  %��  VmU  %��  X�Z  %��  Z ?  %��  \:  %��  ^�I  %��  `E8  %��  b�;  %��  h�;  %��  p�O  %��  xDF  %��  zfV  %��  |�9  %��  ~[9  %��  ��G  %��  �zQ  %��  � h  :   L   	 P  !:   L    {D  %��7  �1  @%��:  �I  %��   6Y  %��  �^  %��  S  %��  )  %��  @3  %��   �0  %��  (4C  %��  0�C  %��  8 aM  %�.:  �I  @%��;  �  %��   _7  %��  )  %��  �O  %��  �n %��  �T  %��  EF  %��  I  %��  �K  %��;  N:  %��;  ,L  %��;  4�E  %�P  :�Z  %�P  ;�Z  %�h  <^  %�h  = P  �;   L    P  �;   L    P  �;   L    eU  %��:  �9  (%7�<  ��  %9�   a@  %:�  b<  %;�  
8  %<�  .  %=�  �H  %>�  �Q  %?�  X  %@�  �.  %A�  �;  %B�  ))  %C�  eH  %D�  I_  %E�  �B  %F�   !3  %G�  " �)  %I�;  �  &I	=  F@ &K�   I�  &L�  K�  &M�   ԃ  &O�<  �b  h&hJ=  `h  &j�   m�  &k�  dh  &lJ=   	=  Z=   L    ��  &n=  �j  0&��=  F@ &��   I�  &��  +def &��  K�  &��  +tag &��   c  &��  ( )�  &�f=  �  &�>  �  &��   c  &��  Cg  &��   �~  &��=  z�   &�^>  `h  &��   m�  &��  L�  &��  dh  &�^>  e  &�d>   �=  >  J�  &�>  �R   'F�>  +tag 'H�   ��  'I�  .� 'J�  �P  'K�>   �  DG  'Mv>  f3   '�?  +Tag '��   Q  '��  .*  '��  �K  '��   gW  '�?  �>  �^   '�?  k@  '�   aE  '�  p0  '�  �>  '�  H  '�  �/  '�  �� 'u2   �F  '?  �<  '0�?  H  '2�   �/  '3�  �� '8u2   qS  ':�?  A9  0'US@  ߣ  'W�   �E  'X�  �^  'Y�  =Y 'ZS@  <  '[�  �=  '\Y@   Jy  ']H  ( �?  �?  rY  '_�?  �1  '~�@  �.  '��   �L  '��   Z  '��@  l@  �V  '��@  ��  '��   f>  '��  Y  '��@   �)  '��@  �A  '/�A    '1P   �  '2P  �N  '3h  o=  '4P  D4  '5P  �^  '6P  `*  '7P  �0  '8P  �G  '9P  �D  ':P  	I:  ';�A  
 P  �A   L    �@  '=�@  �\  '�B  +  '��A   Y�  '��A  �
  '�h  (  '�h  �F  '�h  �C  '�h   <)  '�&B  �A  �,  'sB  �  '�   AK  '�  z8  '�0  V 'sB   yB  P  �R  ',B  	F  '.�B  �  '0�   �P  '1yB   ">  '3�B  x'I�B  l�K 'KB  l`B 'L�B   �[   'EC  �z  'G?   =Y 'N�B   �6  'P�B  O]  'a!.C  4C  U�(  7N  ('��C  >) '�u2   -N  '�u2  V` '�u2  TE  '��  �/  '��   �z  '�?  $ G  '�9C  &8  '� �C  �C  PeS  p'oH  �� 'q   ^  's�>  �
�^  'u�  
[>  'v�   
�W  'w?  (
� 'y�5  0
�=  'z�6  �
�,  '|�<  �
��  '~?  �
�(  '�7  �
AK  '��  0
XL  '�_@  8Jos2 '�!:  h
p�  '��:  �
T  '�u2  0
#9  '��  8
!H '��I  @
�+  '�'J  H
@.  '�zJ  P
�E  '�XJ  X
�P  '�XJ  `
@  '�XJ  h
$S  '�a   p
s  '�a   xJmm '�a   �Jvar '�a   �
Q  '�a   �
<B '��@  �
2Y '��;  �
=  '��  �
=  '�B  �
UV  '�C  �
�(  '��  
=  '�u2   
/:  '��  (
�?  '�u2  0
�]  '��  8Jcvt '��J  @
�R  '�H  H
5$  '��	  P
��  '��  `
HT  '��  h
�*  '��  p
�J  '�?  x
�+  '�?  y
�  '�!C  �
�C  '�U  �
�-  '��  �
j7  '��  �
kN  '��  �
�F  '��  �
#7  '��  �
�(  '�u2  �
rE  '�u2  �
QZ  '��  �
4  '��  �
�@  '��  �
:L  '�u2  �
�G  '�u2  �
�]  '��  �
�W  '��J  �
�/  '��  �
�B  ' �2   
�I  'u2  
s-  '�  
�*  '�  
,  'U  
,  'U   Jbdf '	�C  (
�T  '�  P
#F  '�  X
�U  '�  `
�K  '�  h �=  '�H  #H  �  2H  a    �Q  '�"?H  EH  P�\  x'c�I  �  'e�C   �  'f�K  )�  'g�  �V  'h�  :1  'j�   �^ 'k�  (Jy  'mH  0�  'n�  8�  'p�  <�!  'q  @R0  'r�  `�  's�  duN 't�  h6  'u?  lEpp1 'v�  pEpp2 'w�  �2�  'z�K  �Xc  '{�K  �
�6  '}�K  
)  '~u2  
�8  '�   
�L '�a   (
C  '��  0
��  '��  4Jpp3 '��  8Jpp4 '��  H
y�  '�u2  X
�� '�u2  `
U  '�}
  h �I  '�J  	J  �  'J  �C  �  H  �>    1  '4J  :J  �  XJ  2H  �  �  �   �M  '+eJ  kJ  �  zJ  2H   �<  ':�J  �J  $�J  2H   Zy*  Z   '=�J  4   �^  J  b8  �T   lK  'H�J  �  |T  @'?�K  R�  'A|   �  'B�  n  'C�  
Z�  'D�  �  'E�  Eorg 'G  Ecur 'H  ��  'I   s  'Ku2  ([  'L�0  0c+  'N�  8 R8  'P�J  RG  'T'�K  �K  U[  O  '_ �K  �K  ULL  ͳ  @(@FL  Jy  (BH   �S (C�  ܱ  (D�  .� (E�  ��  (Fh  ��  (G�   
�  (H�  (�P  (J�>  0Ӏ (Ku2  8 ,�  (M�K  L
�  (P�L  ߣ  (R�   x  (S�  .� (U�  ē  (V�L   � (W�L   �  �L   L   � ��  (YRL  ��  ((\M  ߣ  (_�   x  (`�  ē  (b�0  ��  (c�0  Ӷ  (e�   �  (f�  $ r�  (h�L  W�  (mOM  Kw  (t�   7�  (u�2   0�  (w'M  j�  ({�M  ��  (}�   �  (~�  �w  (�   J�  (�[M  1�  (��M  �{  (��M    �M  �  (��M  �   (�N  ��  (��   k  (�N  �q  (��   q  (��  y|  (�N   OM  �M  �  (��M  ��  (�<N  �M  %�  (�!NN  TN  P�  �(M�P  k  (O�   Jy  (PH  R�  (Q|  ��  (R�  �   (S�   �  (T�  $(  (Vh  (|  (Wh  )x�  (Xh  *п  (Z�  ,�J  (\?  0i�  (^FL  8�  (_FL  xC�  (`FL  �= (b�L  �
��  (cM  
p�  (eFL  8
��  (fFL  x
=�  (gFL  �
��  (hFL  �
�  (j�  8
��  (m{2  @
V�  (p�  H
V` (q{2  P
��  (ru2  X
��  (s�  `
/�  (u�V  h
��  (v�  0
��  (w�V  8
j�  (y�V  8
2�  (|	-  X
s  (a0  `
��  (��  h
�  (��V  p
d�  (��  x
|�  (��  �
˽  (��	  �
ʞ  (�$N  �
8�  (��V  � ֥  0(�Q  ��  (�?   �  (�?  v�  (�BN  �  (��  ݺ  (��  ��  (��  c�  (��   +BV (�Q  ( H  �  (��P  ��  (�6Q  "%Q  �P  L��  H(�kS  ��  (��   Ǧ  (��  @�  (��  ��  (��  d> (��  ��  (��  �  (�?  I�  (��   U  (��  (�  (��  0��  (��  8�& (��  <��  (�f	  @?�  (�?  `U�  (��  hw�  (��  p֤  (��  �;�  (�  �ܲ  (��  �w�  (��  ���  (��  ��  (��  ���  (��  �ٛ  (��  ��  (��  �g�  (��  �`�  (��  �x�  (��  ��  (��  �|�  (��  ���  (��   �  (��  n�  (��  ��  (��  ��  (��   `�  (��  (�  (��  0m�  (��  4�m  (��  6A�  (��  8��  (��  @ ��  (�<Q  S�  (�$�S  �S  P��  �(*LT  Ҳ  (,kS   
-�  (-V  H
�  (0Q   
ݺ  (1�  PJNDV (2�  X
�  (<u2  `
K�  (=u2  h
�  (>�  p
��  (?�  t
��  (AFL  x
Z�  (B{2  �
l�  (EU  � LE�  �(��U  ��  (�h   �  (�h  ��  (�h  �  (�h  ��  (��U  �  (��U  x��  (��U  ��  (��U  8��  (��  ���  (��  ���  (��  ���  (��  �
�  ( �  �
R�  (h  �
��  (h  �
V�  (V  �
��  (V   
��  (?  �
6�  (�  �
Ğ  (�  �
"�  (	�  �
��  (
�  �
Т  (�  �
P�  (�  �
W�  (�  �
��  (�  �
��  (�  �
��  (wS  � �  �U   L    �  V   L   	 �  V   L    ��  (LT  ��  (6V  LT  a�   (�V  ߣ  (h   �  (�  �U  (u2  
�  (�  w�  (!�  .�  ("�  �  (#h   �  (%<V  �  (%�V  <V  9�  (G�S  wS  �V   L   � �$  1  8�  `),W  �� ).�   -U )/�  X `�  )1*W  �V  L~�  H)<�W  �� )>�   �� )@?  0��  )A?  1�� )C�  8�� )D�  @ Z�  )F�W  0W  L@�  )Q�W  �  )S�(   ��  )T�W   �(  �W   L   � ��  )V�W  �W  �C  h**0X  �� *,$   �Z  *.�  8�  */?  <X;  *00X  @آ  *1H  ` �  @X   L    �D  *3LX  �W  ��  *?-^X  dX  ۳  `*��X  ��  *�u2   y�  *�		  �� *�		  �� *��  ��  *��   Ǩ  *��  $(2 *�{2  (Ϛ  *��2  0R�  *�|  8_� *��Y  @ ��   *T6Y  �� *WOY   �Y *\`Y  +add *_�Y  �x *e`Y   �  OY  RX  �  |   6Y  $`Y  RX   UY  �  �Y  RX  �  a   �   fY  r�  *g�X  "�Y  �  *�"�Y  �Y  ��  �*�Z  y�  *�u2   2�  *�u2  �� *�u2  � *��  R�  *�|   _� *�.^  ( ��  *�"Z  "Z  ��  *�WZ  �S *�u2   �� *�u2  � *�)[   ��  *�"hZ  "WZ  nZ  ��  0*��Z  9�  *��   �{  *��[  � *��[  ��  *�	\  x  *��  �  *�h  m�  *��   �  *��  $��  *�  ( V��  Z   *�)[  ˟   .�  ��  ��  ��  ��   ��  *��Z  ��  *�"Z  VL�  Z   *��[  ��   ��  Ʊ  ��  ��  g�  �  ��  W�  �  	|�  
K�  ��   8�  *�A[  V��  Z   *��[  c�   ��  p�  �  �  ��  �  ��  ��  }�  	 ��  *��[  ��  *�\  \  $+\  �  �   [�  *nZ  �  h*k�\  �� *n]   �Y *t(]  �? *w(]  �2 *y(]  �! *|=]   �$ *~W]  (�* *��]  0�3 *��]  8k! *��]  @�A *��]  HV- *��]  P�F *�(^  X  *�(^  ` $]  �Y  u2  u2  |   �\  $(]  �Y   ]  �  =]  �Y   .]  �  W]  �Y  �   C]  �  �]  �Y  u2  		  �>  ?   ]]  �  �]  �Y  �  �J   �]  �  �]  �Y  �  �  �   �]  $�]  �Y  Z   �]  $�]  �Y  Z  �  �]   �  �]  �  (^  �Y  cZ  �  �  �>   ^  �  *�8\  ".^  ~�  *�M^  l�  p*J_  R�  *|   �  *�  )�  *�W  ��  *�  2�  *�*   �� *�*  (��  *�_  0��  *�_  8R0  *   @�  *!  H�!  *#�  P��  *$?  X�� *%?  Yb�  *&?  Z��  *(?  [�  *)?  \_� *+�_  ` ګ  *�u_  �� *��_   �Y *��_   $�_  �_  a   ?   @^  u_  $�_  �_   �_  �  *�J_  "�_  �  î  *B�_  2�  *Du2   �� *Eu2  y�  *Fu2   {�  *H�_  ��  *L`  `  �  6`  �C  �  {2  �>   l�  *RC`  I`  $^`  �C  {2  �   P��  �*Wyb  <0 *Y@^   4� *[yb  pJtop *\�  �
O� *^�b   
Xc  *_�b  �
��  *a�  �
�  *b�  �
�  *c�b  �Jcff *eBN  
�  *fwS   
˽  *g�b  (

�  *i�_  0
�  *j?  8
��  *k�  <
z�  *m�  @
�  *n�  D
��  *p�  H
�  *q�  L
~�  *s{2  P
9� *t{2  X
V *v{2  `
�  *w�  h
&  *y	  l
�J *{?  p
�  *}&`  x
��  *~&6`  �
s  *�a0  �
Ğ  *��  �
��  *��2  �
q�  *�7.  �
��  *�f	  �
w�  *��  �
�  *�G(  �
�  *��&  �
�  *��  � �  �b   L   0 �_  �b   L    �_  �  �b   L    �	  x�  *�^`  ջ  *�#�b  �b  �  �*�c  R�  *|   �  *�  )�  *�  ��  *�  2�  *�*   �� *�*  (��  *�  0��  *�  8R0  *�  @�  *�  P�!  *  `��  *�e  ��� *?  �b�  *?  ���  * ?  ��  *"a   �L�  *#a   �_� *%Qe  � ��  *��c  �c  �  d  �b  �   q�  *�d  d  $4d  �b  �  �  h   j�  *�Ad  Gd  �  `d  �b  �  �   ��  *�md  sd  �  �d  �b   *�  *�Ad  �  *��d  �d  $�d  �b   �  @*�,e  �� *�Ke   �Y *��d  �? *�$�c  kI *�$d  rL *�$4d   � *�$`d  (-1 *�$�d  0��  *�$�d  8 $Ke  �b  �  {  �  ?   ,e  T�  *��d  "Qe  Za�  Z   *��e  ��   J�  �  ,�   ה  *�ce  ��  *'�b   �  *F�e  y�  *Hu2   2�  *Iu2  �� *Ju2   ɠ  *L�e  ݬ  *L�e  �e  �  *O/f  f  P��  �*}�g  <0 *�e   4� *��h  �Jtop *��&  �
O� *��h  �
Xc  *��e  x

s  *�a0  �

�  *��  �

V *�{2  �

Ğ  *��  �

��  *��  �

��  *�{2  �

h�  *��2  �

��  *�7.  �

��  *�f	  �

w�  *��  �

��  *��  �

�  *��  �

�  *��b  �

�  *�G(  `
&  *�	  h
�  *��g  p
_� *��h  x
�  *��&  �
�  *��  �
�J *�?  �
˽  *��	  � �   *X�g  �� *[Nh   �Y *f_h  �; *o~h  � *u�h   �  *T�g  h  �  h  f  �   �  Nh  f  �  {  �  {2  G(  ?  	  �g   h  $_h  f   Th  �  ~h  f  u2  �   eh  �  �h  �h  u2  �   �b  �h  X�  *z�g  "�h  �  �h   L   � �e  �h   L    <�  *� �h  ��  �*�i  R�  *|   �  *�C  )�  *�W  ��  *�  2�  *�*   �� *�*  (��  *�  0��  *�  8R0  *�  @�  * �  P�!  *"  `��  *$?  ��� *%?  �b�  *&?  ���  *(?  ��  **a   �L�  *+a   �_� *-jk  � c�  *� j  j  �  j  j  �   �h  ˯  *�-j  3j  $Mj  j  �  �  h   N�  *�Zj  `j  �  yj  j  �  �   Ԝ  *�Zj  h�  *��j  �j  $�j  j   8�  *��j  �j  �  �j  j   p�  @*�Ek  �� *�dk   �Y *��j  �? *�%�i  kI *�% j  rL *�%Mj   � *�%�j  (-1 *�%yj  0��  *�%�j  8 $dk  j  �C  W  �W  ?   Ek  +�  *��j  "jk  !�  *E�k  2�  *Gu2   �� *Hu2  y�  *Iu2   ��  *K|k  Pj�  �*Nsm  <0 *P�h   Ecff *QBN  �4� *Syb  �Jtop *T�  h
O� *Vsm  p
Xc  *W�m  
��  *Y�  
�  *Z�  
�  *[�b  

�  *]�  �
��  *^�  �
��  *`?  �
�  *a?  �
��  *b�  �
�  *c�m  �
z�  *e�  �
�  *f�  �
��  *h�  �
�  *i�  �
~�  *k{2  �
9� *l{2  �
V *n{2  �
�  *o�  �
&  *q	  �
�J *s?  �
�  *uwS  �
�  *w&`  �
��  *x&6`  � �k  �m   L    �k  �  �m   L    1�  *z�k  l�  *�m  �� *�n   >'  *�2n  � *��h   $n  n  �C  W  �W  ?  	  `  6`   �m  �m  �  2n  n  W  �   n  U�  *��m  "8n  :�  *�#Wn  ]n  ,�  (*��n  R�  *�|   Jy  *�Go  � *��3  p�  *��o  o�  *�a     4�  *��n  �� *�	o   �Y *�o  gP *�/o   �  	o  Jn  |  u2  u2   �n  $o  Jn   o  �  /o  Jn    o  \�  *��n  "5o  ١  *�#To  Zo  ��   0�o  y�  2u2   2�  3u2  �� 4u2  % 6�   �  �o  �  		  a    �o  �  *�.�o  p  0�   *�p  ��  *��!   �0 *��!  ک  *��!  �> *��!   "�o  D0 *��o  "p  �  X*��p  b�  *!�p   �  *!�p  E�  *!�p  b�  *!�p  ,�  *q   h�  *q  (�  *2q  0��  *Mq  8c�  *�o  @:�  *!Sq  Hs�  *"Yq  P �Y  ;^  ^e  �h  $q  u2  		  �   �p  U  q  U   q  $2q  �h  a   ?   q  $Mq  �  �&  wS   8q  Bo  En  �G *,p   *"_q  "lq  V�I Z   +-	�q    �7 � � 2* �D  m+;�q  Qs +=�   Qf +>�  Qi +?�  Qu +@�  Qb +A?    D +8r  � +:~q   +u +C�q   t6 +E�q  �E +E/r  �q  OZ   ,�xt  �6  t � #? �2 � X CQ 2 J 	�9 
O 8 � ~1 �> � vH "I \. -( �;  �. !r8 "�K #�- $� %�D &;4 '= (A. 0�: 1�% @m= A�/ Q�" R�5 S�K TV+ U5R Vi, WG X�A `� a�" bY* c�' p�B �W) �C ��D � �FE �� ��# �I ��O �4, �v ��H �> �p ��< �;S �� ��< ��R �JD �NK ��F �� �MM � ' �4 �o# ��% �� �� ��# ��8 �;C �� �[C ��3 ��J �1% �N �> �UH �y �K � �.< ��4 � OZ   (�t  }L  uI & �C  Vs1 Z   �zv  ]F  6B s �@ > �& �1  # . ; 	� 
`6 �& �> D !' Y% �1 $ 83 Y8 �( �( RB �: �I �> � 6 �* $Q b( K7  
# !�9 "E2 #S2 $a2 %Q# &�K '$ (c# ) *�L +�# ,�I -= .nK /(+ 0� 1�O 2X/ 3g 4�L 5i> 6a@ 77 8�5 9iB :0F ;k <+M =S >CF ?W @e APF B� C�P DKG EXG F�R G�) H� I95 J�@ K � �t  �  �v   L   I "�v  !� �v  	�I     A� -%wk  Ak% -(�_  A�) -++&  Ab�  .)�Y  A�  .,;^  AE�  ./^e  Ab�  / �h  � 0&#w  w  �M 80(hw  
H 0*�"   �, 0,hw  P= 0-�.   �  0/�  (V 00nw  0 �  �  A H 06�#  A�= 09�#  =G 0D&�w  �w  e0 (0F�w  
H 0H�"   N� 0I�  .� 0J�  �8  0K�0    AP, 0Q�#  A�M 0_�#  F 1EH  "�w  OZ   ,�Lz  �N  �! �) �E � �Q pF �, �M �P 	�> 
g  C9 ) �0 �: p< }. K? �+ zN �  �) !�D "� #�@ $�5 %�2 &�7 'b& (�9 0� 1*@ @�? AF Qq@ RM S� T�O UY; V�. W, X�- `�9 aO: b�C cwP p�! �%A ��2 �� ��) ��/ ��O �% �Q ��< �n- ��E ��E �� � / �~? �. �n3 ��0 ��7 �,# �C' �� �pR �'P �4 ��' �1J �%> ��8 ��1 ��% �aR ��C �B ��" ��  �/ ��G �?  �� �3 ��6 �� �� �� ��L � �E 21H  V/  Z   2P}z  =M  A! �"  =- 2VXz  �& @33�z  R�  35|   � 36�z   38@   0= 39@   s 3:@    .� 3;@   (WR 3<@   0+ptr 3>a   8 �  �@ 3@�z  �. 3@"{  "{  �z  �'  4.j{  � 40�z   �S 41y  +end 42y  +ptr 43y   � 45({  �R 45�{  ({  D) 5=b  V�- Z   5A�{  '8 7K O �<  e 5L|  +a 5N�w   +b 5O�w  +c 5P�w  +d 5Q�w  +tx 5R�w  +ty 5S�w   �; 5U�{  "|  L�B �6?�}  R�  6A|   � 6B�  �E 6D?  !+ 6E?  l 6F�{  (O 6L|  * 6M|  ,�& 6N|  D:� 6O�w  \�  6RQ  `��  6So  �ݺ  6To  �+NDV 6U�  �8Q 6Wb  �T5 6Y�w  �p5 6Z�w  ��S  6]�  ��3 6^�h  ��J 6_wS  ��Q 6c?   jQ 6d?  ?A 6f?  N 6h0X  { 6k�w  $�m 6l�w  (� 6m�w  ,� 6n�w  0( 6p?  4�  6su�  8��  6u�  �  . 5Z.�}  "�}  "|  h 5[ �}  �=  7v4~  ?1  7xo   �N  7y@   ~S 7{�w  � 7|�w  �� 7}�w   �J 5[.E~  "4~  �}  �: H5f�~  +pt0 5h�   +pt1 5i�  +pt2 5j�   +pt3 5k�  0+op 5mb  @ �7 5oK~  .D 5o�~  "�~  K~  LA 5s,�~  �+ 85|1  30 5~C   �, 5C  I= 5�C  G" 5�C  y( 5�b   R�  5�|  (� 5��z  0 �0 5t-=  �~  �  5xO  U  $e  1  �~   �4 @8��  �� 8��~   �3 8��h  8 *5 8�e  � 8��  e  h�v  9!	�I     h�v  9+	@I     h�v  9A	 I     a�v  9I	�I     a�v  9X	�I     d:�  9gBo  	�I     dc�  9q'p  	�I     a�v  9{	@I     ds�  9�En  	 I     b�6 9�yq  	�I     d  9�&  	`I     \  ��   L    "��  bF5 +��  	�I     atw  �	�I     a�w  �	 I     n�w  	�I     n�w  b	`I     V�8 Z   ,��  �H  � � �J �4 �R F U6 �M ': 	�. 
�" � �6 �I s) � 3 �C �E �  ( �8 	1 �E F* |Q cQ  �D L�  �  ʁ   L    "��  A Pʁ  "�  :!�  �  �  ��  �   �  :$�  �  �  ,�  BN  wS  �  �   �  :*8�  >�  h  R�  �V  �   ��  :.^�  d�  ?  ��  %Q  �  �  �   ��  :4��  ��  �  ��  %Q  �  �  �   9�  (::�  i�  :<$ہ   (�  :=$��  Z�  :>$,�  ��  :?$R�  ��  :@$��    "��  R�  ::�  �  OZ   7VK�  �Q b �  �Q G& �I   OS   7hl�  4-   py�J ���| �P 7���  6/ 7��w   �8 7��w  { 7��w  �J 7��w  M 7�?   �= 7�l�  LGH P7�e�  �� 7��w   .� 7�o  �C 7�?  �! 7�?  	�N 7��w  tS 7��w  � 7��w  {' 7��w  SI 7��}    7��}  @Xc  7�e�  ` ��  u�   L    � 7�ǃ  "u�  G# 7���  "��  ǃ  OZ   ;.��  ` ` " 0;F�  � ;H�z   &K ;J?  N ;K?  	� ;M@   z: ;N@   � ;P�    h  �   L    kG ;R��  c$ ;R;�  "*�  ��  nO ;U��  �6 ;W?   +min ;Y�w  +max ;Z�w  �- ;\�w  HK ;]�w   ; ;_A�  "��  !< ;_��  A�  OZ   ;yȅ  �4 � L: (;~L�  v�  ;��}   l ;�L�  �A ;�{  &K ;�?  �Q ;�?  �� ;��w  .� ;�o   _E ;�o  $c� ;�R�  ( ȅ  �}  b�   L   � �C ;�ȅ  �; ;�L�  "n�  L�D �I;�g�  v�  ;��}   ;2 ;�1  ^7 ;�b�  H ;�b�  8l ;�b�  `0�A ;�{  �H# ;��w  �H�9 ;��w  �H* ;��w  �Hl4 ;��  �HvD ;�?  �H� ;�?  �H?E ;�?  �HN< ;�?  �H ;�{  �H� ;�{  �H�M ;�*�   IV( ;��w  I�  ;�g�  IY@  ;��w  I�K  ;��w  Ic9 ;��w   I1 ;��w  $IjJ ;��  (IR ;��  8I� ;��  HI� ;��  XI�S ;��  hI�$ ;�?  xI-3 ;�b  |I�, ;��  �I�9 ;��  �IO3 ;��  �I�, ;��  �I ��  �H ;��  �' ;���  �  ��  <'��  ��  �  ��  �  ��   Z=  jd  <+È  Ɉ  �  ݈  �  ݈   �  j>  �g  </��  ��  �  �  �  �  �&   �{  <6 �  &�  �  ?�  �  �  �    l  <=��  �n  <B �  �x  <Gc�  i�  �  }�  �  �   1j  <K��  �}  <P��  ��  �  ��  �  �2  ��  ��  ݈   �  ��  <W4  �b  P<Z`�  h  <\��   �v  <]�  ��  <^?�  ��  <_}�  .�  <`��   �  <a�  (V�  <bK�  0��  <cW�  88�  <f��  @��  <gĉ  H "Љ  h�  <Zq�  `�  �4 :��  +j <@    � =�w   v" ?w�  ." ?��  w�  m=1�  Qr =3�w  Qf =4Lz  Qi =5b    =/	�  +u =6��   � =8}z   p =:�  + (==d�  R�  =?|   � =@�z  B� =Ad�  +top =Bd�  �m  =C�    	�  �/ =Ev�  �  OZ   �K�  IO  R1 �G �. �6 q 8& 5 L �- 	�6 
�7 �L J( �B : � ; �9 R& � �8 � � �G Z4 - �" _1 , P! �@  OZ   �D�  ~9  r/ W0 iE �@ J #L �B Q$ YN 	�R 
$; S 88 �H ]L �P �7 �, [O � � �N � ? g: �8  �L �9 nN �< �B  �$ !E "�: #S@ $� %�6 & /� B`�  4� Bj�   5wJ �ύ  4� �j�  .� �b  �� �b  k� �	�  12 �b  8idx �b  8i �b  1tmp *	�    5�' ���  4� �j�  :num �o   5}C �'�  4� �!j�  :idx �!o  :val �!�w   21 ��w  Q�  4� �!j�  :idx �!o   2�Q ��w  o�  4� �"j�   2� �b  ��  4� � j�   5� {��  4� {#j�  :val |#�w   5< kَ  4� k!j�  :val l!b   2�* do  ��  4� dj�   5�N T�  4� Tj�  1R�  X|    22: 5j�  k�  R�  5|  :e 6�z  �m  7�  � 9�  4� ;j�   20 j?  ��  :buf jv{   2�; Pb  ��  :buf P!v{   ,5 � �E     ;/      ���  v�  �1�}  �� `� 7buf �1v{  c� Q� ;2 �11  6� *� �< �1  Ӯ Ǯ �* �1?  h� d� �  �1�w  �� �� �  �1�w  ȯ Ư ��  �1��  �� � 	dN ��  |� j� 	�3 ��h  P� <� 	� ��z  J� 8� 	R�  �|  � � 	* ��w  �� {� 	�P ��w  !� � 	� ��  ô �� 	mP �?  /� 	� 	�/ �?  � Ը !L[ ���  ���~	� ��  x� B� 	V( ��w  μ Ƽ 	u. �j�  �� .� 	�m  ��  �� �� op1 �h  �� ?� !�^ ���  �к~!'7 ���  ���~	�!  U  �� q� !dA {  ���~! ?  ���~	ٶ v{  @� &� 	� b  �� _� ! {  �й~!� {  ���~!�M �  ���~!�N m�  ���~<\� � F     T% I#> F     *       Β  	/� ��  s� o� F F     o�  Uu   %�� ]�  	��  ��  �� �� *�  �F      0�  �  8�  2� *� 8�  2� *� R�  �� �� E�  � � 0� _�  �� �� l�  T� R� y�  }� w� ��  �� �� ��  	� � َ  �F      `� ���  �  O� ?� �  O� ?�  M��  �� �  ��  �� �� ��  c� ]� �e F       � �4�  f �� �� f �� �� � f  � �� #f C� ?�   ��  >F       � �Ȕ  �  �  �� ~� �  �� �� ;َ  BF       BF            ���  �  � � �  � �  B�F     Uu 3�  {   �F     '�  �  Uu T{  F     '�  Uu Tz  �F     ύ  Uu T} s    \��E     4�  Us  \��E     H�  Us  ��E     o�  Uu   # F     }       +�  idx ]o  ^� V� 	.� ^o  �� �� َ  $F       $F            ^ޕ  �  �� �� �  �� ��  JF     '�  ��  Uu Tv  \F     '�  �  Tv �F     Q�  U���~  % � 9�  idx to  $� � 	.� uo  �� �� isX w?  �� �� %�� Ė  v ~�w  �� �� �F     Q�  ��  U���~ �F     '�  Uu T|   َ  �F       P� u��  �  $� � �  $� �  @D�  �F      �F            �R�  �� �� R�  �� ��   %Ц w�  	.� �o  �� �� idx �o  � 	� #�F     �       ��  x1 ��w  �� �� y1 ��w  �� �� x2 � �w  (� &� y2 �$�w  M� K� x3 �(�w  t� p� y3 �,�w  �� �� �F     '�  �  Uu Tvz �F     '�  /�  Tv{ �F     '�  G�  Tv| �F     '�  _�  Tv} �F     '�  w�  Tv~ �F     '�  ��  Tv F     �  U���~R~ Y|   َ  hF      � ��  �  �� �� �  �� ��  D�  �F      �F            �*�  R�  5� 3� R�  5� 3�  TF     '�  H�  Uu Tv  cF     '�  `�  Tv �F     Q�  U���~  %��  �  	�M �b  ^� X� #�F            ͙  val ��  �� �� �F     7�  � RF        � �G�  � �� �� � @� >�  � � i� g� K5 dF       P� �N �� �� B �� ��    �  �F      �� ��  A�  �� �� 4�  ,� *� '�  Y� O� �� N�  �� ��   ��  @	F      @	F     B       ��  ��  7� 5� ��  ]� [� ��  �� �� &@	F     B       ��  �� ��   �F     o�  Uu   %P� ٵ  op2 $h  #<F     	       c�  !K8 -%%�  	@I      #�F     )       ̛  !K8 E%%�  	0I     �F     ��  U T��~Q� R���~X	0I     Y0  %@� �  !K8 ]%%�  	 I     eF     ��  U T��~Q� R���~  #jF            D�  !K8 u%%�  	I      %0� V�  v0 �%�w  �� �� v1 �)�w  7� 1� v2 �-�w  �� �� isV � ?  ��  F       p� �+�  �  �� �� �  � � �  Y� U� ;َ  F       F            ��  �  �� �� �  �� ��  BF     3�  2  ��  GF       �� ���  �  � � �  V� R� �  �� �� ;َ  KF       KF            ���  �  �� �� �  �� ��  B	F     3�  4  �F     ]p ڝ  3�  s  �F     '�  ��  Uu T0 �F     '�  �  T2 F     '�  %�  T4 F     '�  <�  T1 GF     '�  Uu T3  #6 F     %       Ϟ  	}0  �#�w  � � 	i/  �#�w  @� <� > F     Q�  ��  Uu  E F     Q�  [ F     ��  Tt   # F            H�  	}0  �#�w  x� v� 	i/  �#�w  �� ��  F     Q�  &�  Uu  " F     Q�  1 F     ��  Tt   #�F            ��  arg �#�w  �� ��  F     Q�  ��  Uu   F     ��  Tt �  %� ��  		*   �  � �� 	,&  b  �� �� 	�J -b  �� �� 	R0   �  C� ;� 	�  .�  �� �� 	�  �3  � 
� !�R $j{  �л~!�$ $�w  ���~	�: b  a� Y� 	�A b  �� �� ady �  /� !� adx �  � � asb �  �� �� %@� S�  	)�  c'�  � � 	��  d'�  E� A� 	�.  e'  �� ~� 9F     C� �  U���~T2 �F     O� 6�  Us  �F     O� U
w � $ &  \�  F       �� �š  j�  �� �� w�  J� @� w�  J� @� �� ��  �� �� 6��  ��~B=F     T��~   \�  �F       �� �7�  j�  �  � w�  *� (� w�  *� (� �� ��  U� Q� 6��  ��~BF     T��~   �F     o�  O�  Uu  �F     o�  �F     Q�  �F     Q�  �F     Q�  VF     C" ��  U} Tv  cF     C" ��  U} T|  �F     \� �F     -r ��  Tv Q�л~3��  }  �F     ��  0�  U~ T�л~Q���~R�ȷ~X1Y0 �F     -r [�  T| Q�л~3��  ���~ �F     ��  U~ T�л~Q���~R�ȷ~X1Y	s ��~�  #�F     �       0�  	�! �"�w  �� �� 	�! �)�w  �� �� 	<0 �"�_  �� �� �F     Q�  �  Uu  F     Q�  F     Q�  F     Q�   #�F            o�  arg �#�w  � � �F     Q�  Uu   #wF            Ԥ  	� #�w  ?� =� 	/; #�w  f� b� F     Q�  Ƥ  Uu  �F     Q�   #.F            9�  	JB #�w  �� �� 	�! #�w  �� �� 6F     Q�  +�  Uu  =F     Q�   %� ��  	�> &#�w  �� �� 	��  '#�w  =� 5� ZF     Q�  eF     Q�  ��  Uu  pF     h� �F     o�  �F     o�   %� �  arg A#�w  �� �� F     Q�  Uu   #�F            e�  	}0  Q#�w  �� �� 	i/  R#�w  �� �� �F     Q�  C�  Uu  �F     Q�  �F     ��  Tt   %� I�  	0G cb  O� 5� 	�O db  t� V� 	.� eo  �� �� 	P+ fo  �� �� #F     �       ��  idx �!�  �� �� 	8G �!�  �� �� . SF      SF            � l�  �. � � �. @� >� fF     �t U���~#T13�. ���~  �F     �  U���~  %�� a�  	�  #G(  h� d� 	2]  #�  �� �� nn /�  �� �� mm 3�  4� *� 	� #o  �� �� 	�D #o  t� j� %0� C�  tmp ?&�w  �� �� �e nF       `� D#|�  f 3� 1� f X� V� `� f � {� #f �� ��   ��  �F      �� J�  �  �  � �� �  =� 7� ;َ  �F       �F            ���  �  �� �� �  �� ��  BBF     Uu 3�  z   MF     '�  .�  Uu Tz  nF     '�  Uu   �F     ύ  Uu Tx y   #�F     `       ��  idx Y#�  �� �� 	�  Z#G(  � � �F     o�  �F     u�  #uF            �  	� r'�w  6� 4� 	/; s'�w  ]� Y� �F     Q�  �F     Q�   #VF            o�  	JB �'�w  �� �� 	�! �'�w  �� �� eF     Q�  lF     Q�   #&F     0       7�  	6 �'�w  �� �� 	� �'�w  � � �e =F      =F            ��  f >� <� f c� a� &=F            f �� �� #f �� ��   5F     Q�  =F     Q�   #�F     .       ��  	�> �'�w  
� � 	��  �'�w  /� -� F     Q�  F     Q�  F     h�  #wF     P       ��  idx �#b  T� R� 	�  �#G(  y� w� �F     o�  �F     Q�   #*F     M       E�  idx �#b  �� �� 	�  �#G(  �� �� LF     o�   #�F     0       �  	}0  '�w  �� �� 	i/  '�w  � � 	�? '�w  W� S� 	]# '�w  �� �� 	F     Q�  F     Q�  F     Q�   F     Q�   %p� =�  r '�w  �� �� �) �F      �� ((�  * � �  �F     ��  Uu   #�F     <       z�  i 2!�  n� h� 2F     Q�  Uu   َ  qF       @� y��  �  �� �� �  �� ��  D�  	F      	F     	       �  R�    R�     . 3F      3F            �]�  �. ; 9 �. c a FF     �t U���~#T63�. ���~   sF      �� ���   � �  ��  �F      � ���  ��  � � ��  � �   �F      �F            ��      bF     o�  	�  Uu  jF     o�  �F     ��  4�  Uu Tt  F     ��  Tt   #�F     %       ��  val v#�w  E C idx w#b  j h �F     o�  ��  Uu  �F     Q�   #�F            �  idx �b  � � �F     o�  Uu   #mF     ,       ��  	}0  �#�w  � � 	i/  �#�w  � � 	�? �#�w    	]# �#�w  O K uF     Q�  n�  Uu  }F     Q�  �F     Q�  �F     Q�   #5F     8       �  r �#�w  � � W�) GF      Т �* � �   #wF     )       ��  	6 �#�w  ( & 	� �#�w  M K �e �F      �F            ���  f r p f � � &�F            f � � #f  �   F     Q�  ��  Uu  �F     Q�   #�F     F       P�  arg �#�w  D < #�F     /       ;�  	�� �!�  � � 	�N �!�  � � F     h� Uv Ts   �F     Q�  Uu   #�F            ��  arg �#�w   � �F     Q�  ��  Uu  �F     ��  Tt   #�F            �  	}0  �#�w  = 9 	i/  �#�w  w s �F     Q�  ��  Uu  �F     Q�  �F     ��   %p� ֳ  idx 
	b  � � 	�  	o  � � %�� �  	�8 	!o  x t |F     '�  Uu   َ  KF      KF            	��  �  � � �  � �  KF     o�  Uu   #h F     �       j�  idx *	b  	 � 	.� +	b  � � `�  z F      z F     �       3	D�  ��  � � y�  �	 }	 m�  �	 �	 &z F     �       ��  �	 �	 ��  �
 �
 ��    ��   � ;َ  � F       � F            ��  �  d ` �  d `  M��  @� �  ��  � �  @5 2!F       2!F     )       N � � B      p F     o�  \�  Uu  x F     o�   ��  `F      � $#��  ��  zF     Dj Ur   �F     Q�  ��  Uu  �F     Q�  �F     Q�  Uu   #�	F     �       >�  	�! n	�w  A ? 	<0 o	�_  f d �	F     Q�  0�  Uu  �	F     Q�   #F     7      c�  	�: �	b  � � 	�A �	b  � � !�R �	j{  �л~!�$ �	�w  ��~		*  �	�     6�  �F      �� �		�  D�  f d D�  f d Q�  � � B�F     Ts   6�  
F      
F     "       �	h�  D�  � � D�  � � Q�  � � B,F     Ts   F     o�  ��  U  %F     o�  ,F     Q�  8F     Q�  TF     _�  ʷ  U���~Q�л~ �F     ��  �  U~ T�л~Q���~R�ȷ~X1 �F     _�  *�  U���~Tv Q�л~ 
F     ��  U~ T�л~Q���~R�ȷ~X1Y0  %�� |�  !�4 1
b�  �л~!7 2
�  ��~5�  ��E      � 5
�  w�    j�  4 . ]�  � � P�  � � C�      ��  !�E      �� :
#�  ��  Y W ��  �   .�E     ��  C�  U��~T~  Y�E     j�  U�л~T�й~Q���~R��~X0Y0  %�� ƻ  	.� {
o  � � idx |
o  � � #p�E     �       ��  x1 �
�w  � � y1 �
�w  � � x2 �
 �w  � � y2 �
$�w     x3 �
(�w  E C y3 �
,�w  j h z�E     '�  Z�  Uu Ts  ��E     '�  r�  Ts ��E     '�  ��  Ts ��E     '�  ��  Ts ��E     '�  ��  Ts ��E     '�  Һ  Ts ��E     �  U���~R~ Y}   َ  ��E      ��E            {
7�  �  � � �  � �  D�  3F      3F            �
y�  R�  � � R�  � �  '�E     '�  ��  Uu T}  7�E     '�  ��  T} [�E     Q�  U���~  #�E     �       ��  	.� �
o  � � 	�� �
o    idx �
o  } q %p� B�  x1 �
�w    y1 �
�w  Y U x2 �
 �w  � � y2 �
$�w  � � x3 �
(�w  � � y3 �
,�w    � U�E     '�  ��  Uu Tv  g�E     '�  Ѽ  Ty  r�E     '�  �  Tv ��E     '�  �  Tv ��E     �  '�  U���~R| Y|  ��E     '�  Uu Tv   @َ  �E       �E            �
%�  % # �  % #   % � x�  	.� �
o  N H 	�� �
o  � � idx �
o  � � %`� ��  x1 �
�w  � � y1 �
�w  � � x2 �
 �w  � � y2 �
$�w  � � x3 �
(�w   � y3 �
,�w  = 7 Z�E     '�  h�  Uu Tv  z�E     '�  ��  Uu Tv  ��E     '�  ��  Ty  ��E     '�  ��  Tv ��E     '�  ξ  Tv ��E     �  U���~Q~ X| Y}   َ  �E       �E            �
%9�  �  � � �  � �  @D�  Q
F      Q
F             �
R�  � � R�  � �   %�� ��  	.�  o   � 	��  o  T P idx o  � � 	�I ?  ) % %0� u�  x1 �w  g _ x2 �w  � � x3 �w  ` Z y1 #�w  � � y2 '�w    y3 +�w  � � &F     '�  t�  Uu Tz  ?F     '�  ��  Tv  OF     '�  ��  Tx  ZF     '�  ��  Ts  �F     �  ��  U���~Q} Yv  �F     '�   �  Uu Tz  �F     '�  �  Tv  F     '�  0�  Tx  F     '�  H�  Ts  )F     '�  `�  T|  p
F     '�  T|   D�  6�E      � B��  R�  � � R�  � �  @َ  �F       �F             %�  . $ �  . $   %�� ��  v Hb  � � 	eG Jb  � � 	E Kb     ��  ��E      �� Je�  ��  ��E     Dj Ur   ��  ��E      � K��  ��  	F     Dj Uu   �E     ��  Uu Tt   #�	F            ��  v \b  G C �	F     ��  Uu Tt   %@� d�  v ib  � � ��  F      p� oI�  ��  (F     Dj Ut   4F     ��  Uu Tt   %Ч ��  v zb   
 ��  �
F       � ���  ��  �F     Dj Uu   �
F     ��  Uu Tt   %0� G�  v ��w  � � 	eG �U  � � 	E �U  � � 	=F �U  *  &  	�E �U  b  `  ��  �F      p� �+u�  ��  <F     Dj Uu   ��  �F      �� �+��  ��  $F     Dj Us   ��  F      Ш �+��  ��  F     Dj Us   ��  ,F       � �+�  ��  �F     Dj Uu   �F     ��  2�  Uu Tt  �F     ��  Uu   ��  �E      �� -n�  \�  �  �  O�  ! ! B�  c! a! 5�  �! �! (�  �! �! �  6" 0" �  �" �" �  �" �" ��  �" �" ��  # # 5�  ��E      0� QA�  w�  e# c# j�  �# �# ]�  �# �# P�  �# �# C�  �# �#  � @�E      �� L��  � �# �# � $$ "$ � I$ G$ � n$ l$  5�  ��E      �� V��  w�  �$ �$ j�  �$ �$ ]�  �$ �$ P�  
% % C�  /% -%  5�  �E      � [K�  w�  X% V% j�  }% {% ]�  �% �% P�  �% �% C�  �% �%  �E     �� U���~T0Q
�I  ��  ��E      `� � ��  ��   � ��E      Ж ��  � & & � A& ?& � f& d& � �& �&  � 5�E       � /�  � �& �& � �& �& � ' ' � 9' 7'  � ��E      0�  �  � b' `' � �' �' � �' �' � �' �'  ��  ��E      `� &��  ��  �' �' ��   ( (  ��  ��E      �� L��  �  [( G(  ��  ��E       ��E            V �  ��  C) A)  �  �E      �� X��  F�  j) f) <�  �) �) 0�  �) �) �� 6R�  �л~^�  A* 5* $�E     �� ��  U| T(Q�л~ [�E     �� ��  U| T8Q0R} X0Y�л~ �
F     �� U|    & ��E      0� d3�  ? �* �* 3 	+ + �F     L U���~TA  D�  ��E      ��E            �u�  R�  s+ q+ R�  s+ q+  ��  ��E      ��E            ���  ��   5  F      p� ���  N �+ �+ B �+ �+  ��  +�E      �� �F�  ��  , , Wy +�E      �� �� ;, 9, �� � c, a, d�E     ��    y ��E      �� ���  � �, �, �� � �, �, ��E     ��   y ��E       � ���  � �, �,  � � - �, ��E     ��   y 
�E      `� �!�  � &- $- `� � O- M- 3�E     ��   ��  ?�E      ?�E     '       ���  �  t- r- =�  D�E     "       �  �- �- S�E     �� ��  Us  f�E     �� Us T    D�  ��E      ��E            ���  R�  �- �- R�  �- �-  َ  �E      �E            i
/�  �  �- �- �  �- �-  َ  ��E      ��E            P
q�  �  !. . �  !. .  َ  �E       �E            
��  �  n. j. �  n. j.   � F      �� �	��   �. �.  ��  � F      �� �	�  ��  �. �. ��  / /   � F      � F            �	G�   9/ 7/  � 0F      � �	��  � b/ `/ � �/ �/ � 0� C5 8F      8F            �N �/ �/ B �/ �/    َ  �F      �F            K�  �  0 �/ �  0 �/  � IF       IF     T       ��  � =0 70 � �0 �0 &IF     T       � �0 �0 K5 [F       �� �N �0 �0 B 	1 1    َ  �F      0� �	��  �  21 ,1 �  21 ,1  �  �F      `� �		�  �  �1 {1 �F     �r U���~  َ  �F       �F            �	.P�  �  �1 �1 �  �1 �1  Q�E     Q�  h�  Uu  u�E     ��  ��  U���~ ��E     Q�  ��  Uu  ��E     Q�  g�E     ]p ��  U| T��~#�Q R���~X�Y���~3�  ��~ � F     ��  �  U���~ �F     Q�  %�  Uu  WF     yg H�  Uu 3- ���~ �F     '�  e�  Uu T0 F     '�  ��  Uu T0 &F     '�  ��  Uu T0 ,F     ��  ��  U���~Ts  �F     '�  Uu T0  �w  �w  ��   L    �w  ��   L    �w  �   L    @   K  %�   L    "�  /�* ���  �  �!1Q  u. �!j�  ��  �!o  � �o  2�  �o  i �o  j �o  ��  �o  1��  ���  sum ��w    x  ,N; O��E     �      ���  u. Oj�  2 2 �  P��  2 w2 �  Q��  �2 �2 �N Ry�  M3 E3 K8 S��  �3 �3 � T?  4 �3 !�M V��  ��idx Wo  �4 �4 	�< X?  B5 :5 top Yb  �5 �5 i Yb  n6 j6 j Yb  �6 �6 %`� �  	)N o?  �6 �6 	�2 r�w  M7 I7 ~�E     '�  Uu   D�  ��E      ��E            �\�  R�  �7 �7 R�  �7 �7  !�E     '�  z�  Uu T~ ��E     �  ��  U��~ ��E     �  ��  U��~R X~ Y��~� a�E     '�  ��  Uu Ty z�E     '�  Uu   K  �w  �   L    /�J ��  v�   �}  u.  j�  �/  {  ��   ��    ��  3  �w  i  o  .� !o  G "?  _  %�w  T\� H1�? 5��    ?  5�I ���  +�  �&*�  � �&@   8i �@   � �o   5�1 �1�  +�  �$*�  ٶ �$v{  � �$@   8i �@    2 l@   [�  +�  l)*�  � m)@    2�, eu2  y�  +�  e**�   5�K Z��  +�  Z&*�  :val [&?   2	N S?  ��  +�  S+6�   2K L?  ��  +�  L-6�   5^ B�  +�  B$*�  � C$�z   /5$ s�  q' s/y�   ,� p�E     6      �Q�  q' )y�  8 �7 7x1 )�w  n8 d8 7y1 )�w  �8 �8 7x2 )�w  O9 G9 7y2 )�w  �9 �9 7x3 )�w  :  : cy3 )�w  � !�$ !�w  ��!�L !�w  ��!�$ !$�w  ��!:' !.�w  ��XP0 "�  ��P1 "�  v: j: P2 "�  ; ; P3 "�  z; r; E�  ��E       �� 7��  w�  �; �; l�  < < a�  9< 7< V�  ^< \<  ��E     /�  ��  Uu R} X Yy  ��E     /�   �  T| Qv R~ X� �Yy  �E     ��  e�E     ]�  7�  Us TsQ��Y0 ��E     j�  UsY0  ,�, ���E     �      ���  q' �(y�  �< �< 7x �(�w  = �< 7y �(�w  l= d= !Y@  ��w  ��!�K  ��w  ��XP0 ��  ��P1 ��  �= �= 	9 �?  *> (> 5�E     /�  0�  Us R| Xv Yy  �E     j�  M�  UsY0 :�E     ]�  w�  Us TsQ��Y0 E�E     ��   ,%0 ���E     �       �/�  q' �(y�  V> N> 7x �(�w  �> �> 7y �(�w  ?? 1? �  ��E      �� ��  �  �? �? %�E     �r  	�E     j�  Uv Y0  ,/L �`�E     �      ���  9q' �/y�  U7x1 �/�w  @ @ 7y1 �/�w  �@ ~@ 7x2 �/�w  �@ �@ 7y2 �/�w  ZA RA cx �/��  Y7y  /��  �A �A dx �w  	B �A dy �w  �B �B E�  ��E       @x =�  w�  �C �C l�  �C �C a�  �C �C V�   �e �E      �E            .��  f D D f BD @D &�E            f jD hD #f �D �D   �e ��E      px G�  f �D �D f �D �D px f E E #f OE KE   �e �E      �E            Io�  f �E �E f �E �E &�E            f �E �E #f !F F   �e a�E      a�E            c��  f ^F \F f �F �F &a�E            f �F �F #f �F �F   �e  �E      �x |.�  f �F �F zf Ι}�x f 'G #G #f jG fG   @�e y�E      y�E            ~f �G �G f �G �G &y�E            f �G �G #f >H :H    ,R> �0�E     �       �]�  q' �*y�  �H yH �S �*�  �H �H !G  ��~  ��w�E     �g 4�  Us TsQ��R��X| Yv 3��  �� \��E     H�  Tw  ��E     ��  Us   o�F )P�E     `      ���  q' ).y�  0I $I �' *.n�  �I �I B> +.   J �I �Q ,.�  �J �J =9 -.?  �J �J !G  /�~  ��~	�$ 1  �J �J 	�4 2  xK pK 	 4�  �K �K 	E6 5?  M M ��  ��E      �� MB�  ��  �M �M ��  �M �M ��  �M �M ��  �M �M ��  )N #N ��  )N #N �  xN rN �  xN rN �  �N �N �  �N �N �  %O O �  %O O �� 0+�  06�  0A�  L�  �O }O Y�  �O �O �e ��E      Љ ���  f �O �O f P P Љ f DP @P #f �P �P   �e �E      0� ���  f �P �P f 0� f �P �P #f .Q *Q   �e ��E      �� �)�  f kQ iQ f �Q �Q �� f �Q �Q #f R �Q   �e ��E       � �o�  f f  � f BR >R #f �R �R   �e �E       `� ���  f �R �R f S S `� f DS >S #f �S �S   �e O�E      O�E            �3�  f �S �S f T T &O�E            f ?T 9T #f �T �T   �E     h�   ��E     �g ~�  Us Ts�0Q��R��Yy 3��  �� .�E     �g ��  Us T~ Q��R��Yy 3��  �� Q�E     �g ��  Us T~ Q��R��Yy 3��  �� t�E     �g /�  Us T~ Q��R��Yy 3��  �� \��E     D�  T��~ ��E     �g ��  Us T��~Q��R��Yy 3��  �� %�E     �g ��  Us T��~3��  �� g�E     �g Us Ts�03��  ��  ' �?  e�  q' �8y�  )u1 �8  )u2 �8  )v1 �8  )v2 �8   �8  u ��  v ��  w ��  P4  ��w  s ��w   /�/ ���  q' �+y�  �' �+n�  )ppt �+  )x �+�w  )y �+�w  pt ��   /�= ���  q' �*y�   /�; ;j�  q' ;-y�  v�  <-�}  ;2 =-1  * >-�w   @-{  � A-{  �M B-*�  V( C-�w  �  D-��  l4 E-   ,# (`�E     �	      ���  �' ($n�  �T �T  )${  eU QU � *${  RV >V �M +$*�  4W ,W �= ,$�w  �W �W �4 -$?  X �W 	* /u2  ~X fX 	v�  1�}  �Y �Y !(R 2�  ��	� 4@   Z Z i 4@   kZ QZ 	�' 5h  �[ y[ #��E     @       �  !��  j�}  ��~w�  ��E      �� m��  ��  �\ �\  ��E     ��  ��  Us T�Q��~ ��E     ��  Us T��~Q�  %p� i�  !� ��}  ��~!` �&�}  ��~��  ��E       ��E             �w�  ��  �\ �\  ��  ��E       ��E             ���  ��  �] y]  [ `�E      �� ���  � ^ �] z n^ h^ m �^ �^ �� � $_ _ � �_ �_ � ` ` � �` �` � ka _a ��  ��E      �� �]�  ��  �a �a  ��  ��E      0� *��  �  Jb Fb  ��  O�E      O�E            >	��  ��  �b �b  W��  ��E      p� 8	��  �b �b    x�E     ��  �  Uu T��~Qv R X��~� ��E     ��  F�  Uu T��~R X��~� ��E     ��  Us T��~Q��~  #@�E     H       !�  !c� ��}  ��~!MV  ��}  ��~w�  @�E      �� �	��  ��  �b �b  w�  v�E      v�E     
       �	��  ��  -c +c  ��E     ��  Us T��~Q��~  #t�E     g       ��  !� ��}  ��~!` �(�}  ��~��E     ��  ��  Uu T��~Qv R X��~� ��E     ��  ��  Uu T��~R X��~� ��E     ��  Us T��~Q��~  %0� ��  	�? #��  Tc Pc � G�E       G�E     2       $��  � �c �c � �c �c &G�E     2       � d �c K5 Q�E       `� �N &d $d B Md Kd    @��  y�E      y�E             (�  td pd   [�  ��E      ��E             ^��  l�  �d �d  ��  g�E       �� I��  ��  �d �d ��  Ie Ee �� ��  �e �e ��  f f K1�  g�E      �� �
N�  �f �f B�  g g =1�  ��E            N�  Pg Jg B�  �g �g C5 ��E       ��E            rN �g �g B �g �g      ��  �E       � ��  ��  "h h  � ��  �h ~h ��  ~i zi  �E      �� �Z�   �i �i  M��  Ѕ  �  ��  )j j ;�  *�E       *�E             ���  L�  k k  ��  >�E     	 >�E             ���  ��  �k �k  M��  � ��  ��  �l �l ��  =m 1m ��  �m �m ��  �n �n �  uo io �  �p �p �  �q �q (�  �s s 5�   t �s B�  )t #t O�  �t {t \�  �t �t ��  ��E       `� ��  ��  Iu Eu  =i�  A�E     /       6j�  ��~[�E     � T��~   [�E     h� ��E     h�  =z�  ��E     �       0{�  � ��E       �� <��  � �u �u � �u �u �� 0� C5 ��E       ��E             �N �u �u B  v �u    @;�  �E      �E             ML�      y�  3�E      �� 6��  ��  %v #v ��  Kv Iv  ��  =�E       =�E             /�  ��  vv pv  ��  ��E       �� =e�  ��  �v �v ��   w �v  !�E     j�  Qv R��Y1  ,@ Z��E     �      ���  �' Z(n�  Ew 9w � [(4~  �w �w ` \(4~  tx ^x 	tE ^o  ky cy i� a?  	nA b4~  �y �y 	�% c4~  z z #��E     X       ��  	I> ��w  { 	{ 	�L ��w  I{ C{ �e КE      �w ���  f <| :| f b| `| �w f �| �| #f �| �|   КE     ��   %�w �  	�( �o  } } 	�+ �o  } }} 	.� �o  �} �}  ��  ��E       `w �F�  ��  ;~ 3~  �  ��E      ��E             �{�  .�  �~ �~  �E     ��   /�F ���  �' �)n�  i �@   j �@   ]z�  � �?  1sQ ��w  o ��w  �7 ��w  { ��w  �( ��w  AD ��w  � ��w  .K ��w  ��  ��w  P ��w  �) ��w  >I �?  1A? ��     1�N ;��    -9O N�w  p�E           ���  9�' N!n�  U~S O!�w  ? / % w ��  i Yo  � � �e �E      0w w3�  f f 0w f ۀ ׀ #f � �   @�e P�E      P�E            lf [� Y� f �� � &P�E            0f 0#f    @�e 0�E      0�E            Tf Ɓ ā f � � &0�E            f -� '� #f �� �    /� /�  �' /"n�   '�' (?  5�  �' (+z�   /�( ��  �' #n�  v�  #�}  �4 #n�  �A #{  �� #�w   /�  ��  �� 4~   '�+ ?  ��  �� )@~   '�6  ?  ��  ��  &@~   2�* �?  ��  �� �&@~   21N �?  �  �� �#@~   23 �?  ;�  �� �'@~   2� �?  Y�  �� �$@~   2� �?  w�  �� �%@~   5KL ���  �� � 4~   Y�Q Z��E     x      �?�  >�� Z&4~  U.�/ [&{  �� ؂ >�- \&@   Q.v�  ]&�}  L� B� .�= ^&�w  σ �� >�� _&�w  Y>u� `&?  � (��  b�w  �� m� (�+ c?�  ؅ Ѕ N� ӲE      �} h(��  � :� 4� � �� �� �} � �� �� K5 ݲE       �} �N � � B $�  �    N��  `�E      0~ ���  ��  \� Z�  K�e ��E      p~ �f �� � f �� �� p~ f ͇ ɇ #f � �    ��  2�> Eb  ��  :x1 E&�w  :y1 F&�w  :x2 G&�w  :y2 H&�w   /19 
m��  �S  
m#�  �3 
o�h   /P 
_��  �S  
_#�  �3 
a�h   '� 
U�w  ��  �3 
U&�h   '4= 
K�w  �  �3 
K&�h   '�0 
b  \�  �3 
+�h  �M 
+b  )buf 
+v{  idx 
o   /). 
���  �3 
�)�h  )buf 
 )v{  �  
�3  �U  
�	   ' 
��  6�  �3 
�(�h  �^ 
�(�  )buf 
�(v{  ��  
��	  � 
��  �  
��3  �6  
��2  inc 
�#�!  1$ 
�u2  ��  
��    /{G 
�_�  �3 
�'�h  )buf 
�'v{   -�P 
��  �E     �       ���  �3 
�&�h  S� K� � 
�&b  �� �� 7buf 
�&v{  &� � gid 
�b  �� �� !ٶ 
�u2  �PXlen 
��  �X	� 
��  �� �� b W�E       �} 
��  � � � t ;� 7� �} � w� q� � Ŋ �� � �� �� Bv�E     U�T   B)�E     Qw R�X  'y+ 
xb  ��  �3 
x,�h  �M 
y,b  )buf 
z,v{  idx 
|o   '�H 
mb  ��  �3 
m&�h   /4 
`3�  �3 
`)�h  .� 
a)�  �U  
b)3�   �_  /�3 
So�  �3 
S$�h  .� 
T$�  �U  
U$3�   / 
F��  �3 
F#�h  .� 
G#�  �U  
H#3�   /N" 
9��  �3 
9#�h  .� 
:#�  �U  
;#3�   /* 
%�  �3 
%$�h  �N 
&$��  tS 
'$��  � 
($��   '�3 
�w  >�  �3 
�h   '�B 
�w  ^�  �3 
�h   'C+ 
��w  ~�  �3 
��h   'DP 
��  ��  �3 
�)�h  )len 
�*��  )vec 
�*��  �  
��C  mm 
�e�   o  'n9 
��  ��  �3 
�!�h   '�. 
�0N  �  �3 
��h   '<7 
�wS  7�  �3 
� �h   -LJ 
4�  `!F           �! �3 
4/�h  @� "� $ 
5/u2  �� � ��  
6/�  � � 	R�  
8|  G� A� !� 
9�  ��~	v�  
:�}  �� �� 	�  
<?  � � %�� � 	<0 
k�_  �� �� 	K1 
l@X  đ �� 	91 
n?  � � 	�H 
pP  y� q� 		*  
t�  � Ւ Xbuf 
uj{  ��!� 
v|  ��	� 
w�w  �� � 	�Q 
y?  ݓ ѓ 	��  
z?  |� t� A "F      �� 
� O � ؔ � � � v X� T� i �� �� \ ܖ ؖ  ! �"F      �"F             
�#N 3 ,� �  % �"F      � 
�� 6 � � 6 � � B m� g� � N �� �� �"F     h� U�C$   a #F       � 
�d � � ݘ � ͙ �� � �� �� s �� ��  � � P� B� 6� ��~6� ��~� � � ^� �)F     � ;#F      � �A � L� <� � � � � 
 Ȟ Ğ  � � " � �� . e� _� : Ϡ Š F K� ?� R ա ͡ _ =� 1� 6l ��~6y ��~M�  � � � Ѣ ͢ ~�  �,F      @�  � ��  � � ��  8� 2� ��  �� �� @� ��  ޣ ܣ ��  � � B�,F     T��~Q0R��~X0   \-F     � U~� B5-F     T~   ^�  �#F      �#F            F� p�   D� p� � 1� +� � �� �� � ֤ ̤ >�  j$F       � �> P�   � �$F       �$F     +       �	  K� I�  s� q�  �� �� � �� �� � � � � � 	� � &�$F     +       0* 06 0B FN FV F^ �$F     ~z U| Tv Rs�X0   �  �$F      P� �0 0�   �  %F       �� ��  0� .�  X� V�  }� {� � �� �� � ʦ Ȧ � � � � �� 0* 06 0B FN FV F^ [%F     ~z U| Tv Rs�X}    � �%F      �� ��	 �  � � � �� �� �� � D� B�  u� g�  /� !�  ̩ Ʃ ) � � 5 l� d� A ֪ ʪ M d� X� Y � � e ^� V� q ά Ƭ } >� 6� � �� �� � n� b� � � � N��  �%F      `� dL ��  �� �� �  կ ӯ �  �� �� ��  %� #� �%F     h� T�B$  N��  &F      �� i� ��  ��  M� K� ��  w� u�  ;o�  &F      &F            j� }�  ��  �� �� ��  ˰ ɰ  ;9�  '&F      '&F            k G�  a�  �� � T�  � �  ;��  /&F      /&F            lX �  %�  I� G� �  s� q�  ;��  7&F      7&F             �
� ��   M� �� � � �� �� � (� � � � � � D� <� � �� ��  N�e i.F       � �((	 f � � f � �  � f B� >� #f �� ��   N�e �.F      `� �%}	 f ´ �� f � � `� f %� !� #f h� d�   �'F     h� �	 U@<$ p,F     h� �	 U@<$T|  �,F     �� �	 U
��Qv  $ & �-F     h� U@<$T|    � �+F       �� �	�
  �� ��  �� ��  :� 6� � v� p� � ɶ Ŷ � � �� � �� 0* 06 0B FN FV F^ ,F     ~z U| Tv Y0   %F     h� �
 U�?$ �+F     h� �
 U��~T��~ �-F     h�  U��~T��~ 8/F     h� ( U�?$Tw  Z/F     h� U�?$    ��  8)F       8)F            � ��  =� 9� ��  =� 9� &8)F            ��  {� y� K)F     ��   ��  �)F       �)F            *0 ��  �� �� &�)F            ��  ȷ Ʒ �)F     yg ! Uu 3- v  �)F     Ȃ   m)F     ��  Us T��Q} R��~X0Y0   @� �)F       �)F            
�  � �  � � &�)F             R� N�    � +F      � 
`� � �� �� � � �� ��  �*F     �� Uw T
�Q��~  '�5 
)�  A �3 
)#�h   /! 

� �3 

)�h  �� 
)��  �� 
)��  �Q 
)��  ��  
)��   5 % 
�� �S  
�"�  R�  
�"|  � 
�"�z   Y;" 
���E     F      �{ .;2 
�11  � ٸ .G  
�1�~  y� m� (� 
��  � � (�S  
��  \� P� <0 
��_  ;W- ��E      ��E            
�� �- � � v- $�  � i- &��E            �- `� \� �E     �u Us    ;. �E      �E            
� �. �. �� �� �E     �t UsT3  N. !�E      p� 
�� H. �� �� =. �� �� 2. 9� 5� %. p� U. u� q� =b. T�E     )       c. �� �� p. Ҽ м    N. 7�E      �� 
� H. �� �� =. M� G� 2. �� �� %. �� 0U. Db. � c. � � p. � �    K. ?�E      @� 
�H. 9� 5� =. u� q� 2. �� �� %. @� 0U. Db. �� c. � � p. � �     Y� 
�@�E     x       �4 .;2 
�11  =� 3� .G  
�1�~  �� �� (� 
��  � � (�S  
��  H� >� (<0 
��_  �� �� ;W- Z�E      Z�E            
�~ �- � � v- K� G� i- �� �� &Z�E            �- �� �� i�E     �u Us    K�- ~�E       � 
��- �� �� �- 7� 1� �- �� �� � 	. �� �� . ~�E      `� �$ �. � 	� �. Z� X� ��E     �t UsT13�. s   {��E     �t    Y + 
�0�E            �� .;2 
�11  �� ~� .G  
�1�~  �� �� (�S  
��  �� �� (<0 
��_  7� 5� >�E     yg Uu 3- s   5|$ 
k� :ptr 
ka   v�  
m�}  1R�  
r|    5-E 
\% �S  
\#�  ��  
]#�w  �3 
_�h   2@@ 
A�  [ � 
A*[ 8Q 
B*b  �A 
D�w   |  '�Q ��  � v�  �+�}  ٶ �+v{  � �+[ � �+��  dN ��  �< ��  A ��w  2 �?  T\� , 5lM �� v�  �&�}  � �&[ �3 ��h  �@ �?  ʞ  �� �= �?  > ��w  �N ��w  ��  wS  :� �w  C o  � �  ]� ��  �   1� ��w  �m ��w  8Q �b    $N  5�( 45 � 4%�w  :� 5%�w  jS 6%�w  U 7%��  
A 8%�w  ?A 9%?  N :%�]  & n�w  17 n"�w  b o�  e�r �e�r �e�� �18x1 }�  8y1 ~�  8x2 �  8y2 ��  8x3 ��  8y3 ��  8x4 ��  8y4 ��  ]� G� ��  �� ��  8x ��   ] G� ��  �� ��  8x ��   1G� ��  �� ��  8x ��     5�& 	,[ � 	,�z  �\ 	-�   '�R �?  � �  �'��  � �'4~  ` �'4~  �/ ��w  �L ��w  " ��w  � �?  i �o   5) B� �  B��  v�  C�}  �3 F�h  ? H�w  O I�w  �/ J�w  9H L@   �1 M@   E N@   \< O@   �, Q�_  � R�_  s S�_  �R T�_  8i V@   [  W�w   W�w  1j @   �K �w  Q �w  -�  "�w  �  �w    Y�# �@�E     Y       �� .�# �${  b� Z� |ptr �$�  �� �� #V�E            � (x  �@   A� =� (\9 �a   �� |� j�E     u� Tv   ��E     L Us   20 �a   � �# �0{  :idx �0@   \9 �a    2�A �a   � �# �/{   2w0 �@    �# �*{   5WS �& �# �%{   58; �L �# �({  �- �(@    G�M _?  ��E     �       �y .�# _.{  �� �� .�- `.@   H� >� p\� ���E     % y G b� e�  �\(R�  f|  �� �� (|7 h@   � �� ;5 �E       �E            y' N v� t� B �� ��  ��E     �� T1Rv Y�\  K5 ��E       py �N �� �� B �� ��   5`" L� �# L({  R�  N|   5= 8� �# 8${  R�  9$|  � :$�z   ;$@    -Z3 		�  P�E     	      �� �3 		&n  � � �  
	&W  �� �� �^ 	&�  �� �� 	<0 	j  c� Y� cff 	BN  �� �� sub 	wS  � � i� 	�   	��  	�  }� y� <�u  =	��E     #��E     a       5 	n�  	h  �� �� #@�E             	'�  )	{  � � 	�8  *	�W  -� +�  B�E     Us�&T�Q  W� ��E      �� 4	� U� S� � z� x� �� � �� �� =� ��E            � �� �� � �� �� &��E            0�      ,�$ ���E     �       �b �3 �6n  � � �  �6�C  f� b� �  �6W  �� ��  �6�W  �� �� Zy  �6?  2� .� &  �6	  q� k�  �6`  �� �� A: �66`  �� �� cff �BN  � � � \�E      �� �. � L� J� � q� o� �� � �� �� =� ^�E            � �� �� � �� �� &^�E            0�     2�E     2 Us T�TQ�QR�RX�X�  '�B ��  � )cff �.BN  �j �.�  n ��  �  ��  ��  ��   '�; ��  � �& ��  ��  ��  E  ��   o+S ���E     q       �� �3 � f  � � 	R�  �|  [� Y� e6 ��E      �x �s s6 �� ~� �x �6 �� ��   ��E     �� Uv   -�4 ��  ��E           �	! �3 �)f  �� �� �  �)�  Q� G� �  �){  �� ��  �)�  $� � V �){2  �� �� �  �)G(  $� � Zy  �)?  �� �� &  �)	  �� �� �  �)�g  �� �� %�~ �  	s  �a0  � �   	~ �}  K� G� 	�O  ��  �� �� ,�E     Ԃ T	�BH     Q1   S�E     �6 Us T} Q��R~ X �  -y; ~�  p�E     �      �C" 9�3 ~)f  U$ )u2  �� �� ��  �)�  �� �� 	Xc  ��e  ;� 7� ip �u2  �� s� 	�� �u2  �� �� 	<0 ��b  :� 8� <�J vӗE     <��  zӗE     T��  }0v top ��&  k� ]� op ���  %� � 	�\ �H  �� �� �v 	��  2�  9� 1�    } ��  �E     �       ��" .�3 �3�h  �� �� .�j �3�  �  � Rn ��  Z� R� (la �  �� �� (s  �a0  � � �~ (F@ ��  [� Y� ��E     � T}    -�S VU  `�E            ��# yW V+�.  �� ~� ��  W+-#  �� �� 	�  Y�3  �� �� 	s  Za0   � � fm�E     U�UT�T  -�# J�  P�E            �$ yW J,�.  L� H� ��  K,U  �� �� 	�  M�3  �� �� 	s  Na0  �� �� f]�E     U�UT�T  ,(- >@�E     (       ��$ yW >&�.  � � 	�  @�  f� d� 	R�  A|  �� �� W�E     ��  -�F *�   �E     )       �2% yW *&�.  �� �� m  +&�  
� � 	�  -�3  E� C� 	R�  .|  j� h� 	s  /a0  �� �� fI�E     T�UR	�E     X0  -& "�  �E            �t% 9�  ""�3  Ucidx #"�  T G9 �U  ��E     d       ��% .
H �,�w  �� �� >��  �,-#  T(E  ��  � � (��  �U  �� �� <�u  �E      G�3 ��  ��E            �K& >
H �-�w  U.��  �-U  �� �� (E  ��  � �  Y�G �`�E            �x& >
H �'�w  U G� ��  0�E     %       ��& >
H �'�w  U>m  �'�  T(�  ��3  <� 8� (= ��0  w� s�  G� ��  �E     1       ��' >
H �$w  U>m  �$�  TC�) �E      �E     .       ��) �� �� �) �� �� &�E     .       �) � � �) >� <�    G�  {�  ��E     1       �/( >
H {&w  U>m  |&�  TC�) ��E      ��E     .       ��) c� a� �) �� �� &��E     .       �) �� �� �) �� ��    GR cU  ��E     U       �() .
H c'w  � � .��  d'-#  h� ^� (E  f�  �� �� (��  gU  |� n� p�u  t��E     C() ��E      ��E     
       lE) � � 9) <� :� &��E     
       Q) c� _� ��E     �~ Uv Ts     2� ?�  �) 
H ?'w  ��  @'U  E  B�  1� G�  8n G�  la H�  1��  R�     Y(H 5��E             ��) >
H 5!w  U 5> #�) 
H #!w  �0 $!�  �  &�3  s  'a0   'h�  �	U  * )r �	U   ,,�  �	 �E     P       �+ 9B� �	u2  Uss  �			  �� �� ߢ  �	�  �� �� W�Q  �E      �u �	�Q � � �Q @� >� �Q e� c� �Q �� �� �Q �� �� �u �Q (� &� �Q Q� K� R �� �� DR  v R �� �� R � �     ,��  x	@�E     �      �, �  x	!�  G� A� ��  y	!�&  �� �� ��  z	!wS  �� �� 	��  |	)V  � � n }	�  u� Q� 	.� }	�  �� �� #��E     1       �+ !ߢ  �	U  �t @�) h�E      h�E            �	3* �� {�   ,�  5	жE     �      ��, �A 5	!�h  �� �� 9�3 6	!a   T�  7	!?  R� N� #�E     �       �, 	�3 =	f  �� �� �E     �. Us Tt Qq   &зE     �       	 X	n  �� �� ڷE     �. Us Tt Qq    /e? �W- <0 �*�_  �S  ��*  N� ��  1p1 �  p2 �  �i   	u2    '�N ��  �- <0 �(�_  )x �(�  )y �(�  � ��   '� ��  �- <0 �(�_  �S  ��*  � ��   'f7 ��  . <0 �'�_  )x �'�  )y �'�  � ��   /C/ j. <0 j&�_  )x k&�  )y l&�  &| m&h  �S  o�*  1oI t  �i  uu2    ', a�  �. <0 a)�_  .� b)�   ,# U�E     0       ��. 9<0 U!�_  U	)�  W�W  �� ��  ,�& 	 �E     �       ��/ O 	!�_  �� �� 9<0 
!a   T9�  !?  Q%P} a/ 	:0 �b  6� 4�  &��E     .       	L *j  [� Y�   ,�+ �@�E     �       �+0 <0 �,j  �� ~� 	�S  ��*  �� �� 	N� ��  ?� ;� �u p1 �  |� v� p2 �  �� �� 	�i  �u2  � �   'X ��  n0 <0 �*j  )x �*�  )y �*�  � ��   --6 ��   �E     x       ��0 <0 �*j  ]� W� 	�S  ��*  �� �� 	� ��  �� �� |�E     � T0Q1  'J }�  ,1 <0 })j  )x ~)�  )y )�  � ��   /� W�1 <0 W(j  )x X(�  )y Y(�  &| Z(h  �S  \�*  1oI a  �i  bu2    '�? N�  �1 <0 N#j  .� O#�   ,�( B��E     0       �2 9<0 B#j  U	)�  D�W   � �  ,�R кE     8      �3 <0 $j  I� C� �  $�C  �� �� �  $W  �� �� )�  $�W  *� $� Zy  $?  z� v� & �E     u       	��  �  �� �� #L�E     )       �2 	'�  {  �� �� 	�8  �W  � ��  ,�E     ��   ,@N ���E     �       ��3 <0 �)�b  D� :� 	�S  ��*  �� �� 	N� ��  � � `u p1 �  b� \� p2 �  �� �� 	�i  �u2  � �   '"1 ��  �3 <0 �'�b  )x �'�  )y �'�  � ��   -} s�  ��E            �b4 <0 s'�b  d� Z� 	�S  u�*  �� �� 	� v�  k� i� �E     � T0Q1  -gL b�  ��E     T       �J5 <0 b&�b  �� �� 7x c&�  � � 7y d&�  �� �� 	� f�  � � 86 ��E       �� i$5 W6 H� F� J6 p� l� ��E     Ws Us T1  '�E     J5 Us Tv Q| R1  ,`I J��E     �       �86 <0 J%�b  �� �� 7x K%�  �� �� 7y L%�  &�  � &| M%h  v� r� 	�S  O�*  �� �� &ӢE     D       	oI T  � �� 	�i  Uu2  (� $� �E     O� "6 U�T  �E     O� U|    'O A�  e6 <0 A(�b  .� B(�   /a' 5�6 <0 5 �b  )�  7�   ,
6 ���E     $      �K7 <0 �"�b  d� ^� �  �"�  �� �� �  �"{  �� �� )�   "�  E� ?� Zy  "?  �� �� &չE     \       	��  �  �� �� �E     ��   ,^= ���E            �z7 9�  ��Y  U ,gD ��E     �       ��7 9�  ��Y  U92�  �u2  T9�� �u2  Q9R�  �|  R -a! ��  ��E     )       ��8 �  �(�Y  �� �� �? �(�  6� 0� �D �(�  �� �� b�  �(�  �� �� �I ��E      pz ��8 �I (� &� ��E     M Uu Tt   HɨE     �D U�UQ�TR�Q  -�3 ��  ��E     E      �K: �  �(�Y  [� K� �L �(�  
� � �  �(�J  J� B� �I ��E      P| �Y9 �I �� �� ��E     M Uu Tt   WF ��E       �| �LF �� �� ?F � � 2F R� F� %F �� �� �| YF y� w� fF �� �� sF b  Z  ~F �  �  ^�F p�E     D�F �| 6�F ���F   �  (�E     �R -: U��T} Q0 f�E     M Uu Tt      -�$ ��  �E             ��: �  �"�Y  M I b�  �"�  � � �I �E       } ��: �I � � �E     M Uu Tt   H �E     �R U�UQ	�T $ &  -�* d�  ��E     q      ��< �  d"�Y   � Ӏ e"u2  � � �: f"		    ? g"�>  � � 9�= h"?  Xi� j�   cur ku2  � t <�u  ���E     �I ��E      �t n�; �I   ��E     M Uu Tt   W+R ΏE      �t �dR 7 ' WR � � JR Y K =R � � �t oR r j zR � � �R � � �R 	 	 D�R  u �R �	 �	     -z! Z�  p�E            �<= �  Z �Y  >
 :
 �I p�E      p�E     	       \ = �I y
 w
 y�E     M Uu Tt   H��E     pT U�UTt   -  �  @�E     O      ��> �  /�Y  �
 �
 �F /cZ  9 - >�  /�  � � :�  /�  ^ R � /�>  � � !(2 �> ��y	�2 Z  k e !$2 �  ��y	� �  � � 	u�  u2  P J 	��  u2  � � !y> +\  ��y<�u  T��E     ��E     �F �> U T��yQ R��y 0�E     �> U T��yQv R| X0  5[  �>  L    -�F �  ШE     e      �XD �  )�Y  � � �F )cZ  2 $ >�  )�  � � :�  )�   	 � )�>  t p !�2 5[  ��Xcur u2  ��~	�� 	u2  � � 	.� 
�  +  idx �  � � 	� �  � � 	� �[  � � <�0  ��E     <� 6 �E     <@ ]��E     <�u  ��E     %| �@ !�  5[  ��	�4  u2  � � 	��  !u2  � � ��E     �G U T��  %�z :D q Du2  "  val E�  � � 	�� F�    %�{ QA 	R�  t|  � � len u�     ~�E     �� A U��~ ��E     �� <A T ����Q��~ ��E     u� Qv   #��E     f        B !/� �XD ��	�!  ��  X V 	E  ��  } { �E     �D �A U��~Q4R��X0 (�E     O� 8�E     O� I�E     O� Z�E     O�  %{ |C 	R�  �|  � � 	/� ��  � � 	E  ��  � � i ��  � � %P{ �B 	�!  ��  + ' ��E     O� ��E     O� ��E     O� ʪE     O�  ��E     �� �B U��~T8Q0R��~X0Y��~ '�E     �D !C U��~T~ Q} Rs ����3$v "X0 H�E     M ?C Uu T~  �E     �� _C U��~Tv  �E     �� U��~Tv   hD ��E      �{ N�C �D zD g a �{ �D � � �D  �   ��E     M �C Uu Tt  ��E     pT D U��~ �E     �R D U��~Q3 ԬE     �R U��~Q0   �E     �G U��~T��  �  hD  L    '� �S   �D �5 �{2  �� �u2  cur �u2  E  �?   -�K U�  @�E     ]      �F �5 U{2  u g �� Vu2    �? W�  � w �D X�  0   b�  Y�  � � cur [u2    	.� \�  T < c ]h  V N 	�]  ]h  � � <�u  �7�E      z !��  s�  ��	�4 tu2  � � �E     �R �E U��Ts Q��� $ & )�E     M Uu Tt    '�? �  �F �5 {2  �� u2  �L �  �  	�J  cur u2  .� �  c h  �]  h  T�u  H1��  #�  �4 $u2    ,L- �p�E     �       ��G �  �(�Y  I = ? �(Z  � � � �(�  k  e  ? �(�]  �  �  !��  �5[  ��% t �G 	u�  �u2  Q! K! 	��  �u2  �! �! cur �Z  �! �! 	�� �Z  C" =" Pt !�2 �5[  ��(�E     �G U| T��   ��E     �G U| T��  ,�A j��E     �      ��I �  j"�Y  �" �" �2 k"Z  # # cur mu2  m# k# 	�� nu2  �# �# 	�- o�  �# �# �I ƌE      ƌE     	       w�H �I ]$ [$ όE     M Uu Tt   �I ՍE      �s ��H �I �$ �$ ߍE     M Us Tt   �I �E      �E            �	JI �I �$ �$ �E     M Us Tt   �E     �I bI Us  `�E     rL �I Uu Tt  ��E     �J �I U�PT|  �E     �I Us   /H `�I �  `%�Y   ,�2 �`�E     /      ��J �  �'�Y  �$ �$ Xcur u2  �`	�� u2  h% ^% 	� �  �% �% <�u  Ka�E     ��E     M lJ Uu Ts  �E     �K �J U�`Ts  =�E     �J �J U�`Ts  ]�E     rL Uu Tt   -~  ��  0�E     $      ��K �5 �{2  �& �& �� �u2  v' l' cur �u2  �' �' 	�- ��  ( ( 	� ��  �( �( ~end �ʉE     �M  �E     '       �	�K �M �M & �E     '       �M �) �)   q�E     rL �K Uu Tt  �E     �K U�hTz   -GI ��  ��E     c       �rL �5 �{2  �) �) �� �u2  * �) cur �u2  M* K* err ��  t* p* �E     M Uu Tt   -�  O�  ЇE     �       �M 9�5 O#{2  U9�� P#u2  Tcur Ru2  �* �* 	�- S�  0+ $+ 	� T�  �+ �+ i UZ   , , �s c Zh  x, n,   ,�? 1`�E     c       ��M 9�5 1{2  U9�� 2u2  Tcur 4u2  �, �, ��M ��E     "       =�M �M &��E     "       �M *- &-    /I �M �5 {2  ��  u2  cur "u2   ,� 0�E     f       �zN >) RX  h- b- 	R�  |  �- �- X�E     �� MN Uv  k�E     �� eN Uv  �E     �� Uv   Y " �p�E     �       ��O .>) �RX  �- �- (R�  �|  [. Y. b� ��  �\(�5 �u2  �. . ;dP ��E      ��E     8       �]O }P �. �. qP �. �. &��E     8       �P / / �P @/ >/ �P e/ c/   ��E     �� {O Uv Q�\ ��E     u� �O T|  
�E     �� Uv T|   25 ��  P >) �RX  :idx ��  ݰ  �a   ss  ��  1� ��  6^  �		  � �	    20) v�  dP >) v#RX  6^  w#		  R�  y|  �5 zu2  � {�   5�P e�P >) eRX  �5 fu2  � h	  x  i{2  �� j{2   G% G�  ��E     �       ��Q .>) GRX  �/ �/ ..� H�  "0 0 .R�  I|  z0 n0 b� K�  �Le�u  \��E     �� VQ Uv T8Q0R| X0Y�L ؠE     �� nQ Uv  
�E     �� Uv T4Q0R| X0Y�L  '|% .�  +R y�  .${2  �� /$u2  B� 0$u2  )n 1$		  ߢ  2$�0  p 4u2  r 5�  s 6�  1val E�  b F�    '�* ��  �R y�  �&{2  �� �&u2  B� �&u2  )n �&		  p �u2  r ��  w ��  pad ��  1c ��    G�2 ��  0�E           �pT .y�  �{2  1 1 .�� �u2  U2 52 .b�  ��  �3 �3 qp �u2  ��(n �u2  �4 �4 (|A ��  C5 5 (�( ��  7 �6 (�J ��  B8 &8 (�b �?  p9 b9 (��  �?  /: : ( �?  9; ); �Bad a<(�  ee�E     <��  j�E     <�u  [e�E     %�y �S Rc �P  �; �;  %�y 6T 	T�  �  :< 6< !�E     pT U��Tt   ��E     pT UT U��Tt  ��E     h� Uv T|   G�8 ��  ��E     p       �!U .y�  �{2  z< p< >�� �u2  Tqp �u2  �X(n �u2  �< �< Rnum ��  B= >= �E     !U U Uu Tt Q: K�E     !U Uu   Gz* T�  ��E     f      �V >y�  T{2  U>�� Uu2  T.2�  V�  �= x= Rp Xu2  > > Rnum Z�  �> �> (�b [?  3? %? (��  \?  �? �? (�O ^�  \@ V@ (Gs  _P  �@ �@ �Bad ���E     ps Rc }P  �@ �@   -\P ^�  p�E     h      ��] �  ^!Jn  :A .A 	R�  `|  �A �A fi a�3  �A �A 	� b�  5B B key c�   "C C Xlen d		  ��~	�0 e�  ^C XC <�0  �F�E     %P� _] !p$ r�] ��~%В UX n ��  �C �C �` P�E      P�E     (       ��W �` �C �C �` �C �C &P�E     (       6�` ��~j�E     �b Us T��~Q1   W�] x�E       � �^ "D  D �] LD FD �] �D �D @� ^ �D �D 6^ ��~F+^ [4^ ��E            X 5^ E E ��E     �a  ��E     � 7X Us T0 ��E     � Us T��~    �D^ �� �H\ V^ �� c^ 8E 2E p^ �E �E 6}^ ��~F�^ �_ �E      � "0Z �_ �E �E � ` F �E ` gF cF ` �F �F 6&` ��~3` �F �F >` ^G ZG FK` �` .�E      `� V
zY �` �G �G �` �G �G `� 6�` ��~3�E     �b Us T��~Q1   Mt` �� �Y 6u` ��~��E     �a T�E     �b Us T��~Q5  [T` ��E     5       Z Y` H H 6f` ��~��E     �� T(Q0X0Y��~  ��E     � Us T��~   �^ ��E      Б )\ �^ >H 8H Б �^ �H �H �^ �H �H �^ HI DI 6�^ ��~�^ �I ~I �^ �I �I F�^ �` ��E       � �
[ �` "J  J �` LJ JJ  � 6�` ��~��E     �b Us T��~Q1   M&_ P� �[ '_ {J oJ M4_ �� o[ 5_ K K 6@_ ��~T�E     �b Us T��~Q4  �E     �a ��E     �� T|  $ &Q@R	P�E       [_ ��E     5       �[ _ RK PK 6_ ��~��E     �� T@Q0X0Y��~  K�E     � Us T��~   %�E     � 9\ Us T��~ ;�E     �a   �` x�E      x�E     #       x�\ �` xK vK �` �K �K &x�E     #       6�` ��~��E     �b Us T��~Q1   ��E     �a ��E     �b �\ Us T��~Q1 ��E     �b ] Us T��~Q1 ��E     �b >] Us T��~Q1 B�E     �b Us T��~Q4  ��E     � ~] Us T��~ ��E     � �] Us T��~ R�E     �� �] U}  m�E     �� U}   r  �]  L    '�; @�  D^ �  @(Jn  )n A(�  #  B(zv  key D�   len E		  T�0  X1�2 Qzv    '�! �  �^ �  $Jn  � �  key �   len 		  T�0  : '� ��  P_ �  �%Jn  fi ��3  kp �D3  key ��   len �		  n �S   tmp ��  T�0  ]&_ R�  �|  � ��   1�2 �zv  1r ��  p$ ��]    -�% �S   P�E     )       ��_ ca �(�  Ucb �(�  Tkp1 �D3  �K �K kp2 �D3  �K �K 	��  ��  L L 	��  ��  8L 4L  'o2 L�  �` �  L%Jn  fi N�3  tk O�2  key P�   len Q		  n RS   tmp S�  T�0  �]t` R�  `|  � a�   1p$ j�`   r  �`  L    '�$ 8�  �` �  8$Jn  ` 9$�]  val ;r   ,�= . �E            �%a �  . Jn  �L �L 	R�  0|  �L �L 0�E     ��  -; �   �E     g       ��a �   Jn  M �L R�   |  UM OM 2�   u2  �M �M ��  u2  �M �M 	Jy  Go  KN EN !� �  �LH�E     �� Uv T Q�L  -.C �zv  �E     �       �]b 7key ��  �N �N 7len �		  �N �N n �
S   CO 9O 7�E     � T| Q}   'I ��   �b �  �$Jn  + �$?  )len �$�b Jy  �Go  key ��    		  -{M t�  пE     {      �Yd �  t%Jn  �O �O �M u%#r   P P 7n v%�  aP YP 	Jy  xGo  �P �P Xstr y�   ��i z�  TQ NQ � len �		  �Q �Q val �#r  �R �R #��E     B       �c 	R�  �|  
S S !� ��  ����E     � �c T Q�� �E     u� Q��  �E     Yd n�E     pT d U��Tt  ��E     e \��E     =d T ��E     �R U��Q0   G*! ��   `�E     h       �e .Jy  �'Go  1S -S Rstr ��   kS gS %� �d Rch �S   �S �S  K�e `�E      � ��e �S �S � _�e  o�E     Ig Uu     G� z�   �E     x       ��e .Jy  z$Go  T  T Rstr |�   hT dT %P le Rch �S   �T �T  C�e �E      �E            �e �T �T &�E            _�e  �E     Ig Uu     2�? ^S   �e Jy  ^'Go  8ch `
S    2�6  �H  0f :a �H  :b �H  8ret �.  8tmp �.   *�I ��E     	       �mf ?�I UH��E     M Uu Tt   *e6 ��E     0       ��f ?s6 U�6 U U  *,1 �E     H       � g :1 BU >U G1 U {U R1 �U �U ?]1 Rj1 �U �U &�E     -       x1 V V �1 AV ?V   *�) p�E            �Ig * nV dV  *�e p�E     c       �yg ?�e U�e �V �V  *�, P�E     �       ��g - - 	W W "- 2W ,W D/- P� 0- �W |W <- �W �W H- 4X 0X   *e�  `�E     �       �Dj s�  ~X zX ��  �X �X ��  
Y Y ?��  Y��  ��  ��  IY CY �e c�E       �� ��h f �Y �Y f �Y �Y �� f Z Z #f KZ GZ   �e ��E      P� ��h f �Z �Z f �Z �Z P� f �Z �Z #f [ [   �e ��E      �� �?i f f W[ U[ �� f �[ |[ #f �[ �[   �e ��E      @� ��i f  \ �[ f %\ #\ @� f N\ J\ #f �\ �\   �e �E      �� ��i f f �� f �\ �\ #f ] ]   �e $�E      � �)j f P] N] f � f w] s] #f �] �]   ��E     ��  Uu Ty   *��  `�E            ��j ?��  UC5 c�E       c�E            bN �] �] B ^ ^   *��  ��E            �k ?��  U̎  C^ A^ C5 ��E       ��E            pN m^ k^ B �^ �^   *��  ��E     2       �Qk ?��  U?̎  TH��E     �j 3̎  t   *��  ��E     5       ��k ?��  U?��  Tf�E     3��  t   *Q�   �E     h       �	l ?b�  U=o�  p�E            ��  �^ �^ C5 t�E       t�E            �`N �B �^ �^    *'�  ��E     o       ��l ?8�  UD�  _ _ ;َ  ��E       ��E            �yl �  U_ S_ �  U_ S_  ='�  ��E             D�  z_ x_ 8�  �_ �_ C5 ��E       ��E            �N �_ �_ B �_ �_    *ύ   �E     >       ��m ?܍  U�  ` ` ;َ  �E       �E            �Wm �  b` `` �  b` ``  =ύ  (�E            �  �` �` ܍  �` �` C5 ,�E       ,�E            �`N �B �` �`    *� @�E     Q       �Yn � �` �` � ca [a D�  � � �a �a  � 0� D�  � � b b ]�E     �� An Uv  t�E     �� Uv      *�O ��E     �      �]p �O Gb 9b �O �b �b �O �c vc �O -d d D�O 0� �O �d �d �O ie _e �O �e �e �O M�O p� Ap �O Ff Bf �O �f }f P g �f KP 8�E      �� �3P �g �g 'P �g �g �� ?P >h 6h KP �h �h 6WP ��;dP �E      �E     8       ��o }P i i qP ,i *i &�E     8       �P Qi Oi �P vi ti �P �i �i   E�E     �� 
p U��Ts Q�� �E     u� "p T~  ��E     �� U��T~     �E     u� T Q}    *�  p�E     �       �-r '�  �i �i 4�  ij _j A�  �j �j N�  5k -k ?[�  � �  �  h�  �k �k s�  �k �k ��  8l 4l ��  rl nl ^��  �E     َ  p�E      � !5q �  �l �l �  .m $m  M��  P� �q 6��  ����E     '�  iq Uu Ts  ��E     '�  �q Ts ��E     � U} Tw   D�  ��E      ��E     
       F�q R�  �m �m R�  �m �m  ��  3�E       3�E            ,r ��  �m �m  0�E     '�  Uu T0  *��  ��E     j       ��r ��  �m �m ��  Fn <n ��  6��  �`��  �n �n ��  o 	o ��  Go Co �  �o �o [�  ��E            �r �  �o �o '�  �o �o  B��E     T�TQw   *�   �E     i       �Ws �  2p *p <�E     Q�  /s Us  ��E     ]�  Us TsQs��Y1  *86 ��E     '       ��s J6 �p �p W6 �p �p H��E     � Q0  *86 ��E            ��s J6 q q W6 cq ]q H��E     Ws U�UT�T  *�3 @�E     J       ��t �3 �q �q �3 Or Cr �3 �r �r _�3 D�3 Ќ �3 us ks �3 �s �s �3 st it Ќ �3 �t �t l�E     �3 �t Us  H��E     b4 U�UT�TQ�Q    *. ��E     '       ��t �. u u �. H��E     � Q0  *�- ��E     <       ��u �- Nu Ju �- �u �u �- �u �u 0	. @. ��E      ��E     ;       �`H. =. v v 2. Bv >v %. v {v &��E     ;       U. �v �v =b. ��E     %       c. �v �v p. w w     *W-  �E     �       ��w i- 1w 'w v- �w �w �- @x 4x �- �x �x �- �E      � ��v �- !y y � �- �y �y �- �y �y ��E     � T0Q1   @�- d�E      d�E     (       ��- z z �- Az ?z �- fz dz &d�E     (       	. �z �z . d�E      d�E            �^w �. �z �z �. �z �z r�E     �t UsT13�. s   ��E     �t Us T| Q}     *�1 0�E     '       ��w �1 { { �1 P{ L{ HW�E     � Q0  *�1 `�E            �x �1 �{ �{ �1 �{ �{ Hf�E     �w U�UT�T  *�0 ��E     d       ��y �0 3| -| 1 �| | 1 �| �| 1 %} #} �1 ��E       �� ��x �1 J} H} �1 r} n} ��E     �w U| T1  =�0 ��E     D       1 �} �} 1 �} �} �0 $~ "~ &��E     D       01 @,1 ��E      ��E     D       �]1 I~ G~ R1 q~ m~ G1 �~ �~ :1 �~ �~ &��E     D       j1   =�f ��E     (       x1 3 1 �1 X V       *+0 ��E     J       �~z =0 � { J0 � � U0 �� �� _`0  D+0 �� U0 A� 7� J0 �� �� =0 ?� 5� �� `0 �� �� �E     n0 Xz Us  H:�E     �0 U�UT�TQ�Q    *� @�E     �      ��~ � � ق � H� @� � �� �� � � �  �� ��  � 	� ? � * � s� 6 �� �� B � � ^N 6�E     ^V ��E     ^^ P�E     =f ��E     u      g �� �� r B� 6� } ы ǋ � X� N� � ߌ Ռ � f� \� � � � � h� ^� N�e ��E      0� ��{ f f 0� f � � #f A� =�   [� (�E     p       �| � �� |� 0�  �� �� F�E     h� O| Tv  u�E     �� �| U}  $ &T~  $ &Q��� $ & ��E     h� Uw �@$ $ &Tv   N�e ��E      �� �} f 0� .� f U� S� �� f ~� x� #f ֐ А   [ ��E     V       �}  -� )� 0 ( h� d� �E     h� R} Tv  1�E     �� ~} U}  $ &Q
w � $ & ?�E     h� U~  $ &Tv   [� p�E     �       I~ � ޑ ڑ � � � � L� H� ��E     h� �} Tv  ��E     �� $~ U}  $ &Q��� $ & ��E     h� Uw �@$ $ &Tv   ��E     h� i~ T
s 1$ $ & ��E     h� �~ Tv  b�E     h� U���@$ $ &Tv    �()  �E     }       �A 9) Ē �� E) � � _Q)  D]) Џ ^) O� M� j) �� �� t) �� � D�)  � �) @� >� W�E     � T~     *() ��E            �� 9) i� c� E) �� �� _Q)  H��E     �~ U�UT�T  *]b  �E     b       �� ob � � �b H� D� �b �� ~� �b �� �� `|b �E     Yd � Ux  &�E     e Ux   *��  ��E     �       �z� �  '� � �  �� �� �  �� � 0&�  N1�  ��E      �� �
�� N�  F� B� B�  �� |� =1�   �E            N�  �� �� B�  ݗ ۗ C5 #�E       #�E            r`N B �  �    =��  ��E     G       �  �  �  &��E     G       &�  )� %� K��  ��E      �� �$��  d� `� �E     Dj Ut      *o�  ��E     X       �7� ?��  U;5 ��E       ��E            �݁ N �� �� B Ø ��  =o�   �E            ��  � � C5 �E       �E            �`N �B � �    I�X  �X  "~IaG  aG  �g\  \  VI�A  �A  �g5<  5<  ?r�D  �D  > ri0  _0  > I�K  �K  ?vI�6  �6  ?�IF\  F\  ?�gjO  jO  IC  C  `Io+  o+  �gKM  KM  YIBi  Bi  @I],  ],  eI_T  _T  AXI��  ��  @IkA  kA  ?{ d5   �  �  �X $"  �/F     &      �Z X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  	)  �  	5  >   G   �	  	N   	N  �  B"l  r     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  `  -      n�  �  �  `  U    �  �    U   ,  `  -   -   U    �  �"8  >  �   PJ�  2�  L;   �  M@   pos N@   �  P�  SF  Q�   �1 R  (=9 SM  0R�  U`  8y�  V;  @�� W;  H �  ��  �\ �-   m  �U    o  ��  �  �    @   ;  ,  @   ;  @    A  �  	A  2  Z  `  k  ,     :-   �  J�  x Lk   y Mk   )  Ow  	�  B   s�  M   uk   }  uk  V  vk  /  vk   t
  x�  k	  (y  �  N    ��  N   �  	G   B� 
;  L  5    A  s  A  v	  U     �  �  	y  �  (N�  �  P)   Z�  Q)  �  S�  s  T�   [  U�  ?1  WG     �  )    Y�  �  =  N   �K  �   M
  pmoc5  stib	  ltuo|  tolp 	  �  b   "e  k  �  %  <�  x >)   len ?5  *� @A   %  Bp  	�    `�  �  �  G   G   �  U    �  �  q�  �  G     G   G   U    �  %  +  @  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  ��  ()  �  0R   �U   8�  ��  @ �  �  �  �@  	�  �   �  �  G     U      X  �  &  ,  7  X   �  ?D  J  _  X  ;  @    �  Yl  r  G   �  X  @   U    s  ��  �  G   �  X  �   �  W  0�  �  �K   e� ��  �� �7  �� �_  �� ��   �� �  ( �'  ��  �!  lA  �  �@  �  -  �A  	G  S  �  ��   	^  �
  �)  �  �5  �  �G   	�  
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   b   �&	  xx ��   xy ��  yx ��  yy ��   a  ��  	&	  z'  �c	  m  �X   ss  ��   �  �8	    �}	  �	  �	  U    �  ��	  �U  �U      �p	   %  ��	  �  $�	  �	  �   
  �� "�	   �@ #�	  �U  $U    �  7=
  �; 9�	   ��  :�	   L  <
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @	=  ��  	?k   �  	@k  ~  	Bk  �  	Ck  �  	Dk   5  	Fk  (B  	Gk  0�  	Hk  8 �	  	J�  
   	sn  �  	uo   ��  	vo  �  	xk  �
  	zk  (  	{k   �  	}  �  	�#�  �  k  `
�=  R�  
�`   (  
��  |  
��  �  
��  �  
��  �  
��#  v  
�=
  �  
��  (�%  
�=  07&  
��#  8G   
��  X �  	�"J  P  h  
�  �M 
�#   k  
{  R�  
`   �  	�"�  �  %  8
;�  �� 
=�#   �M 
>@    
?=
   r$  
@u  0 5  	�$�  �  %  �
g  �� 
�#   �M 
�#  �  
K   �  
�  (�� 

X  h�� 
�  p�� 
w  x K  	� t  z  �  �	,;  �   	.�   �  	/�  O  	1�  C  	2�  �  	4�   d> 	6�  (A  	7�  0T  	9�  8  	:�  @�  	<�  H�  	=�  PE-  	?�	  X�!  	D�  h:  	F{  �  	Go  ��  	Ho  ��  	Io  ��  	Ko  �  	Lo  �U  	No  ��  	Oo  �)�  	Q�  ��  	R;  ��� 	S�  �K1 	W�  �R�  	X`  �Jy  	Y,  �%  	[=
  ��	  	]�	  �    	^U   ��8  	`+  � L  	 H  N    X	��  �  	�g   E-  	��	  N 	��  �8  	��  P �  	*%�  �  �  0	t�  k  	v{   �  	wg  �@ 	x�  ݖ 	y�  E-  	z�	   N 	|  0�  	}�  pR  	~�  x�  	�  �ߣ  	�K  ��I 	�y  ��  	��  �h  	��  ��S  	��  �4  	��  �8  	��  �  	�U    �  	�-   �  	�k  o  	�k  �L 	�U    �8  	�	  ( �
  	L#�    W  	HL  �  	Jg   = 	K    	L{  d  	M{   �  N   	�  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  	L  (0  	O  #   	g)8  >  �   �
��  =  
�&	   L  
��   $  
��  0�  
��  8m  
�#r!  h�  
�4  pآ  
�A  tG   
��  x ^  n  �  �
  	�)�  �  �   H
�  �  
�U    "  
��  �!  
��   ~	  8	f�  �
  	h{   (  	i{  �� 	k�  �� 	l�    	nk  �  	ok   �  	pk  (�  	qk  0 y  	s    	�$�  �  �  0'	  �N  )�   ?1  *{  }0  +�  i/  ,�  � -&	   �  	�)       H
�  ��  
�u   ?1  
��  (  
�(  4  
�&	  \  
��  0  
�U   @ +!  	�  tag 	�   �U  	�   �  	  �  `  N   	
�  w%   }#  �&  h  �  &     	
�  E   	9
W  � 	;
�   ��  	<
�  �  	=
�  �  	>
�  �#  	?
�   �  	L
(d    �  N   	��  :   �   ^$  1  �!  �!   :  	�j  �  ��  �#  ��  �  �  �  =   I$  ��  �  �  =   �&  �    �    =     �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  ��  @ j  R  �%  	�  x  =}	  H  E#�  	�  �  @JS  �  L�   �  MK  �� O�  .� P�  �  QE   �  R�  (�!  S  08'  Tk  8   W!_  e  -  (l�  k  n{   �M o�  ߣ  pK  �  q�   �  k  )�  �  �  �  S  �   w   .�  �  �  S   �  1�      S       3	  K  6)  /  ?  S  ?   �  �  :Q  W  �  k  S  S   �  >�  "  Y�  �  �  �  �  �  �     �  _�  �  �  �  �  �       $  f�  �  �  �  �  ?   �  l
    �  )  �  �  �   #  x��  �� � �   �  � K  H  � w  P�  � �  X9!  � �  `l� � �  h  � �  p     �)  �  H2�  �S  4�   �  5�  (  6�  04  7�  88  8�  @ �  :�  �  �=u  R�  ?`   �  @�  n  A�  �  B�  1$  C(  2�  E�  �� F�  `�L HU   � �  J�  �  P   �  �  �  �  ,  g  �  �  �   �  &�  �  �  g   �%  *�  �  �  �  ;   �%  -      ;   {  1#  )  �  8  �   �  4D  J  U  �   l  8a  g  �  {  ;  W   �  <�  �  �  �  ;  �   �  @�  �  �  �  �  ;  �  A   �  G�  �  �    g  �  �  �   �'  N    �  '  g  ,   �  S3  9  �  \  g  �  �  A  \   �  &  ��@  �� ��   i'  ��  H   ��  P  ��  X�A ��  `Y ��  h�#  ��  p�  ��  x�  �  �  �8  ���  ��  �U�  ��  ��!  �  ���  �'  ��  �U  �&  �{  � �&  �L  b  �>  �z  'O  �   xC  ��   s/  �R  	z  �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }�  �  U'      m  D   tT   �  v�   A  w�  �  x�  &  y�   !  {   �  �l   r   �  �   �  �  �    c	  �  ��   �   �   �  �    �'  ��   �   �  �   �  �  (  �    T   �!  "!  ��  )`    ��  )�   �  )�    }  �   	"!  O  ;_!  _� =%_!   ݰ  >%�   /!  �  @4!  e!  cA  
�,�!  �!  /  
��!  �� 
�   �M 
��!   ?<  
�,�!  T"  �5  P
�T"  �  
��   �� 
�e"  �Y 
��"  �H 
��"  U@ 
��"   �9 
�#�"  (�A  
�#*#  0�^  
�#U#  8�^  
�#{#  @N7  
�#�#  H 	�!  ��  
��!  (Z  
�q"  w"  �  �"  x!  �   17  
��"  �"  �"  x!   �G  
��"  �"  �  �"  x!  N   %G  
��"  �"  �  �"  x!  �"   N  �@  
�#  #  �  *#  x!  x!  N  N   �;  
�6#  <#  (  U#  x!  N  N   �W  
�a#  g#  �"  {#  x!  `   *;  
��#  �#  �"  �#  x!  `  N   �T  
��#  �  �  
P  �  =  �#  @    �  �#  @    �  
�%  ��  #$  
$  N  $     d�  )%$  +$    :$  �   0�  /%$  K�  6n$  �> 8N   �^ 9�   �  ;F$  Ѽ  >$�$  �$  ў  (@�$  
H BY"   ��  C�  XT D�$    n$  ��  N�$  �$    �$  �  �   B�  V�$  �$  %  �     ��  Z%  !%  �  I%  `  z$  �  �$  �$  �   ��  bU%  [%  �  o%  z$  N   ��  f{%  �%  N  �%  z$  �"   5[ j�%  	�%  ��  @j&  �\ l �#   8` n %  �\ o I%  �_ p o%  �T r $   }�  s :$  (ʬ  t &  0�  u &  8 <  
�  �  �   ?&   @   o 	.&  
5V ?&  0  a&   @    	P&  6Y �a&  0  �&   @   � 	s&  (V ��&  <  �&  @   � 	�&  U )�&  �` J�&  H  �&   @   �� 	�&  vT u�&  !D&  	�J     !f&  	��I     !�&  	��I     !�&  	��I     !�&  	��I     !�&  	�I     N   ��)  �Y  $W �S }Z �W \ �W �S �[ wY 	�\ 
EW !_ �[ M] �\ �` �` �U �V �Z bZ  �Z !a "^ #K[ $eU %,\ &�U '�_ (p] 0,T 1<X @FZ A�] Q�X R�^ S>_ TZ U�] V�Z W�W X<a `t[ a�_ b�X c�` p[ �` ��Y ��V ��Y ��\ ��W �^` ��` �MU ��S �_ ��T �fX ��] ��^ ��_ �.U �'Z �}_ �Y �+] ��] �]T ��W ��\ ��V ��T ��[ ��Z ��T ��^ ��U �mV ��U ��Y ��[ �^_ �8^ �MV �CY �X ��T �W ��V ��U �gY � [  �)  @   	 	�)  "jW ��)  	�I     �   �)  @   T 	�)  "V ��)  	@I     �  �)  @   	 	�)  "O\ ��)  	 I     #T �%  	�I     �  -*  @    	*  #�S A-*  	�I     $"&  e	@I     %k\ H�  P1F     
       ��*  &~ H%=  4� 0� &�1  I%  q� m� 'Z1F     *5  (U	�I     (T�T  %F`    1F     #       ��*  )sid %�  U %�T 	   1F            �7+  &i�  	#�  �� ��  %�_ �N  P0F     �       �),  &>) �'z$  ՙ ϙ *�> �'�"  T+E  ��  )� !� +��  �N  �� �� ,�u  ��0F     -`� .min ��  &�  � .max ��  {� q� .mid ��  � � .map ��$  V� N� +�] �N  �� ��   %\ ��  �/F     �       ��,  &>) �(z$  � � *�> �(N  T.min ��$  @� >� .max ��$  i� c� .mid ��$  �� �� +E  �#�$  � ܝ - � +�] �N  p� l�   %5` <�  4F     �      ��/  &R�  <+`  �� �� &>) =+z$  � � &�  >+�  g� _� &��  ?+�$  Ο Ɵ &VX @+�$  2� .� &��  A+�  r� j� #� C�  ��~#w` E�/  ��~#�^ F�/  ��/0� �/  .n O�  ٠ Ѡ +.� P�  ;� 7� .map Q�$  �� q� +�_ RN  3� /� /`� /  +��  Y  o� i� 00  �� ^z.  1D0  170  1*0  10  -�� 2Q0  �� �� 3�4F     75  (T    0�/  г d�.  1�/  1�/  -г 2�/  (�  �   4�4F     w �.  (U} (Ts  5�4F     �0  �.  (U  45F     ��~�.  (U} (T  3�5F     �0  (U   5�5F     C5  =/  (Ts (Q8(R	�/F      5M6F     O5  W/  (U��~ 3�6F     [5  (U��~(T8(Q| ����(Rs (Y��~  3z4F     [5  (U��~(T8(Q0(R|
����(X0(Y��~  �  �/  @   	 6b^ '	0  7�_ ',N  7yl (,	0  8n *�   �  6]a ]0  7��  +  7)�  +�  7�^ +	0  7yl +	0  8n �   9LT �G   �/F     7       ��0  :a �"�  �� �� ;b �"�  T<`W ��$  ɣ ţ <eW ��$  � � <k[ �N  )� '� <"] �N  V� L�  9�\ ?N  �2F           �n3  =la ?"  � ߤ >�3F     V       �1  <.� M�  b� ^� <�\ NN  �� �� ?p O  �� � - � ?c T�   G� A� ?d UN   �� ��   /�� 2  <.� y�  � � <�\ zN  h� `� ?p {  ͧ ŧ -в ?c ��   1� +� ?d �N   �� }�   -� ?p �  � � ?dot �  "� � @n3  &3F     P� ��2  A�3  [� Y� A�3  �� ~� -P� 2�3  �� �� B�3  B�3  B�3  2�3  � � C�3  �3F     D�3  D�3  303F     =4  (U�U(Tt    En3  83F            �A�3  � � A�3  8� 4� F83F            2�3  s� q� B�3  B�3  B�3  2�3  �� �� C�3  =3F     D�3  D�3  3=3F     =4  (U�U(Tt      G^ /@   74  7F@ /*  7�� 0*  8c 2G   H.� 3G   8min 3"G   8max 3'G   8p 474  I�Y �I�Y WI�S �J4  8mid CG   8q D74  8c2 EG    KHx  wG   8q x74    H  Ln3  `1F     �      �*5  A�3  Ӫ Ū M�3  T2�3  |� p� 2�3  � �� 2�3  �� � 2�3  v� j� 2�3  � �� C�3  �1F     D�3  D�3  N�3  б �4  2�3  Q� G� 24  د �� 24  � �  O4  x2F     _       24  :� 6� 2*4  �� ��   P�*  �*  [QBi  Bi  Q_T  _T  XQF\  F\  �Q�6  �6  � �   ��  �  ~a $"  �6F     �      �e X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  �  B"C  I     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  7  -      n�  �  �  7  U    �  ��  �  U     7  -   -   U    �  �"    �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S  0R�  U7  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��  �  @       @     @      �  2  ,  2  =       :-   B   s�  M   u=   }  u=  V  v=  /  v=   t
  xI  k	  (  �  N    ��  N   �  	G   B� 
  L  0      s    v	  U     �  �  	  =  N   �f  �   M
  pmoc5  stib	  ltuo|  tolp 	  �(  b   "�  �  �  %  <�  x >)   len ?0  *� @   %  B�  	�    `�  �    G   G     U    �  �  q    G   3  G   G   U    �  @  F  [  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  �  ()  �3  0R   �U   8�  ��  @ #  �  �  �[  	�  �       G   .  U   .   s  �  A  G  R  s   �  ?_  e  z  s    @    �  Y�  �  G   �  s  @   U    s  ��  �  G   �  s  �     W  0�6  �  �f   e� �  �� �R  �� �z  �� ��   �� �4  ( �'  ��  �  �  ,G   N   	��	  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �   �  �%6  '  7p8F            ��	  R�  77  � � u8F     �  U�U  �  7  08F     7       �D
   R�  !7  ,� *� !>8F     �  U   "�<  �J  p7F     �       �9  #Jy  �   [� O� #OF  � �	  � � $�� �  P� J� %�7F     �  �
  U�TT	PJ      %�7F     �  �
  Uv T0Q2 %�7F     �    Uv  %�7F     �  $  Uv T0Q0 !8F     �  Uv   &b �@   �6F     V       ��  #Jy  �&  �� �� #x  �&@   "� � #B� �&  �� �� #.� �&@   K� =� $�� �  � � '7F     �  �  U�QT1Q�R !*7F     �  U| Q0  (�a ��6F     &       �>  #Jy  �$  8� 2� )�6F     �   (b }P7F            ��  #R�  }7  �� �� #��  ~U   ŷ �� X7F     �  U�T  &�a cU   `7F            �)  #R�  c7  � �� #f;  d-   ?� ;� #6^  e-   |� x� #��  fU   �� �� k7F     �  U�RT�Q  &�a EU   @7F            ��  #R�  E7  �� � #�  F-   3� /� H7F     �  U�T  *�N �N @*wa wa A*�a �a [*�a �a �*b b �*�a �a Y*�a �a �*�6  �6  B M0   �  �  hb $"  �8F     ]      _i X  ^� �@   �i int �i {S @�   g
  �       	4   v  #	4   �  &	4   |
  )	4    h  ,	4   (�  -	4   0�	  2G   8�  5G   < �   �  	�   �
  8"W   
  K  �   
�  L  
�  M  S  -  �  >   G   �  B"P  V     ��  R   �U    �� ��  �N ��  �6  ��   �  Y�  �  U   �  D  -      n�  �  �  D  U    �  ��  �  U     D  -   -   U    �  �"  "  �   PJ�  2�  L   �  M@   pos N@   �  P�  SF  Q�   �1 R�  (=9 S,  0R�  UD  8y�  V  @�� W  H �  ��  �\ �-   m  �U    o  ��  �  ��    @       @     @    %  �  2  9  ?  J       :-   �  Jz  x LJ   y MJ   )  OV  	z  B   s�  M   uJ   }  uJ  V  vJ  /  vJ   t
  x�  �J  N   �"  �@   �\  0  35  G5  8  >  �[  F;   k	  (�  �  N    ��  N   �  	G   B� 
  L  0    %  s  %  v	  U     �  "  	�  �  (N  �  P)   Z�  Q)  �  S  s  T�   [  U  ?1  WG     z  )    Y�  �  =  N   �s  �   M
  pmoc5  stib	  ltuo|  tolp 	  �5  b   "�  �  �  %  <�  x >)   len ?0  *� @%   %  B�  	�    `�  �    G   G     U    �  �  q!  '  G   @  G   G   U    �  M  S  h  G   G   U    �  `��  �  ��   �% ��  ?1  �G   �&  ��  !  ��   I  �  ()  �@  0R   �U   8�  ��  @ �    �  �h  	  �   !  '  G   ;  U   ;   �  �  N  T  _  �   �  ?l  r  �  �    @    �  Y�  �  G   �  �  @   U    s  ��  �  G   �  �  �     W  0�C  �  �s   e� �  �� �_  �� ��  �� ��   �� �A  ( �'  ��  �!  l%  �  �h  �  -  �%  	o  {  �  ��   	�  �
  �)  �  �0  �  �G   
  �N   �  �-   \#  �@   �   -   �  ,G   \&  7U   �0  D4   b   �V	  xx ��   xy ��  yx ��  yy ��   a  �	  	V	  z'  ��	  m  ��   ss  ��   �  �h	    ��	  �	  �	  U    �  ��	  �U  �U      ��	   %  ��	  �  $
  	
  �   B
  �� "�	   �@ #�	  �U  $U    �  7m
  �; 9�	   ��  :�	   L  <B
  N   ��  �     �    $  K  �%  �%  ,#  �  	   
�$  e#  �  �  [%  A#  z"  6  �  �  �   �"  !Y  "�  #�#  $_"  %�  &�"  'H!  (�  0v  1�  @  Al  Q�   R7  S�$  T�#  U  V   W�  XR  `	  aa  b�"  c�'  p�  ��  �	  ��  �M  ��  �v  ��  �'  �H%  �  �e!  ��  �'%  ��   ��  ��  ��$  ��  �g  �  �P  ��  ��  ��  �  ��$  ��&  �N  ��   �  ��  �;$  ��  �#  ��"  ��  �G  ��  �0  �1  �P  �C&  �:  �_  �A  �^  � �
  @=<  ��  ?J   �  @J  ~  BJ  �  CJ  �  DJ   5  FJ  (B  GJ  0�  HJ  8 �	  J�  
   s�  �  u�   ��  v�  �  xJ  �
  zJ  (  {J   �  }I  �  �#�  �  k  `	�m  R�  	�D   (  	��  |  	��  �  	��  �  	��  �  	�v!  v  	�m
  �  	�  (�%  	�m  07&  	��!  8G   	��  X �  �"z  �  h  	�  �M 	]!   k  	�  R�  	D   �  �"�  �  %  8	;  �� 	=c!   �M 	>^    	?m
   r$  	@�  0 5  �$   &  %  �	�  �� 	c!   �M 	p!  �  	s   �  	�  (�� 	
�  h�� 	�  p�� 	�  x K  � �  �  �  �,k  �   .�   �  /�  O  1�  C  2�  �  4�   d> 6�  (A  7�  0T  9�  8  :�  @�  <�  H�  =�  PE-  ?�	  X�!  D�  h:  F�  �  G�  ��  H�  ��  I�  ��  K�  �  L�  �U  N�  ��  O�  �)�  Q�  ��  Rk  ��� S"  �K1 W�  �R�  XD  �Jy  Y  �%  [m
  ��	  ]�	  �    ^U   ��8  `N  � L   x  ~    X��  �  ��   E-  ��	  N ��  �8  ��  P �  *%�  �  �  0t"  k  v�   �  w�  �@ x�  ݖ y�  E-  z�	   N |<  0�  }�  pR  ~�  x�  z  �ߣ  �s  ��I ��  ��  ��  �h  ��  ��S  �"  �4  ��  �8  ��  �  �U    �  �-   �  �J  o  �J  �L �U    �8  �,  ( �
  L#/  5  W  H|  �  J�   = KA    L�  d  M�   �  N   �A  �   �  bmys=  cinu�  sijsw    bgO  5gibp  snawM  ahoj�    bg�  sijs�    bgq  5gib�  snaw�	  ahoj  BODA4   EBDA�	  CBDA  1tal�  2tal   nmra �	  |  #   g)[  a  �   �	��  =  	�V	   L  	�z   $  	��  0�  	��  8m  	�#W!  h�  	�\  pآ  	�7  tG   	��  x �  �  "  �
  �)�    �   H	�>  �  	�U    "  	��  �!  	��   ~	  8f�  �
  h�   (  i�  �� k�  �� l�    nJ  �  oJ   �  pJ  (�  qJ  0 y  s>    �$�  �  �  0
',  �N  
)�   ?1  
*�  }0  
+�  i/  
,�  � 
-V	   �  �)9  ?     H	��  ��  	��   ?1  	��  (  	�P  4  	�V	  \  	�z  0  	�U   @ +!  �  tag �   �U  �   �  �  �  `  N   
  w%   }#  �&  h  �  &     
�  E   9
z  � ;
   ��  <
�  �  =
�  �  >
�  �#  ?
�   �  L
(�  %  �  N   ��  :   �   ^$  1  �!  �!   :  ��  �  ��  �#  ��  �  �  �  m   I$  �      m   �&  �(  .  �  B  m  B   �   �!  H��  �  ��   S"  ��     ��  �"  ��  �  ��   ;  ��  (%  ��  0�   ��  8��  �  @ �  R  �H  x  =�	  H  E#�  	�  �  @Jq  �  L�   �  Ms  �� O�  .� P�  �  Qc   �  R  (�!  S;  08'  T�  8   W!}  �  -  (l�  k  n�   �M o�  ߣ  ps  �  qz   �  k  )�  �  �  �  q  �   w   .�      q   �  1     5  q  5  /   c	  K  6G  M  ]  q  ]   �  �  :o  u  �  �  q  q   �  >�  "  Y�  �  �  �    �  �  /   �  _�  �  �  �    �  5  /   $  f        �  ]   �  l(  .  �  G    �  �   #  x��  �� � �   �  � s  H  � �  P�  � �  X9!  � �  `l� �   h  � �  p C    �G  �  H
2  �S  
4"   �  
5  (  
6  04  
7�  88  
8�  @ �  
:�  �  �
=�  R�  
?D   �  
@�  n  
A�  �  
B�  1$  
CP  2�  
E  �� 
F  `�L 
HU   � �  
J�    P   �  �  �  �    �  �  �  �   �  &�  �  �  �   �%  *  	  �    k   �%  -$  *  5  k   {  1A  G  �  V  �   �  4b  h  s  �   l  8  �  �  �  k  z   �  <�  �  �  �  k  �   �  @�  �  �  �  �  k  �  7   �  G�    �    �  �  �     �'  N+  1  �  E  �     �  SQ  W  �  z  �  �  �  7  z   �  &  ��^  �� ��   i'  ��  H   ��  P  ��  X�A ��  `Y ��  h�#  ��  p�  �  x�  �5  �  �V  ���  ��  �U�  ��  ��!  �  ���  �E  ��  �s  �&  ��  � �&  �j  �  �  0t�  �  v�   a   w�  �'  x�  !  y�  �#  z�   �  {�  ( �  }p  �  U'�  �  m  D   t9   �  v�   A  w�  �  x�  &  y�   !  {�  �  �Q   W   �  p   �  �  p    �	  �  ��   �   �   �  p    �'  ��   �   �  �   �  �  P  �    9   �!  !  ��  )E    ��  )v   �  )�    }  �   	!  O  ;D!  _� =%D!   ݰ  >%�   !  �  @!  J!  �  �  	�  �  m  �!  @    �  �!  @     �  	�%C  !�b �  (                                        "�9 ,�  @@F     F       �H"  #k  ,�  r� l� #�I -H"  ƹ �� $R�  /D  )� %� %Z@F     0   �  "(c �  �?F     �       ��"  # *�  f� `� & � '�I �  �@$� �  �� �� (�/  �?F       P� �"  )�/  ٺ ׺  *@F     �-  +Ts�+Qw    "R ��  �:F     �      �4'  #k  �(�  � �� #�% �(�  �� �� #�  �(H"  0� $� #P� �(�  ż �� '� ��  �L$R�  �D  � y� ,s  4'  ֽ ̽ ,t 4'  S� E� -p� '$  ,pad �  � � $hc �  t� h� .lc *�  $ �  � 
� *�;F     "0  +T1+Y�L  -�� �$  ,i K�  {� q� &� ,ss R4'  �� �� ,tt S4'  w� g� ,j T�  1� #� /`>F     `       �$  ,val Z�  �� ��  0 ?F     (       ,val n�  � �    /�=F     P       /%  $��  ��  H� F� ,i ��  q� k� *�=F     .0  +T| +Q~   - � �%  ,i ��  �� �� &`� ,ss �4'  A� 7� ,tt �4'  �� �� ,j ��  |� n� /p=F     1       �%  ,val ��  !� �  0(?F     (       ,val ��  [� W�    -�� d&  ,i ��  �� �� &� ,ss �4'  � �� ,tt �4'  �� �� ,j ��  U� M� 0<F            ,val ��  �� ��    0�<F     �       ,i ��  "� � 0�<F     �       ,ss �4'  u� m� ,tt �4'  �� �� ,j ��  c� a� 1:'  �<F      �<F     U       �)L'  �� �� 0�<F     U       2Y'  �� �� 2d'  �� ��      o  3c �o  p'  4#c �8�  5a ��  5l ��   "�b (�  �@F     M      �m,  #k  (#�  r� T� #�I )#H"  �� �� #^b *#J  �� �� #�b +#J  y� m� $� -�  � � ,p .  �� �� ,i /�  �� �� ,x /�  �� �� $�  /�  � � ,y 0�  �� �� $Pb 1�  � 	� $yc 1�  �� �� -ж )  6tmp K�  ��(�/  �AF       � O	�(  )�/  �� ��  7BF     �"  �(  +Q��+R1 **BF     �!  +Uv +Ts   -�� ")  ,tmp �%  ;� 5�  /�AF     3       K)  ,q �  �� ��  8m,  gBF       @� k)�,  �� �� )�,  �� w� )�,  Y� ?� )~,  �� j� &@� 9�,  ��2�,  � q� 2�,  ,� � 2�,  (�  � 2�,  �� �� 2�,  "� � 2�,  �� �� :-  �BF            �*  2-  �� �� 2-  �� �� ;-  �BF     _       2 -  � � 2,-  p� l� 28-  �� �� 2D-  �� �� 2P-  7� /� ;\-  $CF     "       2]-  �� �� *DCF     90  +T0    <�-  0� c+  =�-  2�-  �� �� 2�-  A� 3� 2�-  �� �� 2�-  >� :� 7�DF     .0  +  +U~ +Q��~ 7�DF     90  A+  +U~ | "+T0+Q�� *�DF     90  +U~ +T0+Q��~  :l-  _FF     v       ,  =q-  2}-  �� ~� 2�-  �� �� 2�-  �� �� 2�-  �� �� 7pFF     90  �+  +Uv +T0+Q��~ 7�FF     .0  �+  +Us +Q��~ *�FF     90  +Us | "+T0+Q~   7BDF     "0  T,  +U��~+T ����+Q0+X0+Y�� *EF     0  +U��~    >&b ��  �-  ?R�  �(D  ?�I �(H"  ?`c �(�  ?Xc �(�  @� ��  @�  �N   @Nc �N   Abpp ��  @��  ��  @�  ��  @B� �  Bl-  @Q ��  @Ub ��  C@+ �4'  Aend �4'  @�� ��  @� ��  @.� ��  C@x� �4'     B�-  Alen ��  Ain �  Aout �  @�� �  @� �N    C5len �  5in   5out   .��   .� N     D�b 6�  �8F     �      ��/  Ek  6%�  � � E�% 7%�  �� �� E�  8%H"  �� w� FR�  :D  ;� 5� G� ;�  ��F�  =�  �� �� F�  >�  I� C� F�b @�  �� �� F>b @ �  �� �� -� /  Flc a�  b� Z� F�b b�  �� �� **:F     "0  +T1+R} +Y��  -@� �/  Hp q  � � /�9F     G       �/  Hi }�  1� +� Hs ~4'  �� z� Ht 4'  �� �� *�9F     .0  +Qs   *�:F     .0  +Q}   *}:F     D0  +T} +Q��  I@c ,�/  ?�O  ,H"   J�A "�/  ?�O  "H"   K�/  �8F            �0  L�/  U MF\  F\  �M�[  �[  �N�D  �D   Ni0  _0   MkA  kA  { N    ��  @RF     0SF     z src/gfx/sse2.asm NASM 2.14.02 �@RF              �    ��  �c �c ~c �UF     >       �z �  �  �i -  N   �i �  -  int X  7  B   �c �UF     >       ��c q   �`�c &q   �X}0  5q   �Pi/  Dq   �H d Sq   �@�c bq   ��  �    �  �n �v ~c `�         :{ X  ^� �<   �i S  �
  �  int V   �o V   -  �i u   �  �n 	)   �  -  
<   �  �  
�<   7  �   �  4�   �  �   �   �   	<    
�n -  �n @  �n �q   $  �   �g <l 4  �      �w +�v !  �r ,�p &  �m /sv V   �  V   �  �   o 'm b   �p !�d Nr +k �     gh }q V   �  �   0    Nd \j V   �  0   �   �d k V     std    9t �  �\ �  �l   �l =g ,  P  V  �   �g t ,  n  t  �   T   v       �v �  �\ �  �l   �g �o �  �  �  �   �g Vl �  �  �  �   T   v    �  �s �-  �\ ��  T V   �O  >    ;s �Z  �\ ��  T V   �O  D    v ��q �  v ��e �   t   �d   �  6h �  �   frg 	�
  !/g �  "[r  �  #�t  �  $�q 7   %mi V   ,  &�r  &�( 'hex  (Mq `  )�h {k  *ݰ  |V   +�h ~�q I  O     �h h _    V     ,�s  u �  �  '   ,�s p �  �  '  �   ,�s �v �  �  '  2   ,�s *o �  �  '  8   ,�s *gs �    '  >   ,�s 0dr   &  '  D   ,�s 8�m ;  F  '  V    -Gp =�w J  _  j  '     -�s Qr   �  �  P   -�s T�i   �  �  '   -]h X%d   �  �  P   -p \Xw 2  �  �  P   -p `�k V  �    '   -�o d�g \    $  '   +�� ��s 8  >  '   .wq �   .�r �  T V      ,s 2L  +,s 3�s �  �  b   #m 6Rf e  �  �  b  �   .(m <�   .�m =V   .H� >  .�t ?  .v @  .�r A  .;f B  .�u C  /+s �n (  3  b  V    0,s  i @  b  �    e  
/f J  �f Nqw �  P R  T u   �  u     V   V   V   �    !v xi �  P R  T u   �  u   V   V   V   �    1�d ��m T u   F R  u   e  �    !Dq 
  "�g   2`d Xt .
  +s ECo G  R  �  �    j �	�	  +j �e s  ~  �  �   3j ig �  �  �  �   4Gp 	�j �  �  �  �  �   +j �f �  �  �  V    Cr "	�r �  �  	  �     + i '�h 	  !	  �  �    + i 1~j 5	  @	  �     5#s >�   5A� ?�   5�� @
0   �5m A  �*q 	{l �  �	  �	  T u   �  u    6�m 	3m �  �	  T   �      R  �g H�o R  �	  �	  �   ,�l Mj 
  
  �     5cg Q�    7�n �   8�! <   � t 
*w 2  T
  T V   2  2   nk �Qp {
  F R  u   e  �   nk �Au �
  F R    e  �   9�p 3�k �
  T u   F R  �  �   :'i 3Ee T   F R  �  �    ;�  	J     �     ;�  	8�K           '  <]   =V   <`  =  <  `  <V   V   e  b  >Ln   >uh :  �i Jf ;  	"J     �   &  �  R  �  <�	  <R  ?Z  ?l  @	  �  x`F     �       �	  A�  �  �hBs '�   �d C.
  O`F     (       �F  T V   Ba 2  �hBb #2  �` D]  �^F     �      �r  P R  T u   EH N�  ��E��  N$u   ��Es N1  ��E�s N?V   ��E��  OV   ��EH� OV   ��EZX  O#�   ��F]� P  �XFB� Sr  ��Gk TV   ��H�_F     E       /  Gi aV   �l H�_F     -       R  Gi dV   �h I`F     0       Gi fV   �d  �   �  	<    D�  [^F     U       �  P R  T u   EH x�  �hE��  x!u   �dE�s x-V   �`E��  x8V   �\EH� yV   �XEZX  y�   �TJK�f {	u     D�  �]F     �       �k  T u   F R  Eݰ  �u   �lBfo �/e  �`EH �6�  �X @!	  �  �\F     �       ��  A�  �  �hBstr 1  �` DT
  �\F     J       ��  F R  Eݰ  �!u   �LBfo �8e  �@EH �?�  �� D{
  z\F     *       �G  F R  Eݰ  �   �hBfo �7e  �`EH �>�  �X @�	  f  T\F     &       ��  A�  �  �hE�d M  �` <|   D�
  \F     C       ��  T u   F R  Lݰ  3�  �HLH 3!�  �@ <  D�
  �[F     E       �"  T   F R  Lݰ  3�  �HLH 3!�  �@ M_  0  F  N�  �  O$s �   P"  �u i  �[F     4       �z  Q0  �hQ9  �` MO  �  �  N�  "  N0  ]    Pz  Gk �  �[F            ��  Q�  �h M5  �  �  N�  "   P�  �t   �[F            �  Q�  �h @�  *  T[F     ,       �?  A�  �  �hR  �  @x	  e  ,[F     (       ��  T u   A�  �  �hEݰ  u   �d @�	  �  [F     )       ��  T   A�  �  �hEݰ    �` M�  �  �  N�  �  N0  ]    P�  �t   �ZF            �  Q�  �h @�	  /  �ZF     )       �<  A�  �  �` M�  J  `  N�  -  O�L *>   S<  [q �  vZF     V       ��  QJ  �hQS  �` M&  �  �  N�  -  N0  ]    S�  r �  ZZF            ��  Q�  �h Mk  �  �  N�  -   S�  �d   6ZF     #       �%  Q�  �h TDw F�t YF            �U	k AV   YF            �V�w 9�k �WF           ��  E�f 9&  ��~E�� 9=  ��~E+ 9Pu   ��~E8u :  ��~ �   )   D`  �WF     c       �7  E}m /V   �\E�u /'�  �PE�q /3�  �HF�u 0�   �hFFd 0�   �` D�  WWF     ;       �q  Fp (�   �`Gpid +	b   �l W�  EWF            �D�  WF     6       ��  Bmsg    �h C�  �VF            ��  Em  �   �hE�  *0   �` �   D�  qVF     �       �@  E�  0   �hEm  ,�  �`Xw P  	�J      �   P  	<    @  D�  ;VF     6       ��  E% V   �l Y  2�  �  N�  h  N0  ]    S�  �o �  ZF            ��  Q�  �h <L  Y3  2�  �  N�  h  �   S�  �e   �YF     �       �*  Q�  �hQ�  �` Mr  8  B  N�  h   S*  w e  &YF     \       �n  Q8  �h Z6r kv �   YF            ��  E�  #0   �hBp /�   �` &E �
   %   ȑ  �n �x ~c ,aF     A       ނ X  �i S  �
  �  std  �  9t �   �\ �  �l �  �l =g s   �   �   	�   �g t s   �   �   	�   
T �  v �    Y   �v B  �\ �  �l �  �g �o �       	�   �g Vl �   ,  2  	�   
T �  v �   �   �s �t  �\ ��  
T   �O  D    ;s ��  �\ ��  
T   �O  J    v ��q �  v ��e �   t �  �d f   �   6h �   B  �i �  �  �  -  int   frg 	�  /g +  [r  4  �t  `  �q 7   Mq �  �h {�  ݰ  |  �h ~�q �  �  	,   �h h �  	,  	    �s  u �  �  	2   �s p �  �  	2  +   �s �v     	2  8   �s *o ,  7  	2  >   �s *gs L  W  	2  D   �s 0dr l  w  	2  J   �s 8�m �  �  	2  	   Gp =�w P  �  �  	2  `   �s Qr �  �  �  	V   �s T�i �  �  �  	2   ]h X%d �      	V   p \Xw 8  1  7  	V   p `�k \  P  V  	2   �o d�g b  o  u  	2   �� ��s �  �  	2    wq �m    �r ��  
T    `  !/f JDq 
�  �g �  `d i  s E�x �    	d  �   "j �g Hx   !  '  	d   �l Mox <  G  	d     #cg Q�   $�n �  %�! 4   � &Xt s ECo �  �  	|  �   "j �g H�o �  �  �  	|   �l Mj �  �  	|     #cg Q�   $�n �  %�! 4   �  '9  	�J         �    'R  	@�K     m  `  (  )  (�  )`  (`  �  (    *Ln T  *uh �  �i Jf '�  	�J     +�n N  x �  ,x 
Xx �  �  	N   �g y �  	N      �n -  ,�n �q     	Y   �g <l !  	Y      -�w +�v �  -�r ,�p i   �  N  �  Y  �  .-  $	P�K     i  .=  	%	Q�K     /�  /�  0  �  LaF     !       ��  1�  _  �h2�d )  �` 0�  �  ,aF            �  1�  T  �h2�d (  �` &E �
   q   ��  �n ]} ~c  �         � X  ^� �<   �i S  �
  �  std  �  9t �   �\ �  �l �  �l =g {   �   �   	�   �g t {   �   �   	�   
T �  v �    a   �v J  �\ �  �l �  �g �o �       	�   �g Vl �   4  :  	�   
T �  v �   �   �s �|  �\ ��  
T "  �O  !    ;s ��  �\ ��  
T "  �O  '    v ��q �  v ��e �   t �  �d n   �   6h �   J  �i �  �  �  �  -  int "  frg 	�  /g :  [r  C  �t 	 o  �q 	7�   mi "  ,�  �r  �( hex  Mq �  �h {�  ݰ  |"  �h ~�q �  �  	�    �h h �  	�  	"    !�s  u     	
   !�s p    +  	
  ":   !�s �v @  K  	
  "   !�s *o `  k  	
  "   !�s *gs �  �  	
  "!   !�s 0dr �  �  	
  "'   !�s 8�m �  �  	
  	"   #Gp =�w -  �  �  	
  "�   #�s Qr �      	3   #�s T�i �  '  -  	
   #]h X%d �  F  L  	3   #p \Xw   e  k  	3   #p `�k 9  �  �  	
   #�o d�g ?  �  �  	
   �� ��s �  �  	
   $wq ��   $�r ��  
T "   �  ,s 2�  ,s 3�s     	E   #m 6Rf �  )  4  	E  "o   $(m <o   $�m ="  $H� >�  $�t ?�  $v @�  $�r A�  $;f B�  $�u C�  %+s �n �  �  	E  	"   &,s  i �  	E  "�    �  '/f J9  (�� Nm{ $  
P   
T �  "�  "�  "�  ""  ""  ""  "�   (�f Nqw f  
P �	  
T �  "^  "�  "�  ""  ""  ""  "�   (B~ xR �  
P   
T �  "�  "�  ""  ""  ""  "�   (!v xi �  
P �	  
T �  "^  "�  ""  ""  ""  "�   (*y ��   
T �  
F   "�  "�  "�   )�d ��m 
T �  
F �	  "�  "�  "^    Dq 
9  �g B  `d [	  s E�x t    	t  "�   j �	�  j | �  �  	  "t   *j *{ �  �  	  "�   +Gp 	@� �  �  �  	  "�   j      	  	"   Cr "	�z �  $  /  	  "9    i '�} C  N  	  "�    i 1Wz b  m  	  "�   ,#s >t   ,A� ?d  ,�� @
0   �,m A�  �*q 	z �  �  �  
T �  	  "�   -�m 	�~ �  �  
T �  	  "�      �g Hx   	  	  	t   !�l Mox .	  9	  	t  "�   ,cg Q�   .�n �  /�! <   � Xt c  s ECo |	  �	  	B  "�   j �	�
  j �e �	  �	  	M  "B   *j ig �	  �	  	M  "X   +Gp 	�j ^  �	  �	  	M  "X   j �f 	
  
  	M  	"   Cr "	�r ^  ,
  7
  	M  "9    i '�h K
  V
  	M  "�    i 1~j j
  u
  	M  "�   ,#s >B   ,A� ?d  ,�� @
0   �,m A�  �*q 	{l ^  �
  �
  
T �  	M  "�   -�m 	3m ^  �
  
T �  	M  "�    �	  �g H�o �	    !  	B   !�l Mj 6  A  	B  "�   ,cg Q�   .�n �  /�! <   � 0t 
*w   �  
T "  "  "   (�~ ��| �  
F   "�  "�  "�   (�~ ��} �  
F   "�  "�  "�   (nk �Qp �  
F �	  "�  "�  "^   (nk �Au %  
F �	  "�  "�  "^   1�{ 3�y O  
T �  
F   "|  "�   1xy 3} y  
T �  
F   "�  "�   1�p 3�k �  
T �  
F �	  "|  "^   2'i 3Ee 
T �  
F �	  "�  "^    3H  	�J     �  �  �  �  3a  	H�K     �  �  �  
  4)  5"  4�  5�  4�  �  4"  "  �  E  6Ln \  6uh �  �i Jf 3G  	�J     '�n 
6  x 
�  7x 

Xx �  �  	6    �g 
y �  	6  "�    �n 
  7�n 
�q �  �  	<    �g 
<l 	  	<  "�    8�w 
+�v S  8�r 
,�p [	   �  �  [	  B  �	  M  4�
  4�	  9�  t  :<    S  t      4�  4  ;�  ;�  </  �  �hF     �       ��  =�  �  �h>s '�  �d <7
  �  x`F     �       �  =�  S  �h>s '�  �d ?c  O`F     (       �O  
T "  >a   �h>b #  �` @�  RgF     �      �{  
P   
T �  AH N�  ��A��  N$�  ��As N1�  ��A�s N?"  ��A��  O"  ��AH� O"  ��AZX  O#�  ��B]� P�  �XBB� S{  ��Ck T"  ��DBhF     E       8  Ci a"  �l D�hF     -       [  Ci d"  �h E�hF     0       Ci f"  �d  9�  �  :<    @$  �^F     �      ��  
P �	  
T �  AH N^  ��A��  N$�  ��As N1�  ��A�s N?"  ��A��  O"  ��AH� O"  ��AZX  O#�  ��B]� P�  �XBB� S{  ��Ck T"  ��D�_F     E       t  Ci a"  �l D�_F     -       �  Ci d"  �h E`F     0       Ci f"  �d  @f  �fF     U       �I  
P   
T �  AH x�  �hA��  x!�  �dA�s x-"  �`A��  x8"  �\AH� y"  �XAZX  y�  �TFG�f {	�    @�  [^F     U       ��  
P �	  
T �  AH x^  �hA��  x!�  �dA�s x-"  �`A��  x8"  �\AH� y"  �XAZX  y�  �TFG�f {	�    @�  afF     �       �2  
T �  
F   Aݰ  ��  �l>fo �/�  �`AH �6�  �X <N  Q  �eF     �       �m  =�  �  �h>str 1�  �` @  �]F     �       ��  
T �  
F �	  Aݰ  ��  �l>fo �/�  �`AH �6^  �X <V
  �  �\F     �       ��  =�  S  �h>str 1�  �` @�  FeF     J       �P  
F   Aݰ  �!�  �L>fo �8�  �@AH �?�  �� @�  eF     *       ��  
F   Aݰ  � �  �h>fo �7�  �`AH �>�  �X @�  �\F     J       ��  
F �	  Aݰ  �!�  �L>fo �8�  �@AH �?^  �� @�  z\F     *       �A  
F �	  Aݰ  � �  �h>fo �7�  �`AH �>^  �X <	  `  �dF     &       �|  =�  z  �hA�d M�  �` 4�  @%  �dF     C       ��  
T �  
F   Hݰ  3|  �HHH 3!�  �@ 4�  @O  ndF     E       �  
T �  
F   Hݰ  3�  �HHH 3!�  �@ I�  *  @  J�  �  K$s t   L  �z c  :dF     4       �t  M*  �hM3  �` <!  �  T\F     &       ��  =�  H  �hA�d M�  �` @y  \F     C       ��  
T �  
F �	  Hݰ  3|  �HHH 3!^  �@ @�  �[F     E       �C  
T �  
F �	  Hݰ  3�  �HHH 3!^  �@ I�	  Q  g  J�  S  K$s B   LC  �u �  �[F     4       ��  MQ  �hMZ  �` I�  �  �  J�    J0  )   L�  Gk �  �[F            ��  M�  �h I�  �     J�     L�  �t #  �[F            �,  M�  �h <  K  dF     ,       �`  =�  �  �hN9  �  <�  �  �cF     (       ��  
T �  =�  �  �hAݰ  �  �d <�  �  �cF     )       ��  
T �  =�  �  �hAݰ  �  �` I�  �    J�  �  J0  )   L�  _| (  �cF            �1  M�  �h <�  P  �cF     )       �]  =�  z  �` <
  |  T[F     ,       ��  =�  S  �hN9  �  <�
  �  ,[F     (       ��  
T �  =�  S  �hAݰ  �  �d <�
  �  [F     )       �  
T �  =�  S  �hAݰ  �  �` I�	  #  6  J�  S  J0  )   L  �t Y  �ZF            �b  M#  �h <  �  �ZF     )       ��  =�  H  �` Ik  �  �  J�    K�L *!   O�  [q �  vZF     V       ��  M�  �hM�  �` I�  �    J�    J0  )   O�  r *  ZZF            �3  M�  �h I�  A  K  J�     O3  �d n  6ZF     #       �w  MA  �h P�} ybF           ��  A�f  �  ��~A�� 7�  ��~A+ J�  ��~A8u �  ��~ P2� maF           �5  A�f  �  ��~A�� 7�  ��~A+ J�  ��~A8u �  ��~ Q�  2F  Y  J�  K  J0  )   O5  �o |  ZF            ��  MF  �h 4�  Q�  2�  �  J�  K  "�   O�  �e �  �YF     �       ��  M�  �hM�  �` I�  �  �  J�  K   O�  w   &YF     \       �#  M�  �h R6r kv   YF            �f  A�  #0   �h>p /  �` &E �
   �   ��  �n ـ ~c �iF     �       � ^� �9   �i �O   -   �jF     <       ��   s  �   �Xlen !	-   �h�jF     &       i "-   �`  �   �  	�   �Z a  EjF     �       �a  
S a  �Hsrc 'h  �@
�  3-   ��� t  �Xπ t  �PojF     4       A  i -   �h �jF     E       i -   �`  a  s  h  �   �D  a  �iF     Z       �  
S c  �Hsrc <n  �@
�  H-   ��� t  �`π t  �XjF     4       i -   �h  i0  a  �iF     F       ��  
S a  �Xc �  �T
�  (-   �H� t  �`�iF     )       i -   �h  int  *    ��  �� *kF     {kF     � ~c 2� ��Z   ��  e�n �� ~c p�         � @�� 	5   fint 5   @�� M   S   �  S   @! M   �  k   �  "t  �   �i �   �i �   �  -  X  "�  ��   "g  ~   �   "�  4�   �   "^� ��   �   "*� 	  g  AU� 1  � 5    /rem 5    "V� 	  Aa� e  � �    /rem �    "b� =  A�� �  � �   /rem �   S  "�� q  hfrg �  i�� �	�  On <   pOm <   �P>� �   ߰�jmsb �      �P�� �   ����� 7� '  -  �   ߢ  �� A  L  �  �     �g � �   d  j  �   k_st >�   l�� ?5   �	 B/g �  Q[r  �  m�t  �  n�q 7�   7mi 5   ,�  %�r  %�( Rhex  SMq 3  o�h {>  pݰ  |5   �h ~�q   "  �   C�h h 2  �  5     �s  u S  Y  �   �s p n  y  �  �   �s �v �  �  �  �   �s *o �  �  �  �   �s *gs �  �  �  �   �s 0dr �  �  �     �s 8�m     �  5    &Gp =�w   2  =  �  �   &�s Qr �  V  \     &�s T�i �  u  {  �   &]h X%d �  �  �     &p \Xw �  �  �     &p `�k   �  �  �   &�o d�g   �  �  �   �� ��s     �   wq ��   �r ��  T 5    �  ,s 2  ,s 3�s Y  _       #m 6Rf 8  w  �     �   (m <�   �m =5   H� >�  �t ?�  v @�  �r A�  ;f B�  �u C�  q+s �n �       5    r,s  i      =X    8  D/f J�  8�� N߫ r  P    T �   2#  �   �  5   5   5   S    8C� xZ� �  P    T �   2#  �   5   5   5   S    s�� �� T �   F    �   8  2#    BDq 

�  Q�g 
�  `d 
�  s 
E�x      #  �   j �
	�  j 
| A  L  !#  #   ,j 
*{ `  k  !#  ,#   -Gp 
	@� 2#  �  �  !#  ,#   j 
 �  �  !#  5     Cr 
"	�z 2#  �  �  !#  �    i 
'�} �  �  !#  S     i 
1Wz     !#  �   3#s 
>#   3A� 
?�"  3�� 
@
�   �3m 
A�  � M� 
	�� 2#  e  p  T   !#     T�m 
	�~ 2#  �  T �  !#  �        �g 
Hx    �  �  #   �l 
Mox �  �  #  �   3cg 
Q�   4�n �  t�! �   � UXt B�� 		  uW� 
	   D`� 	  E<	  V� �    F)	  7>� 5   i	  %�r  Rred %d�  l� 0!
  l� � �	  �	  6!   ,l� � �	  �	  6!  A!   -Gp ;� G!  �	  �	  6!  A!   S�    �    ��   )�    �� !   � "D	  ( i	  �� %r
  �� '{� �  T
  T f  e#   WJ� ';� �  T �  N#    f� 5  Xh 8`� 6!  �
  N#   O� =t� N#  �
  N#   �� BͰ N#  �
  N#   n� E� N#  �
  N#   )� I�� N#     N#   �� L7� N#    N#    �� PE� N#  2  8  �#   9#� U�� �  S  N#   9�� Z؟ �  n  N#   � d� �  �  �#   ,� g� �  �  �#  �#   -Gp i;� �#  �  �  �#  �#    N� o�� N#  �  �  �#   � |\� �    �#  N#   c� ���   -  �#  N#  N#   �� ��� B  R  �#  N#  N#   
� �6� g  r  �#  N#   '�� #� �  �  �#  N#   <� � �  �  �#  N#  N#   �� D� �  �  �#  N#  N#   �� x)� �  �  �#  N#   �� �$�      �#  N#   /� �� 6  A  �#  N#   '� u� V  a  �#  N#   ',� #E� v  �  �#  N#   00� 0�� �  �  �  �#   00� 94� �  �  �  �#  N#    �#  �#   :�� �   D 	  T �  ;� �Z  A &
   r
  v� ��  (��  (�  (�-  (��
  (��
  (�  Gr
   '�� �\� h  s  �#  �   '\+  ��� �  �  �#  N#   :�� ��  T �  ;� �Z  L �  A &
   _� 5T  Xh 8� 6!  �  e#   O� =� e#    e#   �� B� e#    e#   n� E2� e#  6  e#   )� I�� e#  P  e#   �� L� e#  j  e#    �� PK� e#  �  �  �#   9#� U� �  �  e#   9�� Zk� �  �  e#   � dg� �  �  �#   ,� g4� �  �  �#  �#   -Gp iI� �#      �#  �#    N� o�� e#  2  8  �#   � |c� M  X  �#  e#   c� �)� m  }  �#  e#  e#   �� ��� �  �  �#  e#  e#   
� �� �  �  �#  e#   '�� U� �  �  �#  e#   <� �� �    �#  e#  e#   �� Dz�   .  �#  e#  e#   �� x�� D  O  �#  e#   �� �Z� e  p  �#  e#   /� �� �  �  �#  e#   '� ;� �  �  �#  e#   ',� #�� �  �  �#  e#   00� 0�� �  �  �  �#   00� 9�� �    %  �#  e#    �#  �#   :�� �   D Y  T f  ;� �Z  XA &
   �  wW� �(�8  (�X  (�}  (�  (�  (�j  G�   '�� �F� �  �  �#  �   '\+  �Q� �  �  �#  e#   :�� ��  T f  ;� �Z  XL �  A &
    E"  V� �    F  �� Y  xclz � 5   Q  �    T �    y"� �$"  7"� 5   ��  %�r  %l� %[�  g  � H�	a  � ��� �  �  N#  g  �   �    ,� �5� �  �  N#  Y#   -Gp �
�� _#  �  	  N#  Y#    Z� �δ �  !  ,  N#     � ��    ��   ss  ��   "� �   �  � ��	  G�   � �E� �  �  e#  �   �   5    ,� ��� �  �  e#  p#   -Gp �r� v#  �  �  e#  p#   �N  �<   Hٖ ��   LU� �|#  P.� �  X f  '� �	�  '� ��� ?  E  |#   ,'� �Ƈ Y  d  |#  �$   -Gp �Ⱥ �$  |  �  |#  �$   ʊ �|#      � �	�  T�g �a� �  �  �#  Y#  Y#    �0   �	  �0  ��� �  �  �#   � �	R!   x� �e#  � �   "�� �  �� �-� <  G  C#  �#   Y�� (z� \  g  C#  �#   zGp *� �#  �  �  C#  �#   &Wd ���   �  �  C#  �    0�6  L��   �  �  C#    �    �N ~�� �  �  C#     � �w�      C#    �    &Y� 1	�� �   9  ?  C#   {J� >
$                         @       H�� @ �   H�� A �    H� H�� �   �  �    r� W�� �   �  �    H�� j<   1� l�   �� o�� �  �  �    1o� |�   1�� �   |� ��    I<� �7� N#  4  ?  C#  �    Ia� �� e#  X  c  C#  5    IP� %j� N#  |  �  C#  �    '`� 7� �  �  C#   '� >� �  �  C#  N#   Э �
�#   A� �R!  "ۧ �'  @� ��  �� �	�    � �`$  (4� "  4v� R!   Y  }0� V  ;� X� K  V  8#  C#   0Wd [!�   p  {  8#  �    � _ʅ �  �  8#    �    �N c�� �  �  8#     0� gε   �  �  8#    �    ~�� lC#   4� "  4v� R!   JG� �+i	  J� �7Y  J� �7	  S#� �  0� �� V  \  p$   0� ׁ q  �  p$  	  "   0� I� �  �  p$  "   Y0� !�� �  �  p$  {$   0� #E� �  �  p$  �$   /� (�� �    p$  5    &Gp -
� �$    %  p$  4   7� 2�� :  @  p$   �� 8�� U  [  p$   &�� >U� �  t  z  p$   &<� Bn� �  �  �  p$  "   F� G	"   �� H�  4v� R!   4  t 
*w �  �  T 5   �  �   8�~ �|�   F    ]  8  2#   8�~ ��} ;  F    �  8  2#   Z� 34� e  T   F    >  2#   Zxy 3} �  T �  F    �>  2#   WU� 
�� �?  T �   �?  �?    �  !� )�� �  )p� �  ) � �  )&�   �  �  �   �  ��   o �
  ��  �std  �  9t �  1�\ �  "�l �   �l =g /  S  Y  �    �g t /  q  w  �   T �  [v �      �v �  1�\ �  "�l �   �g �o �  �  �  �    �g Vl �  �  �  �   T �  [v �   �  �s �0  1�\ ��  T 5   \�O  ]�    ;s �]  1�\ ��  T 5   \�O  ]    ^v ��q �  ^v ��e �   t �  )�d "  �  )6h �  �  <�  	�J     Z   �  =�  <�  	P�K     �  �  �  �  <   K5   3  K�  �  3  5   5   8     _Ln   _uh =  �i X  =F  Jf Q  c  �<�  	J     D�n &!  x �  �x 
Xx �  �  &!   C�g y �  &!  �    `�w +�v �  `�r ,�p �  7� 5      %�r  %q� %� %�� %o�  � b   /it �   /end �  a�s �� �  T   Z   �"   C Z    h� �   /it �"   /end F  a�s 2� �  �   �   �"   C Q   m� 	
<� �  �   T �  �  C   �� 	
� D  �   T D  �  C   6� 	
y� �D   !  T �D  �  C   Uzo  �  6	  6.	  i	  6!  !
  i	  6  -� �!  -� �� s!  y!  "   ,-� � �!  �!  "  "   -Gp �� "  �!  �!  "  "   7� �� �!  �!  "   �� �� �!  �!  "   3n� 5     R!  R!  "  �!  R!  >� l"  �map x� �   @"  K"  l"  �    Cɒ   �� ["  l"  �   �     "  l �"  b� �    �� �   3� �       �   Q  =�"  b   S   �"  !�    E�"  �I� r"   F�"  <�"  
        ���� ��  	`�K     �  #     !#  �     '  8#  Y  C#  �  N#  a  �  f  e#    f    |#  r
  �#    r
  N#  �  �#  	  �#  �  �#  T  �  e#  Y  �#  �  "  "  Y  �   
$  !�    �#  )g� ?  )!� m  )�� {  )K� �  b?� �   �b�� �   �5� �     )݉   �  p$  !�    4  p$  �  K4  4  �    6]  6o  ��� �}F            ��M  Z}F     /       ��$  <  �5   �l  �5   �h 	�  %  �hF     �       �1%  �  '#  �hs 
'S   �d .�  O`F     (       �n%  T 5   a �  �hb #�  �` �  ��F     1       ��%  D� Ze#  �h 	p  �%   �F     �      ��%  �  �#  ��n e#  ��u e#  �Xv e#  �Pw e#  �H 	O  &  `�F     �      �e&  �  �#  ��n �e#  ��u �e#  �Xv �e#  �Pw �e#  �H .3
  Q�F            ��&  T f  D� 'e#  �h .T
  B�F            ��&  T �  D� 'N#  �h 	   �&  ��F     �      �/'  �  �#  ��n N#  ��u N#  �Xv N#  �Pw N#  �H 	�  N'  �F     �      ��'  �  �#  ��n �N#  ��u �N#  �Xv �N#  �Pw �N#  �H S  ��F     1       ��'  D� ZN#  �h 0  (�F     �      ��(  P    T �   H N2#  ����  N$�   ��s N1�  ���s N?5   ����  O5   ��H� O5   ��ZX  O#S   ��~]� P�  �XB� S�(  ��
k T5   ��#!�F     E       �(  
i a5   �l #p�F     -       �(  
i d5   �h ��F     0       
i f5   �d  S   �(  !�    	R  )  ҿF     V      �S)  �  �#  �Xn �N#  �PS� �N#  �h� �N#  �` �  ��F            �~)  j =e#  �h 	.  �)  �F     �      �{*  �  �#  ��n xe#  ��S� {e#  �Ps �e#  �X
� �D	  ��#��F     �       *  x �e#  �H #ݻF     z       0*  x �e#  �@ #��F     Q       W*  0� �e#  �� ҾF     Q       0� �e#  ��  �  ��F     1       ��*  D� Ue#  �h P  ��F            ��*  j Le#  �h 	�  �*  Z�F     H       �+  �  �#  �XD� #e#  �P�� $e#  �h .�  D�F            �H+  j 8e#  �h 	�  g+  �F     V      ��+  �  �#  �Xn �e#  �PS� �e#  �h� �e#  �` 	�  �+  εF            ��+  �  �#  �hD� e#  �` 	A  �+  ��F            �,  �  �#  �hD� N#  �` 	a  6,  f�F     H       �c,  �  �#  �XD� #N#  �P�� $N#  �h �
  I�F            ��,  j =N#  �h 	�  �,  ��F     �      ��-  �  �#  ��n xN#  ��S� {N#  �Ps �N#  �X
� �D	  ��#U�F     �       -  x �N#  �H #q�F     z       @-  x �N#  �@ #�F     Q       g-  0� �N#  �� f�F     Q       0� �N#  ��  8  T�F     1       ��-  D� UN#  �h    6�F            ��-  j LN#  �h .
   �F            �.  j 8N#  �h r  ɮF     W       ��.  P    T �   H x2#  �h��  x!�   �`�s x-5   �\��  x85   �XH� y5   �TZX  yS   �P���f {	�     �  �.  �.  �  T#  +� �g  +� �%�   +�� �6�    *�.  ֭ �.  ~�F     K       � /  �.  �h�.  �d�.  �X�.  �P 	-  ?/  F�F     7      �z/  �  �#  �HS� �N#  �@D� �"N#  ��L� �N#  �X 	  �/  �F     7      ��/  �  �#  �HS� �N#  �@D� �!N#  ���� �N#  �X 	�  �/  ��F     j       �0  �  �#  �hD� |N#  �` y  0  K0  �  k#  +� ��   +�� �)�   +�� �65    *0  �� n0  @�F     d       ��0  0  �h&0  �`20  �X>0  �T 	�  �0  ��F     �      �1  �  �#  ��D� e#  ���  e#  ��S� e#  �X�  e#  �P�� e#  �H 6  ��F            �91  j Ie#  �h 	  X1  4�F     a      ��1  �  �#  ��D� De#  ��0� D$e#  ���� Ee#  �XL� Fe#  �PS� Ze#  �H 	}  �1  ��F     7      �2  �  �#  �HS� �e#  �@D� �"e#  ��L� �e#  �X   ݤF            �=2  j Ee#  �h 	X  \2  ��F     7      ��2  �  �#  �HS� �e#  �@D� �!e#  ���� �e#  �X   ��F            ��2  j Be#  �h 2�  �2  `�F     (       �3  �  �#  �ha �!Y#  �`b �1Y#  �X 	8  '3  ��F     j       �C3  �  �#  �hD� |e#  �` 2j  b3  �F            �o3  �  �#  �h 	�  �3  X�F     �      ��3  �  �#  ��D� N#  ���  N#  ��S� N#  �X�  N#  �P�� N#  �H �
  9�F            �4  j IN#  �h 	�  84  ؝F     a      ��4  �  �#  ��D� DN#  ��0� D$N#  ���� EN#  �XL� FN#  �PS� ZN#  �H �
  ��F            ��4  j EN#  �h �
  ��F            ��4  j BN#  �h 2  5  ��F            �5  �  �#  �h �  �F     �       �q5  T �   F    ݰ  ��   �hfo �/8  �`H �62#  �X 	�  �5  �eF     �       ��5  �  '#  �hstr 
1�  �` 	c  �5  N�F     �       �6  �  I#  �HR� %8�   �@ +�   �Xfra -N#  �P 	%  '6  �F     L       �46  �  v$  �h 	s  S6  �F     �       ��6  �  �#  �XD� �N#  �P�� �N#  �h 	?  �6  ʙF     D      �U7  �  I#  ���N  45   �� 
�   �@Y  �   ���� 	�   �Xslb e#  ��N� |#  �P��F     ^       off �   �H��F     >       ݰ  |#  ��   	  t7  r�F     X       ��7  �  �#  �X�� pe#  �h 	�  �7  ��F     �       �8  �  �#  �HD� e#  �@�� e#  �h� e#  �`&�F     I       �� e#  �X  	�  -8  F     �       �Z8  �  �#  �XD� �e#  �P�� �e#  �h 2	  y8  x�F     I       ��8  �  T#  �Xp �  �P
adr �	�   �h +  �8  �8  �  �#   5�8  �� �8  b�F            ��8  �8  �h 	@  9  �F     O       �9  �  v$  �h 	r  19  V�F     �       ��9  �  �#  �HD� N#  �@�� N#  �h� N#  �`ƖF     I       �� N#  �X  	  �9  ��F     �       ��9  �  I#  �X �6�   �P�� �N#  �h �  �9  �9  �  v$  0  <    *�9  ��  :  f�F     '       �):  �9  �h �  7:  M:  �  v$  +G� "   *):  �� p:  4�F     2       ��:  7:  �h@:  �` �  ��F     }       ��:  F    ݰ  � ]  ��fo �78  ��H �>2#  ��   eF     *       �$;  F    ݰ  � �  �hfo �78  �`H �>2#  �X 	�  C;  ��F     #      �<  �  I#  ��m  L/  ���T  L?�   �� V�   �X�� X4  ��fra YN#  �P#a�F     �       �;  slb _e#  �HY  `
�   �@!� e	  �� �F     �       !� s	  ��  	�  -<  �F     �      �@=  �  I#  ��~ss  �1�   ��~#$�F     �      �<  �N  �5   �\bkt �#  �P� 4  ��ݰ  |#  ��#��F     *      �<  slb 	e#  �H ƏF     �      slb 	e#  �@�� #4  ��  ԑF     �       R� :�   ��fra ;N#  ���� =4  ��~  	�  _=  |�F     h      �>  �  I#  ��~m  ~+  ��~ ��   �X�� �4  ��fra �N#  �Pslb �e#  �Hbkt ��#  �@Y  �	�   ��� �4  ��O� ��  ��ݰ  �|#  ��   ;  7�F     E       �c>  T   F    ݰ  3>  �HH 3!2#  �@ 	�  �>  �dF     &       ��>  �  #  �h�d 
M�  �` �  e  ndF     E       ��>  T �  F    ݰ  3�>  �HH 3!2#  �@ -  �>  ?  �  '#  +$s 
#   5�>  �z 5?  :dF     4       �F?  �>  �h?  �` "  T?  g?  �  �  0  <    5F?  Gk �?  �[F            ��?  T?  �h   �?  �?  �  �   5�?  �t �?  �[F            ��?  �?  �h �   .�  �F     +       �@  T �   a �?  �hb #�?  �` 	�  9@  ܉F     0       �f@  �  >#  �hm  g  �`6^  g)�   �X 	V  �@  ��F     (       ��@  �  >#  �h�  [�   �` 	�  �@  ��F     )       ��@  �  >#  �hm  c  �` �  ��F     �       �mA  �  W0�   ��
tc Y�   �`
e b�   �X
f c�   �P
ip d�   �H
is e�   �@��F     :       
i [�   �l  .�  �F            ��A  idx H6�   ��
tc J�   �h
s O5   �d
ip P�   �X
is Q�   �P
f R�   �H 	F  B  �F     )       �B  T   �  '#  �hݰ  
  �` 	�  >B  dF     ,       �SB  �  '#  �h>�  �  	p  yB  �cF     )       ��B  T �  �  '#  �hݰ  
�  �` �  �B  �B  �  '#  0  <    5�B  _| �B  �cF            ��B  �B  �h 	�  C  �cF     )       �C  �  #  �` M   =C  �   ǅF           ��C  T �  str 	
�  ��� 	
#C  ��Lret 	1��F     w  D  	@,J     s 	�  ��E  	�  �`
dot 	�  ��
end 	�  ��� 	�  ��
tmp 	�  �XM@� 
d 	"�  �@  Z    D  !�    �C  &E �   {�F     L      ��D  T D  str 	
�  ��� 	
#C  ��Lret 	1��F     w  D  	8,J     s 	�  �[E  	D  �l
dot 	�  �P
end 	�  �H� 	�  �@
tmp 	�  �`M� 
d 	"D  �\  �
  �   .�F     M      ��E  T �D  str 	
�  ��� 	
#C  ��Lret 	1F�F     w  D  	0,J     s 	�  �WE  	�D  �h
dot 	�  �H
end 	�  �@� 	�  ��
tmp 	�  �`M� 
d 	"�D  �X  �  �E  �E  �  �  +�L *�   *�E  [q F  vZF     V       �F  �E  �h�E  �` �   F  3F  �  �  0  <    *F  r VF  ZZF            �_F   F  �h >  mF  wF  �  �   *_F  �d �F  6ZF     #       ��F  mF  �h $&� ��D  '}F     3       �
G  �A  �*�  �h� �EC  �`loc �V�   �Xw G  	�,J      Z   G  !�    
G  $�� �5   ^|F     �       ��G  out ��G  �H~� �'�   �@�  �5�   ��p �  �Xw �G  	�,J        Z   �G  !�    �G  $�6  ~  �{F     �       �H  ptr ~  ��~�  ~!�   ��~�A    �h $wa u  �zF     �       �KH  �  u�   ��~�A  v  �h ��N j�yF     �       �}H  ptr j  ��} $�� d�   �yF     3       ��H  �� dM   �hM� d<L  �`]�  dN�   �Xw G  	�,J      $2� L�   xxF     =      �J  wcs L�"  ��mbs L+�  ��g� L7�   ��cc MJ  �hst Nr"  �P�n O   �@-� Pb   ��w G  	�,J     #�xF     N       �I  �  S
�   ���xF     H       e T�  �d  4yF            e Y
�  �`|yF     7       n ]
�   �X    !  $i� G5   JxF     .       �pJ  >� GM   �hwc G"Q  �dw �J  	�,J      Z   �J  !�    pJ  $�� >5   wF     1      ��J  wc > �"  ��~mbs >;�  ��~]�  >G�   ��~w �J  	�,J      $5� /5   vF           ��K  mbs /�  ���� /#�   ��cc 0J  �Xwc 1
Q  �P�n 2   �@-� 3b   ��w �K  	�,J     �vF     Z       e :
�  �T  Z   �K  !�    �K  $;� *	�  �uF     /       �L  ��  *�  �h�� *+�  �`w �K  	�,J      $<� &e  �uF     /       �iL  ��  &�   �h�� &�   �`w yL  	�,J      Z   yL  !�    iL  �div  1  �uF     &       ��L  ��   5   �\��  5   �Xr !1  �h $8� �  fuF     +       �M  ��  �  �hw �K  	�,J      $9� �   ;uF     +       �_M  ��  �   �hw yL  	�,J      �abs 5   uF     *       ��M  ��  5   �lw �M  	�,J      Z   �M  !�    �M  N_T  � tF           ��N  2�  �  ��.� ��   ���  �-�   ��3  �	O  ��tF     �       i  �   �h.tF     �       u 	  �PEtF     �       j �   �`_tF     �       v 
  �H�� 
M   �@�� 	
M   ���tF     V       k 
�   �X�tF     =       /� 
S   ��       �5   O  ]  ]   �N  /� �  sF     �       ��O  key �]  ��2�  �,]  ��.� �9�   ���  �G�   ��3  �	O  ��
i �	�   �h
j �	�   �`w  D  	�,J     TsF     |       
k �
�   �X��  ��  �P
res �5   �L  -� �M   �rF     +       �5P  >M   �hw �J  	�,J      � �5   �rF     +       �zP  �� ��  �hw �J  	{,J      ?V� ��rF     *       ��P  % �5   �lw �P  	p,J      Z   �P  !�   
 �P  ?i� ��rF            ��P  % �5   �l ?\� �orF            �,Q  % �5   �l S� �5   DrF     +       �qQ  �� �sQ  �hw �Q  	`,J      �qQ  Z   �Q  !�    yQ  k �5   rF     )       ��Q  �� �sQ  �h ?� ��qF     #       ��Q  w �K  	V,J      l� �  �qF     V       �BR  .� ��   �X�  �#�   �P
ptr �  �h �� �  MqF     U       ��R  P� ��   �X�  �.�   �P
ptr �  �`
ret �5   �l N-� ��pF     Z       ��R  >�   ��~ N�� ��pF     "       ��R  s ��   �l +� �5   �pF     +       �3S  >�"  �hw �J  	O,J      �� �5   �pF            �B� �?  apF     +       ��S  �� �4�  �hend �NC  �`2�  �W5   �\ �� [�   nF     G      �jT  �A  [.�  ��� [FC  ��2�  [R5   ��p� ]�   �P
s _jT  �h
acc `�   ��
c a5   �d� b�   �H
neg c5   �`
any c5   �\�� c5   �D r   ;� V�  �mF     +       ��T  �� V*�  �hend VDC  �`2�  VM5   �\ �\  0�   �lF     J      �AU  �� 0$�  �Xend 0>C  �P2�  0G5   �Lw �J  	H,J     s ;�  �oE  G�   �` M� -�  llF     9       ��U  �� -,�  �hend -FC  �` �� *D  GlF     %       ��U  �� *%�  �hend *?C  �` �� '�D  lF     3       �V  �� '&�  �hend '@C  �` �� $�  �kF     $       �6V  �� $�  �h �) !�   �kF     $       �hV  �� !�  �h � 5   �kF     $       ��V  �� �  �h *� �D  {kF     -       ��V  �� �  �h 2�!  �V  �F            ��V  �  	"  �h 	�!  W  րF     B       �7W  �  	"  �hw yL  	�,J      .7  ÀF            �`W  x )�   �h v	  nW  xW  �  <!   5`W  �� �W  r�F     Q       ��W  nW  �h 	_  �W  <�F     6       ��W  �  &  �`c 63�  �\�  78  �h c�  2�W  X  �  &  0  <    *�W  �o 4X  ZF            �=X  �W  �h   c  2TX  cX  �  &  =X   *CX  �e �X  �YF     �       ��X  TX  �h]X  �` E  �X  �X  �  &   *�X  w �X  &YF     \       ��X  �X  �h �6r kv   YF            �Y  �  #�   �hp /  �` 2L  >Y  l~F     �      �Z  �  �  �H�#�  Z  �P
res 3�   �X�~F     N      
y -�   �\#�~F     {       �Y  
kk #5   �l�~F     e       
y $�   �d  F     {       
kk (5   �h"F     e       
y )�   �`    �   Z  !�    Z  2-  ?Z  �}F     �       �YZ  �  �  �hs �   �d   gZ  qZ  �  �   *YZ  �� �Z  �}F             ��Z  gZ  �h d�    "df    " �   ��  �n �� ~c  �         � �� e6   �i 6   �� 	
N   �i X  ^� �N   S  �
  �  �  �  t  
6   �  -  int �   g  �   l �   	b� �    	�� �   	3� 6    
std  h  9t m  �\ o  �l h  �l =g   9  ?  }   �g t   W  ]  }   T h  v h    �   �v �  �\ o  �l h  �g �o �  �  �  �   �g Vl �  �  �  �   T h  v h   r  �s �  �\ �o  T �   �O  �
    ;s �C  �\ �o  T �   �O  �
    v ��q o  v ��e o   t h  �d   m  6h   �  frg 	2
  /g �  [r  �  �t  �  �q 7G
   mi �   ,�  �r  �( hex  Mq I  �h {T  ݰ  |�    �h ~�q 2  8  g
   !�h h H  g
  �     "�s  u i  o  r
   "�s p �  �  r
  #�   "�s �v �  �  r
  #}
   "�s *o �  �  r
  #�
   "�s *gs �  �  r
  #�
   "�s 0dr     r
  #�
   "�s 8�m $  /  r
  �    $Gp =�w �
  H  S  r
  #�   $�s Qr h  l  r  �
   $�s T�i h  �  �  r
   $]h X%d h  �  �  �
   $p \Xw }
  �  �  �
   $p `�k �
  �  �  r
   $�o d�g �
      r
    �� ��s !  '  r
   	wq �   	�r �h  T �    �  ,s 2   ,s 3�s o  u  �
   #m 6Rf N  �  �  �
  #�   	(m <�   	�m =�   	H� >�  	�t ?h  	v @h  	�r Ah  	;f Bh  	�u Ch  %+s �n   �
  �     &/f J�� �  "� y� C  I  �
   "� �� ^  i  �
  #A
   "� �� ~  �  �
  #A
  #\    $�U  !� A
  �  �  �
   $d  #U� �
  �  �  �
  #\    $�  '	�� \   �  �  �
   $�� +� h  	    �
  #!   $�� 3�� h  -  8  �
  #!   $I� 7	�� \   Q  a  �
  #L
  #\    $f� ?	j� \   z  �  �
  #L
   $�� G�� !  �  �  �
  #\   #\    	m  XA
   	rs  Y	\   '7�  L
   !  Dq 
�  �g �  `d �	   s E�x     X  #   j �	j	   j | >  I  c  #X   (j *{ ]  h  c  #n   )Gp 	@� t  �  �  c  #n    j  �  �  c  �    Cr "	�z t  �  �  c  #�     i '�} �  �  c  #L
     i 1Wz  	  	  c  #A
   *#s >X   *A� ?z  *�� @
\   �*m Ah  �+�m 	�~ t  ^	  T A
  c  #A
      �g Hx   �	  �	  X   "�l Mox �	  �	  X  #A
   *cg Q   '�n   ,�! N   � -Xt .�~ ��} �	  F   #A
  #N  #t   /xy 3} %
  T A
  F   #Z  #t   � \!!   0�  	�-J     S
  A
  �  L
  0�  	X�K       g
  �  r
  1�   2�   1I  2�  1�  I  1�   �   N  �
  3Ln �  3uh #  �i !  �
  �  �
  1S
  Jf 0�  	�-J     4�n �  x U  5x 
Xx 3  9  �   !�g y I  �  #A
    6�w +�v �  6�r ,�p �	  � �   �  �r  q� � �� o�  � �  7it A
   7end A
  8�s �� h  �  �  �   C S
   �� >  7it �   7end �  8�s x� h  0  6  �   C 6    �h qp  +� r^� u  _  �  #�
  #�    � #�   9zo �  +� 0�� u  �  �  #L
  #�    :�� "5� h  #p      �  6   =   �  >  1p  ;P  <6   �b�  �� ,� �� 7� �  � �� �� �� 	D� 
T� �� P�   =��  �  X    c  1j	  1  >L
  �  ?N    @C  @U  A�  �  �eF     �       ��  B�  i  �hCstr 1A
  �` D�	  eF     *       �  F   Eݰ  � A
  �hCfo �7N  �`EH �>t  �X A�	  >  �dF     &       �Z  B�  ^  �hE�d MA
  �` 1G
  D�	  ndF     E       ��  T A
  F   Fݰ  3Z  �HFH 3!t  �@ G*  �  �  H�  i  I$s X   J�  �z �  :dF     4       �  K�  �hK�  �` G8    #  H�  m
  H0  �    J  Gk F  �[F            �O  K  �h G  ]  g  H�  m
   JO  �t �  �[F            ��  K]  �h A�  �  dF     ,       ��  B�  i  �hL�  �  AC	  �  �cF     )       �	  T A
  B�  i  �hEݰ  A
  �` G�    *  H�  i  H0  �    J	  _| M  �cF            �V  K  �h Ao	  u  �cF     )       ��  B�  ^  �` M�  �  l�F            ��  B�  �
  �XE�L +%!  �@N��F     G       Oi .\   �h  GI  �  �  H�  �
  Pcs  A
   J�   � "  �F     R       �3  K�  �hK�  �` G  A  T  H�  x
  H0  �    Q3  r w  ZZF            ��  KA  �h GT  �  �  H�  x
   Q�  �d �  6ZF     #       ��  K�  �h R#� #)   ��F     *       �  L)   �lSw   	 /J      >S
    ?N      R�� )   ��F     *       �W  L)   �lSw   	/J      R�� �   9�F     Q       ��  Tnc �   �\Ucc �  �hUcp p  �`NM�F     &       Ue 
u  �d  |  �  R�� 
�   ��F     Q       �D  Tnc 
�   �\Ucc �  �hUcp p  �`N��F     &       Ue 
u  �d  Rp� �   ��F     .       ��  L)   �lLB   �`Sw   	 /J      Vr� �
B   ��F     �      ��  Ccs �A
  ��|Os �%
  ��} V�� ��   ��F     H       �7  Cnc �)   �\Occ ��  �hOcp �p  �`N��F     %       Oe �
u  �d  V�� ��   V�F     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`Nj�F     %       Oe �
u  �d  V�� ��   �F     S       �  Cnc �)   �\Occ ��  �hOcp �p  �`N�F     %       Oe �
u  �d  V�� ��   ��F     S       �{  Cnc �)   �\Occ ��  �hOcp �p  �`N��F     %       Oe �
u  �d  VM� ��   ]�F     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`Nq�F     %       Oe �
u  �d  V@� ��   
�F     S       �S  Cnc �)   �\Occ ��  �hOcp �p  �`N�F     %       Oe �
u  �d  VG� ��   ��F     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N��F     %       Oe �
u  �d  V�� ��   d�F     S       �+  Cnc �)   �\Occ ��  �hOcp �p  �`Nx�F     %       Oe �
u  �d  V�� ��   �F     S       ��  Cnc �)   �\Occ ��  �hOcp �p  �`N%�F     %       Oe �
u  �d  Vx� ��   ��F     S       �  Cnc �)   �\Occ ��  �hOcp �p  �`N��F     %       Oe �
u  �d  V�� ��   k�F     S       �o  Cnc �)   �\Occ ��  �hOcp �p  �`N�F     %       Oe �
u  �d  V]� x�   �F     S       ��  Cnc x)   �\Occ y�  �hOcp zp  �`N,�F     %       Oe {
u  �d  V�� l�   ��F     J       �G  Cnc l�   �\Occ m�  �hOcp np  �`N��F     (       Oe o
u  �d  V�� d�   ��F     K       ��  Cnc d�   �\Occ e�  �hOcp fp  �`N��F     (       Oe g
u  �d  V�� \�   -�F     V       �  Cnc \�   �\Occ ]�  �hOcp ^p  �`NA�F     (       Oe _
u  �d  V�� T�   ��F     V       ��  Cnc T�   �\Occ U�  �hOcp Vp  �`N��F     (       Oe W
u  �d  V�� L�   ��F     V       ��  Cnc L�   �\Occ M�  �hOcp Np  �`N��F     (       Oe O
u  �d  V� D�   +�F     V       �c  Cnc D�   �\Occ E�  �hOcp Fp  �`N?�F     (       Oe G
u  �d  V�� <�   ��F     V       ��  Cnc <�   �\Occ =�  �hOcp >p  �`N��F     (       Oe ?
u  �d  V�� 4�   �F     V       �;  Cnc 4�   �\Occ 5�  �hOcp 6p  �`N��F     (       Oe 7
u  �d  VV� ,�   )�F     V       ��  Cnc ,�   �\Occ -�  �hOcp .p  �`N=�F     (       Oe /
u  �d  V�� $�   ��F     V       �  Cnc $�   �\Occ %�  �hOcp &p  �`N��F     (       Oe '
u  �d  VY� �   }�F     V       �  Cnc �   �\Occ �  �hOcp p  �`N��F     (       Oe 
u  �d  V� �   '�F     V       ��  Cnc �   �\Occ �  �hOcp p  �`N;�F     (       Oe 
u  �d  V	� �   ��F     V       �W  Cnc �   �\Occ �  �hOcp p  �`N��F     (       Oe 
u  �d  W�  ��F     0       ��  Cc "*p  �l A�  �  ��F           �8  B�  �  ��Cnc 0L
  ��Cwc 0-�  ��Ouc 1{   �oX�n 7�  �PX-� 8�  �@Ost 9�   ��Sw H  	�.J     N]�F     .       Oe ;u  �h  >S
  H  ?N    8  Y   2^  q  H�  �
  H0  �    QM  �o �  ZF            ��  K^  �h G[  �  �  H�  �
   Q�  w �  &YF     \       ��  K�  �h &E �
   �T   �  ^�n �� ~c p�         q� 1�� 	5   _int 5   1�� M   
X   M   �  X   1! M   ^� ��   p   �i `X  S  �i �   {S @'  g
  M       	p   v  #	p   �  &	p   |
  )	p    h  ,	p   (�  -	p   0�	  25   8�  55   < �
  8"�   1  K?  
'  1�  L?  1�  M?  �
  a�  �  i  �  �  -  �  ��   �  4�  �  bstd  �  9t $  -�\ �  �l �  �l =g �  �  �  �   �g t �      �   T �  Iv �    �  �v �  -�\ �  �l �  �g �o C  g  m  �   �g Vl C  �  �  �   T �  Iv �   )  �s ��  -�\ ��  T 5   J�O  K�%    ;s ��  -�\ ��  T 5   J�O  K�%    � `  � a5  T �D   <� `<  � aM   T �'   Lv ��q �  Lv ��e �  �� j>  �� !|� `  �  T �D  �D   5�� �� �  T M   �'  �'   �� j>(  M/� !�� �  T �'  �'    t �  .�d �  
$  .6h 6  
�  cfrg '$  >�� 	  dW�    ?`� 	  @J  N� �    A7  B>� 5   w  /�r  Ored /d�  l� 0/  l� � �  �  1$   )l� � �  �  1$  <$   *Gp ;� B$  �  �  1$  <$   S� �    �  �   �� �   )�  �   �� !�    � "R  ( w  �� %�  �� '{� �  b  T t  (   MJ� ';� �  T �  �'    f� 5	  Ph 8`� 1$  �  �'   O� =t� �'  �  �'   �� BͰ �'  �  �'   n� E� �'  �  �'   )� I�� �'    �'   �� L7� �'  (  �'   �� PE� �'  @  F  /(   8#� U�� �  a  �'   8�� Z؟ �  |  �'   � d� �  �  /(   )� g� �  �  /(  :(   *Gp i;� @(  �  �  /(  :(   N� o�� �'  �  �  /(   � |\�     /(  �'   c� ��� +  ;  /(  �'  �'   �� ��� P  `  /(  �'  �'   
� �6� u  �  /(  �'    �� #� �  �  /(  �'   <� � �  �  /(  �'  �'   �� D� �  �  /(  �'  �'   �� x)�     /(  �'   �� �$� #  .  /(  �'   /� �� D  O  /(  �'    � u� d  o  /(  �'    ,� #E� �  �  /(  �'   00� 0�� �  �  �  /(   00� 94� �  �  �  /(  �'  �%  F(  F(   2�� ��    D 	  T �  9� �T  A 4   �  Q� ��	  !��  !�  !�;  !��  !��  !�(  C�    �� �\� v	  �	  W(  �    \+  ��� �	  �	  W(  �'   2�� ��  T �  9� �T  L �  A 4   _� 5b  Ph 8� 1$  �	  (   O� =� (  
  (   �� B� (  *
  (   n� E2� (  D
  (   )� I�� (  ^
  (   �� L� (  x
  (   �� PK� (  �
  �
  b(   8#� U� �  �
  (   8�� Zk� �  �
  (   � dg� �
  �
  b(   )� g4� �
    b(  m(   *Gp iI� s(    (  b(  m(   N� o�� (  @  F  b(   � |c� [  f  b(  (   c� �)� {  �  b(  (  (   �� ��� �  �  b(  (  (   
� �� �  �  b(  (    �� U� �  �  b(  (   <� ��     b(  (  (   �� Dz� ,  <  b(  (  (   �� x�� R  ]  b(  (   �� �Z� s  ~  b(  (   /� �� �  �  b(  (    � ;� �  �  b(  (    ,� #�� �  �  b(  (   00� 0�� �  �  �  b(   00� 9�� �    3  b(  (  �%  y(  y(   2�� ��    D g  T t  9� �T  XA 4   �	  eW� �!�F  !�f  !��  !�
  !�*
  !�x
  C�	    �� �F� �  �  (  �    \+  �Q� �  �  (  (   2�� ��  T t  9� �T  XL �  A 4    @0  N� �    A  �� g  fclz � 5   _  �    T �    g"� �$0  B"� 5   ��  /�r  /l� /[�  u  � H�	o  � ��� �  �  �'  u  �  p    )� �5� �  �  �'  (   *Gp �
�� (      �'  (   Z� �δ �  /  :  �'  �    � ��    ��  ss  �|   "� �A!   �  � ��	'  C�   � �E� �  �  (  �  p   5    )� ��� �  �  (  (   *Gp �r� (  �  �  (  (   �N  �<   Hٖ ��   LU� �$(  P.� �A!  X t  '� �	�  '� ��� M  S  $(   )'� �Ƈ g  r  $(  4)   *Gp �Ⱥ :)  �  �  $(  4)   ʊ �$(    ,  � �	�  R�g �a� �  �  L(  (  (    �0   �	)  �0  ��� �    �(   � �	M$   x� �(  � �)   �� �N!  �� �-� J  U  �'  �(   S�� (z� j  u  �'  �(   hGp *� �(  �  �  �'  �(   Wd ��� �   �  �  �'  p    0�6  L�� �   �  �  �'  �   p    �N ~�� �    �'  �    � �w�   .  �'  �   p    Y� 1	�� p   G  M  �'   iJ� >�(                         @       D�� @ �   D�� A �    H� H�� p   �  �    r� W�� p   �  p    D�� j<   -� l|   �� o�� �     �    -o� ||   -�� |   j� �|    E<� �7� �'  B  M  �'  �   Ea� �� (  f  q  �'  5    EP� %j� �'  �  �  �'  p     `� 7� �  �  �'    � >� �  �  �'  �'   Э �
�(   A� �M$  ۧ �[!  @� ��  �� �	p    � �)  (+� %  +v� M$   g  k0� V  ;� X� Y  d  �'  �'   0Wd [!� �   ~  �  �'  p    � _ʅ �  �  �'  �   p    �N c�� �  �  �'  �    0� gε �   �  �  �'  �   p    l�� l�'   +� %  +v� M$   >/g   T[r  $  m�t  P  n�q 7�%   Bmi 5   ,u  /�r  /�( Ohex  :Mq �  o�h {�  pݰ  |5   �h ~�q �  �  �%   F�h h �  �%  5     �s  u �  �  �%   �s p     �%     �s �v !  ,  �%  �%   �s *o A  L  �%  �%   �s *gs a  l  �%  �%   �s 0dr �  �  �%  �%   �s 8�m �  �  �%  5    Gp =�w �%  �  �  �%  u   �s Qr �  �  �  �%   �s T�i �      �%   ]h X%d �  '  -  �%   p \Xw �%  F  L  �%   p `�k �%  e  k  �%   �o d�g �%  �  �  �%   �� ��s �  �  �%   wq ��   �r ��  T 5    u  ,s 2�  ,s 3�s �  �  �%   #m 6Rf �  
    �%  P   (m <P   �m =5   H� >u  �t ?�  v @�  �r A�  ;f B�  �u C�  q+s �n �  �  �%  5    r,s  i �  �%  �R    �  ?/f Jm  5�� Nm{   P �  T �   �'  �   �  5   5   5   X    5B~ xR B  P �  T �   �'  �   5   5   5   X    s*y �� T �   F �  �   �  �'    :��   � y� �  �  &   � �� �  �  &  {%   � �� �  �  &  {%  p    �U  !� {%  �  �  &   d  #U� &      &  p    �  '	�� p   6  <  &   �� +� �  U  `  &  m   �� 3�� �  y  �  &  m   I� 7	�� p   �  �  &  X   p    f� ?	j� p   �  �  &  X    �� G�� m  �  �  &  p   p    m  X{%   rs  Y	p   +7�  X    m  Q�� u   �� "=� F  V  $&  /&  p    2A� &/&   2V� '	p    #  >Dq 	
z  T�g 	�  `d 	�  s 	E�x �  �  e'  Q&   j �		7  j 	| �  �  p'  e'   )j 	*{      p'  {'   *Gp 		@� �'  #  .  p'  {'   j 	 B  M  p'  5    Cr 	"	�z �'  e  p  p'  z    i 	'�} �  �  p'  X     i 	1Wz �  �  p'  {%   3#s 	>e'   3A� 	?�'  3�� 	@
p   �3m 	A�  ��� 		� �'      T #  p'  #   R�m 		�~ �'  +  T {%  p'  {%    �  �g 	Hx �  T  Z  e'   �l 	Mox o  z  e'  {%   3cg 	QQ&   +�n Q&  t�! �   � uXt :��  
<!  ��  
��� �  �  �'  5   ��  
?� �  �  �'  �'   ��  
$U�     �'  �'   #� 
�f� #  .  �'  5    Gp 
+
� �'  G  R  �'  �   �# 
��� �'  k  v  �'  �'   �# 
��� �'  �  �  �'  �'   � 
4"� �'  �  �  �'  �'   � 
8+� �'  �  �  �'  �'   Gpop 
��� M   �    �'   ��  
Dy�     �'   �U  
J� _'  5  ;  �'   �U  
Nj� �'  T  Z  �'   �  
R	�� p   s  y  �'   �4 
V&� �  �  �  �'   6 
Z�� _'  �  �  �'   6 
^>� �'  �  �  �'   Gend 
b�� _'  �  �  �'   Gend 
f�� �'        �'   �  
j�� �'  -   3   �'   �  
m�� �'  L   R   �'   0  
q1� �'  k   q   �'   0  
t�� �'  �   �   �'   d  
x�� �'  �   �   �'  p    d  
{�� �'  �   �   �'  p    �� 
��� �   �   �'  p    ?� 
�5   '2 
�_'  V� 
�	p   �� 
�	p   T M   +E� 5   �  HG� �+w  H� �7g  H� �7	  :#� �"  0� �� �!  �!  )   0� ׁ �!  �!  )    %   0� I� �!  �!  )  %   S0� !�� �!  �!  )  ")   0� #E� 
"  "  )  ()   /� (�� *"  5"  )  5    Gp -
� .)  N"  Y"  )  h!   7� 2�� n"  t"  )   �� 8�� �"  �"  )   �� >U� �  �"  �"  )   <� Bn� �  �"  �"  )  �$   F� G	�$   �� H�  +v� M$   h!  t 
*w �%  !#  T 5   �%  �%   5�~ ��| H#  F �  �   �  �'   ;�{ 82� w#  T �   F �  �?  �  �'   ;�~ � �#  F �  #  �  �'   5�~ ��} �#  F �  {%  �  �'   ;�� 3\� �#  T #  F �  rE  �'   ;xy 3} $  T {%  F �  �E  �'   � \!m   6  6<  
w  1$  /  w  6"  -� �$  -� �� n$  t$  �$   )-� � �$  �$  �$  	%   *Gp �� %  �$  �$  �$  	%   7� �� �$  �$  �$   �� �� �$  �$  �$   3n� 5     M$  
M$  �$  �$  M$  >� f%  vmap x� �  :%  E%  f%  p    Fɒ   �� U%  f%  �  p     
%  <)  	�/J     
_   {%  <B  	`�K     
�  �%  
u  �%  <   75   �  7u  u  
�  5   
5   
�  �%  ULn �  Uuh �  �i 
m  &  
  &  _   Jf 
#  $&  
5&  w<�  	�/J     ?�n �&  x �&  xx 
Xx s&  y&  �&   F�g y �&  �&  {%    V�w +�v �  V�r ,�p �   
Q&  @"'  y�� *'  W�� O�&  $   W�� <�&  $  {%  �   zX� -{� ('�'  |� p   $    A�&  %M   :'  &�     <�&  	@�K     }�  _'  	 �K     
M   
�  e'  
�  p'  7  �  %X   �'  &�    
5  �'  
g  �'  
�  �'  <!  7�  �  M   S   7M   
S   
<!  �'  ~Z  �   
�  �'  o  �  
t  (  '  t  
,  $(  
�  /(  	  �  �'  
�  L(  
	  W(  
�	  b(  b  �	  (  
g  (  
�  %  0  g  %|   �(  &�    �(  .g� M  .!� {  .�� �  .K� �  X?� �   �X��     5�      .݉   %�  )  &�    
h!  )  �"  7h!  h!  �  ,  6<  6N  '�"  O`F     (       ��)  T 5   a �%  �hb #�%  �` �
  ��F     1       ��)  D� Z(  �h �  RgF     �      ��*  P �  T �   H N�'  ����  N$�   ��s N1�  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P{%  �XB� S�*  ��k T5   ��#BhF     E       �*  i a5   �l #�hF     -       �*  i d5   �h �hF     0       i f5   �d  %X   �*  &�    `  +  ҿF     V      �E+  �  5(  �Xn ��'  �PS� ��'  �h� ��'  �` <  d+  �F     �      �B,  �  h(  ��,n x(  ��	S� {(  �Ps �(  �X	
� �R  ��#��F     �       �+  x �(  �H #ݻF     z       �+  x �(  �@ #��F     Q       ,  	0� �(  �� ҾF     Q       	0� �(  ��  ~  a,   �F     �      ��,  �  h(  ��,n (  ��u (  �Xv (  �Pw (  �H ]  �,  `�F     �      �-  �  h(  ��,n �(  ��u �(  �Xv �(  �Pw �(  �H �
  ��F     1       �9-  D� U(  �h �	  ��F            �d-  j =(  �h 'A  Q�F            ��-  T t  D� '(  �h 'b  B�F            ��-  T �  D� '�'  �h .  �-  ��F     �      �..  �  5(  ��,n �'  ��u �'  �Xv �'  �Pw �'  �H   M.  �F     �      ��.  �  5(  ��,n ��'  ��u ��'  �Xv ��'  �Pw ��'  �H a  ��F     1       ��.  D� Z�'  �h   �fF     U       �R/  P �  T �   H x�'  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �TY��f {	�     �  `/  �/  �  �'  $� �u  $� �%�  $�� �6p    "R/  ֭ �/  ~�F     K       ��/  `/  �hi/  �du/  �X�/  �P ;  �/  F�F     7      �,0  �  5(  �HS� ��'  �@D� �"�'  ��L� ��'  �X   K0  �F     7      ��0  �  5(  �HS� ��'  �@D� �!�'  ���� ��'  �X �  �0  ��F     j       ��0  �  5(  �hD� |�'  �` �  �0  �0  �  (  $� ��  $�� �)p   $�� �65    "�0  ��  1  @�F     d       �A1  �0  �h�0  �`�0  �X�0  �T �  `1  ��F     �      ��1  �  h(  ��D� (  ���  (  ��	S� (  �X	�  (  �P	�� (  �H   �1  4�F     a      �?2  �  h(  ��D� D(  ��0� D$(  ��	�� E(  �X	L� F(  �P	S� Z(  �H ^
  ��F            �j2  j L(  �h �  �2  Z�F     H       ��2  �  h(  �XD� #(  �P	�� $(  �h D
  ��F            ��2  j I(  �h '�	  D�F            �3  j 8(  �h �  +3  �F     V      �c3  �  h(  �Xn �(  �PS� �(  �h� �(  �` �  �3  εF            ��3  �  h(  �hD� (  �` O  �3  ��F            ��3  �  5(  �hD� �'  �` o  �3  f�F     H       �'4  �  5(  �XD� #�'  �P	�� $�'  �h �  I�F            �R4  j =�'  �h �  q4  ��F     �      �O5  �  5(  ��,n x�'  ��	S� {�'  �Ps ��'  �X	
� �R  ��#U�F     �       �4  x ��'  �H #q�F     z       5  x ��'  �@ #�F     Q       +5  	0� ��'  �� f�F     Q       	0� ��'  ��  F  T�F     1       �z5  D� U�'  �h   6�F            ��5  j L�'  �h '�   �F            ��5  j 8�'  �h B  afF     �       �'6  T �   F �  ݰ  ��   �lfo �/�  �`H �6�'  �X q  F6  N�F     �       ��6  �  �'  �HR� %8p   �@	 +�  �Xfra -�'  �P �	  �6  �F     �       ��6  �  ](  �XD� ��'  �P	�� ��'  �h M  �6  ʙF     D      ��7  �  �'  ���N  45   ��	 
�  �@	Y  �   ��	�� 	p   �Xslb (  ��	N� $(  �P��F     ^       off p   �H��F     >       	ݰ  $(  ��   (  �7  r�F     X       ��7  �  h(  �X�� p(  �h �  �7  ��F     �       �]8  �  h(  �HD� (  �@	�� (  �h	� (  �`&�F     I       	�� (  �X  �  |8  ��F     7      ��8  �  h(  �HS� �(  �@D� �"(  ��L� �(  �X *
  ݤF            ��8  j E(  �h f  9  ��F     7      �<9  �  h(  �HS� �(  �@D� �!(  ���� �(  �X 
  ��F            �g9  j B(  �h �  �9  `�F     (       ��9  �  R(  �ha �!(  �`b �1(  �X F  �9  ��F     j       ��9  �  h(  �hD� |(  �` x
  :  �F            �:  �  h(  �h �  3:  X�F     �      ��:  �  5(  ��D� �'  ���  �'  ��	S� �'  �X	�  �'  �P	�� �'  �H �  9�F            ��:  j I�'  �h �  �:  ؝F     a      �=;  �  5(  ��D� D�'  ��0� D$�'  ��	�� E�'  �X	L� F�'  �P	S� Z�'  �H �  ��F            �h;  j E�'  �h �  ��F            ��;  j B�'  �h Y"  �;  �F     L       ��;  �  )  �h (  �;  ��F            ��;  �  5(  �h !#  FeF     J       �<<  F �  ݰ  �!�   �Lfo �8�  �@H �?�'  �� �  [<  �F     �      �n=  �  �'  ��~ss  �1p   ��~#$�F     �      (=  �N  �5   �\bkt �(  �P	� h!  ��	ݰ  $(  ��#��F     *      �<  slb 	(  �H ƏF     �      slb 	(  �@	�� #h!  ��  ԑF     �       	R� :�   ��fra ;�'  ��	�� =h!  ��~  �  �=  F     �       ��=  �  �(  �XD� �(  �P	�� �(  �h   �=  x�F     I       �>  �  �'  �Xp ��   �Padr �	�   �h 9  >  >  �  *(   (>  �� =>  b�F            �F>  >  �h t"  e>  �F     O       �r>  �  )  �h �  �>  V�F     �       ��>  �  5(  �HD� �'  �@	�� �'  �h	� �'  �`ƖF     I       	�� �'  �X  )  ?  ��F     �       �<?  �  �'  �X �6�  �P	�� ��'  �h "  J?  ]?  �  )  0  <    "<?  �� �?  f�F     '       ��?  J?  �h �!  �?  �?  �  )  $G� %   "�?  �� �?  4�F     2       ��?  �?  �h�?  �` �   H#  ��F     N       �B@  T �   F �  ݰ  8�?  �H,fo 8-�  �@H 84�'  �� p  a@  �hF     �       �{@  �  v'  �hs 	'X   �d �  �@  �eF     �       ��@  �  v'  �hstr 	1{%  �` d  �@  ��F     (       ��@  �  �'  �h�  [p   �` �  A  |�F     h      ��A  �  �'  ��~m  ~+�   ��~	 ��   �X	�� �h!  ��fra ��'  �Pslb �(  �Hbkt ��(  �@	Y  �	p   ��	� �h!  ��	O� ��  ��	ݰ  �$(  �� w#  ��F           �iB  F �  ,� '#  ��,fo <�  ��H C�'  ��p iB  �`��F     �      i p   �h�F     �      c 	i  �_   
p  �#  eF     *       ��B  F �  ݰ  � {%  �hfo �7�  �`H �>�'  �X �   �B  ��F     �       �\C  �  �'  ���� 
�4p   ���� 
�	p   �H4� 
�_'  �@#�F     ^       <C  i 
�p   �X y�F            i 
�p   �P  �  {C  ��F     )       ��C  �  �'  �hm  c�   �` �  ��F     �       �'D  �  W0p   ��tc Y�   �`e b�   �Xf c�   �Pip d�   �His e�   �@��F     :       i [�   �l  '�  �F            ��D  idx H6�   ��tc J�   �hs O5   �dip P�   �Xis Q�   �Pf R�   �H 5  'l  ��F            ��D  T �D  x *�D  �h �  �D  �D  �  &  Zs  {%  $ss  *p    (�D  �� E  ��F     *       �7E  �D  �h�D  �`�D  �X Z  VE  �dF     &       �rE  �  k'  �h�d 	M{%  �` u  �#  M�F     I       ��E  T #  F �  ݰ  3rE  �HH 3!�'  �@ �%  �#  ndF     E       �F  T {%  F �  ݰ  3�E  �HH 3!�'  �@ �   F  6F  �  v'  $$s 	e'   (F  �z YF  :dF     4       �jF   F  �h)F  �` �  xF  �F  �  �%  0  <    (jF  Gk �F  �[F            ��F  xF  �h �  �F  �F  �  �%   (�F  �t �F  �[F            ��F  �F  �h �  G  �F     I       �6G  �  �'  �X��  
�M   �h �  ��F     O       ��G  T M   x �'  �Xy �'  �P/� M   �h '�  ��F            ��G  T �'  x *�'  �h Z  �G  ��F            ��G  �  �'  �h R   �G  l�F     %       �
H  �  �'  �h �   )H  J�F     !       �EH  �  �'  �h�N  
{p   �` v  dH  ��F     �       ��H  �  �'  �H��  
�#�'  �@m  
�_'  �X R  �H  L�F     w       ��H  �  �'  �X��  
�(�'  �Pm  
�_'  �h   �H  �F     4       �$I  �  �'  �X �F            i 
Ep   �h    CI  �F            �PI  �  �'  �h   ^I   ~I  �  �'  0  <   Y�i 
�p     "PI  Z� �I  ��F     C       ��I  ^I  �X�pI  �I  �qI   �pI  ��F            �qI  �h  �  �I   �I  �  �'  $@� 
�(5   "�I  T� "J  r�F     P       �3J  �I  �X�I  �P <  RJ  l�F            ��J  �  &  �X�L +%m  �@��F     G       i .p   �h  �  �J   �F     r       ��J  �  &  �X�� G&p   �P�  G3p   �H M  �J  dF     ,       �K  �  v'  �h�z  �  �  2K  ��F     6       �NK  T #  �  v'  �hݰ  	#  �P   mK  ��F            �zK  �  &  �h �  �K  ��F            ��K  �  &  �h   �K  �cF     )       ��K  T {%  �  v'  �hݰ  	{%  �` .  �K  	L  �  v'  0  <    (�K  _| ,L  �cF            �5L  �K  �h <  TL  �cF     )       �aL  �  k'  �` �  �L  R�F     S       ��L  �  &  �Xc 7X   �T�� 7#p   �Hc�F     9       i 8p   �h  �  �L  �L  �  &  Zcs  {%   (�L   � M  �F     R       �M  �L  �h�L  �` L  -M  CM  �  �%  $�L *�%   "M  [q fM  vZF     V       �wM  -M  �h6M  �` �  �M  �M  �  �%  0  <    "wM  r �M  ZZF            ��M  �M  �h �  �M  �M  �  �%   "�M  �d �M  6ZF     #       �N  �M  �h =#� �5   ��F     >       �:N  F@ �{%  �X =%� x5   ��F     �      ��N  F@ x{%  ��}�\ x*{%  ��}�� x55   ��}� y$  ��~s z	p   �X�� �M   ��}4w �N  	�DJ      %_   �N  &�    �N  =c� m5   I�F     �       �DO  �� m{%  ��� n$  �@s o	p   �X4w �N  	�DJ      =�  bM   �F     �       ��O  F@ b{%  ��k c�   �h� g$  �@s h	p   �`4w �N  	�DJ      �&  �F     r      �P  F@ O)$  �@��  P�'  �X4w P  	�DJ     k S�   �P %_   P  &�    P  �&  ��F     ?      ��P  F@ <'$  ���� <9{%  ���� <F�  ����  =�'  �X4w �P  	�DJ     k @�   �P %_   �P  &�    �P  �&  �F     �       ��P  ��  .�'  �`E�F     P       i 5p   �h  '  ��F     o       �.Q  ��  ).�  	`�K      '  ��F     �      ��Q  F@ ,$  ��}�F     o      i p   �X9�F     <      � $  ��~s 
p   �P   1  �Q  �Q  �  *&  [B� "/&  [�  "(p    (�Q  � �Q  (�F     *       �R  �Q  �h�Q  �`�Q  �X �  5R  <�F     6       �_R  �  �%  �`c 63P  �\�  7�  �h \}  2pR  �R  �  �%  0  <    "_R  �o �R  ZF            ��R  pR  �h �  \�  2�R  �R  �  �%  �R   "�R  �e �R  �YF     �       �	S  �R  �h�R  �` �  S  !S  �  �%   "	S  w DS  &YF     \       �MS  S  �h �6r kv �   YF            ��S  �  #p   �hp /�   �` �$  �S  �F            ��S  �  %  �h �$  �S  րF     B       ��S  �  %  �h4w T  	�DJ      %_   T  &�    �S  'E  ÀF            �:T  x )�   �h �  HT  RT  �  7$   (:T  �� uT  r�F     Q       �~T  HT  �h &E �
  ]�  A!  "]t  A!  " q    ��  �n � ~c q� �� 4   
       �int �� Q   	��K     W   �  ! Q   	��K      �u   ��  x�n � ~c �         �� 7�� 	5   yint 5   7�� M   S   !�  S   7! M   ^� �|   k   !�i |   z!X  !S  !�  !�  !�i �   !�  !-  �  �|   �  4�   �   ]� �   {S @l  g
  M       	k   v  #	k   �  &	k   |
  )	k    h  ,	k   (�  -	k   0�	  25   8�  55   < �
  8"�   7  K�  l  7�  L�  7�  M�  d �   !�
  {�  |std  �  9t 7  4�\ �  �l �  �l =g �    	  �   �g t �  !  '  �   T �  [v �    �  �v �  4�\ �  �l �  �g �o V  z  �  �   �g Vl V  �  �  �   T �  [v �   <  �s ��  4�\ ��  T 5   \�O  .�'    ;s �  4�\ ��  T 5   \�O  .�'    ]�� l]	 ~� `>  � a�  T �0   �� j>*  �� `k  � a5   T �'   �
 `�  � a�0  T T   � [�  � \�c  T �c   F	 [�  � \�b  T �b   ^v ��q �  ^v ��e �  �� j>x  � !�� �    T T  T   A� �&  <  T �b  �U   �� j>�  � q� �'  i  T �'  �V   �� j>W  A� '  �  T �c  �V   �� j>�   !t �  5�d �  7  56h I  �  }frg 	�'  B/g �  _[r  �  ~�t  
  �q 7�'   <mi 5   ,/  #�r  #�( `hex  aMq �  ��h {�  �ݰ  |5   �h ~�q k  q  �'   C�h h �  �'  5     �s  u �  �  �'   �s p �  �  �'  �   �s �v �  �  �'  �'   �s *o �    �'  �'   �s *gs   (  �'  �'   �s 0dr =  H  �'  �'   �s 8�m ]  h  �'  5    'Gp =�w �'  �  �  �'  /   '�s Qr �  �  �  �'   '�s T�i �  �  �  �'   ']h X%d �  �  �  �'   'p \Xw �'      �'   'p `�k �'  !  '  �'   '�o d�g  (  @  F  �'   �� ��s Z  `  �'   wq �<   �r ��  T 5    /  ,s 2p  ,s 3�s �  �  (   #m 6Rf �  �  �  (  
   (m <
   �m =5   H� >/  �t ?�  v @�  �r A�  ;f B�  �u C�  �+s �n K  V  (  5    �,s  i d  (  �t    �  D/f Jn	  6� N�� �  P �	  T 5   m1  5   �  5   5   5   S    6�� Nm{ 	  P �	  T �   m1  �   �  5   5   5   S    6@  x� B	  P �	  T 5   m1  5   5   5   5   S    �� �i� T 5   F �	  5   �  m1    BDq 	
n	  _�g 	w	  `d 	�  s 	E�x �	  �	  Q1  T(   j �		U  j 	| �	  �	  \1  Q1   /j 	*{ �	  �	  \1  g1   0Gp 		@� m1  
  "
  \1  g1   j 	 6
  A
  \1  5    Cr 	"	�z m1  Y
  d
  \1  n	    i 	'�} x
  �
  \1  S     i 	1Wz �
  �
  \1  �'   #s 	>Q1   A� 	?�0  �� 	@
k   �m 	A�  ��
 		�� m1  �
    T S   \1  S    Q� 		� m1  #  .  T 5   \1  5    M�m 		�~ m1  I  T �'  \1  �'    �	  �g 	Hx �	  r  x  Q1   �l 	Mox �  �  Q1  �'   cg 	QT(   �n T(  b�! |   � Xt 	�  s 	ECo �  �  �1  �(   j �		3  j 	�e     �1  �1   /j 	ig &  1  �1  �1   0Gp 		�j �1  I  T  �1  �1   j 	�f h  s  �1  5    Cr 	"	�r �1  �  �  �1  n	    i 	'�h �  �  �1  S     i 	1~j �  �  �1  �'   #s 	>�1   A� 	?�0  �� 	@
k   �m 	A�  �M�m 		3m �1  '  T �'  �1  �'    �  �g 	H�o �  P  V  �1   �l 	Mj k  v  �1  �'   cg 	Q�(   �n �(  b�! |   � B�� 	�  �W� �   D`� 	�  E�  N� �    O�  <>� 5     #�r  `red #d�  l� 0�  l� � "  (  �/   /l� � <  G  �/  �/   0Gp ;� �/  _  j  �/  �/   S� �    �  �   �� �   )�  �   �� !�    � "�  (   �� %
  �� '{� �  �  T �  �2   cJ� ';� �  T *  �2    f� 5�  dh 8`� �/  0  �2   O� =t� �2  J  �2   �� BͰ �2  d  �2   n� E� �2  ~  �2   )� I�� �2  �  �2   �� L7� �2  �  �2   �� PE� �2  �  �  �2   F#� U�� �  �  �2   F�� Z؟ �    �2   � d�      �2   /� g� 4  ?  �2  �2   0Gp i;� �2  W  b  �2  �2   N� o�� �2  z  �  �2   � |\� �  �  �2  �2   c� ��� �  �  �2  �2  �2   �� ��� �  �  �2  �2  �2   
� �6� �  
  �2  �2   $�� #�   *  �2  �2   <� � @  P  �2  �2  �2   �� D� f  v  �2  �2  �2   �� x)� �  �  �2  �2   �� �$� �  �  �2  �2   /� �� �  �  �2  �2   $� u� �  �  �2  �2   $,� #E�     �2  �2   (0� 0�� �  3  9  �2   (0� 94� �  S  m  �2  �2  �'  �2  �2   G�� ��    D �  T *  =� �u  A �   
  P� �Z  )��  )��  )��  )�J  )�d  )��  >
   $�� �\�      3  3   $\+  ���    +  3  �2   G�� �3  T *  =� �u  L 3  A �   _� 5�  dh 8� �/  �  �2   O� =� �2  �  �2   �� B� �2  �  �2   n� E2� �2  �  �2   )� I�� �2  �  �2   �� L� �2    �2   �� PK� �2       3   F#� U� �  ;  �2   F�� Zk� �  V  �2   � dg� j  p  3   /� g4� �  �  3  &3   0Gp iI� ,3  �  �  3  &3   N� o�� �2  �  �  3   � |c� �  �  3  �2   c� �)�     3  �2  �2   �� ��� *  :  3  �2  �2   
� �� O  Z  3  �2   $�� U� o  z  3  �2   <� �� �  �  3  �2  �2   �� Dz� �  �  3  �2  �2   �� x�� �  �  3  �2   �� �Z� �    3  �2   /� ��   )  3  �2   $� ;� >  I  3  �2   $,� #�� ^  i  3  �2   (0� 0�� �  �  �  3   (0� 9�� �  �  �  3  �2  �'  23  23   G�� ��    D �  T �  =� �u  XA �   Z  eW� �)��  )��  )�  )��  )��  )�  >Z   $�� �F� L  W  83  3   $\+  �Q� l  w  83  �2   G�� �3  T �  =� �u  XL 3  A �    E�  N� �    O�  �� �  fclz � 5   �  |    T |    �"� �$�  <"� 5   �%  #�r  #l� #[�     � H�	�  � ��� K  `  �2     �   k    /� �5� t    �2  �2   0Gp �
�� �2  �  �  �2  �2   Z� �δ �  �  �  �2  �    � �%    ��   ss  �w   "� �\#   *  � ��	�  >*   � �E� &  ;  �2  �   k   5    /� ��� O  Z  �2  �2   0Gp �r� �2  r  }  �2  �2   �N  �<   Hٖ ��   LU� ��2  P.� �\#  X �  '� �	.  '� ��� �  �  �2   /'� �Ƈ �  �  �2  4   0Gp �Ⱥ 4       �2  4   ʊ ��2    �  � �	e  M�g �a� �  T  3  �2  �2    �0   �	�  �0  ��� �  �  C3   � �	�/   x� ��2  � ��   �� �i#  �� �-� �  �  ~1  I3   g�� (z� �     ~1  O3   �Gp *� U3    %  ~1  O3   'Wd ��� �   >  I  ~1  k    (�6  L�� �   c  s  ~1  �   k    �N ~�� �  �  ~1  �    � �w� �  �  ~1  �   k    'Y� 1	�� k   �  �  ~1   �J� >k3                         @       Q�� @ �   Q�� A �    H� H�� k   >  �    r� W�� k   X  k    Q�� j<   4� lw   �� o�� �  �  �    4o� |w   4�� w   �� �w    H<� �7� �2  �  �  ~1  �    Ha� �� �2  �  �  ~1  5    HP� %j� �2    #  ~1  k    $`� 7� 8  >  ~1   $� >� S  ^  ~1  �2   Э �
I3   A� ��/  ۧ �v#  @� �x  �� �	k    � ��3  (� d0  v� �/   �  �0� V�  ;� X� �  �  s1  ~1   (Wd [!� �       s1  k    � _ʅ .  >  s1  �   k    �N c�� T  _  s1  �    (� gε �   y  �  s1  �   k    ��� l~1   � d0  v� �/   D�$ �"  B;	 K� 9  � � �  �  �0   	 $�0  �@ �   �  &�0  �    C �  �� �0  �  �0   �L R�"   SN�  E>  hh %7� 	1  n  y  1  y   S�  "6   ��  *	�   R�"   hh -	� 	1  �  �  /1  y   ��  2F �  �  /1  y   p 5�  y  �  �  :1   �� 9*� �        :1  E1   �� <&� �  4   ?   :1  E1   �
 @: K1  W   ]   /1   �
 D� �  u   �   /1  5    �� Ky    �  � N�� �  �   �   1  y   b� S�� �   �   1   �  V� �  �   �   1  �    S	 !4�  � g�� �  !  $!  1  �    \+  x �  <!  L!  1  �  �    �4 �� �  d!  j!  1   �  ��	 y  �!  �!  1   0  �h� y  �!  �!  1   Y
 �  �   �!  �!  1   � ��� �   �!  �!  1    ��� �   �!  "  1  �   	 ��� "  )"  1  �  1   6 �E� �  A"  G"  1   iend �� �  _"  e"  1   �  ��    /  �y  T L)  q� �"    A� �"  �g l� �0  �"  �"  �0  �0   T L)  H �  =� �u  X �� 
#  R�"   fget 
�
 �0  
#  1   Tag �  T �"   �� \#  �	 �� �0  B#  �0   T L)  �� �0  �  �0   TG� �+  T� �7�  T� �7�  a#� %  0� �� �#  �#  �3   0� ׁ �#  �#  �3  �  ^0   0� I� �#  �#  �3  ^0   g0� !�� $  $  �3  �3   0� #E� %$  0$  �3  �3   /� (�� E$  P$  �3  5    'Gp -
�  4  i$  t$  �3  �#   7� 2�� �$  �$  �3   �� 8�� �$  �$  �3   '�� >U� �  �$  �$  �3   '<� Bn� �  �$  �$  �3  M0   F� G	M0   �� H�  v� �/   �#  �� ��  t 

*w �'  H%  T 5   �'  �'   6�~ �� o%  F �	  5   �  m1   6nk �Au �%  F �  �'  �  �1   6�~ ��} �%  F �	  �'  �  m1   0 
E �0  �%  Tag �  T �"  1   I�� 3� &  T S   F �	  ,(  m1   I~� 3�� ;&  T 5   F �	  �'  m1   I'i 3Ee e&  T �'  F �  nQ  �1   Ixy 3} �&  T �'  F �	  nQ  m1   A� 4  �&  T |-  E� �  J�O  �&  .�'  .�b   KU  �'  �&  8�b   A8� 4  #'  T |-  E� �  J�O  '  .�'  .�c   KU  �'  '  8�c   6 � �� N'  T L)  E� �  KU  �0   U� 

�� Y  t'  T |   Y  Y   c# 
	
l� Y  T |   Y  Y    2�  	 EJ     Z   �'  2�  	h�K     <  �'  /  �'  <   85   �  8/  /  �  5   5   �  (  jLn �  juh �  !�i Z   !Jf 2|	  	EJ     D�n j/  x �(  kx 
Xx v(  |(  j/   C�g y �(  j/  �'    �n �(  k�n �q �(  �(  p/   C�g <l �(  p/  �'    l�w +�v �	  l�r ,�p �  <y� 5   
!)  #��  #]� #��  <�
 5   L)  #��  # #=� #�  m�� pL)  C-  >�   ��� `4   �� 0K� �)  �)  �0  )4   /��  �)  �)  �0  q4   0Gp x� �0  �)  �)  �0  q4   �> @@� L)  �)  �)  �0  5    � L�� *  *  �0   �=9 #G� 5   L)  /*  5*  �0   �1 V 5   M*  b*  �0  M   k   G4   x� ��	 5   z*  �*  �0  �'  k   G4   �� �� �*  �*  �0  S    g� ��� 5   �*  �*  �0  !)    ��� �*  �*  �0   i� �w 5   +  	+  �0   b �X 5   !+  ,+  �0  M4   H� �� 5   E+  U+  �0  �  5    ?,	 2�� 5   L)  v+  �+  �0  ;4   ?�� 3; 5   L)  �+  �+  �0  A4   ?� 41� 5   L)  �+  �+  �0  M   k   G4   ?u� 5�� 5   L)  ,  ,  �0  �'  k   G4   ?� 6�  5   L)  :,  O,  �0  �  5   M4   (u� �� 5   i,  o,  �0   (�� )�� 5   �,  �,  �0   (�� 3< 5   �,  �,  �0   (k� U� 5   �,  �,  �0   (�� f�� 5   �,  �,  �0   
� wF� -  -  �0   � B�(  H�� C!)  L� D%)4  P� H(%  X L)  Et-  NM $�   m !9  �f 'Z-   OH-  m�� xKL)  d/  >L)   n�� �
 �-  �-  4  4   n��  �-  �-  4  #4   $�� �v� �-  �-  4  5   )4   �fd ��� 5   	.  .  4   �=9 ��  5   |-  1.  7.  4   @,	 ��� 5   |-  Y.  d.  4  ;4   @�� ��� 5   |-  �.  �.  4  A4   @� �� 5   |-  �.  �.  4  M   k   G4   @u� �z 5   |-  �.  �.  4  �'  k   G4   @� �c
 5   |-  !/  6/  4  �  5   M4   �_fd \5   p��� *  |-  X/  4  5     |-   T(  �(  9�  9�    �/  �    9�  -� H0  -� �� �/  �/  M0   /-� � �/  �/  M0  X0   0Gp �� ^0  �/  0  M0  X0   7� �� 0  0  M0   �� �� 30  90  M0   n� 5     �/  �/  M0  H0  �/  >� �0  imap x� �   �0  �0  �0  k    Cɒ   �� �0  �0  �   k     d0  L)  �0  �  �0  %S   �0  &|    9M-  �  �"  �0  L)  �"  �"  J  9  1  9  2f-  	��K     �  /1  �   :1  �   �  �	  Q1  �	  \1  U  �	  �  s1  �  ~1  �  �1  �  �1  3  �  E%2  Ky �|-  K� �|-  K: �|-  P� �	2  �� ��1  �1  \2   �K �2  \2  5     K� ��1   ���1  2�1  	��K     2�1  	@�K     2�1  	��K     �1  \2  22  	8�K     Ux  �	�K     U�  �	�K     U�  �	�K     *  �2  �  *  �  �2  �  �  �  �2  
  �2  �  
  �2  3  3  �  3  Z  3  �  Z  �2  �  83  e  d0  �  �  %w   k3  &|    [3  5g� �  5!�   5��   5K� X  o?� f   �o�� �   �5� �     5݉ �  %e  �3  &|    �c  .d  �b  �b  �#  �3  %  8�#  �#  .  �  |-  4  8|-  d/  /4  �;4  �0   �(  !)  k   �  �5   `4  � f4  ��� S4  C-  �Z  �   9�  9�  �� �G            ��M  �G     �       ��4  	<  w5   �l	  w5   �h VE/  K�4  5  �  4  0  <     �4  � '5  �G     +       �05  �4  �h  �4  V� S5  �G     -       �\5  �4  �h d
  {5  �hF     �       ��5  �  b1  �hs 	'S   �d ""%  O`F     (       ��5  T 5   a 
�'  �hb 
#�'  �` ;  ��F     1       ��5  D� Z�2  �h �  G     �      �)7  P �	  T 5   H Nm1  ����  N$5   ��s N1�  ���s N?5   ����  O5   ��H� O5   ��ZX  O#S   ��]� P�'  �XB� S)7  ��k T5   ���G     E       �6  i a5   �l JG     -       	7  i d5   �h wG     0       i f5   �d  %S   97  &|    �  RgF     �      �e8  P �	  T �   H Nm1  ����  N$�   ��s N1�  ���s N?5   ����  O5   ��H� O5   ��ZX  O#S   ��]� P�'  �XB� S)7  ��k T5   ��BhF     E       "8  i a5   �l �hF     -       E8  i d5   �h �hF     0       i f5   �d    �8   �F     �      ��8  �  !3  ��3n �2  ��
u �2  �X
v �2  �P
w �2  �H �  �8  `�F     �      �19  �  !3  ��3n ��2  ��
u ��2  �X
v ��2  �P
w ��2  �H "�  Q�F            �c9  T �  D� '�2  �h "�  B�F            ��9  T *  D� '�2  �h �  �9  ��F     �      ��9  �  �2  ��3n �2  ��
u �2  �X
v �2  �P
w �2  �H �  :  �F     �      �a:  �  �2  ��3n ��2  ��
u ��2  �X
v ��2  �P
w ��2  �H �  ��F     1       ��:  D� Z�2  �h �  �:  ҿF     V      ��:  �  �2  �Xn ��2  �PS� ��2  �h� ��2  �` �  ��F            �;  j =�2  �h �  -;  �F     �      �<  �  !3  ��3n x�2  ��S� {�2  �P
s ��2  �X
� ��  ����F     �       �;  
x ��2  �H ݻF     z       �;  
x ��2  �@ ��F     Q       �;  0� ��2  �� ҾF     Q       0� ��2  ��     ��F     1       �6<  D� U�2  �h 	  ~G     �       ��<  P �	  T 5   H xm1  �X��  x!5   �T�s x-5   �P��  x85   �LH� y5   �HZX  yS   �D�G     ;       �f {	�   �l  �  ��F            �=  j L�2  �h I  %=  Z�F     H       �R=  �  !3  �X	D� #�2  �P�� $�2  �h "g  D�F            �}=  j 8�2  �h :  �=  �F     V      ��=  �  !3  �Xn ��2  �PS� ��2  �h� ��2  �` )  �=  εF            �>  �  !3  �h	D� �2  �` �  />  ��F            �L>  �  �2  �h	D� �2  �` �  k>  f�F     H       ��>  �  �2  �X	D� #�2  �P�� $�2  �h 0  I�F            ��>  j =�2  �h v  �>  ��F     �      ��?  �  �2  ��3n x�2  ��S� {�2  �P
s ��2  �X
� ��  ��U�F     �       Q?  
x ��2  �H q�F     z       u?  
x ��2  �@ �F     Q       �?  0� ��2  �� f�F     Q       0� ��2  ��  �  T�F     1       ��?  D� U�2  �h �  6�F            �@  j L�2  �h "   �F            �A@  j 8�2  �h 7  O@  }@  �  �2  *� �   *� �%�   *�� �6k     A@  ֭ �@  ~�F     K       ��@  O@  �hX@  �dd@  �Xp@  �P �  �@  F�F     7      �A  �  �2  �HS� ��2  �@D� �"�2  ��L� ��2  �X �  :A  �F     7      �uA  �  �2  �HS� ��2  �@D� �!�2  ���� ��2  �X �  �A  ��F     j       ��A  �  �2  �hD� |�2  �`   �A  �A  �  �2  *� ��   *�� �)k   *�� �65     �A  �� B  @�F     d       �0B  �A  �h�A  �`�A  �X�A  �T z  OB  ��F     �      ��B  �  !3  ��	D� �2  ��	�  �2  ��S� �2  �X�  �2  �P�� �2  �H �  ��F            ��B  j I�2  �h �  �B  4�F     a      �YC  �  !3  ��	D� D�2  ��	0� D$�2  ���� E�2  �XL� F�2  �PS� Z�2  �H B	  �G     �       ��C  T 5   F �	  ݰ  �5   �lfo �/�  �`H �6m1  �X �  �C  �\F     �       ��C  �  �1  �hstr 	1�'  �`   
D  ��F     7      �ED  �  !3  �HS� ��2  �@D� �"�2  ��L� ��2  �X �  ݤF            �pD  j E�2  �h �  �D  ��F     7      ��D  �  !3  �HS� ��2  �@D� �!�2  ���� ��2  �X �  ��F            ��D  j B�2  �h 1@  E  `�F     (       �;E  �  3  �ha �!�2  �`b �1�2  �X �  ZE  ��F     j       �vE  �  !3  �hD� |�2  �` 1  �E  �F            ��E  �  !3  �h *  �E  X�F     �      �!F  �  �2  ��	D� �2  ��	�  �2  ��S� �2  �X�  �2  �P�� �2  �H ~  9�F            �LF  j I�2  �h P  kF  ؝F     a      ��F  �  �2  ��	D� D�2  ��	0� D$�2  ���� E�2  �XL� F�2  �PS� Z�2  �H d  ��F            ��F  j E�2  �h J  ��F            �!G  j B�2  �h 1�  @G  ��F            �MG  �  �2  �h �
  lG  �eF     �       ��G  �  b1  �hstr 	1�'  �` "�"  �G            ��G  p 
%1  �h �  �G  �G     <      �sH  �  �1  ��	m  �1�   ��	�  �Ak   �� �|   �X
slb ��2  �P
bkt �C3  �HY  �	k   �@� ��#  ��O� ��  ��ݰ  ��2  �� �  �H  N�F     �       ��H  �  �1  �H	R� %8k   �@ +�   �X
fra -�2  �P t$  �H  �F     L       ��H  �  �3  �h   I  �F     �       �GI  �  3  �X	D� ��2  �P�� ��2  �h �  fI  ʙF     D      �J  �  �1  ��	�N  45   �� 
�   �@Y  |   ���� 	k   �X
slb �2  ��N� �2  �P��F     ^       
off k   �H��F     >       ݰ  �2  ��   �  ;J  r�F     X       �WJ  �  !3  �X�� p�2  �h Z  vJ  ��F     �       ��J  �  !3  �H	D� �2  �@�� �2  �h� �2  �`&�F     I       �� �2  �X  H%  NG     J       �&K  F �	  ݰ  �5   �Lfo �/�  �@H �6m1  �� o%  z\F     *       �vK  F �  ݰ  � �'  �hfo �7�  �`H �>�1  �X W  �K  F     �       ��K  �  >3  �X	D� ��2  �P�� ��2  �h 1�  �K  x�F     I       �
L  �  �2  �Xp ��   �Padr �	|   �h �  L  "L  �  �2   ,
L  �� EL  b�F            �NL  L  �h �$  mL  �F     O       �zL  �  �3  �h 
  �L  V�F     �       ��L  �  �2  �H	D� �2  �@�� �2  �h� �2  �`ƖF     I       �� �2  �X  �  M  ��F     �       �DM  �  �1  �X	 �6�   �P�� ��2  �h 0$  RM  eM  �  �3  0  <     DM  �� �M  f�F     '       ��M  RM  �h �#  �M  �M  �  �3  *G� ^0    �M  �� �M  4�F     2       ��M  �M  �h�M  �` �%  eF     *       �9N  F �	  ݰ  � �'  �hfo �7�  �`H �>m1  �X 1�"  XN  4G            �rN  �  �0  �hx �0  �` �%  G            ��N  Tag �  T �"  p 
1  �h   �N  �G     1       ��N  �  y1  �h	m  _�   �`	�  _(k   �X �%  �G     G       �AO  T S   F �	  	ݰ  3,(  �H	H 3!m1  �@ �  `O  pG     0       �|O  �  51  �hptr -y  �` 1�  �O  NG     "       ��O  �  @1  �h�L 9$E1  �` %  �O  �F     �      ��P  �  �1  ��~ss  �1k   ��~$�F     �      �P  �N  �5   �\
bkt C3  �P� �#  ��ݰ  �2  ����F     *      oP  
slb 	�2  �H ƏF     �      
slb 	�2  �@�� #�#  ��  ԑF     �       R� :|   ��
fra ;�2  ���� =�#  ��~  &  
G     C       �3Q  T 5   F �	  	ݰ  3�'  �H	H 3!m1  �@ V  RQ  T\F     &       �nQ  �  �1  �h�d 	M�'  �` �'  ;&  �[F     E       ��Q  T �'  F �  	ݰ  3nQ  �H	H 3!�1  �@ �  �Q  �Q  �  �1  *$s 	�1   ,�Q  �u R  �[F     4       �R  �Q  �h�Q  �` s  5R  |�F     h      ��R  �  �1  ��~	m  ~+�   ��~ �|   �X�� ��#  ��
fra ��2  �P
slb ��2  �H
bkt �C3  �@Y  �	k   ��� ��#  ��O� ��  ��ݰ  ��2  �� x  S  �dF     &       �$S  �  W1  �h�d 	M�'  �` e&  ndF     E       �nS  T �'  F �	  	ݰ  3nQ  �H	H 3!m1  �@ �	  |S  �S  �  b1  *$s 	Q1   ,nS  �z �S  :dF     4       ��S  |S  �h�S  �` �  �S  �S  �  51  *�� 2y   ,�S  X� T  �G            �T  �S  �h�S  �` �0  "�  �G            �TT  T T  x *T  �h W  sT  �G     0       ��T  �  1  �hptr %y  �` "(#  �G            ��T  �5  �0  �h q  �T  �T  �  �'  0  <    ,�T  Gk �T  �[F            �U  �T  �h W  U  U  �  �'   ,U  �t BU  �[F            �KU  U  �h �  �&  SG     �       ��U  T |-  E� �  J�O  �U  .�'  .�b   @� KU  ��p+�U  �'  �&   m  �   �H�	 +�'  �� 	 +�&  �� <  "  EG            �V  T �b  x .�U  �h �&  �
G     �       ��V  T |-  E� �  J�O  XV  .�'  .�c   @� KU  ��p+{V  �'  '   m  �   �H�	 +�'  �� 	 +'  �� i  "H  �G            ��V  T �'  x .�V  �h �  "u  �
G            �W  T �c  x .�V  �h #'  JG     G       �aW  T L)  E� �  @� KU  �hm  (�0  �` �
  �W   G     *       ��W  T S   �  b1  �hݰ  	S   �d 1�  �W  G            ��W  �  @1  �h ?   �W  �G     2       ��W  �  51  �h    X  �G     (       �6X  �  @1  �h�L <$E1  �` G"  UX  �G     #       �bX  �  1  �X )"  �X  \G     3       ��X  �  1  �X �  �X  ��F     (       ��X  �  y1  �h	�  [k   �`   �X  4G     (       �Y  T 5   �  b1  �hݰ  	5   �d �   "N'  �F     +       �OY  T |   a 
Y  �hb 
#Y  �` "t'  	G     +       ��Y  T |   a 
	Y  �hb 
	#Y  �` s  �Y  T[F     ,       ��Y  �  �1  �hLn	  �    �Y  [F     )       �Z  T �'  �  �1  �hݰ  	�'  �` T  Z  #Z  �  �1  0  <    ,Z  �t FZ  �ZF            �OZ  Z  �h 8  nZ  �ZF     )       �{Z  �  �1  �` �!  �Z  *G     �      ��Z  �  1  ��it ��  ���@ ��   �H� �y  �P�� ��   �X �   [  �G     a       �[  �  1  �Xptr N&y  �P >  >[  ��F     )       �[[  �  y1  �h	m  c�   �` >  ��F     �       ��[  �  W0k   ��tc Y|   �`e b|   �Xf c|   �Pip d|   �His e|   �@��F     :       i [�   �l  "$  �F            �Z\  idx H6�   ��tc J|   �hs O5   �dip P|   �Xis Q|   �Pf R|   �H A
  y\  dF     ,       ��\  �  b1  �hLn	  �  .  �\  �cF     )       ��\  T �'  �  b1  �hݰ  	�'  �` "
  �\  �\  �  b1  0  <    ,�\  _| ]  �cF            �]  �\  �h Z  <]  �cF     )       �I]  �  W1  �` !  h]  ,G     �      ��]  �  1  �H��  g#�   �@�
 iy  �X �  �]  �]  �  �0   ,�]  �� �]  G     *       ��]  �]  �h �   �]  �]  �  1   ,�]  j ^  �G     "       �^  �]  �h   )^  ?^  �  �'  *�L *�'    ^  [q b^  vZF     V       �s^  )^  �h2^  �` H  �^  �^  �  �'  0  <     s^  r �^  ZZF            ��^  �^  �h �  �^  �^  �  �'    �^  �d �^  6ZF     #       �_  �^  �h q t~
G     5       �D_  	�S t�  �X�� u�0  �h - n5   <
G     B       ��_  3c n5   �\	�S n�  �P�� o�0  �h qe� h�	G     R       ��_  	�S h�  �X�� i�0  �h -� N5   �G           ��`  	�S N�  �H	B� N$M   �@	�� N05   ��	�  N=k   ���� P�0  �h	G     @       o`  
e R
5   �d N	G     9       �`  
e W
5   �` �	G     9       
e \
5   �\  -� J5   �G            ��`  	�S J�  �h -� D5   nG     I       �,a  	�S D�  �X�� E�0  �h -b :�   G     i       ��a  	�S :�  �H�� ;�0  �h/ <�  �X+G     =       
e =	5   �d  -�a 15   �G     r       �$b  	�S 1�  �X	x  1!�   �P	�� 1-5   �L�� 2�0  �h�G     >       
e 3	5   �d  -�a &5   G     �       �vb  	�S &�  �X�� '�0  �`
e (5   �l -�� �  uG     �       �tc  3fd 5   ��~	�� "�'  ��~e� #r�� �b  �b  �3  5    s�g  c  G     *       �c  �b  o� Lc  �h	�� #�0  �` t� )4  @c  dG            �Rc  �  Lc  �h�3   u� DG            �L�0  �h   -�a ��  �G     Q      ��d  	xF ��'  ��}	�� �+�'  ��}?1  �5   �l`� ��  �k
fd 5   ��}P� �d  r�� d  d  �3  5    s�g 3d  nG     *       �Pd  �c  o� d  �h	�� �0  �` t� )4  sd  �G            ��d  �  d  �h�3   u� �G            �L�0  �h  �G     C       
e 	5   �d  -�� �5   SG            ��d  	�S ��  �h -�� �5   G     4       �?e  	�S ��  �X�� �4  �h �1  Me  �e  �  b2  0  <   Wvit ��0  X�� 1  X0 �  X; �  Wve �5      �?e  �e  6G     �       �@f  Me  ��~w_e  �e  :`e  :le  :ue  :~e  ��e  :�e    Y_e  HG     �       ;`e  �`;le  �h;ue  ��~;~e  ��~Y�e  �G     [       ;�e  �\   �1  Nf  Xf  �  b2   �@f  xf  *G            ��f  Nf  �h �.  �f  �G     E       ��f  �  4  �X	x  ��  �P	�� �(5   �L	2� �7M4  �@�G     '       
e �	5   �l  �.  g  �G     U       ��g  �  4  �X	B� �#�'  �P	]�  �2k   �H	/ �DG4  �@
s �
�   �`�G     (       
e �	5   �l  �.  �g  8G     U       �h  �  4  �X	B� �M   �P	]�  �+k   �H	/ �=G4  �@
s �
�   �`PG     (       
e �	5   �l  d.  0h  D G     �       ��h  �  4  ��~	�� �-A4  ��~+w �h  	�bJ     � G     �       
e �	5   �l  %Z   �h  &|    �h  7.  �h  ��F     h       ��h  �  4  �X	� �*;4  �Px  ��  �`
e �5   �l .  i  B�F     �       �>i  �  4  ��~��F            
e �	5   �l  1�-  ]i  0�F            �ji  �  4  �h �-  xi   �i  �  4  �fd �5   �� �!)4    ji  � �i  ��F     E       ��i  xi  �h�i  �d�i  �X �,  �i  t�F     u       �(j  �  �0  �X+w 8j  	�bJ     
ptr |�   �h %Z   8j  &|    (j  �,  \j  ��F     �       ��j  �  �0  �X+w �j  	�bJ     ��F            
e g	5   �l  %Z   �j  &|    �j  �,  �j  ��F            �Uk  �  �0  ��~��F             k  
e V
5   �l ��F     �       2� Z	�  ��~{ [�   �`��F     �       
e \5   �\   �,  tk  ��F     �      �@l  �  �0  �H+w Pl  	xbJ     ��F            �k  
e 4	5   �l ��F     Z       �k  2� =	�  �X��F     J       
e >
5   �h  ��F     �       I� H
k   �P��F     i       
e I
5   �d   %Z   Pl  &|    @l  o,  tl  �F     �       ��l  �  �0  �h+w �l  	hbJ      %Z   �l  &|    �l  O,  �l  ��F            �m  �  �0  �X+w m  	XbJ     ��F     0       
e #	5   �l  %Z   m  &|   
 m  ,+  <m  |�F           �n  �  �0  �H	x  �  �@	�� +5   ��2� 	�  �P+w 'n  	ObJ     ��F            �m  
e 	5   �l ��F     e       �m  { �   �`��F     D       
e 
5   �\  B�F     @       
e 
5   �X  %Z   'n  &|    n  	+  Kn  �F     n       ��n  �  �0  �X/ � M4  �P{ ��  �`�F     3       e �	5   �l  �*  �n  ��F     h       �o  �  �0  �X��F            �n  e �5   �l ��F            e �
5   �h  1�*  "o  f�F     ?       �/o  �  �0  �h �*  No  �F     T       �}o  �  �0  �h�� �/!)  �d+w �o  	@bJ      %Z   �o  &|    }o  �*  �o  ��F     m       ��o  �  �0  �hc � S   �d+w �o  	:bJ      %Z   �o  &|    �o  b*  p  ��F     �      �-q  �  �0  ��~B� �&�'  ��~]�  �5k   ��}/ �GG4  ��}+w �o  	4bJ     s �|   ��~% ��  �oc�F     �       �p  I� �
k   ��~��F     Y       e �
5   �h  W�F             �p  e �
5   �d w�F             q  e �
5   �` ��F     @       nl �M   �X  5*  Lq  @�F     �      �xr  �  �0  ��~B� VM   ��~]�  V.k   ��~/ V@G4  ��~+w 'n  	/bJ     s �|   �X��F     �       �q  I� \
k   ��~��F     Y       e ]
5   �l  ��F           I� x
k   ��~��F             4r  e q
5   �h �F             Wr  e s
5   �d @�F     a       e y
5   �`   �)  �r  �F     /       ��r  �  �0  �h �)  �r   �r  �  �0  0  <   W�it H�     �r    �r  ��F     +       ��r  �r  �h  �r   "s  ��F     �       �Zs  �r  ��~w�r  :s  :�r   Y�r  �F     �       ;�r  ��~  n)  hs   ~s  �  �0  *� 0%)4    Zs  � �s  $�F     �       ��s  hs  �hqs  �` 10  �s  �F            ��s  �  S0  �h 0  �s  րF     B       �t  �  S0  �h+w 'n  	*bJ      "�  ÀF            �Ft  x )|   �h   Tt  ^t  �  �/   ,Ft  �� �t  r�F     Q       ��t  Tt  �h V9  2�t  �t  �  (  0  <     �t  �o �t  ZF            ��t  �t  �h p  VV  2�t   u  �  (  �t    �t  �e #u  �YF     �       �4u  �t  �h�t  �` �  Bu  Lu  �  (    4u  w ou  &YF     \       �xu  Bu  �h �6r kv �   YF            ��u  �  #k   �hp /�   �` !&E !�
  ZL)  %  "Z*  \#  "Z�  \#  " �   �  t�n �H ~c ��         �) E�� 	5   uint 
5   E�� M   X   FM   +�  
X   E! M   $�$ (|   v�# �   -�   �   1�     +�i 
�   wZ  �   J�7  �    JF(  �   J�=  �   JFD  �    +�i 
�   x$�$ cp   $^� ��   
�   $]�   +X  {S @�  g
  M       	�   v  #	�   �  &	�   |
  )	�    h  ,	�   (�  -	�   0�	  25   8�  55   < $�
  8"  $HP 9�   
�  E  K�  �  F�  E�  L�  E�  M�  +�  
�  +�  +�  +-  $F �  $�  ��   $�@ /  $�  4  
0  +S  K�� e�   $:G  �  +�
  y�  zstd  `  9t �  =�\ g  $�l `  .�l =g �  �  �  u   .�g t �  �  �  u   T `  av `    
x  �v a  =�\ g  $�l `  .�g �o 	  -  3  �   .�g Vl 	  K  Q  �   T `  av `   
�  �s ��  =�\ �g  T 5   L�O  M=2    ;s ��  =�\ �g  T 5   L�O  MC2    �� `�  $� a5   T U2   � �  =�\ �g  T 5   L�O  M72    ,S �;  =�\ �g  T 5   L�O  MU2    �H `\  $� a`  T Ik   Nv ��q g  Nv ��e g  Nv � Y g  Nv �9+ g  �A 
K �  T `  Ik  Ik   $�� j>H  '�% 
!�' �  �  T Ik  Ik   � 
�)   T 5   U2  U2   '� 
q� U2  6  T U2  �   $�� j>�  W�9 
!�, 6  T U2  U2    +t 
`  B�d �  �  B6h �  a  {frg �0  X�� 	
�  |W� �   Y`� 	�  Z�  b� g    [�  O>� 5   �  %�r  cred %d�  l� 0�  l� �   %  �0   ?l� � 9  D  �0  �0   @Gp ;� �0  \  g  �0  �0   S� �    �  �   �� �   )�  �   �� !�    � "�  ( 
�  �� %  'J� ';� `  �  T &  [:   W�� '{� `  T �  r:    f� 5�
  dh 8`� �0  -  [:   'O� =t� [:  G  [:   '�� BͰ [:  a  [:   'n� E� [:  {  [:   ')� I�� [:  �  [:   '�� L7� [:  �  [:   .�� PE� [:  �  �  �:   P#� U�� `  �  [:   P�� Z؟ `    [:   � d�     �:   ?� g� 1  <  �:  �:   @Gp i;� �:  T  _  �:  �:   .N� o�� [:  w  }  �:   � |\� �  �  �:  [:   c� ��� �  �  �:  [:  [:   �� ��� �  �  �:  [:  [:   
� �6� �  	  �:  [:   2�� #� 	  '	  �:  [:   ,<� � =	  M	  �:  [:  [:   ,�� D� c	  s	  �:  [:  [:   ,�� x)� �	  �	  �:  [:   ,�� �$� �	  �	  �:  [:   ,/� �� �	  �	  �:  [:   2� u� �	  �	  �:  [:   2,� #E� 
  
  �:  [:   C0� 0�� `  0
  6
  �:   C0� 94� `  P
  j
  �:  [:  U2  �:  �:   A�� ��    D �
  T &  Q� ��  A �   
  <� �W  5�}  5��  5��  5�G  5�a  5��  \   2�� �\� �
    �:  /   2\+  ���   (  �:  [:   A�� �/  T &  Q� ��  L /  A �   _� 5�  dh 8� �0  }  r:   'O� =� r:  �  r:   '�� B� r:  �  r:   'n� E2� r:  �  r:   ')� I�� r:  �  r:   '�� L� r:  �  r:   .�� PK� r:      �:   P#� U� `  8  r:   P�� Zk� `  S  r:   � dg� g  m  �:   ?� g4� �  �  �:  �:   @Gp iI� �:  �  �  �:  �:   .N� o�� r:  �  �  �:   � |c� �  �  �:  r:   c� �)�     �:  r:  r:   �� ��� '  7  �:  r:  r:   
� �� L  W  �:  r:   2�� U� l  w  �:  r:   ,<� �� �  �  �:  r:  r:   ,�� Dz� �  �  �:  r:  r:   ,�� x�� �  �  �:  r:   ,�� �Z� �    �:  r:   ,/� ��   &  �:  r:   2� ;� ;  F  �:  r:   2,� #�� [  f  �:  r:   C0� 0�� `  �  �  �:   C0� 9�� `  �  �  �:  r:  U2  �:  �:   A�� ��    D �  T �  Q�  �  XA �   
W  IW� �5��  5��  5�  5��  5��  5��  \W   2�� �F� I  T  �:  /   2\+  �Q� i  t  �:  r:   A�� �/  T �  Q�  �  XL /  A �    Z�  b� g    [�  �� �  }clz � 5   �  �    T �    ~"� �$�  O"� 5   �!  %�r  %l� %[�  
�  � H�	�  � ��� G  \  [:  �  0  �    ?� �5� p  {  [:  f:   @Gp �
�� l:  �  �  [:  f:   .Z� �δ `  �  �  [:  �    � �!    �<  ss  �  "� �%*   
&  � ��	�  \&   � �E� "  7  r:  0  �   5    ?� ��� K  V  r:  }:   @Gp �r� �:  n  y  r:  }:   �N  �<   Hٖ ��   LU� ��:  P.� �%*  X 
�  '� �	*  '� ��� �  �  �:   ?'� �Ƈ �  �  �:  �;   @Gp �Ⱥ �;      �:  �;   ʊ ��:    
�  � �	a  e�g �a� `  P  �:  f:  f:    �0   �	�  �0  ��� �  �  �:   � �	�0   x� �r:  � ��   $�� �2*  �� �-� �  �  p9  �:   f�� (z� �  �  p9  �:   Gp *� ;       p9  �:    Wd ��� �   9  D  p9  �    C�6  L�� �   ^  n  p9  �   �    ,�N ~�� �  �  p9  �    ,� �w� �  �  p9  �   �     Y� 1	�� �   �  �  p9   �J� >;                         @       ]�� @ �   ]�� A �    'H� H�� �   9  �    'r� W�� �   S  �    ]�� j<   =� l  '�� o�� `  �  �    =o� |  =��   �� �   ^<� �7� [:  �  �  p9  0   ^a� �� r:  �  �  p9  5    ^P� %j� [:      p9  �    2`� 7� 3  9  p9   2� >� N  Y  p9  [:   Э �
�:   A� ��0  $ۧ �?*  @� �s  �� �	�    � �m;  (� �1  v� �0   
�  �0� V�  ,;� X� �  �  e9  p9   CWd [!� �       e9  �    ,� _ʅ )  9  e9  �   �    ,�N c�� O  Z  e9  �    C� gε �   t  �  e9  �   �    !�� lp9   � �1  v� �0   X/g 
�  g[r  �  ��t  �  ��q 72   Omi 5   ,  %�r  %�( chex  RMq {  ��h {_  �ݰ  |5   �h ~�q =  C  2   _�h h S  2  5     �s  u t  z  &2   �s p �  �  &2  �   �s �v �  �  &2  12   �s *o �  �  &2  72   �s *gs �  �  &2  =2   �s 0dr     &2  C2   �s 8�m /  :  &2  5     Gp =�w I2  S  ^  &2      �s Qr `  w  }  O2    �s T�i `  �  �  &2    ]h X%d `  �  �  O2    p \Xw 12  �  �  O2    p `�k U2  �  �  &2    �o d�g [2      &2   �� ��s ,  2  &2   wq �   �r �`  A= %�( h  s  U U2  &2  U2   T 5    
  ,s 2h  ,s 3�s �  �  a2   .#m 6Rf �  �  �  a2  �   (m <�   �m =5   H� >  �t ?`  v @`  �r A`  ;f B`  �u C`  +s �n C  N  a2  5    �,s  i \  a2  �    
�  Y/f J�#  � N�� �  P (  T 5   �3  5   `  5   5   5   X    �� Nm{ �  P (  T �   �3  �   `  5   5   5   X    B~ xR :  P (  T �   �3  �   5   5   5   X    @  x� w  P (  T 5   �3  5   5   5   5   X    *y �� �  T �   F (  �   �  �3   � �i� �  T 5   F (  5   �  �3   $M N�7   P �5  T �2  �B  �2  `  5   5   5   X    �N N�G W  P �5  T �   �B  �   `  5   5   5   X    =. N� �  P �5  T   �B    `  5   5   5   X    / N~/ �  P �5  T �   �B  �   `  5   5   5   X    U N�1   P a4  T �2  �K  �2  `  5   5   5   X    }F N�> _  P a4  T �   �K  �   `  5   5   5   X    � N�' �  P a4  T   �K    `  5   5   5   X    ! N<5 �  P a4  T �   �K  �   `  5   5   5   X    �. NG8 %  P 5  T �2  fP  �2  `  5   5   5   X    :Z NO0 g  P 5  T �   fP  �   `  5   5   5   X    a N� �  P 5  T   fP    `  5   5   5   X    �O N�@ �  P 5  T �   fP  �   `  5   5   5   X    rL N�' -  P �3  T �2  mU  �2  `  5   5   5   X    �M N�F o  P �3  T �   mU  �   `  5   5   5   X    �- N�0 �  P �3  T   mU    `  5   5   5   X    #' N�J �  P �3  T �   mU  �   `  5   5   5   X     x[ 0   P �5  T �2  �B  �2  5   5   5   X    �, x�F m   P �5  T �   �B  �   5   5   5   X    C x�U �   P �5  T   �B    5   5   5   X    � x�% �   P �5  T �   �B  �   5   5   5   X    gG xYY $!  P a4  T �2  �K  �2  5   5   5   X    � x�* a!  P a4  T �   �K  �   5   5   5   X    �@ x�3 �!  P a4  T   �K    5   5   5   X    �% x�* �!  P a4  T �   �K  �   5   5   5   X    L x�G "  P 5  T �2  fP  �2  5   5   5   X    LF x[ U"  P 5  T �   fP  �   5   5   5   X    ! xkB �"  P 5  T   fP    5   5   5   X    `* xR1 �"  P 5  T �   fP  �   5   5   5   X    �1 x�A #  P �3  T �2  mU  �2  5   5   5   X    �+ x I#  P �3  T �   mU  �   5   5   5   X    � x�> �#  P �3  T   mU    5   5   5   X    �3 xj+ P �3  T �   mU  �   5   5   5   X     �A ��#  ��  �
�     O~5 5   �$  %�  %�H %�H %
#  R�� �%  � y� )$  /$  �2   � �� D$  O$  �2  �1   � �� d$  t$  �2  �1  �     �U  !� �1  �$  �$  �2    d  #U� �2  �$  �$  �2  �     �  '	�� �   �$  �$  �2    �� +� `  �$  �$  �2  $    �� 3�� `  %  %  �2  $    I� 7	�� �   7%  G%  �2  X   �     f� ?	j� �   `%  k%  �2  X     �� G�� $  �%  �%  �2  �   �    m  X�1   rs  Y	�   7�  X    
$  R�Q n'  � �3 �%  �%  �2   � �Q �%  &  �2  �2   � !D &  *&  �2  �2  �     �U  DL �2  C&  I&  �2    d  #=* �2  b&  m&  �2  �     �  '	�$ �   �&  �&  �2    �� +KK `  �&  �&  �2  �%    �� 3� `  �&  �&  �2  �%    I� 7	j- �   �&  �&  �2  �2  �     f� ?	� �   '  !'  �2  �2    �� G�K �%  :'  J'  �2  �   �    m  X�2   rs  Y	�   7�  �2   
�%  <�� �'  2�� "=� �'  �'  �2  �2  �    AA� &�2   AV� '	�    
s'  XDq 	

�'  g�g 	�'  `d 	*  s 	E�x (  (  �3  3   j �		�)  j 	| 1(  <(  �3  �3   ?j 	*{ P(  [(  �3  �3   @Gp 		@� �3  s(  ~(  �3  �3   j 	 �(  �(  �3  5    .Cr 	"	�z �3  �(  �(  �3  �'    i 	'�} �(  �(  �3  X     i 	1Wz �(  �(  �3  �1   /#s 	>�3   /A� 	?{3  /�� 	@
�   �/m 	A`  �.�
 		�� �3  U)  `)  T X   �3  X    .�� 		� �3  )  �)  T s'  �3  s'   e�m 		�~ �3  �)  T �1  �3  �1    
(  .�g 	Hx (  �)  �)  �3   �l 	Mox �)  �)  �3  �1   /cg 	Q3   �n 3  ��! �   � hXt ��$ KG� �+�  K� �7�  K� �7�
  R#� �+  0� �� n*  t*  };   0� ׁ �*  �*  };  �  �1   0� I� �*  �*  };  �1   f0� !�� �*  �*  };  �;   0� #E� �*  �*  };  �;   /� (�� +  +  };  5     Gp -
� �;  2+  =+  };  L*   7� 2�� R+  X+  };   �� 8�� m+  s+  };    �� >U� `  �+  �+  };    <� Bn� `  �+  �+  };  ~1   F� G	~1   �� H`  v� �0   
L*  't 
*w 12  ,  T 5   12  12   �~ ��| ,,  F (  �   �  �3   �~ �� S,  F (  5   �  �3   (�{ 82� �,  T �   F (  ~\  �  �3   (�� 3� �,  T X   F (  �2  �3   (6X ��O �,  F �5  �B  X   �  �#  �7   (�H qE -  F �5  �B  X   �  �#  �7   (VX 'B B-  F �5  �B  X   �  �#  �7   (�~ � j-  F (  s'  �  �3   �~ ��} �-  F (  �1  �  �3   (�V ��< �-  F a4  �K  X   �  �#  �7   (t. q�8 �-  F a4  �K  X   �  �#  �7   (R' '�C '.  F a4  �K  X   �  �#  �7   (d$ �P= Y.  F 5  fP  X   �  �#  �7   (,K qM; �.  F 5  fP  X   �  �#  �7   (�! 'Z( �.  F 5  fP  X   �  �#  �7   (DO �� �.  F �3  mU  X   �  �#  �7   (� q]D !/  F �3  mU  X   �  �#  �7   (qO ' S/  F �3  mU  X   �  �#  �7   �8  i� n/  I2  I2   (�� 3\� �/  T s'  F (  ��  �3   (xy 3} �/  T �1  F (  K�  �3   �T �3@ �/  A {9  {9  �1  �7   �5 �'C 0  A �8  �8  �1  �7   '# 	
l� #�  60  T �   #�  #�   uX �� ]0  A �7  �7  �1  �7    �& �0  A �6  �6  �1  �7   WU� 
�� #�  T �   #�  #�    D�  D�  �  
�0  �  �  D�  -� y1  -� �� �0  �0  ~1   ?-� � 1  1  ~1  �1   @Gp �� �1  +1  61  ~1  �1   7� �� J1  P1  ~1   �� �� d1  j1  ~1   /n� 5     
�0  �0  
~1  y1  �0  >� �1  �map x� 0  �1  �1  �1  �    _ɒ   �� �1  �1  0  �     �1  `�  	%cJ     _   
�1  F�1  `�  	p�K       
2    
&2  <   )5   {  )    {  5   5   �  
a2  SLn s  Suh �  +�i $  
�2  �%  
�2  _   �%  
�2  �2  F�2  +Jf 
�2  n'  
�2  �2  s'  
�2  �2  �`�'  	7cJ     Y�n o3  x I3  �x 
Xx '3  -3  o3   _�g y =3  o3  �1    i�w +�v �'  i�r ,�p *  h��  3  i3  -X   �3  1�    �'  
�3  (  
�3  �)  (  �5 DV4  �5 E�W �3  �3  V4  �    i HnE �3  �3  V4  X     i M 4  4  V4  �1    i R6 +4  ;4  V4  �1  �    Jy  W�   .� X	�    �3  
V4  z [
5  z \$? �4  �4  
5  M     i _iN �4  �4  
5  X     i d�J �4  �4  
5  �1    i l�O �4  �4  
5  �1  �    B� tM    .� u	�    a4  

5  �@ x�5  �@ y�H 65  F5  �5  M   �     i |@: Z5  e5  �5  X     i ��> y5  �5  �5  �1    i ��* �5  �5  �5  �1  �    B� �M    �� �	�   .� �	�    5  
�5  {W ��6  {W �� �5  6  �6   �@ �^ 6  6  �6    i �w3 06  ;6  �6  X     i �_M O6  Z6  �6  �1    i ��= n6  ~6  �6  �1  �    B� �M    �� �	�   .� �	�    �5  
�6  Z�6  ��   �
%'I  %�6 %}M %�N %M? %�, %� %4   [��6  �5 �7  � N% 7  ,7  �7  V4  �7   �g �< @7  K7  �7  X    �g �D _7  o7  �7  �1  �    �g �& �7  �7  �7  X   �  �#   /H @V4   /9 A�7  F �3   �6  
�7  �#  �P �8  � �E �7  �7  �8  �5  �7   �g � 8  8  �8  X    �g �@ 18  A8  �8  �1  �    �g ?A U8  j8  �8  X   �  �#   /H @�5   /9 A�7  F 5   �7  
�8  HS Z9  � �6 �8  �8  Z9  
5  �7   �g f) �8  �8  Z9  X    �g x9 �8  9  Z9  �1  �    �g �? !9  69  Z9  X   �  �#   /H @
5   /9 A�7  F a4   �8  
Z9  �  
e9  �  
p9  �4 <:  � 4 �9  �9  <:  �6  �7   �g \7 �9  �9  <:  X    �g �C �9  �9  <:  �1  �    �g R4 :  :  <:  X   �  �#   /H @�6   /9 A�7  F �5   {9  
<:  S�3 �  SAG   &  
[:  �  &  �  
r:  �  �  �  
�:    
�:  �
    [:  /  
�:  �
  
�:  W  
�:  �  W  r:  �  
�:  a  �1  �  �  -  ;  1�    
;  Bg� �  B!�   B��   BK� S  j?� a   �j�� �   �5� �     B݉ �  -a  };  1�    L*  
};  �+  )L*  L*  *  �  D\  Dn  D�  D�  y  G     �      ��<  P (  T 5   H N�3  ����  N$5   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   ���G     E       �<  i a5   �l JG     -       �<  i d5   �h wG     0       i f5   �d  -X   �<  1�    �  RgF     �      �">  P (  T �   H N�3  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   ��BhF     E       �=  i a5   �l �hF     -       >  i d5   �h �hF     0       i f5   �d  �  �fF     U       ��>  P (  T �   H x�3  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �T34�f {	�     :  ~G     �       �Y?  P (  T 5   H x�3  �X��  x!5   �T�s x-5   �P��  x85   �LH� y5   �HZX  yX   �D�G     ;       �f {	�   �l  w  afF     �       ��?  T �   F (  ݰ  ��   �lfo �/�  �`H �6�3  �X �	  �?  ��F     �      �@  	�  �:  ��n [:  ��u [:  �Xv [:  �Pw [:  �H �	  5@  �F     �      �|@  	�  �:  ��n �[:  ��u �[:  �Xv �[:  �Pw �[:  �H �  T�F     1       ��@  D� U[:  �h -  I�F            ��@  j =[:  �h 6�  B�F            �A  T &  D� '[:  �h 6�  Q�F            �6A  T �  D� 'r:  �h   UA   �F     �      ��A  	�  �:  ��n r:  ��u r:  �Xv r:  �Pw r:  �H �  �A  `�F     �      �B  	�  �:  ��n �r:  ��u �r:  �Xv �r:  �Pw �r:  �H 8  ��F     1       �-B  D� Zr:  �h �  �G     �       ��B  T 5   F (  ݰ  �5   �lfo �/�  �`H �6�3  �X 6�+  O`F     (       ��B  T 5   a 12  �hb #12  �` �5  �  ��G     �      ��C  P �5  T �2  H N�B  ����  N$�2  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       �C  i a5   �l E�G     -       �C  i d5   �h r�G     0       i f5   �d    ^�G     �      �E  P �5  T �   H N�B  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   ��N�G     E       �D  i a5   �l ��G     -       �D  i d5   �h ��G     0       i f5   �d  W  ��G     �      �KF  P �5  T   H N�B  ����  N$  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       F  i a5   �l ��G     -       +F  i d5   �h +�G     0       i f5   �d  �  �G     �      �wG  P �5  T �   H N�B  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ���G     E       4G  i a5   �l V�G     -       WG  i d5   �h ��G     0       i f5   �d  ,  FeF     J       ��G  F (  ݰ  �!�   �Lfo �8�  �@H �?�3  �� 7  �G  �F     V      �H  	�  �:  �Xn �r:  �PS� �r:  �h� �r:  �` �  6�F            �JH  j L[:  �h �	  iH  f�F     H       ��H  	�  �:  �XD� #[:  �P�� $[:  �h {  9�F            ��H  j I[:  �h 6   �F            ��H  j 8[:  �h �  I  ҿF     V      �CI  	�  �:  �Xn �[:  �PS� �[:  �h� �[:  �` �	  bI  ��F            �I  	�  �:  �hD� [:  �` &  �I  εF            ��I  	�  �:  �hD� r:  �` F  �I  Z�F     H       �J  	�  �:  �XD� #r:  �P�� $r:  �h }  ��F            �2J  j =r:  �h �  QJ  �F     �      �/K  	�  �:  ��n xr:  ��S� {r:  �Ps �r:  �X
� ��  ����F     �       �J  x �r:  �H ݻF     z       �J  x �r:  �@ ��F     Q       K  0� �r:  �� ҾF     Q       0� �r:  ��    ��F     1       �ZK  D� Ur:  �h �  ��F            ��K  j Lr:  �h 6d  D�F            ��K  j 8r:  �h a4  �  f�G     �      ��L  P a4  T �2  H N�K  ����  N$�2  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ��_�G     E       �L  i a5   �l ��G     -       �L  i d5   �h ��G     0       i f5   �d    ��G     �      �N  P a4  T �   H N�K  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   ����G     E       �M  i a5   �l �G     -       �M  i d5   �h 3�G     0       i f5   �d  _  �G     �      �:O  P a4  T   H N�K  ����  N$  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ���G     E       �N  i a5   �l g�G     -       O  i d5   �h ��G     0       i f5   �d  �  w�G     �      �fP  P a4  T �   H N�K  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ��p�G     E       #P  i a5   �l ��G     -       FP  i d5   �h ��G     0       i f5   �d  5  �  ��G     �      ��Q  P 5  T �2  H NfP  ����  N$�2  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       UQ  i a5   �l �G     -       xQ  i d5   �h D�G     0       i f5   �d  %  0�G     �      ��R  P 5  T �   H NfP  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   �� �G     E       �R  i a5   �l o�G     -       �R  i d5   �h ��G     0       i f5   �d  g  ��G     �      ��S  P 5  T   H NfP  ����  N$  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       �S  i a5   �l ��G     -       �S  i d5   �h ��G     0       i f5   �d  �  ��G     �      �U  P 5  T �   H NfP  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       �T  i a5   �l (�G     -       �T  i d5   �h U�G     0       i f5   �d  ,,  NG     J       �mU  F (  ݰ  �5   �Lfo �/�  �@H �6�3  �� �3  �  8�G     �      ��V  P �3  T �2  H NmU  ����  N$�2  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ��1�G     E       \V  i a5   �l ��G     -       V  i d5   �h ��G     0       i f5   �d  -  ��G     �      ��W  P �3  T �   H NmU  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��]� P�1  �XB� S�<  ��k T5   ����G     E       �W  i a5   �l ��G     -       �W  i d5   �h �G     0       i f5   �d  o  ��G     �      ��X  P �3  T   H NmU  ����  N$  ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ����G     E       �X  i a5   �l 9�G     -       �X  i d5   �h f�G     0       i f5   �d  �  I�G     �      �#Z  P �3  T �   H NmU  ����  N$�   ��s N1`  ���s N?5   ����  O5   ��H� O5   ��ZX  O#X   ��~]� P�1  �XB� S�<  ��k T5   ��B�G     E       �Y  i a5   �l ��G     -       Z  i d5   �h ��G     0       i f5   �d  �  ��G     W       ��Z  P �5  T �2  H x�B  �h��  x!�2  �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�2    0   ��G     U       �G[  P �5  T �   H x�B  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �T34�f {	�     m   ��G     �       ��[  P �5  T   H x�B  �X��  x!  �P�s x-5   �L��  x85   �HH� y5   �DZX  yX   �@%�G     ?       �f {	�   �h  �   ��G     W       �~\  P �5  T �   H x�B  �h��  x!�   �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�     �   S,  ��F     N       ��\  T �   F (  ݰ  8~\  �Hfo 8-�  �@H 84�3  �� �(  �\  �hF     �       �]  	�  �3  �hs 	'X   �d �(  7]  �eF     �       �S]  	�  �3  �hstr 	1�1  �` "3  a]  �]  �  a:  &� ��  &� �%0  &�� �6�    7S]  ֭ �]  ~�F     K       ��]  a]  �hj]  �dv]  �X�]  �P   �]  ��F     7      �-^  	�  �:  �HS� �r:  �@D� �"r:  ��L� �r:  �X �  L^  ��F     7      ��^  	�  �:  �HS� �r:  �@D� �!r:  ���� �r:  �X �  �^  ��F     j       ��^  	�  �:  �hD� |r:  �` �  �^  F�F     7      �_  	�  �:  �HS� �[:  �@D� �"[:  ��L� �[:  �X a  ��F            �G_  j E[:  �h �  f_  �F     7      ��_  	�  �:  �HS� �[:  �@D� �![:  ���� �[:  �X G  ��F            ��_  j B[:  �h 8<  �_  `�F     (       �`  	�  �:  �ha �!f:  �`b �1f:  �X }  1`  ��F     j       �M`  	�  �:  �hD� |[:  �` "�  [`  e`  �  �:   *M`  �� �`  b�F            ��`  [`  �h "  �`  �`  �  x:  &� �0  &�� �)�   &�� �65    7�`  �� �`  @�F     d       �a  �`  �h�`  �`�`  �X�`  �T 8�  0a  �F            �=a  	�  �:  �h w  \a  ��F     �      ��a  	�  �:  ��D� r:  ���  r:  ��S� r:  �X�  r:  �P�� r:  �H �  ��F            ��a  j Ir:  �h �  b  4�F     a      �fb  	�  �:  ��D� Dr:  ��0� D$r:  ���� Er:  �XL� Fr:  �PS� Zr:  �H �  ݤF            ��b  j Er:  �h �  ��F            ��b  j Br:  �h 8�  �b  ��F            ��b  	�  �:  �h �   P�G     W       �zc  P a4  T �2  H x�K  �h��  x!�2  �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�2    $!  ��G     U       �d  P a4  T �   H x�K  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �T34�f {	�     a!  \�G     �       ��d  P a4  T   H x�K  �X��  x!  �P�s x-5   �L��  x85   �HH� y5   �DZX  yX   �@��G     ?       �f {	�   �h  �!  �G     W       �Ce  P a4  T �   H x�K  �h��  x!�   �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�     �!  ��G     W       ��e  P 5  T �2  H xfP  �h��  x!�2  �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�2    "  Y�G     U       �gf  P 5  T �   H xfP  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �T34�f {	�     U"  ��G     �       �g  P 5  T   H xfP  �X��  x!  �P�s x-5   �L��  x85   �HH� y5   �DZX  yX   �@��G     ?       �f {	�   �h  �"  c�G     W       ��g  P 5  T �   H xfP  �h��  x!�   �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�     �,  �G     G       ��g  T X   F (  ݰ  3�2  �HH 3!�3  �@ �"  �G     W       �zh  P �3  T �2  H xmU  �h��  x!�2  �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�2    #  ��G     U       �i  P �3  T �   H xmU  �h��  x!�   �d�s x-5   �`��  x85   �\H� y5   �XZX  yX   �T34�f {	�     I#  �G     �       ��i  P �3  T   H xmU  �X��  x!  �P�s x-5   �L��  x85   �HH� y5   �DZX  yX   �@?�G     ?       �f {	�   �h  8m&  �i  �G            ��i  	�  �2  �h "�%  �i   j  �  �2  Gcs  �2   *�i  � #j  ��G     Y       �4j  �i  �h�i  �` 8�$  Sj  ��F            �`j  	�  �2  �h "/$  nj  �j  �  �2  Gcs  �1   *`j   � �j  �F     R       ��j  nj  �hwj  �` �#  T�G     W       �Ik  P �3  T �   H xmU  �h��  x!�   �`�s x-5   �\��  x85   �XH� y5   �TZX  yX   �P34�f {	�     `  �  
�G     J       ��k  T `  x 
Ik  �Xy 
Ik  �P/� 
`  �o 6�  ��G            ��k  T Ik  x 
*Ik  �h �  ��G     J       �l  T 5   x 
U2  �Xy 
U2  �P/� 
5   �l �,  K�G     d       ��l  F �5  H ��B  �ht �*X   �d�@ �<�  �X7* ��#  �`vsp �%�7  �P �,  ��G     �      �r  F �5  H q�B  ��t q(X   ���@ q:�  ��7* r�#  ��vsp r%�7  ����G           %m  ��  x  �X # � ?m  �u �?m  �@ <i  ��n  �� �+ ^m  um  cm  ?m  nm  )?m   �� �7 �m  �m  cm  �m  �m  
?m   9�� $H �m  �m  cm   �� i �m  �m  cm  5    !�@ �r   !H ��B  :@Y �4  n  `�G     �       �^n  jO �   jO �   	�  ,n  �X
"r  ��  ��   �T�@ r  �XH �B  �X# ;`> �! �n  ��G     �       �jO �   jO �   	�  ,n  �X��  ��   �P�@ r  �XH �B  �X#  #0� �n  �u ��n  �� <c. �np  �� �  o  o  o  �n  o  )�n   �� �: +o  Ao  o  5o  ;o  
�n   9�� ; Ro  Xo  o   �� *R io  to  o  5    !�@ �r   !H ��B  :@Y T �o  �G     �       �p  �M �   �M �   	�  �o  �X
r  ��  ��   �T�@ r  �XH �B  �X# ;`> � 4p  6�G     �       ��M �   �M �   	�  �o  �X��  ��   �P�@ r  �XH �B  �X#  #`� �p  �u ��p  �� I<? ��� �P �p  �p  �p  �p  �p  )�p   �� # �p  �p  �p  �p  �p  
�p   9�� � �p  �p  �p   �� !6 
q  q  �p  5    !�@ �r   !H ��B  :@Y �B fq  ��G     �       ��q  �M �   �M �   	�  rq  �X
r  ��  ��   �T�@ r  �XH �B  �X# ;`> �M �q  ��G     �       ��M �   �M �   	�  rq  �X��  ��   �P�@ r  �XH �B  �X#   �  �p  ;o  �m  -  ��G     �      �Dt  F �5  H '�B  ��~t ')X   ��~�@ ';�  ��~7* (�#  ��~vsp (%�7  ��~��G     0       �r  i 85   �l ��G     �      �s  s A	�1  �`ss  E5   �\p�G     J       s  i J5   �X ��G     0       =s  i L5   �T ��G     ,       as  i O5   �P �G     R       i Q5   �L  h�G     �      s V	�2  �@ss  Z5   ��]�G     V       �s  i _5   �� ��G     0       �s  i a5   �� ��G     ,       !t  i d5   �� �G     V       i f5   ��   B-  ��F           ��t  F (  ,� 's'  ��fo <�  ��H C�3  ��p �t  �`��F     �      i �   �h�F     �      c 	�  �_   �  j-  eF     *       �>u  F (  ݰ  � �1  �hfo �7�  �`H �>�3  �X �  ]u  N�F     �       ��u  	�  v9  �HR� %8�   �@ +0  �Xfra -[:  �P T  �u  F     �       ��u  	�  �:  �XD� �r:  �P�� �r:  �h =+  v  �F     L       �v  	�  �;  �h   1v  �F     �       �^v  	�  �:  �XD� �[:  �P�� �[:  �h �  }v  ʙF     D      �3w  	�  v9  ���N  45   �� 
0  �@Y  �   ���� 	�   �Xslb r:  ��N� �:  �P��F     ^       off �   �H��F     >       ݰ  �:  ��   X+  Rw  �F     O       �_w  	�  �;  �h �  ~w  r�F     X       ��w  	�  �:  �X�� pr:  �h W  �w  ��F     �       �x  	�  �:  �HD� r:  �@�� r:  �h� r:  �`&�F     I       �� r:  �X  8�  7x  x�F     I       �`x  	�  a:  �Xp ��   �Padr �	�   �h "�*  nx  �x  �  �;  0  <    7`x  �� �x  f�F     '       ��x  nx  �h "�*  �x  �x  �  �;  &G� �1   7�x  �� �x  4�F     2       �y  �x  �h�x  �` �-  G�G     d       �wy  F a4  H ��K  �ht �*X   �d�@ �<�  �X7* ��#  �`vsp �%�7  �P �-  ��G     �      ��~  F a4  H q�K  ��t q(X   ���@ q:�  ��7* r�#  ��vsp r%�7  ���G           z  ��  x  �X #p� -z  �u �-z  �@ <i  ��{  �� �2 Lz  cz  Qz  -z  \z  )-z   �� �T tz  �z  Qz  ~z  �z  
-z   9�� pK �z  �z  Qz   �� gV �z  �z  Qz  5    !�@ �r   !H ��K  :@Y i {  \�G     �       �L{  jO �   jO �   	�  {  �X

  ��  ��   �T�@ r  �XH �K  �X# ;`> / }{  ��G     �       �jO �   jO �   	�  {  �X��  ��   �P�@ r  �XH �K  �X#  #�� �{  �u ��{  �� <c. �\}  �� �W �{  |  �{  �{  |  )�{   �� �6 |  /|  �{  #|  )|  
�{   9�� ]: @|  F|  �{   �� �U W|  b|  �{  5    !�@ �r   !H ��K  :@Y 7I �|  �G     �       ��|  �M �   �M �   	�  �|  �X
  ��  ��   �T�@ r  �XH �K  �X# ;`> Q" "}  2�G     �       ��M �   �M �   	�  �|  �X��  ��   �P�@ r  �XH �K  �X#  #�� w}  �u �w}  �� I<? ��� �; �}  �}  �}  w}  �}  )w}   �� � �}  �}  �}  �}  �}  
w}   9�� � �}  �}  �}   �� �9 �}  ~  �}  5    !�@ �r   !H ��K  :@Y T T~  ��G     �       ��~  �M �   �M �   	�  `~  �X
�~  ��  ��   �T�@ r  �XH �K  �X# ;`> �/ �~  �G     �       ��M �   �M �   	�  `~  �X��  ��   �P�@ r  �XH �K  �X#   �}  )|  �z  �-  ��G     �      �,�  F a4  H '�K  ��~t ')X   ��~�@ ';�  ��~7* (�#  ��~vsp (%�7  ��~ɴG     0       �  i 85   �l ��G     �      j�  s A	�1  �`ss  E5   �\l�G     J       �  i J5   �X ��G     0       %�  i L5   �T �G     ,       I�  i O5   �P �G     R       i Q5   �L  d�G     �      s V	�2  �@ss  Z5   ��Y�G     V       ��  i _5   �� ��G     0       �  i a5   �� ߸G     ,       	�  i d5   �� �G     V       i f5   ��   '.  C�G     d       ���  F 5  H �fP  �ht �*X   �d�@ �<�  �X7* ��#  �`vsp �%�7  �P Y.  ��G     �      �%�  F 5  H qfP  ��t q(X   ���@ q:�  ��7* r�#  ��vsp r%�7  ��ݪG           :�  ��  x  �X #�� T�  �u �T�  �@ <i  �ރ  �� �- s�  ��  x�  T�  ��  )T�   �� g? ��  ��  x�  ��  ��  
T�   9�� �E   Ȃ  x�   �� �I ق  �  x�  5    !�@ �r   !H �fP  :@Y .< 5�  X�G     �       �s�  jO �   jO �   	�  A�  �X
1�  ��  ��   �T�@ r  �XH fP  �X# ;`> �L ��  ~�G     �       �jO �   jO �   	�  A�  �X��  ��   �P�@ r  �XH fP  �X#  #� ��  �u ���  �� <c. ���  �� w �  /�  �  ��  (�  )��   �� U @�  V�  �  J�  P�  
��   9�� AJ g�  m�  �   �� Z& ~�  ��  �  5    !�@ �r   !H �fP  :@Y �8 ڄ  �G     �       ��  �M �   �M �   	�  �  �X
+�  ��  ��   �T�@ r  �XH fP  �X# ;`> �2 I�  .�G     �       ��M �   �M �   	�  �  �X��  ��   �P�@ r  �XH fP  �X#  #@� ��  �u ���  �� I<? ��� �$ ��  Ѕ  ��  ��  Ʌ  )��   �� OP �  ��  ��  �  �  
��   9�� e �  �  ��   �� �R �  *�  ��  5    !�@ �r   !H �fP  :@Y �X {�  ��G     �       ���  �M �   �M �   	�  ��  �X
%�  ��  ��   �T�@ r  �XH fP  �X# ;`> � �  ިG     �       ��M �   �M �   	�  ��  �X��  ��   �P�@ r  �XH fP  �X#   �  P�  ��  �.  ��G     �      �S�  F 5  H 'fP  ��~t ')X   ��~�@ ';�  ��~7* (�#  ��~vsp (%�7  ��~ŠG     0       ч  i 85   �l ��G     �      ��  s A	�1  �`ss  E5   �\h�G     J       (�  i J5   �X ��G     0       L�  i L5   �T �G     ,       p�  i O5   �P �G     R       i Q5   �L  `�G     �      s V	�2  �@ss  Z5   ��U�G     V       �  i _5   �� ��G     0       �  i a5   �� ۤG     ,       0�  i d5   �� �G     V       i f5   ��   6)  y�   G     *       ���  T X   	�  �3  �hݰ  	X   �d �.  ?�G     d       ��  F �3  H �mU  �ht �*X   �d�@ �<�  �X7* ��#  �`vsp �%�7  �P �.  ��G     �      ���  F �3  H qmU  ��t q(X   ���@ q:�  ��7* r�#  ��vsp r%�7  ��ٖG           ��  ��  x  �X #P� ��  �u ���  �@ <i  �G�  �� �N ܊  �  �  ��  �  )��   �� �) �  �  �  �  �  
��   9�� �= +�  1�  �   �� � B�  M�  �  5    !�@ �r   !H �mU  :@Y 7! ��  T�G     �       �܋  jO �   jO �   	�  ��  �X
��  ��  ��   �T�@ r  �XH mU  �X# ;`> � �  z�G     �       �jO �   jO �   	�  ��  �X��  ��   �P�@ r  �XH mU  �X#  #�� b�  �u �b�  �� <c. ��  �� �# ��  ��  ��  b�  ��  )b�   �� �( ��  ��  ��  ��  ��  
b�   9�� W Ќ  ֌  ��   �� 
2 �  �  ��  5    !�@ �r   !H �mU  :@Y � C�  �G     �       ���  �M �   �M �   	�  O�  �X
��  ��  ��   �T�@ r  �XH mU  �X# ;`> �S ��  *�G     �       ��M �   �M �   	�  O�  �X��  ��   �P�@ r  �XH mU  �X#  #�� �  �u ��  �� I<? ��� �Y "�  9�  '�  �  2�  )�   �� f J�  `�  '�  T�  Z�  
�   9�� nQ q�  w�  '�   �� �, ��  ��  '�  5    !�@ �r   !H �mU  :@Y �0 �  ��G     �       �"�  �M �   �M �   	�  ��  �X
��  ��  ��   �T�@ r  �XH mU  �X# ;`> 6U S�  ڔG     �       ��M �   �M �   	�  ��  �X��  ��   �P�@ r  �XH mU  �X#   Z�  ��  �  !/  ��G     �      ���  F �3  H 'mU  ��~t ')X   ��~�@ ';�  ��~7* (�#  ��~vsp (%�7  ��~��G     0       :�  i 85   �l ��G     �      ��  s A	�1  �`ss  E5   �\d�G     J       ��  i J5   �X ��G     0       ��  i L5   �T ގG     ,       ِ  i O5   �P 
�G     R       i Q5   �L  \�G     �      s V	�2  �@ss  Z5   ��Q�G     V       O�  i _5   �� ��G     0       t�  i a5   �� אG     ,       ��  i d5   �� �G     V       i f5   ��   �  ۑ  d�G     ;       ��  	�  ,2  �h 6  6  �G            ��  T U2  x 
.�  �h S/  g�G     �       ���  N� iI2  �H�5 i.I2  �@ÉG     0       |�  tmp o5   �\ �G     0       tmp s5   �X  �9  ��  ��G     �      �,�  	�  B:  ��}t X   ��}�@ /�  ��}7* J�#  ��}w <�  	��J     X�G     |       p 4	[2  �X  -_   <�  1�   
 
,�  �9  `�  f�G     )       �z�  	�  B:  �hc X   �d �9  ��  4�G     1       ���  	�  B:  �hc �1  �`n )�   �X �)  ߓ  �dF     &       ���  	�  �3  �h�d 	M�1  �` �'  n/  M�F     I       �K�  T s'  F (  ݰ  3��  �HH 3!�3  �@ 2  �/  ndF     E       ���  T �1  F (  ݰ  3K�  �HH 3!�3  �@ "(  ��  ��  �  �3  &$s 	�3   *��  �z �  :dF     4       ��  ��  �h��  �`    �  �F     �      �%�  	�  v9  ��~ss  �1�   ��~$�F     �      ߕ  �N  �5   �\bkt �:  �P� L*  ��ݰ  �:  ����F     *      ��  slb 	r:  �H ƏF     �      slb 	r:  �@�� #L*  ��  ԑF     �       R� :�   ��fra ;[:  ���� =L*  ��~  9  D�  \�G     �      ���  	�  `9  ��}t X   ��}�@ /�  ��}7* J�#  ��}w <�  	��J     $�G     |       p 4	[2  �X  �8  Җ  2�G     )       ��  	�  `9  �hc X   �d �8  �   �G     1       �2�  	�  `9  �hc �1  �`n )�   �X A8  Q�  (}G     �      ���  	�  �8  ��}t X   ��}�@ /�  ��}7* J�#  ��}w <�  	��J     �G     |       p 4	[2  �X  �7  ߗ  �|G     )       ���  	�  �8  �hc X   �d 8  �  �|G     1       �?�  	�  �8  �hc �1  �`n )�   �X o7  ^�  �xG     �      �͘  	�  �7  ��}t X   ��}�@ /�  ��}7* J�#  ��}w <�  	��J     �{G     |       p 4	[2  �X  "L  �  ��  U U2  �  ,2  &�\ %U2   7͘  �A "�  �xG     N       �3�  U U2  �  �X�  �P :  R�  |xG     )       �o�  	�  ,2  �h�L =   �` "�  }�  ��  �  ,2  &ݰ  72   7o�  �5 ��  .xG     N       �Ǚ  }�  �X��  �P ,7  �  xG     )       � �  	�  �7  �hc X   �d K7  �  �wG     1       �F�  	�  �7  �hc �1  �`n )�   �X 6B  �wG            �v�  T U2  x 
*U2  �h "C  ��  ��  �  !2  0  <    *v�  Gk ��  �[F            �Ú  ��  �h ")  њ  ۚ  �  !2   *Ú  �t ��  �[F            ��  њ  �h �/  �pG     �      ��  A {9  ;= �{9  ��~s �)�1  ��~vsp �7�7  ��~8qG     �      �@ ��  ��7* �#  �`FqG     c       ��  n ��   �h 5tG     ~       Λ  w �5   �d �uG     �       �\ 	5   ��   "�9  �  #�  �  B:  &H �6  Gvsp ,�7   *�  F, F�  �pG     *       �_�  �  �h
�  �`�  �X �(  ~�  dF     ,       ���  	�  �3  �h�'  �  `)  ��  ��F     6       �՜  T s'  	�  �3  �hݰ  	s'  �P �)  ��  �cF     )       ��  T �1  	�  �3  �hݰ  	�1  �` "~(  %�  8�  �  �3  0  <    *�  _| [�  �cF            �d�  %�  �h �)  ��  �cF     )       ���  	�  �3  �` �  ��  ��F     (       �̝  	�  k9  �h�  [�   �` 9  ��F     �       �[�  �  W0�   ��tc Y�   �`e b�   �Xf c�   �Pip d�   �His e�   �@��F     :       i [�   �l  6  �F            �˞  idx H6�   ��tc J�   �hs O5   �dip P�   �Xis Q�   �Pf R�   �H �/   jG     �      ���  A �8  ;= ��8  ��~s �)�1  ��~vsp �7�7  ��~BjG     �      �@ ��  ��7* �#  �`PjG     c       o�  n ��   �h ?mG     ~       ��  w �5   �d �nG     �       �\ 	5   ��   "�8  ş  �  �  `9  &H 
5  Gvsp ,�7   *��  � 
�  �iG     *       �#�  ş  �hΟ  �`ڟ  �X �   60  	G     +       �f�  T �   a 	#�  �hb 	##�  �` 60  
cG     �      �R�  A �7  ;= ��7  ��~s �)�1  ��~vsp �7�7  ��~LcG     �      �@ ��  ��7* �#  �`ZcG     c       
�  n ��   �h IfG     ~       -�  w �5   �d �gG     �       �\ 	5   ��   "�7  `�  ��  �  �8  &H �5  Gvsp ,�7   *R�  �" ��  �bG     *       ���  `�  �hi�  �`u�  �X k�# %5   tHG     �      �k�  H V�  �$ %��  ��yV�  fmt %-�1  ��y��  %Ak�  ��y&G &	5   �l�HG     t      S 8�   �`��  B5   �\� [�   �X2�  \�   �T#�� ��  c 3X   ��~ # � â  res �$�2  �Hc �X   �G #0� �  res �$�2  ��c �X   �� #`� �  res �$�2  ��c �X   �� #�� R�  S �M   ��~c �X   ��.� �5   �� #�� ��  S 	M   ��~c 
X   ��.� 5   �� #�� �  ��  5   ���M q�  ��zS 5M   ��~.� 65   ��c 7X   ��hSG     F       c /#X   ��  �TG     @      R�  res F$�2  ��c GX   ��~S _��  ��~ H � S d[2  ��~   �   -X   ��  ��     �   ]0  \G     �      �u�  A �6  ;= ��6  ��~s �)�1  ��~vsp �7�7  ��~V\G     �      �@ ��  ��7* �#  �`d\G     c       -�  n ��   �h S_G     ~       P�  w �5   �d �`G     �       �\ 	5   ��   "7  ��  ��  �  �7  &H V4  Gvsp ,�7   *u�  �. ȥ  �[G     *       ��  ��  �h��  �`��  �X kP %5   �:G     �      ���  H e�  �$ %�  ��ye�  fmt %-�1  ��y��  %Ak�  ��y&G &	5   �l�:G     t      S 8�   �`��  B5   �\� [�   �X2�  \�   �T#P� ��  c 3X   ��~ #�� �  res �$�2  �Hc �X   �G #�� �  res �$�2  ��c �X   �� #�� :�  res �$�2  ��c �X   �� #� u�  S �M   ��~c �X   ��.� �5   �� #@� ��  S 	M   ��~c 
X   ��.� 5   �� #p� .�  ��  5   ���M q�  ��zS 5M   ��~.� 65   ��c 7X   ���EG     F       c /#X   ��  �FG     @      u�  res F$�2  ��c GX   ��~S _��  ��~ H�� S d[2  ��~   6�0  �F     +       �˨  T �   a #�  �hb ##�  �` "�  ٨  �  �  ,2  &�L *=2   7˨  [q �  vZF     V       �#�  ٨  �h�  �` 8}  B�  �[G            �O�  	�  ,2  �h "  ]�  p�  �  ,2  0  <    7O�  r ��  ZZF            ���  ]�  �h "_  ��  ��  �  ,2   7��  �d ש  6ZF     #       ��  ��  �h tC aM   �:G     2       �/�  M   �h5   �d�  �Xw ?�  	�J      -_   ?�  1�    
/�  �% ,�   H8G     ;      �R�  B� ,$�2  ��|�  ,3�   ��|.� ,@�   ��|�S ,M�  ��|�� -u3  �P�8G     �       ��  d� 4
�   �hH�� s 6�   ��}  {9G     �       i G�   �`�9G     �       d� H�   �XH � s J�   ��}      ��   6G     ;      �`�  B� ��   ��|�  �,�   ��|.� �9�   ��|�S �F�  ��|�� �u3  �P�6G     �       �  d� �
�   �hH�� s �   ��}  @7G     �       i �   �`Y7G     �       d� �   �XH�� s �   ��}    �P �5   �5G     D       ���  Jy  ��  �Xd ��  �o T�N �5   �5G            �֬  �S ��  �h T� �5   �5G            �
�  �S ��  �h l�$ ��5G            �:�  �S ��  �h � �5   05G     [       �g�  �  ��~ m�* ��4G     [       ���  �  ��~ m,X �z4G     [       ���  �  ��~  �5   �3G     �       �.�  out �.�  ��ߣ  �'�1  ����  �>k�  ��vs ��#  �@p ��5  �� M    �5   +3G     �       ���  out �.�  ��~ߣ  �&�1  ��~0��  �
�   ��~E  �5   ��~ TD �		  �2G     6       ��  + �.�  �hn �'�  �`WD �.5   �\�S �;�  �Pw (�  	��J      �   -_   (�  1�    
�  9J �		  61G     �      ���  + �.�  ��~n �&�  ��~�S �/�  ��}B� �M   �X�� �	�   �Pk �	�   �H �9 �5   �0G     �       ���  �� ��1  �X� �5   �l T>0 �5   �0G            �(�  �S ��  �h Tb? �5   �0G            �\�  �S ��  �h l� �u0G            ���  �S ��  �h ~> ~5   F0G     /       ��  Jy  ~�  �h_  ~)�  �`w ��  	ЋJ      �  -_   ��  1�    
�  L y5   0G     /       �U�  Jy  y�  �h_  y9[�  �`w ��  	ȋJ      �  FU�  3Z u�   �/G     2       �ı  B� u�2  �h�  u*�   �`.� u8�   �X�S uE�  �P �a q�   �/G     2       �(�  B� q�   �h�  q#�   �`.� q0�   �X�S q=�  �P >( oH  �/G     .       �o�  H  �l�  �`w ��  	��J      �, nH  [/G     *       ���  �2  �lw (�  	��J      $R mH  -/G     .       ���  �2  �l�  �`w �  	��J      -_   �  1�    
��  �  lH  
/G     #       �A�  w (�  	��J      {  kH  �.G     +       ���  �  �hw �  	��J      �* j5   �.G     .       �ǳ  �  �h5   �dw �  	��J      � i5   �.G     /       ��  �2  �h�  �`w �  	��J      -_   �  1�    
�  #R hH  T.G     .       �j�  �2  �l�  �`w �  	��J      '! g
��  ".G     2       ���  ��  �h5   �d�  �Xw �  	}�J      �2  F��  z  fH  �-G     +       ��  �  �hw �  	v�J      �I M5   -G     �       ���  �� M�1  ���� Nu3  �`d� P	�   �hlen Q	�   �X2 ^	�   �Pp-G     O       s S
�   �H  > I5   -G            �̵  c I5   �l Y+ F5   �,G     $       ���  c F5   �l eO B5   �,G     "       �@�  c B5   �lJy  B�  �` �9 <5   t,G     I       ���  c <5   �\Jy  < �  �Pd =X   �o neZ 85   \,G            �n;F 45   D,G            � 05   *,G            ��  Jy  0�  �h �P ,5   ,G            �6�  Jy  ,�  �h �I (5   �+G     %       �z�  �� ("2  �hJy  (;�  �` � #5   �+G     P       ���  �� #+2  �hJy  #D�  �` dO 5   y+G     "       � �  c 5   �lJy  �  �` �9 5   .+G     K       �P�  c 5   �\Jy  !�  �Pd X   �o _ �M   Y*G     �       ���  B� �S   �X]�  �-�   �PJy  �H�  �Hw �  	p�J     �*G     �       i ��   �h�*G     �       c �5   �d    �5   *G     D       �I�  Jy  ��  �Xc �X   �g� ��   �h �I �5   �)G     /       ���  �2  �hk�  �`w ��  	h�J      .! �5   �)G     /       �׹  �2  �hk�  �`w (�  	X�J      �S �5   ?)G     x       ��  �2  ��~0w �  	P�J      G0 �5   �(G     x       �Y�  �2  ��~0w ��  	H�J       �5   �(G     7       ���  ��  �h�   �`�2  �Xk�  �Pw (�  	8�J      -* �5   Y(G     7       ��  ��  �h�   �`�2  �Xk�  �Pw �  	(�J      -_   �  1�   	 
�   �5   �'G     x       �o�  ��  ��~�   ��~�2  ��~0w ��  	 �J      .* �5   i'G     x       �»  ��  ��~�   ��~�2  ��~0w (�  	�J      �S �5   6'G     3       ��  �  �h�2  �`k�  �Xw (�  	 �J      E0 �5   'G     3       �`�  �  �h�2  �`k�  �Xw �  	��J      �S �5   �&G     x       ���  �  ��~�2  ��~0w ��  	�J      F0 �5   &G     x       ���  �  ��~�2  ��~0w (�  	؊J      �H �5   �%G     3       �[�  B� �$2  �hߣ  �C2  �`��  �Zk�  �Xw ��  	ЊJ      �V �5   U%G     �       �н  B� �S   ��ߣ  �>2  ����  �Uk�  ��vs ��#  �@p �a4  �� \) �5   s$G     �       �W�  B� � S   ��~]�  �/�   ��~ߣ  �2  ��~��  �1k�  ��~vs ��#  ��p �5  �� � �5   D$G     /       ���  ߣ  �#2  �h��  �:k�  �`w �  	��J      �8 �5   $G     /       ��  ߣ  �$2  �h��  �;k�  �` � �5   �#G     `       ���  Jy  ��  �Hߣ  �=2  �@��  �Tk�  ���� �u3  �h��	��  U2G n�  �  s�  V�  5    U3G ��  ��  s�  ��  )V�   U3G ��  ��  s�  ��  ��  
V�   U3G Ϳ  ӿ  s�   o�M �X   ��  �"G     b       �%�  	�  X�  �Xc �	X   �o/ ��   �` o�9 �X   L�  Z#G     [       �|�  	�  X�  �X
s�  c �	X   �o/ ��   �` !�� �u3   !�C �5    �$ �V�  �P R �5   z"G     }       ��  Jy  ��  ��ߣ  �>2  ����  �Uk�  ��vs ��#  �@p ��3  �� �H �5   �!G     �       ���  B� �#2  ��}ߣ  �B2  ��}0��t�  V2G ~�  ��  ��  e�  5    V3G ��  ��  ��  ��  )e�   V3G ��  ��  ��  ��  ��  
e�   V3G ��  ��  ��   p�M �X   �  ^!G            ��  	�  O�  �h p�9 �X   C�  r!G     0       �U�  	�  O�  �h
��   AB� ��1   A�C �5    �$ �e�  ��~��  ��   ��~E  �	5   ��~  z5   � G     �       ��  B� zS   ��~ߣ  z=2  ��~0��  {
�   ��~E  }5   ��~ ]) s5   �G     �       ���  B� sS   ��~]�  s.�   ��~ߣ  sO2  ��~0��  t
�   ��~E  v5   ��~ � o5   zG     x       ���  ߣ  o"2  ��~0w �  	��J      �"S �G     �       �#�  S �   �h�  0�   �di I�2  �X >T �5   G     �       �w�  ߣ  �#2  ��~0��  �
�   ��~E  �5   ��~ >� �5   eG     �       ���  Jy  ��  ��~ߣ  �<2  ��~0��  �
�   ��~E  �5   ��~ >S �5   �G     �       �?�  Jy  ��  ��~ߣ  �=2  ��~0��  �
�   ��~E  �5   ��~ �[? �G     2       ���  Jy  ��  �hB� �7S   �`w �  	��J      >jL ��  LG     3       ���  `  �&2  �h�� �G2  �`Jy  �^�  �Xw ��  	��J      >XM �M   !G     +       �8�  B� �M   �hw �  	x�J      >�M ��  �G     #       �n�  w ��  	p�J      >� �5   �G     5       ���  6A �5   �ltF �(�1  �`�M �65   �h�) �L�1  �Xw (�  	`�J      >�- �5   /G     �       �S�  xF ��1  �X�) �*�1  �Pw �  	V�J     �G     ;       e �	5   �l  >�� �5   G     +       ���  `  ��1  �hw �  	O�J      Z6  ��  �[G     O       ���  	�  �6  �Xstr ��1  �Pn �&�   �H�[G     8       i ��   �h  ;6  �  4[G     S       �Y�  	�  �6  �Xstr ��1  �PD[G     @       i ��   �h  6  x�  �ZG     L       ���  	�  �6  �hc �X   �d 6  ��  �YG     	      ��  	�  �6  �Hw �  	��J     ZG     �       P( �	�   �h"* �	M   �P  "�5  �  �  �  �6   *�  mZ <�  �YG     .       �E�  �  �h �5  d�  `YG     O       ���  	�  �5  �Xstr ��1  �Pn �&�   �HtYG     8       i ��   �h  e5  ��  YG     S       ��  	�  �5  �Xstr ��1  �PYG     @       i ��   �h  8F5  %�  �XG     Q       �?�  	�  �5  �hc |X   �d ""5  M�  o�  �  �5  &B� yM   &�� y&�    *?�  �D ��  �XG     6       ���  M�  �hV�  �`b�  �X 8�4  ��   XG     c       ��  	�  5  �Xstr l�1  �Pn l&�   �H0XG     P       i n�   �h  8�4  1�  �WG     g       �l�  	�  5  �Xstr d�1  �P�WG     X       i f�   �h  8�4  ��  |WG     <       ���  	�  5  �hc _X   �d "n4  ��  ��  �  5  &B� \M    *��  q' ��  VWG     &       ���  ��  �h��  �` 4  �  WG     M       �E�  	�  \4  �hstr R�1  �`n R&�   �X �3  d�  �VG     e       ���  	�  \4  �Xstr M�1  �P �3  ��  ZVG     H       ���  	�  \4  �hc HX   �d "�3  ��  ��  �  \4  &Jy  E�   *��  cS  �  4VG     &       ��  ��  �h��  �` "�'  �  C�  �  �2  qB� "�2  q�  "(�    *�  � f�  (�F     *       ��  �  �h(�  �`5�  �X �  ��  <�F     6       ���  	�  g2  �`c 63�  �\�  7�  �h r2  2��  ��  �  g2  0  <    7��  �o �  ZF            ��  ��  �h h  rN  2/�  >�  �  g2  �   7�  �e a�  �YF     �       �r�  /�  �h8�  �` "�  ��  ��  �  g2   7r�  w ��  &YF     \       ���  ��  �h �6r kv �   YF            ���  �  #�   �hp /�   �` 8P1  �  �F            �&�  	�  �1  �h 61  E�  րF     B       �e�  	�  �1  �hw u�  	؋J      -_   u�  1�    
e�  6�  ÀF            ���  x )�   �h "  ��  ��  �  �0   *��  �� ��  r�F     Q       ���  ��  �h +&E +�
  s&  %*  "s�  %*  " ~   �  �n [ ~c ��G     �      �� ^� �9   �i �� 	L   int �� _   j   _   �  j   ! _   �i 	-  
�Z 4_   6H     H       ��   S 4e   �Xsrc 4<�   �Pn 59   �h q   �   
i[ 0�   �H     7       �C  S 0�   �hsrc 0'C  �`len 03-   �X I  
�[ 'L   �H     ]       ��  e 'L   �\B� '_   �P�Z ',-   �Hs (_   �h [ 
_   b
H     @      ��  e 
L   �\s �   �h 
�Z 
9  0
H     2       �9  9  �hD  �d-   �Xw `  	��J      D  9  Jf D  q   `  9    P  
�[ -   
H     +       ��  �  �hw �  	ՕJ      K  �  q   �  9    �  �[ �
9  �	H     f       �@  s �!�  �Xc �,D  �T�  �6-   �H�[  �  �`�	H     H       i -   �h  �Z �
9  l	H     3       ��  ?  �h�  �`�  �Xw �  	ΕJ      9  �  y[ �
9  =	H     /       ��  �  �h�  �`w �  	ǕJ      \ �-   	H     /       �%  �  �h�  �`w �  	��J      �Z �
9  �H     .       �k  �  �hD  �dw `  	��J      Z[ �
9  �H     /       ��  �  �h�  �`w `  	��J      �[ �-   �H     /       ��  �  �h�  �`w `  	��J      b[ �
9  TH     .       �=  �  �hD  �dw �  	��J      �Z �L   !H     3       ��  �  �h�  �`-   �Xw `  	��J      \ �L   �H     3       ��  ?  �h�  �`-   �Xw `  	��J      q[ �L   �H     3       �'  �  �h�  �`-   �Xw `  	��J      \ �L   �H     /       �m  �  �h�  �`w `  	��J      �[ �L   ]H     /       ��  �  �h�  �`w �  	x�J      �Z �
9  *H     3       �  ?  �h�  �`-   �Xw `  	p�J      �[ �
9  �H     /       �G  ?  �h�  �`w �  	i�J      �Z �
9  �H     3       ��  9  �h�  �`-   �Xw �  	`�J      q   �  9    �   \ �
9  �H     3       ��  ?  �h�  �`-   �Xw `  	X�J      �Z �
9  bH     3       �F  ?  �h�  �`-   �Xw `  	P�J      �Z �
9  3H     /       ��  ?  �h�  �`w �  	I�J      �Z ��  H     2       ��  �  �h�  �`L   �\w �  	@�J      �i �[ �9   �H     2       �/	  �  �h�  �`L   �\w `  	8�J      [ �}	  �H     2       �}	  �  �h�  �`L   �\w `  	0�J      S  [ ��	  kH     2       ��	  �  �h�  �`L   �\w �  	(�J      X  �Z �
  <H     /       �
  �  �h�  �`w `  	 �J      �
  �Z �l
  H     /       �l
  �  �h�  �`w �  	�J      &E �Z ��
  �H     /       ��
  �  �h�  �`w �  	�J      �
  �Z �_   �H     \       �
  s ��   �Xc �$L   �Ti �	-   �h �[ �_   VH     ,       �_  s �e   �hG[ �9�   �`\ �_   	@�K      Q[ �_   ,H     *      ��  s �!e   �Xdel �;�   �Pm �R�  �Hw �  	�J     tok �_   �hp �_   �` _   �  �+  �_   yH     �       ��  s ��   �H�Z �)�   �@�H     �       i �-   �h�H     x       ;�  ��  �g�H     a       j �-   �X    t �[ �-   H     m       ��  s ��   �X[ �*�   �Pn �	-   �h �\  �_   �H     p       �A  s ��   �Xc �"L   �Tss  �	-   �`�H     J       i �-   �h  (\ �_   .H     n       ��  s ��   �X[ �*�   �Pn �	-   �h �[ }-   � H     m       ��  s }�   �X[ }+�   �Pn ~	-   �h �[ r_   X H     i       �#  s r�   �Xc r!L   �Ti s	-   �h �[ k�   ��G     Y       ��  s kC  �Xc k!L   �T�  k+-   �H�[ l�  �` H     ;       i m-   �h  �  �  �  �[ f-   ��G     3       �  S f!e   �hsrc f>�   �`]�  fJ-   �Xw `  	 �J      ��  UL   E�G     �       ��  a U�   �Xb U(�   �P]�  U2-   �Hi V	-   �h]�G     k       �[ Z�  �g�[ [�  �f  �[ PL    �G     %       ��  a P�   �hb P(�   �` Bi  @L   ��G     r       �R  a @�   �Xb @'�   �Pi A	-   �h��G     Z       �[ C�  �g�[ D�  �f  �  5L   <�G     r       ��  a 5C  �Xb 5'C  �P�  51-   �HL�G     [       i 6-   �h^�G     B       �[ 7�  �g�[ 8�  �f   �[ (_   ��G     �       �i  S ( e   �Hsrc (=�   �@]�  (I-   ��� )_   �hπ *�   �`i ,	-   �X �S  $_   �G     ;       ��  S $e   �hsrc $<�   �` �9  _   ��G     �       �&  S  e   �Hsrc 2�   �@]�  >-   ��� _   �hπ �   �`i 	-   �X ;�  _   ��G     S       �S e   �Xsrc 1�   �P� _   �hπ _   �`  �   ��  �n �\ ~c ~H           �� �  �  �i -  N   �i �  -  int X  �  �N   7  B   �  4q   ^� �N   ]� j   d j   �n �  0\ @p\ c   �   �  c    ;\ ;] c   �   c    �\ 0V\ c   "  �  c      ] �\ c   K  c   �   c   |   M\ $] c   t  c     �      �\ �\ c   c   }  �       	�  �  
�  �   =H     C       ��  `  @�  �X�� @+c   �Tret Ac   �l �   H     :       �  fd ;c   �l 	c   �   �H     W       �|  `  0�  �X?1  0)c   �Tfd 05  �H_fd 1c   �l 	�   "  EH     g       �  fd c   �\x  �   �P�� )c   �X2� 8|  �Hoff  	�   �h�\ !c   ret #}   �` 	�   K  �H     a       �}  fd c   �\buf   �P.� )�   �H� 9  �@ret c   �l�\ c    	�  t  ~H     f       �fd c   �\B� $}  �P.� 3�   �HE\ C  �@ret c   �l  �   ��  �n �h ~c `�         �� ^� �:   )   �i X  S  �
  �  std  ?  9t 	�   �\ 	F  �l 	?  	�l 	=g �   �   �   
T   	�g 	t �   �   �   
T   T ?  v ?    f   �v 	O  �\ 	F  �l 	?  	�g 	�o �     !  
c   	�g 	Vl �   9  ?  
c   T ?  v ?   �   �h 	`u  � 	a   T �   �` 	[�  � 	\Y  T Y   �] 	`�  � 	av  T    �� 	j>�  G` !b �  �  T      �c �` �    T Y      �� 	j>�  c �e �  2  T �     �� 	j>a   t ?  �d s   �   6h �   O  �  �  �i w  �  -  int �  �  
�:   �  4�  �  frg 	5  �� 	�  W� �   `� 	�    � F    �  >� �  .  �r  red d�  l� 0�  l� � O  U  
?   l� � i  t  
?  E   Gp ;� K  �  �  
?  E   S� Q   �  Q  �� Q  )�  Q  �� !Q   � "	  ( .  �� %f� 5�   h 8`� ?    �   O� =t� �  4  �   �� BͰ �  N  �   n� E� �  h  �   )� I�� �  �  �   �� L7� �  �  �   	�� PE� �  �  �  
�   !#� U�� ?  �  �   !�� Z؟ ?  �  �   � d�   
  
�   � g�   )  
�  �   Gp i;�   A  L  
�  �   	N� o�� �  d  j  
�   "� |\�   �  
�  �   "c� ��� �  �  
�  �  �   "�� ��� �  �  
�  �  �   "
� �6� �  �  
�  �   #�� #� 	    
�  �   $<� � *  :  
�  �  �   $�� D� P  `  
�  �  �   $�� x)� v  �  
�  �   $�� �$� �  �  
�  �   $/� �� �  �  
�  �   #� u� �  �  
�  �   #,� #E� �    
�  �   %0� 0�� ?    #  
�   %0� 94� ?  =  W  
�  �  	       &�� �Q   D �  T �  '� �  A �   �  (� �D  )�j  )��  )��  )�4  )�N  )��  *�   #�� �\� �  �  
  v   #\+  ��� 
    
  �   &�� �v  T �  '� �  L v  A �   _� 5�   h 8� ?  j  �   O� =� �  �  �   �� B� �  �  �   n� E2� �  �  �   )� I�� �  �  �   �� L� �  �  �   	�� PK� �  	  
	  
&   !#� U� ?  %	  �   !�� Zk� ?  @	  �   � dg� T	  Z	  
&   � g4� n	  y	  
&  1   Gp iI� 7  �	  �	  
&  1   	N� o�� �  �	  �	  
&   "� |c� �	  �	  
&  �   "c� �)� �	  �	  
&  �  �   "�� ��� 
  $
  
&  �  �   "
� �� 9
  D
  
&  �   #�� U� Y
  d
  
&  �   $<� �� z
  �
  
&  �  �   $�� Dz� �
  �
  
&  �  �   $�� x�� �
  �
  
&  �   $�� �Z� �
  �
  
&  �   $/� ��     
&  �   #� ;� (  3  
&  �   #,� #�� H  S  
&  �   %0� 0�� ?  m  s  
&   %0� 9�� ?  �  �  
&  �  	  =  =   &�� �Q   D �  T �  '� �  XA �   D  +W� �)��	  )��	  )��	  )��  )��  )��  *D   #�� �F� 6  A  
C  v   #\+  �Q� V  a  
C  �   &�� �v  T �  '� �  XL v  A �    �  � F    �  ,"� �$�  "� �  ��  �r  l� [�  �  � H�	�  � ���     
�  �  �  )    � �5� .  9  
�  �   Gp �
�� �  Q  \  
�  �   	Z� �δ ?  t    
�  Q   � ��    ��  ss  �5   "� ��   �  � ��	l  *�   � �E� �  �  
�  �  )   �   � ��� 	    
�  �   Gp �r� �  ,  7  
�  �   �N  ��  Hٖ �w  LU� ��  P.� ��  X �  -'� � �	�  .�g �a� ?  �  
  �  �    �0   �	�  �0  ��� �  �  
N   � �	X   x� ��  � ��   �� ��  "�� �-�   #  
Y  �   /�� (z� 8  C  
Y  d   0Gp *� j  \  g  
Y  d   1Wd ��� Q  �  �  
Y  )    %�6  L�� Q  �  �  
Y  Q  )    $�N ~�� �  �  
Y  Q   $� �w� �  �  
Y  Q  )    1Y� 1	�� )       
Y   2J� >�                         @       3�� @ ~  3�� A ~   H� H�� )     w   r� W�� )   �  )    3�� j�  � l5   �� o�� ?  �  w   o� |5   �� 5   4� �5    5<� �7� �      
Y  �   5a� �� �  4  ?  
Y  �   5P� %j� �  X  c  
Y  )    #`� 7� x  ~  
Y   #� >� �  �  
Y  �   Э �
�   A� �X  ۧ ��  @� ��  �� �	)    � ��  (6�    6v� X   �  70� V�  $;� X� '  2  
  Y   %Wd [!� Q  L  W  
  )    $� _ʅ m  }  
  Q  )    $�N c�� �  �  
  Q   %� gε Q  �  �  
  Q  )    8�� lY   6�    6v� X   9f 3  �^ <g     
�   B� �   '�V  :   '�^ :    :�c �  ;get  �^ �  Z  `  
�   <�^ %)�   "�^ Hc �  �  =�O  
�   T     >G� �+.  >� �7�  >� �7�  ?0c �	  �^ (f �  �  
�   B� �   @�V  :   �'�^ :    A�d �|  ;get  �_ j  1  7  
�   <�^ %)�   "=_ �^ i  t  B�O  i  C�   
�  �   T �   9�^ �  �^ �b �  �  
   B�    '�V  :   '�^ :    D#b ;get  ld *  �  �  
0   <�^ %)|   "xc �] !  ,  B�O  !  CY   
0  �   T     E�  E�  .  F�  F.  GE�  -�   -� �� y    
	   -� � �  �  
	     Gp ��   �  �  
	     7� �� �  �  
	   �� �� �  �  
	   Hn� �    X  X  	  F  FX  >� q  Imap x� �  E  P  
q  )    Jɒ   �� `  
q  �  )        q  bb %>  �  �  K�n -�  �  L�  �  M:     F   3  �  �  F�  F�  �  Fl  F�  q  �  �  F�  F�  F�  F�  v  �    D  &  F�  FD  F�  �  C  �  N  �  Y  F�  F�  L5   �  M:    p  g�   !� I  �� W  K� �  ?� �  �� �  5� �  ݉ �  L�  �  M:    �  �  L�  �  N:   � 	  �      |    L�  *  M:    F  �  0  O@	  I  S  P�  ,   Q;  cg v  �H            �  RI  �h O!  �  �  P�  I  S�� �v   T  X_ �  �H     $       ��  R�  �hR�  �  O�  �  �  P�  �   Q�  Qf   �H            �  R�  �h Fv  U�  H     
       �R  T   Vx *  �h O�  `  j  P�  T   TR  Ah �  HH     7       ��  R`  �h O�  �  �  P�  !  S�� �v   T�  .e �  $H     $       ��  R�  �hR�  �  O  �    P�  
  S�� X+Y   Q�  d 7  
H            �H  R�  �hR  �` O�  V  `  P�     QH  e �  �H            ��  RV  �h O  �   �  P�  _  Wѭ �-�   T�  g] �  xH     {       ��  R�  �XR�  �P O�  �  �  P�  �   Q�  >]   RH     %       �(  R�  �h O�  6  @  P�  �   Q(  ^^ c  @H            �l  R6  �h X�  �  2H            ��  Y�  6  �h ZY  O�  �  �  B�O  �  CY   P�  6  [�    T�  �a   �H     P       �   B�O    CY   R�  �X\  ]�   R�  �P F  U�  �H            �V  T Y  Vx .   �h X  u  �H            ��  Y�  �  �h OE  �  �  B�O  �  C�   P�  �  [�    T�  4a �  vH     P       �  B�O  �  C�   R�  �X\�  ]�   R�  �P F2  U  hH            �:  T �  Vx .  �h XA  Y  ZH            �f  Y�  �  �h On  y  �  =�O  P�  �  ^ Tf  �a �  .H     ,       ��  =�O  Ry  �h^ _P  �  �H     R       �  Y�  w  �h`  (�  �``ss   8)   �Xaw +  	{�J      L�  +  M:      b-  R  tH     Q       ��  Y�  w  �X`ss  ()   �Pcptr Q  �haw �  	w�J      L�  �  M:    �  drb �d   �H     �       �  e�c (3  	`�K     e�^ "	  	��K     e�h '�  	P�K      F|  Oe  "  ,  P�     Q  %g O  H            �X  R"  �h f6r kv Q  YF            ��  `�  #)   �hVp /Q  �` �i &E �
  g�  �  "g�  �  " �   t�  �n �n ~c  �         t� ^� �5   �i �  �  t  V   �i V   �  -  int p   X  g  J   frg S  /g �   [r  �   	�t  �   
�q 7Y   Mq !  �h {,  ݰ  |p   �h ~�q 
    t   �h h    t  p     �s  u A  G  z   �s p \  g  z  �    �s �v |  �  z  �   �s *o �  �  z  �   �s *gs �  �  z  �   �s 0dr �  �  z  �   �s 8�m �    z  p    Gp =�w �     +  z  �    �s Qr �  D  J  �   �s T�i �  c  i  z   ]h X%d �  �  �  �   p \Xw �  �  �  �   p `�k �  �  �  z   �o d�g �  �  �  z   �� ��s �  �  z   wq ��    �r ��  T p    �   /f JDq 
.  �g 7  `d Xt  e  S  �  ^  S  �
  �  std  �  9t 	�  �\ 	�  �l 	�  �l 	=g �  �  �  
   �g 	t �  �  �  
   T �  v �    �  �v 	q  �\ 	�  �l 	�  �g 	�o   =  C     �g 	Vl   [  a     T �  v �   �  �s 	��  �\ 	��  T p   �O   �    ;s 	��  �\ 	��  T p   �O   �    !v 	��q �  !v 	��e �   t �  "�d �  �  "6h   q  #�   	��J     #�   	x�K     l 
r  b� 
i    �� 
i   3� 
V    $�   �   %w   &p   %!  &�   %�   !  %p   p   'Ln �  'uh �  �i �  Jf �  #<  	��J     (�n �  )�w +�v H  )�r ,�p M  *� p   I  +�r  +q� +� +�� +o�  � �  ,it S   ,end S  -�s �� �  �  �  �   C e   �� �  ,it �   ,end �  -�s x� �  �  �  �   C V    h� -  ,it �   ,end �  -�s 2� �    %  �   C �   �h q_  .� r^�   N  �  �  �    � #�   �j 	j  ]s 	  ]s �m �  �  �   d� �q �  �  �  �   5� 7q �  �  �  �   �g �n   �  �  �  �   /c� 5p    /4� 6_   s 9	M  .�g <�l   <  �    	    0}j 
�  0ol �    �j �  ,it '   ,end S  -�s �m �  �  �  -   C ^   �h 	  ,it �   ,end �  -�s 
r �  �  �  !   C ]    �m N	  ,it �   ,end �  -�s )i �  @	  F	  8   C �   1Om Q�
  �
  2�
   3�q or v	  �	  L  W   3�q %l �	  �	  L  ]   �q Rk �	  �	  L   48� UEi   N	  �	  �	  L  �  c  i   4�j q�l   N	  
  !
  L  �  o  i   4Vk ��p   N	  A
  V
  L  �  u  i   4gq ��n   N	  v
  �
  L    {  i   5�q <j N	  �
  �
  L  p    G k   N	  1zo ,�
  x  3zo �j �
  �
  �  �   6to �   7�p ,j �
  
    �  p    � 0��   -  =  �  ^  �   �i D%s   U  e  �  ^  �   zo WJr y  �  �  �  �   48� Z�k   �
  �  �  �  �  c  i   4�j ]ok   �
  �  �  �  �  o  i   4Vk `�o   �
    (  �  �  u  i   4gq cBp   �
  H  ]  �    {  i   }j g�  ol j�  	 �
  8j �&r �  8�o �i �   I  �  V   ]   �  �  �  �  �  -  �  %_  x  �  jl %I    �  %j  %�  "�m M  "�j [  �  ^  j  -  	  8  9Z  r  N	  L  &N	  %�
  %�  %=  %�  )   %	  �
  �  %x  :p   �  ; �  <�� �  %�  =�  =�  >(	  �  NH            ��  ?�  >  �h >�    .H            �  ?�  3  �h >  4  H            �A  ?�  �  �h >�  `  �H            �m  ?�  �  �h >o  �  �H            ��  ?�  �  �h @V
  �  vH     X      �h  ?�  R  ��A�n �3  ��A-� �R{  ��Bst �i  ��Cw x  	��J     D�l �j  �PEes �  �OF H     �       Ecp �_  �HEcps ��  ��G�� Ee �  �l   He  x  I5    h  @!
  �  bH           �&  ?�  R  ��A�n �@�  ��Bn �Nu  ��Bst �i  ��Cw 6  	��J     D�n �I  �PEds �x  �HF�H     !       Ee �  �l  He  6  I5    &  @�	  Z  H     G      ��  ?�  R  ��A�n q9�  ��A-� qRo  ��Bst ri  ��Cw x  	�J     D�n uI  �PEds vx  �HF�H     $       Ee z  �l  @�	    �H     K      ��  ?�  R  ��A�n U.�  ��A-� UIc  ��Bst Vi  ��Cw �  	"�J     D�n YI  �@Eds Zx  ��FeH     $       Ee ^  �\  He  �  I5    �  J�
  Q�  �  K�  R  K0  w    L�  �r �  �H     +       ��  M�  �h L�  Dn   tH     -       �#  M�  �h N�	  1  ;  K�  R   L#  �o ^  <H     7       �g  M1  �h O}  �H            ��  D�h �-  	x�K      P:  ��  �H            ��  ?�  �  �hBnc �/�  �dBwc �>�  �X Q�  #H     g       �  Dn �5N	  	`�K      N�
  $   7  K�  �  K0  w    L  �r Z  �H     +       �c  M$  �h R   n �  �H            ��  M$  �h @(  �  �H     |       ��  ?�  �  �XA�n <.  �PA-� <O	  �HEwc =	V   �lCw 
  	ȗJ      He  
  I5   
 �  @�  .  6H     �      �k  ?�  �  �XBseq 4�  �PEuc 	<   �oCw 
  	 �J      S�  V   �  $H            ��  ?�  �  �h S�  p   �  H            ��  ?�  �  �h N�  �  �  K�  �   R�  yq   �H             �  M�  �h Ne    ?  K�  �  T�q W�  T�i W8�   R  �i b  �H     =       �{  M  �hM&  �dM2  �` &E �
   (   ��  �n �t ~c @�         	� X  ^� �<   �i S  �
  �  �  �  t  p   �i p   �  -  int �   g  	d   std    9t 
  	�\ 
!  �l 
  
�l 
=g �   �   �   /   
�g 
t �   	    /   T   v     �   �v 
�  	�\ 
!  �l 
  
�g 
�o >  b  h  >   
�g 
Vl >  �  �  >   T   v    $  �s 
��  	�\ 
�!  T �   �O  �	    ;s 
��  	�\ 
�!  T �   �O  �	    v 
��q !  v 
��e !   t   �d �     6h 1  �  frg 	�	  /g R  [r  [  �t  �  �q 7�	   mi �   ,�  �r  �( hex  Mq �  �h {  ݰ  |�   �h ~�q �  �  �	    �h h �  �	  �     !�s  u   #  �	   !�s p 8  C  �	  "R   !�s �v X  c  �	  "�	   !�s *o x  �  �	  "�	   !�s *gs �  �  �	  "�	   !�s 0dr �  �  �	  "�	   !�s 8�m �  �  �	  �    #Gp =�w �	  �    �	  "�   #�s Qr      &  �	   #�s T�i   ?  E  �	   #]h X%d   ^  d  �	   #p \Xw �	  }  �  �	   #p `�k �	  �  �  �	   #�o d�g 
  �  �  �	   �� ��s �  �  �	   $wq ��   $�r �  T �    �  ,s 2�  ,s 3�s #  )  
   
#m 6Rf   A  L  
  "�   $(m <�   $�m =�   $H� >�  $�t ?  $v @  $�r A  $;f B  $�u C  %+s �n �  �  
  �    &,s  i �  
  "<      '/f J�  (�� Nm{ <  P �  T p   "�  "p   "  "�   "�   "�   "�	   (B~ xR y  P �  T p   "�  "p   "�   "�   "�   "�	   )*y �� T p   F �  "p   "  "�    Dq 
�  �g �  `d �  s E�x �  �  �  "S
   j �	a  j |     �  "�   *j *{ *  5  �  "�   +Gp 	@� �  M  X  �  "�   j  l  w  �  �    
Cr "	�z �  �  �  �  "�    i '�} �  �  �  "�	    i 1Wz �  �  �  "�	   ,#s >�   ,A� ?�  ,�� @
0   �,m A  �
*q 	z �  /  :  T p   �  "p    -�m 	�~ �  U  T �	  �  "�	    �  
�g Hx �  ~  �  �   !�l Mox �  �  �  "�	   ,cg QS
   .�n S
  /�! <   � 0Xt 1t 
*w �	  �  T �   "�	  "�	   (�~ ��| 	  F �  "p   "  "�   (�~ ��} ?	  F �  "�	  "  "�   2�{ 3�y i	  T p   F �  "�  "�   3xy 3} T �	  F �  "  "�    4`  	0�J     �	  �	  �  �	  4y  	��K     �  �	  �  �	  5�   6�   5�  6�  5�  �  5�   �     
  7Ln �  7uh �  �i Jf 4�  	B�J     '�n �  x �
  8x 
Xx u
  {
  �    �g y �
  �  "�	    9�w +�v �  9�r ,�p �  � #�   ��  �  
�u .u   �
  �
  �   
�s �s       �  "�
   
�o Uu   )  4  �  "�
   
�u t   L  W  �  "�
   
�s �t   o  z  �  "�
   
�u �u   �  �  �  "�
   
�s bt   �  �  �  "�
   
�s js   �  �  �  "�
   
3 �s   �    �  "�
   
�u �s     )  �  "�
   
�t t   A  L  �  "�
   
t (t   d  o  �  "�
   
u �t �
  �  �  �  "�
   -�u u �
  �  �  "�
    :�u �
Et �   S
  �
  �  �  �  �  �  5a  5�  ;�	    <<    =�  =  >�  /  �hF     �       �I  ?�  �  �h@s '�	  �d A�  O`F     (       ��  T �   @a �	  �h@b #�	  �` B�  RgF     �      ��  P �  T p   CH N�  ��C��  N$p   ��Cs N1  ��C�s N?�   ��C��  O�   ��CH� O�   ��CZX  O#�	  ��D]� P�	  �XDB� S�  ��Ek T�   ��FBhF     E       o  Ei a�   �l F�hF     -       �  Ei d�   �h G�hF     0       Ei f�   �d  ;�	  �  <<    B<  �fF     U       �T  P �  T p   CH x�  �hC��  x!p   �dC�s x-�   �`C��  x8�   �\CH� y�   �XCZX  y�	  �THI�f {	p     By  afF     �       ��  T p   F �  Cݰ  �p   �l@fo �/  �`CH �6�  �X >�  �  �eF     �       ��  ?�  �  �h@str 1�	  �` B�  FeF     J       �7  F �  Cݰ  �!p   �L@fo �8  �@CH �?�  �� B	  eF     *       ��  F �  Cݰ  � �	  �h@fo �7  �`CH �>�  �X 5w   B?	  �dF     C       ��  T p   F �  Jݰ  3�  �HJH 3!�  �@ >�  �  �dF     &       �  ?�  �  �hC�d M�	  �` 5�	  Bi	  ndF     E       �b  T �	  F �  Jݰ  3  �HJH 3!�  �@ K�  p  �  L�  �  M$s �   Nb  �z �  :dF     4       ��  Op  �hOy  �` K�  �  �  L�  �	  L0  �    N�  Gk �  �[F            �  O�  �h K�      L�  �	   N  �t B  �[F            �K  O  �h >  q  �cF     (       ��  T p   ?�  �  �hCݰ  p   �d >w  �  dF     ,       ��  ?�  �  �hP�  �  >:  �  �cF     )       �  T �	  ?�  �  �hCݰ  �	  �` KX    $  L�  �  L0  �    N  _| G  �cF            �P  O  �h >f  o  �cF     )       �|  ?�  �  �` K�  �  �  L�  �	  M�L *�	   Q|  [q �  vZF     V       ��  O�  �hO�  �` K�  �  �  L�  �	  L0  �    Q�  r   ZZF            �!  O�  �h K  /  9  L�  �	   Q!  �d \  6ZF     #       �e  O/  �h A�  �'H            ��  Dru ��
  	y�K      R�  ��  'H     �       ��  ?�  �  ��~@c �'�
  ��~ Ro  v�  d&H     �       �  ?�  �  ��~@c v'�
  ��~ RL  m5  �%H     �       �Q  ?�  �  ��~@c m"�
  ��~ R)  ds  �$H     �       ��  ?�  �  ��~@c d"�
  ��~ R  [�  6$H     �       ��  ?�  �  ��~@c ["�
  ��~ R�  R�  X#H     �       �  ?�  �  ��~@c R"�
  ��~ R�  I-  �"H     �       �I  ?�  �  ��~@c I"�
  ��~ R�  @k  �!H     �       ��  ?�  �  ��~@c @"�
  ��~ Rz  1�  �H           ��  ?�  �  ��~@c 1"�
  ��~ RW  (�  �H     �       �  ?�  �  ��~@c ("�
  ��~ R4  %  H     �       �A  ?�  �  ��~@c #�
  ��~ R  c  JH     �       �  ?�  �  ��~@c "�
  ��~ R�
  �  ~H     �       ��  ?�  �  ��~@c "�
  ��~ S�
  �  nH            ��  ?�  �  �h T�  2�    L�  
  L0  �    Q�  �o 3  ZF            �<  O�  �h 5�  T�  2S  b  L�  
  "<   QB  �e �  �YF     �       ��  OS  �hO\  �` K  �  �  L�  
   Q�  w �  &YF     \       ��  O�  �h U6r kv D  YF            �  C�  #0   �h@p /D  �` &E �
   �   ��  �n _v ~c  �         �� X  ^� �<   �i S  �
  �  a  b   �  �  t  |   �i �  -  x  �   int �   Qv )   �  �<   h  	�   �   8  	�     	V   g  	p   �  	4�   std  z  9t 
  	�\ 
�  �l 
z  
�l 
=g '  K  Q  �   
�g 
t '  i  o  �   T z  v z      �v 
�  	�\ 
�  �l 
z  
�g 
�o �  �  �  �   
�g 
Vl �  �  �  �   T z  v z   �  �s 
�(  	�\ 
��  T �   �O  L
    ;s 
�U  	�\ 
��  T �   �O  R
    v 
��q �  v 
��e �   t z  �d     6h �  �  �  frg 	�	  /g �  [r  �  �t  �  �q 7

   mi �   ,  �r  �( hex  Mq b  �h {m  ݰ  |�   �h ~�q K  Q  *
    �h h a  *
  �     !�s  u �  �  5
   !�s p �  �  5
  "�   !�s �v �  �  5
  "@
   !�s *o �  �  5
  "F
   !�s *gs �    5
  "L
   !�s 0dr   (  5
  "R
   !�s 8�m =  H  5
  �    #Gp =�w X
  a  l  5
  "   #�s Qr z  �  �  ^
   #�s T�i z  �  �  5
   #]h X%d z  �  �  ^
   #p \Xw @
  �  �  ^
   #p `�k d
      5
   #�o d�g j
     &  5
   �� ��s :  @  5
   $wq �   $�r �z  T �      ,s 2N  ,s 3�s �  �  p
   
#m 6Rf g  �  �  p
  "�   $(m <�   $�m =�   $H� >  $�t ?z  $v @z  $�r Az  $;f Bz  $�u Cz  %+s �n *  5  p
  �    &,s  i B  p
  "�    g  '/f J	  (�w N0y �  P T  T <   "�  "<   "z  "�   "�   "�   "
   (ww x�u �  P T  T <   "�  "<   "�   "�   "�   "
   )�x ��v T <   F T  "<   "g  "�    Dq 
	  �g   *`d Xt 0	  s ECo I  T  �  "�
   j �	�  j �e u  �  �  "�   +j ig �  �  �  "�   ,Gp 	�j �  �  �  �  "�   j �f �  �  �  �    
Cr "	�r �  �    �  "	    i '�h   #  �  "
    i 1~j 7  B  �  "
   -#s >�   -A� ?*  -�� @
0   �-m Az  �
M� 	x �  �  �  T �  �  "�   .�m 	3m �  �  T 
  �  "
    T  
�g H�o T  �  �  �   !�l Mj 	  	  �  "
   -cg Q�
   /�n �
  0�! <   � 1t 
*w @
  V	  T �   "@
  "@
   (nk �
w }	  F T  "�
  "g  "�   (nk �Au �	  F T  "
  "g  "�   2�x 3�y �	  T �  F T  "�  "�   3'i 3Ee T 
  F T  "�  "�    4�  	��J     
  
  �  
  4�  	��K       *
    5
  5�   6�   5b  6  5  b  5�   �   g  p
  7Ln   7uh 5  �i Jf �
  84  	J     '�n $  �n   9�n �q �
  �
  $    �g <l �
  $  "
    :�w +�v #  :�r ,�p (   �
  ;
  :  <<    =�  >�u ?Å �   @7� f  l  �   @�� |  �  �   $w !
�    $G� $�     A	:  BH  ?  �  (  �  T  �  5�  5T  BU  Bg  C    x`F     �       �  D�  �  �hEs '
  �d F0	  O`F     (       �X  T �   Ea @
  �hEb #@
  �` G_  +H     �      ��  P T  T <   HH N�  ��H��  N$<   ��Hs N1z  ��H�s N?�   ��H��  O�   ��HH� O�   ��HZX  O#
  ��~I]� P
  �XIB� S�  ��Jk T�   ��K�+H     E       A  Ji a�   �l KM,H     -       d  Ji d�   �h Lz,H     0       Ji f�   �d  ;
  �  <<    G�  �*H     W       �&  P T  T <   HH x�  �hH��  x!<   �`H�s x-�   �\H��  x8�   �XHH� y�   �THZX  y
  �PMN�f {	<     G�  *H     �       �}  T <   F T  Hݰ  �<   �hEfo �/g  �`HH �6�  �X C#  �  �\F     �       ��  D�  �  �hEstr 1
  �` GV	  �)H     }       �  F T  Hݰ  � �
  ��Efo �7g  ��HH �>�  �� G}	  z\F     *       �[  F T  Hݰ  � 
  �hEfo �7g  �`HH �>�  �X C�  z  T\F     &       ��  D�  �  �hH�d M
  �` 5�  G�	  M)H     E       ��  T �  F T  Oݰ  3�  �HOH 3!�  �@ 5

  G�	  �[F     E       �6  T 
  F T  Oݰ  3�  �HOH 3!�  �@ Pa  D  Z  Q�  �  R$s �   S6  �u }  �[F     4       ��  TD  �hTM  �` PQ  �  �  Q�  0
  Q0  �    S�  Gk �  �[F            ��  T�  �h P7  �  �  Q�  0
   S�  �t   �[F            �  T�  �h C�  >  T[F     ,       �S  D�  �  �hU	  �  Cz  y  $)H     )       ��  T �  D�  �  �hHݰ  �  �` C�  �  [F     )       ��  T 
  D�  �  �hHݰ  
  �` P�  �  �  Q�  �  Q0  �    S�  �t   �ZF            �$  T�  �h C�  C  �ZF     )       �P  D�  �  �` P�  ^  t  Q�  ;
  R�L *L
   VP  [q �  vZF     V       ��  T^  �hTg  �` P(  �  �  Q�  ;
  Q0  �    V�  r �  ZZF            ��  T�  �h Pm      Q�  ;
   V�  �d 0  6ZF     #       �9  T  �h Wux <1�(H     .       �v  Eptr <Nv  �XI�� =�  �h �   Xax 00�   �(H     J       ��  Eptr 0Mv  �XI�� 1�  �h Yy +1F(H     f       �Zl  �  ,(H            �  D�  �  �h CV  "  �'H     J       �<  D�  �  �XJv �   �l C�  [  <�F     6       ��  D�  v
  �`Ec 63�  �\I�  7g  �h [  2�  �  Q�  v
  Q0  �    V�  �o �  ZF            ��  T�  �h 5N  [5  2�  �  Q�  v
  "�   V�  �e   �YF     �       �/  T�  �hT�  �` Pt  =  G  Q�  v
   V/  w j  &YF     \       �s  T=  �h \6r kv �  YF            ��  H�  #0   �hEp /�  �` &E �
   %U   :;9I  $ >  $ >  & I  :;9   :;9I8   :;9I8  	   
 I  :;9n  I  ! I/  ;   .?n4<d   I4  4 :;9I?<   :;9I  I   I    :;9   :;9I8   :;9I8  :;9   :;9I  >I:;9  (   (    <  :;9    :;9I8  !4 :;9I?  "4 :;9I?  #:;9  $.?:;9n2<d  %.?:;9nI2<d  & :;9I82  ' :;9I82  (/ I  ).?n42<d  *4 I?4<  +. 4@�B  ,.Gd   - I4  .  /4 :;9I  0.1nd@�B  1 1  21  34 1  41  54 1  6.4@�B  7 :;9I  8.Gd@�B  9 I4  : :;9I  ;4 :;9I  <  =4 :;9I  >.Gd@�B  ?.G:;9d   @.1nd@�B  A  B.?:;9I@�B  C4 :;9I  D4 :;9I  E.?:;9n@�B  F.?:;9nI@�B  G I   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   4 :;9I  !.?:;9'I@�B  " :;9I�B  #4 :;9I�B  $��1  %�� �B  &��1  '1R�BXYW  ( 1�B  )  *4 1  +4 1�B  ,�� 1  -.?:;9'@�B  . :;9I�B  /4 :;9I�B  0.?:;9'   1 :;9I  24 :;9I  34 :;9I  4.1@�B  5. ?<n:;9  6. ?<n:;9   �� �B   1�B  4 1�B   :;9I8   :;9I�B  4 :;9I�B   I   I  	 :;9I8  
(   U  ��  ��1   :;9I  4 :;9I   :;9I  ��1  1R�BUXYW   :;9I  4 1  .?:;9'I@�B   :;9I8   :;9I�B  4 :;9I�B  4 :;9I�B  'I  .1@�B  1R�BXYW  :;9   :;9I  4 :;9I    1  ! :;9I  "4 :;9I�B  #1R�BUXYW  $:;9  %4 :;9I  &  'U  (4 :;9I  ).?:;9'I@�B  *4 :;9I  + 1  ,���B1  -
 :;9  .& I  /1R�BUXYW  0�� 1�B  1I  2! I/  3(   44 1  5'  6.?:;9'@�B  71R�BUXYW  81R�BXYW  9��  :  ; :;9I�B  <1  =.:;9'I   >
 :;9  ?  @���B  A :;9I  B :;9I�B  C.:;9'I@�B  D1U  E4 :;9I  F :;9I8  G
 1  H.?:;9'   I.?:;9'I   J4 1  K�� 1  L. ?<n:;9  M4 :;9I  N1R�BXYW  O :;9I  P4 :;9I  Q$ >  R>I:;9  S :;9I  T.:;9'   U :;9I8  V.:;9'I@�B  W.?:;9'I   X <  Y.?:;9'   Z.:;9'I   [4 :;9I  \
 1  ] :;9I8  ^>I:;9  _:;9  ` :;9I  a.:;9'   b.?:;9'@�B  c4 :;9I?<  d.?:;9'I@�B  e
 :;9  f�� �B1  g���B1  h.:;9'@�B  i:;9  j :;9I  k :;9I  l(   m :;9I  n4 :;9I  o1U  p.?:;9'I@  q.:;9'@�B  r1R�BXYW  s���B  t1  u.1@�B  v. ?<n:;  w. ?<n:;9  x%  y$ >  z   {&   |>I:;9  }4 :;9I?<  ~5 I  :;9  �4 :;9I
  �.?:;9'@�B  �4 :;9I  �
 :;9  �1UXYW  �.:;9'I@�B  �
 :;9  � :;9I  ����B  �4 1   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   :;9   :;9I8  I  ! I/  4 :;9I?<  .?:;9'I    :;9I  !4 :;9I  "  #.?:;9'I@�B  $ :;9I�B  %4 :;9I  &  '4 :;9I�B  (���B  )�� �B   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  >I:;9  I  ! I/   4 :;9I?<  !.?:;9'I@�B  " :;9I  #.?:;9'@�B  $ :;9I   %   :;9I  $ >  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I  # :;9I8  $:;9  % :;9I8  & :;9I8  '(   (4 :;9I  )4 :;9I  *4 G:;  +4 G:;9  ,.:;9'I   - :;9I  .4 :;9I  /4 :;9I  0.:;9'   1
 :;9  2.:;9'I@�B  3 :;9I�B  44 :;9I�B  5
 :;9  6  74 :;9I�B  8��1  9�� �B  :��  ;��1  <.:;9'I@�B  = :;9I  > :;9I�B  ?4 :;9I�B  @4 :;9I�B  A.:;9'I   B :;9I  C4 :;9I  D
 :;9  E  F4 :;9I  G�� �B1  H.:;9'@�B  I :;9I  J1R�BXYW  K 1�B  L  M4 1�B  N1R�BUXYW  OU  P�� 1  Q4 :;9I  R  S��  T.:;9'@�B  UU  V1XYW  W 1  X4 1  Y1R�BUXYW  Z4 1  [
 1  \1UXYW  ]1  ^1U  _ :;9I  `.:;9'@�B  a.?:;9'I@�B  b :;9I�B  c1R�BXYW  d�� 1�B  e
 1  f :;9I  g :;9I  h4 :;9I  i. :;9'   j���B1  k.:;9'   l>I:;9  m1U  n1  o.:;9'I@�B  p4 :;9I  q
 :;9  r1R�BUXYW  s���B1  t.1@�B  u 1  v���B  w4 1  x. ?<n:;9  y. ?<n:;9  z. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  #:;9  $ :;9I  % :;9I8  &>I:;9  '4 :;9I  (4 :;9I  )4 G:;9  *.:;9'I   + :;9I  ,4 :;9I  -
 :;9  .  /4 :;9I  0  1.:;9'   2 :;9I  34 :;9I  4.:;9'I   54 :;9I  6
 :;9  7
 :;9  8.:;9'I@�B  9 :;9I�B  :4 :;9I�B  ;4 :;9I�B  <��1  =�� �B  >��1  ?.:;9'@�B  @ :;9I  A.:;9'I@�B  B4 :;9I�B  C :;9I�B  D
 :;9  EU  FU  G�� 1  H.:;9'@�B  I.:;9'I@�B  J  K  L :;9I  M :;9I�B  N�� 1�B  O��  P4 :;9I�B  Q1R�BUXYW  R 1�B  S4 1  T
 1  U��  V4 1�B  W
 1  X1U  Y1  Z.:;9'   [.:;9'I@�B  \4 :;9I  ]1R�BUXYW  ^.:;9'@�B  _���B1  `4 :;9I  a1R�BXYW  b 1  c1R�BXYW  d1U  e :;9I  f :;9I  g :;9I  h.1@�B  i 1  j1  k4 1  l.1@  m.1@�B  n. ?<n:;9  o. ?<n:;9  p. ?<n:;   %   :;9I  $ >  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  # :;9I8  $:;9  % :;9I  &4 G:;  '>I:;9  (4 :;9I  )4 G:;  *4 :;9I  +.:;9'@�B  , :;9I  -.:;9'I@�B  .4 :;9I�B  /.:;9'@�B  0 :;9I�B  1  24 :;9I�B  31R�BUXYW  4 1�B  5U  64 1�B  71R�BXYW  8��1  9�� �B  :��1  ;  <��  =
 :;9  >U  ?��  @4 1  A1U  B
 1  C1  D�� 1  E1R�BUXYW  F 1  G1R�BXYW  H.:;9'   I :;9I  J4 :;9I  K  L4 :;9I  M.:;9'I   N.:;9'I@�B  O :;9I�B  P�� 1�B  Q.:;9'I@�B  R :;9I�B  S4 :;9I�B  T4 :;9I�B  U
 :;9  V.:;9'@�B  W :;9I  X.:;9'@�B  Y�� �B1  Z.:;9'I   [ :;9I  \4 :;9I  ]
 :;9  ^  _1  `���B  a :;9I  b :;9I�B  c :;9I  d4 :;9I  e4 :;9I  f
 :;9  g
 :;9  h.:;9'   i
 :;9  j1R�BUXYW  k :;9I  l4 :;9I  m4 :;9I  n4 :;9I  o���B1  p���B1  q.1@�B  r 1  s4 1  t
 1  u.1@  v1R�BXYW  w1U  x. ?<n:;9  y. ?<n:;9  z. ?<n:;   %   :;9I   I  :;9   :;9I8  'I   I     	$ >  
'  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I  $ >  & I  4 :;9I?<   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  # :;9I8  $:;9  % :;9I  & :;9I8  '>I:;9  (4 :;9I  )4 :;9I  *4 G:;  +.:;9'I@�B  , :;9I�B  -���B1  .�� �B  / :;9I  0 :;9I  14 :;9I  24 :;9I�B  34 :;9I�B  4.:;9'   5 :;9I  6  74 :;9I  8.:;9'I   9 :;9I  :4 :;9I  ;4 :;9I  <
 :;9  =  >! I/  ?.:;9'@�B  @ :;9I  A.:;9'I@�B  B4 :;9I�B  C.:;9'I   D
 :;9  E4 :;9I  F.:;9'@�B  G  H��1  I��1  J :;9I�B  K�� 1�B  L��  M.:;9'   N.:;9'I@�B  O  P
 :;9  Q :;9I�B  R4 :;9I�B  SU  T��  U�� 1  VU  W1R�BUXYW  X 1  Y 1�B  Z4 1�B  [1R�BXYW  \1R�BXYW  ]
 :;9  ^1R�BUXYW  _1R�BXYW  ` :;9I  a.1@  b.1@�B  c1  d4 1  e1U  f
 1  g4 1  h
 1  i1  j1U  k1R�BUXYW  l. ?<n:;9  m. ?<n:;9  n. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I8  #4 G:;9  $4 :;9I  %4 :;9I  &.:;9'I   ' :;9I  (4 :;9I  )
 :;9  *  +4 :;9I  ,  - :;9I  ..:;9'   /.:;9'   0 :;9I  1 :;9I  24 :;9I  34 :;9I  4.:;9'I@�B  5 :;9I�B  64 :;9I�B  7
 :;9  8U  9U  :4 :;9I�B  ;  <��1  =�� �B  >��1  ?  @1R�BUXYW  A 1  B 1�B  C4 1�B  D1R�BXYW  E1R�BUXYW  F�� 1  G
 1  H
 1  I1  J1U  K1U  L4 1  M1UXYW  N1UXYW  O1  P.:;9'@�B  Q.:;9'I@�B  R :;9I�B  S4 :;9I�B  T1R�BUXYW  U4 1  V4 :;9I�B  W1R�BUXYW  X1R�BXYW  Y1R�BXYW  Z��  [ :;9I�B  \.:;9'I   ]
 :;9  ^�� 1�B  _���B1  ` :;9I  a
 :;9  b.:;9'@�B  c.1@�B  d. ?<n:;9  e. ?<n:;9  f. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/   :;9I   4 :;9I?<  !:;9  " :;9I8  #4 :;9I  $4 G:;9  %:;9  & :;9I  ' :;9I8  (>I:;9  ).:;9'   * :;9I  +4 :;9I  ,.:;9'I   -
 :;9  .  /4 :;9I  0  1.:;9'@�B  2 :;9I�B  34 :;9I�B  44 :;9I�B  5
 :;9  6  7��  8�� �B  9��  :��1  ;4 :;9I  <U  =��1  >.:;9'@�B  ? :;9I�B  @4 :;9I�B  A.:;9'I   B :;9I  C.:;9'   D :;9I  E4 :;9I  F
 :;9  G�� �B1  H.:;9'I@�B  I�� 1  J :;9I�B  K :;9I  L.:;9'I@�B  M1R�BUXYW  N 1�B  OU  P4 1  Q4 1�B  R
 1  S1R�BUXYW  T1U  U1U  V1  W4 :;9I  X.:;9'I@�B  Y���B1  Z :;9I  [4 :;9I�B  \.1@�B  ] 1  ^1  _ 1  `  a4 1  b. ?<n:;9  c. ?<n:;9  d. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I8  #4 :;9I  $4 :;9I  %4 :;9I  &4 G:;9  '.:;9'I@�B  ( :;9I�B  )���B1  *�� �B  + :;9I  ,4 :;9I�B  -4 :;9I�B  .
 :;9  /U  0  1��1  2.:;9'I   3 :;9I  4 :;9I  5��1  61R�BUXYW  7 1�B  8 1  9U  :4 1  ;4 1�B  <
 1  =1U  >�� 1  ?1R�BUXYW  @4 1  A1U  B.:;9'   C
 :;9  D  E  F4 :;9I  G.:;9'I   H :;9I  I4 :;9I  J.:;9'@�B  K :;9I�B  L4 :;9I�B  M.1@�B  N4 1  O1  P  Q
 1  R. ?<n:;9  S. ?<n:;9  T. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I  #:;9  $ :;9I8  % :;9I8  &4 :;9I  '4 :;9I  (4 G:;9  ).:;9'   * :;9I  + :;9I  ,  -4 :;9I  ..:;9'I@�B  / :;9I�B  04 :;9I�B  1
 :;9  2U  3��1  4�� �B  5�� 1�B  6��1  71R�BUXYW  8 1�B  9U  :4 1  ;4 1�B  <1U  =1  >�� 1  ?
 1  @1U  A4 1  B.:;9'I   C :;9I  D4 :;9I  E4 :;9I  F :;9I  G
 :;9  H4 :;9I�B  I  J.:;9'I   K4 :;9I  L.:;9'@�B  M :;9I  N���B1  O1R�BXYW  P :;9I�B  Q4 :;9I  R1R�BXYW  S  T  U.:;9'I@�B  V :;9I�B  W :;9I  X4 :;9I�B  Y4 :;9I�B  Z
 :;9  [.:;9'@�B  \.1@�B  ] 1  ^
 1  _. ?<n:;9  `. ?<n:;  a. ?<n:;9   %   :;9I  $ >  & I  $ >     :;9   :;9I8  	 I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  ! :;9I  ":;9  #:;9  $ :;9I8  % :;9I8  &! I/  '4 :;9I  (4 :;9I  )4 :;9I  * :;9I8  +4 :;9I  ,4 :;9I  -:;9  . :;9I8  /4 G:;9  0.:;9'I@�B  1 :;9I�B  2���B1  3�� �B  4 :;9I  54 :;9I�B  6
 :;9  71R�BUXYW  8 1�B  9U  :4 1  ;��1  <4 :;9I�B  =4 :;9I  >��1  ?.:;9'I   @ :;9I  A :;9I  B4 :;9I  CU  D1R�BUXYW  E1R�BXYW  F  G  H4 1  I4 1�B  J1R�BXYW  K 1  L1R�BUXYW  M1U  N1  O�� 1  P
 1  Q��  R.:;9'@�B  S.:;9'I   T :;9I  U4 :;9I  V  W4 :;9I  X.:;9'I@�B  Y :;9I�B  Z :;9I  [4 :;9I�B  \4 :;9I�B  ]
 :;9  ^.:;9'@�B  _.:;9'   `
 :;9  a�� 1�B  b
 1  c :;9I�B  d :;9I  e.1@�B  f4 1  g1  h1U  i 1  j 1  k. ?<n:;9  l. ?<n:;9  m. ?<n:;   %  $ >   :;9I  $ >  & I     :;9   :;9I8  	 I  
4 :;9I?<  I  ! I/   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   5 I  >I:;9  :;9    :;9I8  !4 :;9I?<  ":;9  # :;9I  $ :;9I8  %:;9  &4 :;9I  '4 :;9I  (4 G:;  )4 :;9I?  *4 :;9I?  +4 G:;9  ,.:;9'I@�B  - :;9I�B  . :;9I�B  / :;9I  04 :;9I�B  1  21R�BXYW  3 1�B  4  54 1�B  6
 1  71  8��1  9�� �B  :U  ;��1  <�� 1  =1R�BUXYW  >U  ?4 1  @.:;9'I   A :;9I  B :;9I  C4 :;9I  D4 :;9I  E
 :;9  F  G4 :;9I  H4 :;9I�B  I
 :;9  J 1  K4 1  L1U  M1R�BUXYW  N��  O4 :;9I  P :;9I  Q.:;9'   R���B1  S.:;9'@�B  T.:;9'I@�B  U :;9I�B  V4 :;9I�B  W
 :;9  X4 :;9I�B  Y��  Z
 :;9  [  \
 1  ]1  ^1U  _.:;9'I   ` :;9I  a4 :;9I  b4 :;9I  c.:;9'@�B  d4 :;9I  e
 :;9  f�� �B1  g :;9I�B  h1R�BUXYW  i :;9I  j :;9I  k.:;9'   l���B  m1R�BXYW  n���B1  o���B  p1XYW  q.:;9'I@�B  r :;9I  s1R�BXYW  t.1@�B  u 1  v.1@�B  w1XYW  x4 1  y. ?<n:;9  z. ?<n:;9  {. ?<n:;   4 1�B  (   �� �B   1�B  4 :;9I�B  4 :;9I   :;9I8  (   	4 :;9I?<  
 :;9I8   I  4 G   I   :;9I  U  4 :;9I?<  ��1  4 G:;9   :;9I   :;9I  ��1  4 :;9I  4 :;9I  4 :;9I�B   :;9I�B    4 1   1  1R�BUXYW  4 :;9I�B  :;9   U  ! :;9I  "4 1  #  $  %& I  &'I  '1U  (I  )4 G:;9  *4 :;9I  + :;9I�B  ,:;9  -! I/  .1U  /(   0'  1 :;9I8  2 :;9I8  3  4 :;9I  51  6 :;9I8  7.:;9'   8�� 1�B  94 :;9I  :4 :;9I�B  ;1R�BUXYW  <.1@�B  =.:;9'@�B  >. ?<n:;9  ? :;9I8  @.:;9'I@�B  A4 :;9I  B
 1  C1R�BUXYW  D :;9I  E.:;9'I   F1R�BXYW  G :;9I�B  H1  I
 :;9  J
 :;9  K>I:;9  L$ >  M1R�BXYW  N :;9I  O���B1  P.:;9'I   Q!   R4 G:;  S.:;9'I@�B  T. ?<n:;9  U:;9  V.:;9'@�B  W�� 1  X��  Y:;9  Z.:;9'   [
 :;9  \ 1  ] <  ^>I:;9  _4 G:;  ` :;9I  a :;9I�B  b.?:;9'I   c
 1  d :;9I  e>I:;9  f(   g:;9  h4 1  i1XYW  j1XYW  k1R�BXYW  l%  m$ >  n   o:;9  p&   q4 :;9I?  r1R�BUXYW  s.?:;9'I@�B  t.?:;9'   u��  v.:;9'I  w4 :;9I  x1UXYW  y.:;9'  z
 :;9  {.:;9'@�B  |4 :;9I  }1R�BXYW  ~ 1  . ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   :;9  ! :;9I8  ">I:;9  #(   $4 :;9I  %4 :;9I?  &.:;9'   ' :;9I  (.:;9'@�B  ) :;9I�B  *4 :;9I  +4 :;9I�B  ,4 :;9I�B  -1R�BXYW  . 1�B  /  04 1  1��1  2�� �B  3 :;9I  41R�BXYW  5�� 1  6.:;9'I   74 :;9I  8  94 :;9I  :
 :;9  ; :;9I  <.:;9'I@�B  = :;9I�B  >
 :;9  ?U  @1R�BUXYW  A4 1�B  B4 1  C
 1  D
 1  E1R�BXYW  F1  G1R�BUXYW  H1U  I�� 1�B  J4 :;9I  K1U  L 1  M  N.:;9'I@�B  O :;9I�B  P4 :;9I�B  Q.:;9'I   R :;9I  S4 :;9I  T.:;9'@�B  U1R�BUXYW  V :;9I�B  W4 :;9I�B  X
 :;9  Y.:;9'   Z :;9I  [4 :;9I  \
 :;9  ] :;9I  ^1R�BXYW  _1R�BUXYW  `��1  a1  b  cU  d.?:;9'I   e.1@�B  f 1  g4 1  h���B1  i1UXYW  j�� �B1  k. ?<n:;9  l. ?<n:;9   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I   :;9I8  :;9   :;9I8  >I:;9  (   (    <   :;9I8  '   I  'I  &   :;9   :;9I  >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !4 G:;9  "4 G:;  #.:;9'I@�B  $ :;9I�B  %4 :;9I  &4 :;9I�B  '
 :;9  (��1  )�� �B  *��  +��1  ,.:;9'@�B  -���B1  ..:;9'I   / :;9I  04 :;9I  1���B  2��  3.:;9'I@�B  4 :;9I�B  54 :;9I�B  64 :;9I  7  84 :;9I�B  91R�BUXYW  : 1�B  ;U  <4 1�B  =1R�BUXYW  >! I/  ? :;9I  @.:;9'@�B  A.:;9'   B :;9I  C.:;9'I   D4 :;9I  E4 :;9I  F1U  G 1  H
 1  I
 1  J1  K4 1  L1U  M4 1  N1R�BXYW  O4 :;9I  P
 :;9  Q  R :;9I�B  S
 :;9  T  U :;9I  V :;9I  W  XU  Y�� 1  Z.:;9'I@�B  [
 :;9  \.1@�B  ]4 1  ^. ?<n:;9  _. ?<n:;9   %  $ >   :;9I  $ >  5 I     :;9   :;9I8  	 I  
& I  4 :;9I?<  I  ! I/   :;9I   :;9I8  >I:;9  (   :;9   :;9I8  'I   I  >I:;9  (    <   :;9I8  '  &   :;9   :;9I  >I:;9  :;9    :;9I8  !4 :;9I?<  "4 :;9I  #4 G:;9  $4 G:;  %.:;9'I@�B  & :;9I�B  '���B1  (�� �B  ).:;9'I@�B  * :;9I�B  +4 :;9I  ,4 :;9I�B  -
 :;9  .U  /4 :;9I�B  0��  1��1  2��1  34 :;9I�B  4��  5.:;9'@�B  6.:;9'I   7 :;9I  84 :;9I  9
 :;9  :���B  ; :;9I  <.:;9'@�B  =4 :;9I  >4 :;9I�B  ?U  @1R�BXYW  A 1�B  B  C4 1�B  D1U  E! I/  F.:;9'   G :;9I  H4 :;9I  I  J :;9I�B  K  L�� 1�B  M :;9I  N
 :;9  O
 :;9  P�� 1  Q.1@�B  R 1  S4 1  T4 1  U
 1  V1R�BUXYW  W4 1  X1  Y. ?<n:;9  Z. ?<n:;9  [. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<   :;9I8  :;9  :;9   :;9I  (    I  !! I/  "4 :;9I  #4 :;9I  $! I/  %:;9  & :;9I8  ' :;9I8  (.?:;9'I@�B  ) :;9I�B  *4 :;9I  +4 :;9I�B  ,��1  -�� �B  .��1  /4 :;9I�B  0
 :;9  1U  21R�BUXYW  3 1�B  4U  54 1�B  61R�BUXYW  74 1  8�� 1  9
 1  :.:;9'I   ; :;9I  <4 :;9I  =.:;9'I@�B  >���B1  ?.:;9'@�B  @ :;9I  A  B :;9I�B  C��  D.:;9'   E
 :;9  F.:;9'I@�B  G :;9I�B  H4 :;9I�B  I  J4 :;9I�B  K.:;9'@�B  L :;9I�B  M1R�BXYW  N1R�BUXYW  O.:;9'   P :;9I  Q.:;9'I   R4 :;9I  S4 :;9I  T.:;9'I@�B  U1R�BUXYW  V1R�BXYW  W1U  X��  Y1R�BXYW  Z :;9I  [  \4 :;9I  ].:;9'@�B  ^ :;9I  _4 :;9I  `.1@�B  a.1@�B  b 1  c 1  d4 1  e 1  f
 1  g1U  h1  i1R�BXYW  j  k. ?<n:;9  l. ?<n:;9  m. ?<n:;  n6    %  $ >   :;9I  $ >     :;9   :;9I8   I  	4 :;9I?<  
 :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I  & I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<  >I:;9  I  ! I/  :;9   :;9I8    :;9I8  ! :;9I8  "! I/  #.?:;9'I@�B  $ :;9I�B  %4 :;9I�B  &
 :;9  '
 :;9  (U  )4 :;9I  *4 :;9I  +��1  ,�� �B  -��1  .4 :;9I�B  /1R�BUXYW  0 1�B  1U  24 1�B  34 1  4.?:;9'@�B  5 :;9I�B  64 :;9I�B  71R�BUXYW  8 :;9I  91R�BXYW  :.?:;9'   ; :;9I  <.:;9'I   =4 :;9I  >.:;9'I@�B  ?4 :;9I  @4 :;9I�B  A1R�BUXYW  B4 :;9I  C1R�BUXYW  D
 1  E.:;9'I@�B  F
 1  G1U  H1U  I.:;9'@�B  J :;9I  K
 :;9  L  M4 :;9I  N  O4 :;9I  P.:;9'   Q
 :;9  R
 :;9  S.1@�B  T 1  U. ?<n:;9  V. ?<n:;9  W. ?<n:;   �� �B   1�B  (    :;9I8   :;9I8   I   I  4 1�B  	4 :;9I�B  
 :;9I8   :;9I  ��1  ��1   :;9I   :;9I�B   :;9I  4 :;9I�B  1R�BUXYW   :;9I8  4 :;9I  'I  �� 1  U   :;9I  :;9  :;9   1  4 :;9I  4 :;9I  1R�BXYW  I   ! I/  !4 :;9I  "& I  #  $'  %U  &  '.:;9'I   (4 :;9I�B  ) :;9I  *.1@�B  + :;9I8  ,.:;9'@�B  -.:;9'I@�B  . :;9I�B  /.:;9'   04 1  1  2.:;9'I   3�� 1�B  4(   5.:;9'   64 1  7 :;9I�B  84 :;9I  9 :;9I  : :;9I  ;1R�BXYW  <
 :;9  =1  > :;9I  ? 1  @1R�BXYW  A4 :;9I?<  B��  C1R�BXYW  D1U  E :;9I8  F
 1  G.:;9'I@�B  H���B1  I. ?<n:;9  J :;9I8  K1R�BUXYW  L:;9  M1U  N1R�BUXYW  O>I:;9  P:;9  Q :;9I  R4 :;9I�B  S$ >  T
 :;9  U <  V>I:;9  W1R�BUXYW  X4 :;9I  Y.:;9'@�B  Z>I:;9  [1  \��  ]  ^
 1  _4 1  ` 1  a4 G:;  b4 :;9I  c :;9I  d4 :;9I?  e
 :;9  f���B  g. ?<n:;9  h4 G:;9  i4 :;9I  j:;9  k :;9I  l :;9I  m:;9  n4 G:;  o.:;9'@�B  p
 :;9  q4 :;9I  r. ?<n:;  s%  t$ >  u   v&   w4 :;9I?<  x:;9  y(   z 1  {�� �B1  | :;9I�B  }.:;9'I@�B  ~
 :;9  1XYW  �1XYW  �
 :;9  �
 :;9  �1UXYW  �.1@�B   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   ! I/  !4 G  "4 :;9I  #4 :;9I  $4 G:;  %.:;9'I@�B  & :;9I�B  '���B1  (�� �B  ) :;9I  * :;9I  +4 :;9I�B  ,
 :;9  -U  .4 :;9I�B  /U  01UXYW  1 1  24 1�B  3��1  4���B  5��1  6.:;9'   7 :;9I  84 :;9I  9.:;9'I@�B  : :;9I�B  ; :;9I  <4 :;9I�B  = :;9I�B  >  ?4 :;9I�B  @1R�BUXYW  A 1�B  B4 1  C
 1  D
 1  E1XYW  F  G.:;9'I   H4 :;9I  I
 :;9  J  K  L.1@�B  M 1  N1U  O1  P. ?<n:;9  Q. ?<n:;9   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<  .?:;9'@�B   :;9I�B  ���B1  �� �B  .?:;9'I@�B   4 :;9I�B  !��1  ".?:;9'I@�B  # :;9I�B  $4 :;9I�B  %��1  &.:;9'I@�B  '���B1  (.:;9'@�B  )�� 1  *. ?<n:;9   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !4 :;9I
  ".?:;9'I@�B  # :;9I�B  $4 :;9I�B  %�� 1  &U  '4 :;9I  (1R�BUXYW  ) 1�B  *��1  +�� �B  ,4 :;9I�B  -U  .4 :;9I  /  0  11R�BXYW  24 1�B  3.:;9'I   4 :;9I  54 :;9I  64 :;9I  7��1  81R�BUXYW  94 1  :1  ;1  <1U  =4 1  >.:;9'I   ? :;9I  @4 :;9I  A4 :;9I  B  C  D.?:;9'I@�B  E :;9I�B  F4 :;9I�B  G4 :;9I  H4 :;9I�B  I.?:;9'  J.?:;9'   K.1@�B  L 1  M. ?<n:;9  N. ?<n:;   %  . @   %  $ >   :;9I  $ >  .?:;9'@�B   :;9I   %U  $ >   :;9I  ;   $ >  & I     I  	! I/  
9:;9  :;9  .?:;9n<�d   I4  .?:;9n<d   I  4 :;9nI?<  .?:;9nI<  . ?:;9nI<  . ?:;9n�<  .?:;9n<  .?:;9n�<  9:;   :;9I?<l   .?:;9nI<d  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I   9:;9  ! :;9  "4 :;9I<l  #9:;9  $4 :;9I<l  %m>I:;9  &(   '(   (:;9  ):;9  * :;9I  +.?:;9n<d  ,.?:;9n2<d  -.?:;9nI2<d  . :;9I8  /.?n4<d  0.?n4<d  1.?:;9n<  2 <  3.?:;9n<�d  4.?:;9nI<�d  5 :;9I82  6.?:;9nI<d  7/ I  80 I  9.?:;9n<  :.?:;9n<  ;4 G  < I  =B I  >4 nG  ?4 G  @.Gd@�B  A I4  B :;9I  C.G@�B  D.G@�B  E :;9I  F4 :;9I  G4 :;9I  H  I  J  K4 :;9I  L :;9I  M.Gd   N I4  O :;9I  P.1nd@�B  Q 1  R I  S.1nd@�B  T. ?:;9n@�B  U. ?:;9I@�B  V.?:;9n@�B  W. G@�B  X4 I4  Y.G:;9d   Z.?:;9nI@�B   %  $ >  ;   9:;  :;9   :;9I?<l    :;9I  .?:;9nI<d  	 I4  
/ I  0 I  & I  ��  / I  4 :;9nI?<l   4 nG   I  $ >  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  :;9  :;9   :;9I  .?:;9n<d  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d    :;9I8  !9 :;9  " <  # :;9I82  $/ I  %0 I  &:;9  '4 G  ( I  )B I  *4 nG  +9:;9  ,.?:;9n<�d  -4 :;9nI?<  .4 G:;9  /4 G  0.G:;9d@�B  1 I4  2 :;9I   %U  $ >   :;9I  ;   9:;  :;9   :;9I?<l   .?:;9nI<d  	 I4  
/ I  0 I  & I  ��  / I  4 :;9nI?<l   4 nG   I     $ >  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  *.?:;9n<�d  +.?:;9nI<�d  , :;9I82  -.?:;9nI<d  ./ I  /0 I  0.?:;9nI<  1.?:;9n<  2.?:;9n<  34 G  4 I  5B I  64 nG  7.?:;9n<�d  84 :;9nI?<  9I  :! I/  ;4 G  <.Gd@�B  = I4  > :;9I  ?.G@�B  @.G@�B  A :;9I  B4 :;9I  C4 :;9I  D  E  F  G4 :;9I  H :;9I  I.Gd   J I4  K :;9I  L.1nd@�B  M 1  N I  O.1nd@�B  P.?:;9@�B  Q.G:;9d   R.?:;9nI@�B   %   :;9I  $ >  .?:;9I@�B   :;9I  4 :;9I     I  	& I  
 :;9I  4 :;9I       7 I  &   $ >    %    I   I4   :;9I  4 :;9I  / I  & I   :;9I   I4  	.Gd@�B  
4 :;9I  4 :;9I   :;9I8   I   I   :;9I  4 :;9I   1    .G@�B  .?:;9n2<d  4 I4  :;9   I4  .?:;9n<d  .?:;9I@�B  .?:;9nI<   :;9I  $ >  .?:;9n2<d  I  .Gd    .?:;9nI<d  !! I/  " :;9I  #  $.?:;9I@�B  %(   &.?:;9nI2<d  '.?:;9n<d  ( :;9  )4 nG  *.1nd@�B  + :;9I  ,.?:;9n<�d  -.?:;9nI<�d  ..G@�B  / :;9I8  0.?:;9nI2<d  1 :;9I?<l   2.Gd@�B  3 :;9I82  4/ I  5.1nd@�B  64 G  7m>I:;9  8.?:;9n<  9.?:;9nI2<  : :;9I82  ;0 I  <4 G  =7 I  > I  ?.?:;9�@�B  @4 :;9I?<  A:;9n  B :;9  C.?:;9n<d  D9:;9  E9  F: :;9  G I8  H :;9I?<l   I.?:;9nI<d  J :;9I  KB I  L
 :;9  MU  N.?:;9@�B  O :;9I?<l   P :;9I?<l   Q4 :;9I<l  R(   S:;9  T.?:;9nI<d  U <  V4 :;9I<l  W.?:;9nI<  X.?:;9nI2<  Y.?:;9n2<�d  Z.?:;9n<  [0 I  \��  ]/ I  ^4 :;9nI?<l   _4 nG  `4 :;9nI?<  a.?:;9nI<cd  b4 nG  c.G:;9d   d IJ  e%U  f$ >  g   h9:;9  i:;9  j :;9I?<l   k :;9I82  l :;9I82  m9:;9  n4 :;9I<l  o:;9  p :;9I  q.?n4<d  r.?n4<d  s.?:;9n<  t0 I  u4 :;9I<
l  v:;9  w:;9  x.?:;9nI<  y:;9  z.?:;9nI2<�d  { :;9I?<
l   | :;9I?<l   }:;9  ~ :;9I8  4 Gn  �! I/  �;   �9:;  �&   �.?:;9n<�d  �.?:;9nI<d  �4 :;9I<  �4 :;9I?  �4 nG  �. 4@�B  �.4@�B  �  �4 :;9I  �.?:;9@�B  �.?:;9I@�B  �.?:;9I@�B  �I  �   �. ?:;9I@�B  �.?:;9nI@�B  �4 :;9Il   %U   :;9I  $ >  & I   :;9I  ;   $ >  :;9  	 :;9I8  
9:;   :;9I?<l   .?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I  9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I   .?:;9n<d  !.?:;9n<d  ".?:;9n2<d  # I  $.?:;9nI2<d  %.?n4<d  &9 :;9  '/ I  (.?:;9n<�d  ).?:;9nI<�d  * :;9I82  +.?:;9nI<d  ,0 I  - <  ..?:;9n<  /.?:;9n<  04 G  1 I  2B I  34 nG  49:;9  5.?:;9n<�d  64 :;9nI?<  7 :;9I8  8.?:;9nI<cd  9<  :.?:;9nI<  ;9  <>I:;9  =: :;9  >I  ?! I/  @4 G  A.Gd@�B  B I4  C :;9I  D.G@�B  E :;9I  F :;9I  G.Gd   H I4  I :;9I  J.1nd@�B  K 1  L I  M.Gd@�B  N  O4 :;9I  P :;9I  Q.1nd@�B  R.?:;9I@�B  S4 I4  T :;9I  U4 :;9I  V.?:;9I@�B  W.G@�B  X4 :;9I  Y.G:;9d     I   I4   :;9I  / I   I4  & I   :;9I8  .Gd@�B  	4 :;9I  
 I  .?:;9nI2<d   I   1  .?:;9n2<d  4 :;9I  .G@�B  4 :;9I   :;9I  4 :;9I   I4  :;9   :;9I  .?:;9n<d    .Gd   .?:;9nI<  $ >  .?:;9n2<d  .Gd@�B   :;9I  .?:;9nI<d   .?:;9n<d  ! :;9  ".1nd@�B  #  $ :;9I  %I  &! I/  '.G@�B  (.1nd@�B  ).?:;9n<�d  *.?:;9nI<�d  +/ I  , :;9I  - :;9I?<l   .4 nG  /(   0.?:;9nI2<d  14 :;9I?<  2 :;9I82  3 :;9I82  44 I4  5.?:;9n<  64 G  7B I  8.?:;9nI2<  90 I  ::;9  ;.?:;9n<  <4 G  =.?:;9I@�B  > :;9  ?9:;9  @9  A: :;9  Bm>I:;9  C I8  D :;9I?<l   E.?:;9nI<d  F.?:;9n<d  G.?:;9nI2<d  H :;9I  I0 I  J��  K/ I  L4 :;9nI?<l   M.?:;9nI<  N4 :;9I<l  O(   P.?:;9nI2<  Q:;9  R.?:;9nI<d  S.?:;9n2<�d  T4 :;9I<l  U4 nG  V4 :;9nI?<  W.:;9<  X4 nG  Y  Z :;9I  [ :;9I  \.G:;9d   ] IJ  ^%U  _$ >  `   a;   b9:;  c9:;9  d4 :;9I<
l  e:;9  f.?:;9nI<  g:;9  h.?:;9nI2<�d  i :;9I?<
l   j :;9I?<l   k:;9  l :;9I8  m9:;9  n4 :;9I<l  o:;9  p :;9I  q.?n4<d  r.?n4<d  s.?:;9n<  t0 I  u <  v.?:;9nI<d  w&   x.?:;9n<�d  y4 :;9I<  z. :;9<  {. :;9I<  |.:;9I<  }4 :;9I?  ~4 I?4<  4 nG  �4 :;9I  �4 :;9I  �1  �4 1  �1  �4 1  � I  �.?:;9nI@�B   %  4 :;9I?  $ >   I  $ >    I   I4  / I   I4   :;9I  .Gd@�B  & I  4 :;9I  	 :;9I  
4 :;9I   I   :;9I8   I   1  .?:;9nI<d     I4  :;9   :;9I  .?:;9n<d  4 :;9I  .G@�B  4 :;9I    .?:;9n2<d   :;9I  .Gd   .?:;9nI<  / I   :;9I82  .?:;9n2<d   .1nd@�B  !$ >  ".G@�B  #(   $.?:;9n<d  %I  &! I/  '.?:;9nI2<d  (.?:;9nI2<d  ) :;9  * :;9I  +4 I4  ,.1nd@�B  -.?:;9I@�B  ./ I  /.?:;9n<�d  0.?:;9nI<�d  1.Gd@�B  24 G  3 :;9I  4 :;9I?<l   54 nG  6.?:;9n<  74 :;9I?<  8B I  94 G  :4 1  ;4 1  <m>I:;9  =0 I  > I8  ?.?:;9nILM2<d  @.?:;9nILM2<d  A.:;9I<  B :;9  C.?:;9n<d  D9:;9  E9  F.?:;9nI2<  G :;9I82  H.?:;9nI<d  I.?:;9n<  J��  K4 :;9I<  L I  M.?:;9nI<d  N4 :;9I<l  O: :;9  P:;9  Q :;9I?<l   R I82  S :;9I2  T :;9I  U4 G:;9  V.G:;9d   W  X4 I4  Y1  Z IJ  [0 I  \��  ]9 :;9  ^4 :;9nI?<l   _4 :;9I<l  `(   a:;9  b0 I  c.?:;9nI<  d.?:;9nI2<  e:;9  f.?:;9nI<  g.?:;9n2<�d  h.?:;9nI2<d  i.?:;9nI<d  j4 nG  k.?:;9n<�d  l4 :;9nI?<  m:;9  n.?n4<�d  o4 nG  p��:;9  q.?:;9@�B  r.4<d  s.4d@�B  t.I4d@�B  u.4@�B  v4 :;9I  w1  x%U  y$ >  z   {;   |9:;  }9:;9  ~9:;9  4 :;9I<l  �:;9  � :;9I  �.?n4<d  �.?n4<d  �.?:;9n<  �4 :;9I<
l  �:;9  �.?:;9nI2<�d  � :;9I?<
l   � :;9I?<l   �:;9  � :;9I8  �:;9  � I84  �.?:;9nL<d  �.?:;9nILM<d  �4 :;9I<  �.?:;9nI<d  �.?:;9nILM<d  � :;9I82  �.?nL4<d  �.:;9<d  �.:;9<d  �: :;9  �4 nG  �  �I  �   � I  �4 I?4<  �. 4@�B  �.4@�B  �.1d@�B  �1  �.1d@�B  � :;9I  � :;9I  �4 :;9I  �.?:;9nI@�B    I   :;9I   I4  / I   :;9I  4 :;9I  4 :;9I  4 :;9I  	 I4  
& I  4 I4     I  .G@�B     :;9I  4 :;9I  .Gd@�B  .?:;9I@�B   :;9I8   I   1  / I   I  .?:;9n<d  .?:;9n<   :;9I  .?n4<d  :;9   I4  .?:;9n2<d   .?:;9nI2<d  ! :;9I8  ".Gd   #U  $ :;9I  %(   & :;9I  '.?:;9nI<  (.?:;9n<  )B I  *.1nd@�B  +$ >  ,.?:;9n2<d  -I  ..?:;9nI<d  / :;9I82  0   1! I/  2.?:;9n<d  3  44 :;9I  5 :;9  6.G@�B  7.1nd@�B  8.Gd@�B  9.?n4<�d  :.?n4d@�B  ;.?n4d@�B  <:;9  = :;9I?<l   >.?:;9I@�B  ?.?:;9n<�d  @.?:;9nI<�d  A :;9I82  B4 nG  C.?:;9nI2<d  D4 G  E4 :;9I?<  F7 I  G :;9I  HU  I:;9  J :;I8  K :;9I  L��  M/ I  N4 :;9nI?<l   Om>I:;9  P.?:;9nI2<  Q0 I  R:;9  S4 nG  T.?:;9I@�B  U.4<d  V.42<d  W.?:;9nI<  X :;9  Y9:;9  Z9  [: :;9  \ I8  ] :;9I?<l   ^.?:;9nI<d  _.?:;9n<d  `4 G  a0 I  b4 :;9I<l  c(   d.?:;9nI2<  e.?:;9nI<d  f.?:;9n2<�d  g4 :;9I<l  h <  i4 :;9nI?<  j4 nG  k.:;9I@�B  l.?:;9@�B  m.?:;9@�B  n. ?:;9I@�B  o.:;9Id@�B  p.:;9I2d@�B  q :;9I  r.G:;9d   s IJ  t%U  u$ >  v I  w:;  x   y;   z9:;  {9:;9  |4 :;9I<
l  }.?:;9nI<  ~:;9  .?:;9nI2<�d  � :;9I?<
l   � :;9I?<l   �:;9  �9:;9  �4 :;9I<l  �:;9  � :;9I  �.?n4<d  �.?:;9n<  �0 I  �9 :;9  �.?:;9nI<d  �&   �.?:;9n<�d  �>I:;9  �4 nG  �! I/  �:;9  �:;9  �.:;9@�B  �.?:;9@�B  �.?:;9nI@�B   %   :;9I  $ >  4 :;9I?<  $ >   I  7 I  & I  	   
.?:;9I@�B   :;9I   :;9I  4 :;9I  &   .?:;9I@�B   I  4 I4  I  ! I/  .?:;9I@�B   :;9I   :;9I  4 :;9I    .?:;9I@�B  4 :;9I  4 :;9I  .?:;9I@�B   %  $ >   :;9I  $ >  9:;9  .?:;9nI<   I  .?:;9nI<  	 I  
& I  .G@�B   :;9I  4 :;9I   :;9I  4 :;9I     &   .G@�B   %U   :;9I  & I  $ >  ;   9:;  :;9   :;9I?<l   	.?:;9nI<d  
 I4  / I  0 I  .?:;9nI<   I  4 nG   I  $ >  9:;9   :;9  4 :;9I<
l  9:;9  9  4 :;9I<l  : :;9  m>I:;9  (   (   .?:;9n<d  .?:;9n<�d  .?:;9nI<�d   :;9I8   .?:;9nI2<  !.?:;9nI2<  ".?:;9n2<d  #.?:;9n<d  $.?:;9n2<d  %.?:;9nI2<d  & :;9I82  '0 I  (:;9  ) :;9  * I8  +:;9  ,:;9  - <  ..?:;9nI<d  /.?:;9n2<�d  0.?:;9nI2<�d  1.?:;9nI2<d  2 :;9I?<
l   3 :;9I?<l   4 :;9I?<l   5.?:;9nI<d  6/ I  7:;9  8 :;9I8  9�:;9  :�:;9  ;.?:;9nI2<d  < :;9I�8  =��   > :;9I  ?�:;9  @0 I  A�:;9  B��  C/ I  D�:;9  E4 G  F I  G   H :;9I82  I.?:;9nI<d  J.?:;9n<d  K9 :;9  LI  M! I/  N! I/  O.Gd   P I4  Q.1nd@�B  R 1  S :;9I  T.1nd@�B  U.G@�B  V :;9I  W :;9I  X.Gd@�B  Y I4  ZB I  [��:;9  \��:;9  ] 1  ^�� :;9  _.G:9d@�B  ` :;9I  a4 I4  b.G:;9d@�B  c4 :;9I  d.?:;9nI@�B  e4 :;9I  f.?:;9nI@�B  g IJ   %U   :;9I  $ >  & I  $ >  9:;9   :;9  4 :;9I<l  	9:;9  
4 :;9I<l  :;9  :;9   :;9I  .?:;9n<d   I4  .?:;9n<d  .?:;9n2<d   I  .?:;9nI2<d   :;9I8  / I  9 :;9   <   I  ;   9:;  :;9   :;9I?<l   .?:;9nI<d  0 I  ��   / I  !4 :;9nI?<l   "4 nG  #4 G  $   % I  &B I  '4 nG  (9:;9  )4 :;9nI?<  *m>I:;9  +(   , :;9I8  -.?:;9nI<cd  ..?:;9nI<d  / :;9I82  0 :;9I?<l   1:;9  2 I8  3.?n4<d  4.?:;9nILM<d  5.?nL4<d  6 I84  7.?:;9nL<�d  8. ?:;9nI<  94 I?4<  :I  ;   < I  =4 G  >.Gd@�B  ? I4  @.Gd@�B  A :;9I  B :;9I  C4 I4  D4 :;9I  E4 :;9I  F  GU  HI  I! I/  J.G:;9d   K I4  L.1nd@�B  M 1  N.Gd   O.G@�B  P.G:;9d@�B  Q.G@�B  R.1nd@�B  S.GId@�B  T :;9I   %U  $ >   :;9I  ;   & I  $ >  9:;  :;9  	 :;9I?<l   
.?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I     9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  *.?:;9n<�d  +.?:;9nI<�d  , :;9I82  -.?:;9nI<d  ./ I  /0 I  0 <  1.?:;9nI<  2.?:;9n<  3.?:;9n<  44 G  5 I  6B I  74 nG  8.?:;9n<�d  94 :;9nI?<  :. ?:;9nI<  ;I  <! I/  =4 G  >.Gd@�B  ? I4  @ :;9I  A.G@�B  B.G@�B  C :;9I  D4 :;9I  E4 :;9I  F  G  H  I4 :;9I  J :;9I  K.Gd   L I4  M :;9I  N.1nd@�B  O 1  P I  Q.1nd@�B  R.G:;9d@�B  S.G:;9d@�B  T.G:;9d   U.?:;9nI@�B   %U  $ >   :;9I  ;   $ >  & I  9:;  :;9  	 :;9I?<l   
.?:;9nI<d   I4  / I  0 I  ��  / I  4 :;9nI?<l   4 nG   I     9:;9   :;9  4 :;9I<l  9:;9  4 :;9I<l  m>I:;9  (   (   :;9  :;9   :;9I  .?:;9n<d   .?:;9n<d  !.?:;9n2<d  " I  #.?:;9nI2<d  $ :;9I8  %.?n4<d  &.?n4<d  '9:;9  (.?:;9n<  ).?:;9n<  * <  +.?:;9n<�d  ,.?:;9nI<�d  - :;9I82  ..?:;9nI<d  // I  00 I  1.?:;9nI<  2.?:;9n<  3.?:;9n<  44 G  5 I  6B I  74 nG  8&   9.?:;9n<�d  :4 :;9nI?<  ;I  <! I/  =9  >:;9  ? :;9I<l   @.:;9<d  A: :;9  B4 G  C.Gd@�B  D I4  E :;9I  F.G@�B  G.G@�B  H :;9I  I4 :;9I  J4 :;9I  K  L  M  N4 :;9I  O :;9I  P.Gd   Q I4  R :;9I  S.1nd@�B  T 1  U I  V.1nd@�B  W.?:;9@�B  X.?:;9I@�B  Y. ?:;9@�B  Z.Gd@�B  [.G:;9d   \.?:;9nI@�B      �  �      /home/computerfido/.local/share/lemon/sysroot/usr/include/gfx /home/computerfido/.local/share/lemon/sysroot/usr/include/gfx/window /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/sysroot/usr/include/bits /home/computerfido/.local/share/lemon/sysroot/usr/include/lemon /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include/freetype/config /home/computerfido/.local/share/lemon/sysroot/usr/include/freetype  graphics.h   window.h   main.cpp    list.h   types.h   stdint.h   fb.h   stddef.h   surface.h   types.h   stdio.h   ipc.h   unistd.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h    G 	�@     
�ff!.  tt!.�  	:@     �*  	]@     � 	�'
�' t �	�K t��+��<tKxfftK� ot�>	�'
� t�K
�+�( t ���<tKK +mt%����'��= jt�>Zt<ZK
�H<
t&$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�.K�k�<60B�4�B �8R:�<(.*�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9%$/AtK/Z/��T���.��u	,(!>�X
K
(�
g(�-<=	��, t � / �kv>f��f���u,fftJg,fftJg�& J( t��& J( t�tf � ��"u%�* f�/f�, �9 fG �; �  .Y �f fM �t �� f� �� �h .���u�<f5 J; t& <K+f �7.Df9�J�trX�t<K'f�J='f�JZ'f�)J<='f�)J<">4<;tf6K�K- g.�� J	�w  �" t f�	u*ut �* f �8 �H fY �J �, .k �{ f_ �� �� f� �� �} .�!u�<f: J@ �( <�t���<K)f�J=)f�JZ)f�+J<=)f�+J<! >3 <: t f8 K � K0���t � t�tJ" X' t <Y$�)t/<�h$�(t�.L�K00tg\+tgZy.mh $X4 tg t f eClRfIfY<<4.t��*[� f�}���<J  	l@     ����  	�@     � 
�u  	�@     � �  	�@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K  	�@     �  	@     )�#���tY��Y����  	�@     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	t@     �	 � t J / �   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftinit.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftmodule.h   stdlib.h   fterrors.h     	�@     �o oX	JrX�
BzJZ	x<
XX �tXtXtY�<�
�m	 Z  t F�	fNL��	K	�	 Z  � F�	fN���	K	�	 Z  � F�	t\�JJ7 J\� R. J J3������<v
�Y	X�X=M�~J	[�
BzJZ	x<X���.yf��qJfJ<�[y'?[�/ utX B�   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  fthash.c   ftobjs.c   ftutil.c   ftcalc.c   ftcalc.h   ftrfork.c   fttrigon.c   ftadvanc.c   ftoutln.c   ftgloadr.c   ftstream.c   ftpsprop.c   ftsnames.c   stddef.h   stdio.h   setjmp.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   autohint.h   ftserv.h   ftincrem.h   fttrigon.h   fthash.h   ftstream.h   ftlist.h   ftoutln.h   ftvalid.h   ftrfork.h   tttables.h   tttypes.h   psaux.h   svprop.h   svsfnt.h   svpostnm.h   svgldict.h   svttcmap.h   svkern.h   svtteng.h   ftsnames.h   <built-in>    string.h   stdlib.h   ftfntfmt.h   fterrors.h     	`@     3=2Ju/<JJ<IJ��"=	=t0<	<=t(f=I0J	<=th0	<?�x��Kz^�<	XK�<Z
�M
K
	Y!fyJ<X� .�f�H>Y<1�YZ�xJJYXJ���x�f  �x.. 	�@     �LX	JL	vJZ
<	�=J%u.J
<�JKX?X	zf	u��$�u<�
�u<�
X�uJ<<�
v�� �.�jL��j�
JK
w	���j�
F�J��jL
w	��J��jL�
�j�K
1	�N�J��jL�
�j�K
1	��J��j�W
�j��<<� z 
 L+ W ]�  =?t.w;>r=7�Dt	�J	=	=2r<<f�>
�	ZJ	=	=2y<<f==a.�<?q=7�t�=.�=?t��
�>
V<	JJ	=	=2y<<f�>
�		XJ	=	=2r<<fYN8N= U.	
w.	Z;u<	=	t�&�&:	K<,tZ:fJ>= �~t=>X�ZZ&Y;=&�u=;==�%X�)tmttjJ�J�M�JY<%<<
�M�<t`v_Y)@_�yJCy C ...y.wJ)LlX"XX ....HJ8X�?Gi  ...+�H��Y�<�L<]�t�pJXJJN�~IY� <XJY�<�~JI[�J�<�~X��pX	<<�	J�>
Z	v	IKLJw<$�.�>
�[/���xVX	`Xt�+Y	<	�l�
X		f	K!M=F	?	L;	@�=uvKut!u	JX=KKLaX;;-.=KKL�t	�|L	�t�| 
�K
�J
wL
K	=
�M	��|L
	�<�| 
GML"	^<
�<
GM	��|	�.m	�|�J 	^<�J 	�.y^
vJWKJ>�[X�JZ  �XnX�{���JX(�5X!X�.myJZ:�,h<L^zJ=<Le<fJw'!M'9?!t=I=!h	'g�	=h:	>w9	?x<X<m<tW
Z�X J.<IY�zXz DHu�Y!tu!���X	<t�M����YZ�e�J��lX�y
t�xYt����J�y<	L�>YNKG>K �	=LYNY�>[K� Ju	=>K
	Y��}�<�vXu�X��}J3 =�'t=mg� �=>w	X X < Y X < . < X < . < � J = - < =>�	X=>w	X X < Y X < . < X < . < � = - K>��L<
<K
w	� J
.(>xn X < g X f <% � < K% - < =>�� #�|L�t.�|f�J�| �J�| 
�!
K;J�	L
��L
?
GM��|LL��|LL
	=�
��|<	K�J
�F
�J�|fIK
�	�|<
��J	�|<Z
�J�|<<	
�M��|LL
?
GM�	�|���	�| �J
�J�|<
�Jd@,	<
u 	J
C
wJR
yJQ����|tL��|�<
<K<
<K�L
M	��J�|X Jf�<i�|>�J�%iK.�<u�|�JL�v�|�J��=�|�J��Lu�|�<K�%fKZ�K�|�J<����|XJ�J��L�|�J'�f�|�J�<�L�|<<%iK.�<u�|�J�J<J<J<�L�|Jf%fKZ�xJ<�=�|�Jt��z [G1Bw
	Ȑ<��
�Z�
�Z�0
�Z[
yVNT^8LT
<
yR
zQJ��	�z�[G1Bw
	J�<XZ�>
>i
B
<O  .��=Kf=0 J < gym J �
��`!f � . />)=X<-=).)<<�>�	g	1 � < .
.v � "  = - K& ; K ; =  3  " < <" J J	 < �! t	 I Y L	   >�%<<�=%..�6J7O2<<ttY� X])	.A.)	.3�X	K;gx<
	KJ� � H� < . � . /�	J=	/	.#�M	+1.1f&M?+J?$fJ0.
tg<KLt<�< � J u  � < � < X J u  X < � < < X �  <3 <' J � yX � J t Y J t
�xX�uv,��G?<Y<<
@I�;Yf
AI�:Yf
BI�9Yf
CI�8Yf
D n�UwVv���v^�X %�?Y"
\t$J
\< $ .
 	�3@     S���.�~(X!�Ju!��~(=IK(KHAEK.(XJM0ABw%Gw%t��~0*<�t��['JFK)'H-L�� K/  < :]��~�W[�=Kt	 �  K<  Yf	 1# s J�IY�3�fJf� �luJ[=t�Bzef[=t��~ S��<*tJ<	Z�LKX foJ..o�.nKK=u��yQ@XX 	p6@     � W�~f�tM�~Y.�
	K�� �  �.��   .J8�t, X <W&��~�X�~�<<���n r�tKI=uGMtY1�t[
t^�}���  .	z 
�|<�t	� �~��usJt X��=JA	� ��KYYUKKYGKYYZ:3f�KGKKKM;$?=8KL<K<L �TuvuugggX <X��;� � JJ=_X��Z�!�ZW�
<	�IKI	K`
<	h	KOi.� �KJK�O	F�KI	Kt�KIKI	K� ��ZvX �.�"iK{ytK	ZJ	�J�	<nXfofMtY0��|�J�|J�f �| f ��f�o=NYt.kWt\�z�Xt��JY[J�3XY[�yt�~X�X�yJ[�~YX�
����Z�xX���x�f  �xff	� ��	� �f[vv
X"��!v`!��!KcX%u%8�%�%�& ��#�#���[	tL~]C x� R tZt�
-J	m��l	K�EZ
f�	N�m�fJX�k���z 4 �e Xe�X� ��u
�=�u��k	u�EZ
f�\�l�ftX�kt�
�r�.f�`J X..	u�s	�Yi Xd<�"�j���&X�NPzfZtCY���vJ3JLJH'�J;'=3;2=sK2fK( %JIu+K4I;JJY4;JJZ��jvY�%<%J<=X�L�j�%<M%+<?>�
JM�jt�%<%J<=��L�jYV�#8��,:K,-�,KL�jJ�<��j֐�MsJ�jf�%<K%-<=�<J
<MX 	�@@     �tLkctt� ����	��"�s	�<	=��? � &  �   ?
 	��i��%<%�<f<�	L��i���L�
X	K�	K	K�	4��itL<
<K
KfM
	K��J	��iLJ�1KL8cKIYZX<x.	��&t t.	=	=�	ua	�Ks	K	K7��iY�%<%t<�-�J	K�<yfK�<�i��%<<%J<=<�%<<%J<=��%<<%J<=����j�%<%�<f��Y 0 D�.�   Xi J[��Zt�z%XX��jJkX-.`[ X! t u /4 VwXJq	J4t�v�Z0,XD<<XH�
�'�	f�}NW���
M�`f$�V�� �zP
ZwJ
Lt]z<uYKZYq�)Yf�<..zP
L]�H�^]z<uY�YX���vu�Jtp�.<n<�.2
	��5�gtLJ
JK
1	�JJJ
$J<�K�gL
1	�J f�L�%Xg�fJ��K<<�N�L%Xg�fJ��K<<�N�KIKIKJ <.�J� .  J��� .Bf>XE�X�g�X��w�f���[[t u� X X u � < u J .   [BzJ�  .z.zxJ`  ..q ��`�[Q�	K[JLZ
<	Z	u.
<VJqXXd�
��X8< X <#[<K
Jt
J4 s .�5w �J X tT wt	<=
qX. l�."�� X �  XvK i	   J �Z$ f fq-.YLtJN��� � t  XvY	J.=
	Y�	�mtK
xJ.Yvf*��'$tm<�	��Z)/'�IJZ
<	��Z/-tIJwX4X'c�-n�?�a X��% Y�� uf � u J X  J	YFj � w�  t  <��t  wX X .  X��t���>
.ii� lf t l J X  <YE] ��G[  nXXt<w� �  t  < � X J .  ��et�[� tf J X  <	YA S  t  <��< v. t  X��v�t�� Xht y� C X y Q < y Q .  
 	YNF\ �f  �� Xit y� 5 X y Q < .   [!  ..-z.�[ ...9[
�W Xit v� 
� X v 
J < v 
J .   [/X ..JG[  ..�[C X <[t< v� 
  � < v 
J .   Z
�MKXJvJ
. v�
.� zX � <[t< � t   Z
�MYXvf�
J�z<[x	RK�
<�iXLZ
t
VJ
Xr X .�o X	z�	�3  .k.X�n�tX q<	 toJ&�JZ
<�@W	h@X tsJ.  s .�X Y9 sY�[f�J<Y
	Z		J�y m y.t . .	�T�zPJ<[
	Z		J�<X _ X.!<�TPt[
	ZJ�t. W�T�zPJ<[
	Z	J�E3 Jf  ��T�zPJ<[
	Z	J�zJ4 z Jf  ���[
= X�v.z�_u<�[	vZ
<	YKwZM
�M
`JsqX	fY�
� ��~[	vZM
�M
`JsqX .�  � �fz�	Xo���~�	vJsZM
���9 J
J�}t[	v
	YNX�JsZM
f�Xu(z�~XX�f.. �~J�.  ..�~ �.�@ X J[vJX�X��z��;tL�JY<$<J
�Q�<.<sJ.�zPZ5 X < K5�/���w	t
t	Y.h
	�	K	K,<	M�<ZtZY!wX	JXm%.f.t[X�%.n�Z(;K(<M	Z	�VJXYoXo.o<�=K�KIK�~X=�t��}K<X�NNJY[�\��#�E3 <..�~��d�zJ�XJ�f��_	��EZ
f� wJM
��`���^t�!�B	�JsZM
�<f�t��{fCI	�$	J<�~X��� 	�X@     � 	�X@      	Y@     [vF]=�ZKK?Y>Y>Y/n�-;��� ��.gx��uftl�X	@�!J	<ZY,= Y> �N
fJZ�J�J!o	<X�$�g�XJ�W��(I/. ���c� � f��(.�mZzP�
	Z	�Y.i�.if.� Y p5 [Y�5pf�,.�?@b/uJ=J=",�q	�V���c!F=Kh�
v�

��"Z:i"-HJ"vH>�Wg;=;Y<ZJYc=AzJ=V>=w
�
���
M0��<	RX	K	L<�kSAS�"u����~.oX=	<�#=0;=;KI=;=;Y	\	KJ"t=#��(Y^2yXCX2y<�Y2�2zX<Zu��X�KUK>�<Y�Z����q;<]��<OfJ@ �cK=I�>H�=I���RxXDxX�{yXCyX�uj�J<�<<W=8
 � �~ �X �~f < �J J �~ <L���
�=�~�YIY�TX� �~��X �eXog� tZ#K#K
i.�
�J+	�	M	 �  J x.X<��Y�� v� 
' � t�}�<�.�}�[=>�t�}����}J���y�}.���}����}<���������h<?�;Y�� �J\
�
����6 ��(�!J�yJ��JN�M!J�yJ<��JN�J��
X	M�!�eJ�ftKwXYN	v�Js�M
X	�e"&MU	��	�}XJ�4 Jh4f�[
< 0 .�
<	/mJ< m�	��XJXX��}J�X����J;W��9�7��
4 f$�
�4 XiJ	�	� �t�uf	�fvJ#O	[#}
J	j#	"	�	���~�J/�VIKV]KzPL<LxXR<J�I�f�X�y��Xv<�w�Xv<�� 	�e���	�|�t	�|�	v��*>=?K
F��LZ\zJZEK
J7K>HLX9�  	�5 y�	� 	uXG  �	
fAv?������ �	�}X� �5 f�z�w��tX	��.�&Xf��
t�X�<�</
�
�W�u/��<	f�:JyJZ�
N��`$X	f.�f�_J!.JJbJ�r,XW�)�֐....X 	 j@     ���v�sJ
t� XZX�</
M
OX .. r� <�I�  .-p�X	y<�� ff..�i���T{xRtY�	J>:/X<�kIY Y	�z��VjuX�rJX^J\9?9@ZI/  ff��v�o��f��Qy�h�}JY<	�I��}Yf	�I��}Yf	�h,�X rX�X�[<��&�	�[	VLX Z*  > =  ? K
  F^5��0� )�< \)Ju; 8	@)J	=Z<KIH��zX	J	K	?�=>KGK=wX,XJ(<XJJ+�K	<��t��q u"vLZJ<K
 J	J�	v
	YNX�JsZM
�	�c<�
J..a iiXn X�]wJGK5:�5���s�X�������w	.=v<	.KvJ	.=v<	.=v<	fY;Y�.��� tJ�Z
K
W�� .��	�[GL�<k�X[@x�f=)M��[$�t��mz'<>V'Jt<=I=IYYX>X		�X	:.�"�< � �	�f�W�	Z��MU_�zLX
f�L
�
<K
Yw	�	H"�`< J	�<?�\�=Twt"!y<A�zY Y	�Z�y<X	��M�yL
fK
K�L
M	�	���]�yL
�u
Iw Y	�	�J�.��&G�H. � � � f X J � < � � �9��zY Y	�9[Y� �z��XXX�� X�~t� 	ps@     � X4.�w�	twX	�wX	f.��

� =X # J	 zJ	X .	K-X	#X.P
=
K
 � L- M�
 v�9 
J
z�H'	J�-�� Y Y Y Y Y Y Y Zu�X� �
��t	J
	��oX.XK"� �Y�J
J�t
JtL
		�>�Z�S
	J%#J�	Vf ;C�"�		�%	!�A�A.�
Jf
JfLY0XoK0�hJ/uuuuuuv�Y���	�|JZ
�X���1$JuJh�
	[��}���JxJf�...�|JH tH fu�=K����� X JY/��JZ
fXMG1  
sJfoJX  �WN\]J#JW<Zt
.XJrJ.  
h�fG[  q[AK��J	X�Y<
<hJ.L
XX ..x�F\mt=ft�`XfJX 	�y@     5�JJ[�Y<<<
<Nu=w<f<<X#� = XvH</XRJ<<7u l��
zXq�.!��~��~J�X�~J<Y
	��F@	�x<>
	Z�Y�	� 3FZ'K	8u'KX 
�~���~tU4�J�	'K�~<.�'KJX Jmf^J
"X Y/ ;X%fK'=';K�� .�	�~���~t� ��YL!JM��X � �
t tX<0�~<�X�~J<<�t�� �I/g(�?�K0Jgt�L�K0Jg��L�K0Jg��KAK0Jg.J./K3K0Jg.KKl�Ha[JZ
�fuI/  �u��	X p�
	gt<x�hJJht
	Z��	^��	X z�uI/.	m�m
.f�|�wy{J�..<<
.�LP��(X.TK� � W�W�e�W@{cyJ%U>1yXN%.X%<1S@%;1%W.X%<1S2%;?%I<f%J:B��!
f
�%�JMd"�JM;#�F<0JM:#�-<M;�B>JK���
f�L-nJ�T�hX.K�W]�YYtEm.lCW�J�..
��f
� ~N
XJ
JL[9�<J�
�XL� =tX.
�X�� �J� X t.F<!
f:��J� X t.
�f�
��
�tx�hJJht
	Z��	^��	X z�uI/.	m�m
.f�x�hJJht
	Z��	^���	X z�uI/.	m m
.f�x�hJJht
	Z��	^J3�	X z�uI/.	m m
.f��j
<XXJLK%Xt<]t
�JN�zW�J�
��J
�~�
XJL[J�zt
�XJ�	�%pJ��
J�
	X�zJWJJ
Xf��yJ�X X
�z��	��<�+�	�<	L�}�yCu[<X�]�yCu[<X���x�hJJht
	Z��	^3�	X zJuI/.	m�m
.f��w�0:�t�JvL�<��X� Y�{v�~J�X�~J�J�����f..	R��	�
�
	Y/?<.2'K	I=�	<@J�J	� �	Ks�	�	Yx.	/-	Lx�/-J.	/x���W	=x�t�W	=xf	=W	L]�	�	�	K	i� �	/�	/�	=��k�R��X� -J=.��f��fJ�|�J><<XEJ0<<XSJ"<<Xa��X>X<YX<.<X%W<%J<=Z�>�	�zfy	J	VK	;Y<Y�Yn��#xn���<<Ye/Y�}J`.��t?�}XL��}`.�?tL��0<wg;KI5</5;=;=5J�}�.��t?�}XL<��}Z.�?tL<�
�K(=;=(LX���u`�
\�.sJ<s <wJ��;/Z�|J`.�?tL�M*./*I//o��oX��|t.�?tL<�K&<[G0<10<ihX.�}f	NK	:ZY��f1v��w�<<<Y;=Z�|J`.�?tL� XgV>K��|�.�?tL<�: X X�[=:���i�e�e��|.k�Z<=
mX�Z=� 
fwu�=��X
z�OS�
�JL=Lf  ��
v<O�/X</<Y
 ��X=Z!:!h>1HH[)g��� ..x��kJ.<...�~�w 	<wX	�<Y[K,vX JzJ^  T�w 	<wX	�<Z[K,vX JzJ^  ��y)_y<�qX)_Z
��
XJ
J�...yX�;=�=�
.y)_y<�qX)_Z
��
XJ
J�...yX׫=�=��#��
JrXJr
J�<JM	w�	<Lv�LX [J%X�X�z�v���
XX<�[L.M�~JL�KK���LM� .J
b.
PJ0 ��J�2
xJRK@* �IK JJEJ<fD..�� OJ1fL 4fuX���y�YXV�X/M�}X[���}X.��{Z�~J�M�~YX�	��	� �t��}JX�..�<x
XvX6><Z[�Z��{��Mf...oOX ...�vJ
X....J�x
XvX6><Y[�Z��{��Mf...oOX ...�vJ
X....�~�x	XwX6=<Y[�Z��|��Mf...oOX ...�vJ
X....���s�u�X�P�rZY�[3. t �lt  Z�~�X[�~�XJ�
	���	� J��kJXJg�XF�[wJZ8�uYy�_�n��Npu<K�}tY<<��g� .�� ��tu��pJLJ�<X
<J
JY�X Jh�Z�}
	w�u�KIK
L:L
���
<<[��[�K
Q�v
	�
JX .._�!X\�
�|�� 
�~
XJJ��K	��|�	�
�|�W=>���J���w	fKM
sX
JJ<s<
�X
J<�uTuJw/�
JJ�x-��# J	v�01IGX!H��OoOK��
J	YY�vY��	�vY��	�X ..ut�}X�f<X� 
Ji�tK� JLK�X?
JJfX
J
J	�K�v�t��tn��kJGvw
�<X
J<J�kY��JX ...7 cf4  7 J4 <J�kY��L
 �LJYXMLK�K�lX�
J�aX&XT<������Wof�X�8�< GZ=<<
�	MKW	ۭxUKX�5
tJN
z<K;K@	JKwLJ��XK
�*<.fXJ. ���.f�|K
JJ�?#u;K?
u;�	[�	K	�4�	��K�`�t�RB	vX�Js�M
�
,TJ,t�_�� �<K
f�|�_X� �K<Z
JE X�EI	Z&	J<�[��$���=��|Xt�`�� AZ=�/ 
xfw�/ u%<)Jx�)R�!X=�
_J
�&Z&VX
\J<�<>,JL:=s�#L4.�<<JJZ<:=J s JWf�
D)xU�X>
J�K�..7<�
>� A�Of
<JL.g(X"JK*(e<=I>JgJ(KH><Am<y<.L"XM]B(x<AOoMBtX <)JLtJ=�'.0X+JI=).>�X<.Lt<>
�
'J
J �= � K= I�
�+XE@=).<>�JL
��
�MMY�.(XuIK(KHA(GHK0ABw%Gw%t� ��XX�OJ1X X�	W��JJ	N�@$J� �;?WYfX/Jt<.Xi<<FtZ@
 ��(�~�tK(�~K�JZ�~(=IK(�MABw%Gw%�tzf(�~�<K(�~I��Z�~K(IK(JM�	�X(�~�tK(�~KJ�Z�~(A~IK(�M��#	fg#;x<=�/u.Ju�=sW=�t
�M0�� <>�*�  X �.oJ<X<r��aJ=v	wX��XL�����=X	LX	�J- r . X �`<�@G[XJXP$X<J�5E<%O7JZXY5%?qRZ�M��YZ�e��/X ...x�t��(   <���<X<X
<JL[HL
M	Z�	KO
+O(J,tNYLf....t\J$X����YZ�e
�f�d<<�� xJ	�e<#%�Ws�
X�p
t.pJJ
<p
J�
JJ
K;��	K�JX .J�e�
�;��YKL�[<����:�Y�==Xjt<Jkt 
JL>=L
<Q	��O
Zu�K�K-=h
t�Mr�<�
J	Z	�J+7J	XY�sJ	� �	� �t� �X 	��@     	0X 	Щ@     �j8\Y�~J��~X�..<<
.�L
� ~�
XJ
J"J�. �) � K) WL)��
 qX <Z
<� Jt
�~����� �	��rXsXJ;	�J	��~J�
�X��~XL�8	���X	<�<�~�
��J���XJ<��~JWJJ�
�XJ�	� � i  X t J �  g	 <Z�JJL�~W�J
���	8��~Y�	�
�~��
�	�	t�	� �3 + <3 X+ J	 W Y J	 I[Y�	=ZX�X&���;`XyXKX>&Jt^J.�J�.�@  �1<[U[�<uu�JrJX�pJ�..<
X�
�J�p���
�
X<���.]o<Oj�p�J�pJ�
��
�J�p ��
�
X<�q�� �pX��pt<�Kkeg39�pXu���
	��h�}J��}���o�Jf�rJ
�XL��X
X�
!�2X!X6;�XfJ�>�r�J�rJ
Xf��rXf��qY���
	�
�p���9�p���	�~
�rX���X
�
��8j0VZ
Z.����r�
�L��
X�

�J
<�
7�
	f\
	�XJ	�3$;	K3$J	Y3$t	Y3$t	Z	�J	�	ZH>	Y	g	g	g�
)�J��q�J�q<��K
J�X�>�q�J
�����q��X[�� �q��sf �f� �pX
���
�pX��X�
�r�	�<�� X�NJ� 9�pX��<�<���GYhZ/ ;K/~N bY/ tY/>/, JL�X�� �q��t�<X��J�Yh�t!.a<!.a<�e<�!JfJ�(M �  X J  X K ��<2 �+ J�
<	��K	M$,	L<�<� 
<��nX�tM�n�X���K
	� 	K	�X�
JL
�	Y�
	K"��J  "5 t t < s	�<Y	YJY	uJY	wZ//�K=���~��<
X:�X�nZ�~�JM�~���
	���	� �
ZXY��~�
�
]��U�K<L��� �KM�L�<! Y <( � <I �K<�RJ	�fZ�;�I�X�~��mXJZ
������XP�m.X��^F	<<�~�~��oJ�
��1c����p����'�>'����Jt��
t
<%JJLXX� 
<����	KX��n��~�JM�~YX�
	���	� ��	����oX��;j�	�X�X;���~X� ��~
s�=tf	f�[z.!5.f�`X
�"��6���Y
J�
P��pXZ�~�JM�~��t�J�	�fJ	� �
�!�TJh�rpCy.��
�rX���X��b�w%nfu%�%�%�#�#�v#RgX�6�|f�;� ��E�X�
J	Y�ot	��G�X�5�	��~�XX���~X�~X� ��nX��~�JM�~YX�
	���	� J��w [xJc[8u�Yy�_� <O�.
i.X\c<
X��<J��t��tX=K������YZe�XXhKJ�J  ...zt�sJ�X<<��t��X ...�Y<�u��J....Y��u�
� X� �xn<
�<<.`Y<L�s
�JX�tJ��
XJL�� �&	�rJ�
���	�J<�If	Kt:&
��
�tL�sJWJJ�
����sJJ
��J�e<thX.f<X<w�	�
t"h�<�
<�s�JWJJ�
��J�(��AWKA;(�%��
	�	K	K	K��
�st
��
��	�	K	K	K�.*&��X<%xJ�
�%<%X<��s�J�sJ�
��L
���
<��s� �st.�K43J.
�s�t��sY����	��~fS�b\9[7u�Yxf`��� 	p�@     �n/� �h
t3L.	�.3J	@�& X	�	u	�	�KK:	K.gtuw�XJJ zJ Q sJ   Z
��Lp+JT�(�XUEI
fo�� Y��!-�!�fo�/� �h
�
W1
X �D e�	�9J	O.�& X	�	=	Zk�uw�XJJ BJ ?J �J   Z
�XL(sJ�p�XEI�)Y�S!-�!�
I�f'Y�'� �wJ	<`<r��iJ=vT��XL	�d�Y���� �.Z<<=
X � <YK� .
��wfc�� �tX>% W < YM�  -X 	��@     f<� f <LJJ=^
>�wfB
,>g.[	=Z
�
iEc. `���>sK[>=S����=UPLY@;uK=<z���y��sX&F\^	�_t� �_t�EZ
f� Z��X]EZ�
QX �XJ(.  JI^J"X.r�HvLXb�(X�_���x	(>��MY
Q  .ti . .o�X
�� �   `  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftfntfmt.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h     	p�@     Yt � � �   |  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftlcdfil.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftlcdfil.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fterrors.h     	��@     �
K
K�� I�     �      /home/computerfido/Desktop/freetypetest2/freetype/src/truetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  ttdriver.c   ttgload.c   ttgxvar.c   ttinterp.c   ttobjs.c   ttpload.c   ftcalc.h   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   tttables.h   ftmm.h   tttypes.h   ttgxvar.h   ttinterp.h   ttobjs.h   sfnt.h   svmm.h   svmetric.h   svtteng.h   svttglyf.h   svprop.h   ttdriver.h   fterrors.h   ftmemory.h   string.h   <built-in>    ftlist.h   ftoutln.h   stdlib.h     	��@     �wu�xX	JfZ<;.b�<�; YO swX <p&JK�&7K&K�&GY[
M
OG�=�
	0	K<X�3�uWJ�"ggg�/��r���	fK4*�u�  u/  u+ u' r J u #  �nt t Z  , � v, H >   �  u  �4 0 X .4 t�.�}�5�	<tXb9	<t<tp�	<t�u.�	
<tft�	�tf\> � �Xt�	*tXtX<tX<tXz<Y	AtftX�X�0 � �^x6 � �Yw	. � �zX � �u � �u � �o � t ty�y5 � �Xt�tv�tn�/ � ��X#<<Oy	�K�<u��X�X��X
f�][J=# wt�>H�=�ftj�J=2 yt�
��<Ju6<J� <Z��<Xx��-/	&J	u� $Jt�<i6<fJJ�LIsuud�.�<�	\J"<"o.Jo<	u� t�<g$w� <�<�	d�"�	u;��x&��=<IKKw��J1��w&��=<IKKw��J1�A�A��
�!��)J=K)J@IB=�
���
���q���!f���Stz�z��g<
�	�	�]f(ty�	�	�����rt�ZtJh"tg
Q<
<]u	u�J	Z2'X<ti<
<Y4�Xm.*�=t+ t�
 J/ st
 J3 I�q�suX�
�p@
<���$��;-i;s?;qM�Y�=t�p@0<�J�
	�/�[��Z
	�t9w:s$�v���XX�~�
	��tv�~
�z�� ��]<Z<J	�"��]f<�(�p�<g
M�H.fX	iXL$rt	>
�	�t<> WX J
Z�H� Y
	� f��~�J�~t�XK X�t=JJ=-K� �<� f�t<� <
f$J<���K	d��	u-	�� K X.. k.�K �*�% �I � I  �QXWuwx.���!	t��v�t<�
	2=I	=1c	/>�tZg.	i�2.	=?G�L	=>Y��	Lzt	=AX[*
J XMJ
�.� .1z.B�<.<��
k?�}vZU�2 �# J���wJ
�K
<M	� �J��w
�K
w	�!�J��w��
�wtK
w	��J�-�/fP�vXf
XK!u:u!Z�v��� �k�K!ve�u!Xp�?<?tJ6�JrL?<�w���M�w
�K
1	�#�J�x� ==v	fqMi
	K� n�Zv�. ��zPJXZ���0�37+-�S.	-�+�+ �H �-�( �� JZ	

�^#
�_
`
	X:J8 Y> �XZ(��� J�X� X�...sJ
t�J� .J...� � X2.��^�]X ..t��<�]}yY�<X�f..��j�X
�
���[
�+ f	��X�X>f.% ^�		��< X+ ��.z
	yxt�
�XX�JJ���<-�L	J<�
�	>
X
Y;=
<LI/  Jkt
X�<t.�;��
	�u.KtJX.f.�	�yt�$�� J
Jut@P3�	��6U�
� �KX$ �. ��_!J
	Jwt>P3�$g�<� J�'/JJ.JK
t	Z�u?X .f	�J�3�i,
f	���Z
	Z�9Ks�+� t5�	\�M�21�M<<<
fK
K<w	�2�M
M	�2�M���2J�M<�2J?@<��	s� XA5t)	\�M�2?�M<<<<$�2<
�M<K
K<w	�2�M
M	�2�M��2	�M<��2�?@.X�	s$`� <t�MX�NF�<X���X���X�zf��vXX 	��@     �~g?Zt<X���������r�f�f �>rvZY�����X1p�wZ���X � ����X �t A[u ���FuZf	 � / d	 L   K ; �  �  �^��JZt	 u 1 e	 = �  �[��XX<.hw�zvr0X������H�
	Z� �  � �	 IZ��
J	Z��K;��K;�X�
J	Z��K;��K;�X�
J	Z+	I��K;�X����e� r� �c�
Cy.`sf_y<'yt'J<yXQJ�
�L@X .�y�=L�m�jJy�glz�g����usuIuI׹u�!j�g!i�!qh	r!�	t!�w�uyx��voyuztLv��FN���	KJ [G	WY0p���X lJg �q�Y]�M���p���X ��6x<�=
v<<Y�v$y�x����z*u*t��z*�*���
v.kz��z �|�fz]o�t}v�|�����|���� �|�g�f�|t�� �|th�f�|tg�fL�|httt�X .W��yu��y<u�����~�.�8�w�Y��JtZ	�3<JK%Iu%y�/KNX�#ttJ���fp.t  .M�p�"u%�zt*"�t*�z�u�"�z��t"�Xv�}�|u�������vr<�������f�
t J�&f;�
 � t
 i.�  .��%��%��{�
.u<�M
<XQ  .& yt# �M�Mv .�JX 	��@     �~zlKa�	Y��Nm<	�
�J�>//��.<
J	�nJn<JX<	/	Z� JZ=;�/K_�Q�d�)��	yJ;�X	/	[� JZ=;X/K]�
>
�K	;K
?<� �
.v.�K�Y�
�X<X
J<�/��v
�		J� � 2 ; K X <	 ��1
hX!J	m.J � 2 ; K X <	 �zJ K  <2 - K	 ��	��	;X]��	�tZ
t	Y0ttp�#�	Ytjf	JfZV	>	Z:!@Xw �  �=X��  .lJ�=XtfJX=..l ��uX�
�ut.�
JX
�u K
1	��
J/g� =�uX�
t�u 
.K
1	��
J�v�&UuuK&= ���YJ8M#t<��0YL�xJRZ��Y
�J�=
� 3* x JX�Y
Jf A�	MG����zJ�
f
�u"jqIY�t�
�!J
M-:
v!Uu!v
	/��S><L�
J�JJ=
�T
J�JJ=
z�XYtK�^�	�J	[	=K;<><!f)JJ<f�?
	J	LJ	[JJJ<J<��~#FY�XZf...�~�z<B�0 rt � �  � <. 	� � Y 
� �	�J	�	g<	� �  J	 ; XKX�XX� <V	
�J	�	=K;<L<!f)JJ<fZ?
	J	LJ	�JJJ<J<X	g,h��	�����zfy�
�vJouuwYt0Y��|/�t�}���~��X�����Y�8��Y�X JX���vtK�`�6f�fKqJ���}9:=��������~�
P
Y;�
X���~<���}:�<[�}84�
�
J<�J�}<�<[�}8
 7<; �
 K; I�J�}<�<[�}
4�;��J
�~<;;�Y;gE�U?&�A�<<
�b����� <���H.�;YX0
�.X		��
�"
X�JZV�X�
		�� J � �
 K!�	/�(Q�h�(�<�7J[�h(�fu�h
K
w	�4�JJ	 uJX����J/ �~X X J X�<X[q 
	������ �   �, -  =/   �	 J�� �  �, - =-  	 � �@��<[�}��	�X	�	Q�J	. �  �, - =,  	 �>>�(�	�#��#0r v  �h   
 f K 
  w	  �/ �J J+ 	 f ���	�XYVJXVZd>h8Z��ZS?
JvX<ZXM��[�i 
.v<�KX�KL�+�'X<\� 
Z <v
�M
fNut[	 Y  ; K X I X��Ft.oX�uv�qXK;gfK� JX<.D�
M�;=X�5��X<.PX,X._
J�
J�NjrY;K)
� �H ��	 �0  �. X0 � ;?  	 �0 . X0 J?  	 �  z JJ-bXJJ	�<	X�JJf �  � �	 I[��%�=u
zr<L
XJ	Jt�<�� ..
 �~�# ��h�
�XJ
 K1 �
 Y1 s�	J
�
X<��L�
JX
<- � tm
<�
�
XX
 �3 �
 K3 s�7JX� J��X
�
XJi ��
1X
<jLdLf	v�JX �% � K% W�%�	 �$  h J/ t J$ J J/ t$ 
< L! tJ$ 
X	 K$ 	 �  t �/uXX
�
XJi t�$>$rJL
��
�X
f g6 � Y6 sh6�Y6sk
	�

�
�X
JjL	�X�X<	i2 � < JJ�
 X
Jl+ . �L^GX �   J, wJ  	� J, w J	 J- A� J� X�X� Jf4w 	JJ4w<	 < �_�	Jw<�uuK	�B
<�
X	��XgIg�
	�~
<@�	K<y<K�� <KKL�f
�
J[-JJv��KySA)1
=-=
�	�@
<��Zt .�	�K
vJ	<�WK;	Kv�
<JJ	h�<�$XgIg$g��X=��	�KZIV��K=�	K;K=V	KK;	K�Jh�=$XJ�B;
Y; $%:tXFJ2%X5z�'=��{@�.�JYp�O0Y.�#	t.X
��2�=�<.�Ny�4�=�f"	./-w.#
Xv.�zJA"Y8#X\]FX:�?�!tX�=�
�MZXmJ=YgV=f0K@X .../��y�<2
 �L V �	 Z   �  � xX/�o�
XnLX�	��~!���	��y�- gt��tZ
	Y(./
	Y(J=
	Y(J=
	Y(J<wt
	Yg
	Yu
	Yw�n��t
Xt^x)uuhv uu�u�.�%eu JM$�JZ
- X	ht-�&?q	t-hd	v	/&	N*	K	�	L�Q<X�	�.	��um u�Q u��JZ<XJJz<Xtt�ZMULJJj<tXZ�JJ��<tttJZ<XJJz<Xtt�JZ<XJJz<Xtt��ZJ?<��=���ZF=.;M<JNX�=��	�< Xz� /B s6L:�@ImvklJu�
�	�v���
�	i!
	Y��
�	k!"
	Y<t< jX+����
m.�3�tt���uM8=t�<tY0t2I0[2e\%J	���
	��.,<,t<tfwu���X�<
	�� ��^<�f�� 	�t��uM0tp=�
J	��R�->�R<<<<
<K
K<w	�-�R
M	�-�R���-J�R<�-J>?.<��_<�� 	E�	��Rt
.K
1	��-J<�jtȬ.�ft.)<9=>)JJ/�
�(�t�	x(F�<�	\(<<	jf�gX��BJ<	uJZ>ZY@�	uJ�dJ+�X<Jbf
	v&	w	��g��g.
.Y
w	��J.<&tXx<=&Cv<=&	<f<f<�fujttp�K�z. � t, /1 : J
	f�.X
<X
�XbX������u�}�
 �/ � b�
 �/ W
�/�
�/I�
t.
 �? ��
pJN
X
tX
 �; �
 u; W
�;�_t
"�;W��;g�pM&�A�<<
�i<>� &  � I['� ��~�� �'� 1����;YX0
�.X		��
�#J
X�hJ>
		�.w�J7^r�<\f]!f7�!< �	� � �  =  � J	 G^	.�d�	�<Z".w[Z�dX��dJX�
�d<K
Kw	��J=�d
w	��J( uJ	 <��|@;"&�K/X"</X"�tJ	�;K6<LX	�:"Jg"J% w <	 JZ�K;K
Xk��6 ��$J�
	��� ��@ �~ X �� �����}Ȏ����}.��"��?		L�fX.qJ�h�ff.	��. g   �, -  =/   �	 < t��� �  �, - =-  	 � � � ��~
��~<%�t���~J9� �X/ ��$J��~	�X	t	Q�<	<J< u  �, - =,  	 � �6 ��  �}�~, !Xg!����=JG^�KJGX��4 �  	�6"�"X	 wJ �>�d
XK
w	�XJ��d
K
w	�>J�
X3��6 ��$</ n�$<6 �4 � ��~���~X	�XTH�d> X J L  � [  [  H > � J�o<�I9�Y
+�L-�Lv�K�ntYJZ@J<�Jw
���{.�st�JX0I�X� <[J��� X  �� ��	t��u
���yK#bjX<#JK#�#�#�!�!�!�!�
F@:�jiJX_
�	Y!:X�
	Y#<X�
�
�<�+L	&!LSJ-<!JKL	�<v�y!�<
�yJK
w	��Ju�y
JK
w	��J	q	X
fM�
�
��.��u
����|f%���K;�L�\	wJxJ-f�
t��w
M�u
���Yt�J8J<��|��T���Xu
%�y
4 �:�
	��sX
JK
1	��J	g�s
tK
1	��J	��s
tK
1	�\�J	��s
tK
w	��J	��s
tu
M	��J	��s
tK
w	��J�����  �|X8 s	�	���|��u
rX	/�k��Jj�	�	�
Jv�	�	�	�	�	�	�	�	�	�	�X	x	��"x���L�yvJw"��sf	K"u}	u	u	uY*	g�,�
;h
t�}��t#XktZ�}Z
�J
�&
O7X�
�	�	���z	��
	�	�ڐ���yX�~d	f9~�~�uVuuVuu��~J��M� �	�	�.�.-
K	�AS	�u�gI	�$q!^#tz�	z#	g�
��1t;�{J2Z#�Xusu,�{J;,N;F.�2f�,6w,Gtu.-uK<u�*uuu��/�";�M>��X�u
�}X�<	 � ( I J\�
X	
�
J5\58KIY5[tu
�w9[u
4 �	�(X(u 	j�F�kF�Cy�	�	�Xt< �9 % �9 Wh9%t�J	Zn�	<	v �! . }! O K!  �  Y  J	 xJ�"J	��	="J	K
9	Y"q	L�	="t	K	Y"q	L
	=
7�	="t	K	Y	L"Jt�	="t	K	w<	Y	L�z.	�	�	�Xt	�	�&hg. o J	 J	X�&V=NTI	K&=I	u	v&=I	u	u&X=Jxo	ug*	gg,	�X���X��X	r��
J	��rXJ
XK
w	��J	u�r
tK
w	��J	��r
tK
w	��J	��r
tK
w	��J	��r
tu
w	��J	��r
tu
w	��J�
	�[G	uz<	>	YJ	M[�~��{�X�J�{tX��tu	f;K
��!)X/;K
I=
>	=I=	J� ���	 CJ�M�uwE9XxJ[xyJ_HyX	Xv.K`w<uuYZZXx�MU?JZZVMZTsK]TsvWu�KwZ	��xK5
<5v<��7���t�
	�
<
X4�
J	�)	��x
JK
w	�N
FJ�	=�x
w	��J	>��p<tgJLJJX	�~	�.'/J 'XX�����X�X�~	��	�W	K��X�	�� X�^��X	�X	K	w	�. �@�yM��X,Jf,tK,�,�,�*�*X�*X�*X�K
X	�t	� 	" VZ	��x�X�xX.
K
J�
	K���	=�x�<X	�	�	�	��yX�w��O�t�{��|�o#.o.#.oJ�JK;*.J;J�t�.�5J>5bJJNy�		f%JJ$�1I�(<(<J(K��0<G�	 �z!�7�J.X�z�X?I7J�zX
JK
w�	�z��J1<E� ��JJJetZ</�X��%J�U*��@J?.�- o./n<.oJ<nJ�JKL<<H?IHKK=:K=>��@�<<z	<h<hJX	>%f	M[Y	<h<hJXJ <..Mt	Z%f	M�	Dr<rJ	Z%f	M[�J_�K�4�K<�4<�K<
.K
w	�4��Kf�4JX&�W�&;=WXX��n
����	�sgJY�Y�Z�=9L�&:�0�/'�/X4t"<4 �" .	�;K*<K�& ���
 ��
t	�{� X��sgY�#X	>:	>J�~�
-JXX���.�tJXv<h�~�-M<�tJ	X\$I�~<M
-J����K�~<[
-J�X���~X
�Jf��~��	�<I[	K"-=��J	��y�L�y
�<ht�0
	�X��
<ft<M<��
	LL	$7�	\.|t .	^f�"^J." X�
�sLqX<�FX	j�(dJJX>F[
��<
J	Yt(jJ�tjJX<!XJ%tI[
X:	Xh"X:2h.5t2�J�25tJ3�	J*V0JJfff	[�fXȞ58*wJ0J	J(�BWSCqz�^��>� t�tYuY�-��� X�<� <p<XXpJJZJ�.�.t�����
t�	mZwX>	^	zJZ9LM>%�	 �& 	 =% J 9^1�>�_���	 � 	 K
  qJ	ZG	?�xJ	|
qJXX<t�}t�f
t	N�	J
����@X
t�y 
.�v
�v��.��1�~xXJ\1�1x[yXQ�
t�	U	OlXt	_>lJOm�>xNLMXL.%M	 �& 	 =% J 9^1��>	 � 	 =  J G`�
X�
ti	�K	hf	��	K,�E	K�	K�	K	�
<	/,
J,<J	=,
J,<J	=
<	u
<	L�	ZJ" fiK	M	
I	KV�-�
.�
!�.
	�	vJ	��K	i�L.�$XJLGKv= � 3 I. J K I X�wutp�L�u�
��[
X.
tJ
��
Gw&
J
�Jj
<
�<:�
�:;
h:�
�:Wj�G�]G�x�
"�
�Jj
<
�J��*�;K<J�0�;=Y;YZVZ
.�9<3=G�!z�JtX�, �$ t�YIK=U�9�G[�k 	#<	��;	u	Z	= � * ; K X	 I\w	 �2 l�	 J8 lJ	 J �  :	 Z! iX � � X��
Xt
t	;�	�9	?Z ���tu)��X�x	���&K;KJ?0�
	Y<J!zJX�|trnt�L	�L�L%
��%
� �X ��KX5X	fJ�	�	"�% � . <Vz�<
X	�CNJ<	��	���	HX
	�	�J�JK�� � J �z<         �.<=JJIwtJ�tI[��J	JhJH.Z1<.�J .1tJ3�	<#VJJX�JLl..	g�r��rX<
<K
w	��J<t zJJL
�	Y�r�X��XJ <��z�5F(@IERX�����Z	%�	��X	K�JJ	�z��	��	��1�	J<���t
J� Je 	� �	K�X
"��
%�o��x�
c�
Jc�
X�J	��
�
Y��C8JX	�Y/WJ=e
�*W*g)J�#0L
_vfu
x�K
0y<
_Jy�
�<�
 �	�1 �t/..W/=IftJ[J�J�
J?�
W��{.X�<.vV3eȂ�x
�	�1 �t.-A=/��	�
)�
t�K���<J.i	.�+�Y / ;=6-;J9H?K	Q,v<.�<X�Xwtp��LxJ��dֺ<
J	h	KX E�	.
t�?	��	�JhKXEX�
�JMt���KMK3�KX<.Z�	�K	�JZ=/S*JJ��tt
JJ
fJ
Jh<�d.� t� fx`t�MM xJ% R JZ'y.u':JZt�
JX x��6/I>C�vXm��[�M[
�Z.
X��z&t����K�	 <"  J J I 	X t J   t I[/�.xJ	 �  t Ib�
t��
�~fz&t����K�	 <,  J J I 	X t J   t I[/�.xJ	 �  t Ib�
t��
Bf$T/�YMK.X �q�=u�LZL�.<J� X�f��L�.<M^
�M
X�
 Y �) sNf�
J
 �+ �
 Y+ ;��ZX�
J�XN�X
t	Z!z<	P!	�!z<	P!xMXX�
J�~�t���~�J
�~<u<Z
Xf� J� 
�~�*�
K*;
L*�
K*sN�
|�
�M
%z�/,V<Y3;
<*w<=-.n�7
.	�XJ	�$xJ`<x�$x<J`.xX.0
	�J>:>8J
J	�&VJ*J<�J� 
���y5 x�! � t�L
�
�XJXM
UF.f\
	�#.!X�
�^JZ"=[GM=<��J� .X�	H�	Yo<	Yz�#X!X� X� 	`kA     vt 	pkA     ��.�{&YIKJ>fZ��=&I]
	Z,J!gJJX
	�h&���;��;�3F��FzX!0F�lFz.!X�Fx  f*fs�1��-�),)0���y�u.	�vuXJJY
��
X.�<1P+v���iu�tFm�XN�/� J�t�~J<�}JY
������~��z�"fdWW\�ft"J)+fX*'��
X	gY
X	uY
X	uY
c�"rXXnJiXt��	�<h�<�h����`x�KfKJX�� 
J�
t��
 J��}u�����~u��-��
t�~�J�w.� � � � � .�}�~�
 �U.
#f
]X��y��Xn ;KX-��,�)s=,<.;�� "�[=X"�`gX�� 
X�uu�n�J)<%�'Ig�
!X_f!J
�
�t_�&JZX&<
�<
J�&#fKz<	XWgsuJ6J�6�� X�~�����	:�{�
��
t	��uV��h
�ytX!AJL
-�

�X
�|�1	� .	��|..X	��	/	��X�}Y�uX1�
 ���
�t�t�Y�uX1�
 ��{����,WW��}
�yt�	�/ ��~��=?��
	��+zfJ�Jh
��	�{	
.	.'�q#BzX	?!J	>#	YT-
X�w!X<J<%	JX	^ZAKAWJuX	��� ��.'Hu.!��	�	K@� ���pXpXXX=XJ .oXZY]�Z<K
	YjJ*. 	�wA     �{gwX	 wX	J.�'JY�tZ<
	
J.

�`f.	v�%
<f.	`X(Xt�Jr	�K	:ZZKW�;K�>�J- ��<JuJv	=I=	JC	y<C^�i�r<�Xaf
	��cXtJX*/Xi ;<�r.���"[#*.V.
% ��zt4z��Z�<f�Z
�����#�V�D�!I	t�Z!�u���������U���X�!�*�|<f�t)Ji<.t)�
t�.
<�<�<Jf<N
f
J	�4<BJ"�<O
�%[J�	$�	K�J�ZL��
6���<;�L
�
J�t
t
��	�z�J	�2'fJ����eJ!��;L	t	�zJ��6$.J	J
�}��X��J	�zJ	�K f , �( �, < .	 �Z�J'!�# ����� �f, s#�,*�%#��U��s��[�wX�S�wX�X�X�/�
	��-su(JM%�J�  f�t�'1u*qJv'/1N'*K'�'L�J<Ȃ�5�.�~��~��l�
����	3tr.��J����4�Z����$�U�J�(�t
LUK-*
Py�-Qw -
J
�tJXJMc[G�L�L�zwX?q[g�BS�z<=z^�]X Z�>vX
Xv�
f
X�
XuJ<
�<ut3�X<�	�	uH�J�?	H��O��
�d�����d�!�IK��d�!�IK��e�]J
tK
w	�"�!J���eJ ���VJJ�)�VKKIKJ��)�V��)�V��(�c%</-KZZ�������X��dHK�q� pLJXX��dHK�q��pLJX�X��d
f���d
f�u;u���WM
�	��J�'�XM
����'�z��nJ�m.Z �u�	<�n<J��J���^t��<
Jv���Iu��#;L�|X�\� t	�suI<JK.J�
JX�#uU=#WIKKr�Yt�� �	x	���!�_
sK
f�!su�.JL	�I!�<X�t�!rCy<Jv/#u#�LHK,v�m<JJ��X� �vJ���>���
�e����rt3�.mt	6�j ��$L
	
�	60�<	<t���nL
�3�
����G�9?9y��������l,t�
=�=
X>	(� �� ��$L
� �
�(�	�IX�G�&�!�E��X���l���lJ��
%�-[-�$���	��G�
#���eJ���f����f����[J���$�iJ8��~�����iJD.��iJD���iJ8���`
sK
f�!su�.JL	�I!�<X�t��#rCy<Jv/%�KKIK,v�m<Ȃ��!
	�J
�{��<qf
��	�	K.�$�`!
vr��R�u�I[����n*J<t�1Js�)tW<)Xt>JJX>�<t<�Xut	J�,<JJ,<<�����k
%�	_�j �$I�L
	��f��a!
vr��xJRv�t��k�#K1W8<�.��;����U�� fJ�)�U�J�(�e��e��e��U�J�*�U�J�*�X�)��V��'�d���d���T
��tJ�*�T���,�X;9t��'�V��)�VX�*�XKGKKgJ�'�c����c����fKJ�J<v
S
A�.u��
�	�'%J���c����Z��%�dJ����VJ�)�VJ�t�)�V ��)�VJ��+��T��)�V��)�V��)�cJ����c��WJ�J�'�V��)�V�sX�)��VJ��+<��y���Z
��
��	�	uJX�%�V>����)�U6�><���)�U��+�^t�su<JLY&J
J�
JWJ\[
��N�sK!ZpK;KJY������eL
��
J	�t<J����XM����(�h
��K
L/0)D�;=����h
��t�	�	�o ��$L
		�<t<f��WJ��%�tK�*L��t:�H>)=;u)<fJ���WM��it
JK�
�itw	��Jf�(�dJ����w?U
uNE=	oJ
��H�	Y
	
�L$�<J	>
�	��>�=;JJ?9Kt>t���X;9�v��<XJX�2�eL�*M	�%<%u;KI=%=%t?9?�=
Cy<C
��?�m��uw��
>:>
�<h?�m����fL�)M	�<t
J	�&<JX��eL�	#(Jf(t<x����XM�֐�&�ZJf�
�����{'%J[J�	$�	K���y/
t�u�f.=�JI���w$?
��X�	CX�		<X�		< X�	C#���
#X	�D	

$�	�� f���gJ�+ ��h
��K
L/0)D�;=����gJ>
��5X#�K�#X��#X��5X#�K�$X��$���������^
>rZ
<�.I�	�f��KX�		�X�J	=vX	KX�
	��W��J�gX�&\���!���J�VX
	��	�5����lX
� �����{X�	�c�	���n<XxX��
������	L�	"	�t�s
%�����	��G�
#�&�}��J�
	��W��J�TX���8XaDXaDXa8X���R���&���f�o&<JJ��n.<Ȃ�	�	���
�X� 
�X	� 	��	�� ���� ��	�cXt<MX�x��	�!�L!�.!<>�JJ<����\X	J2K,<�X����t��<��q	J2K,J�X�X.Xi-X.X�	�2NX	�1���fX�X�p > �<�	V>\!J!J��-�.X��_
h���L���k�#K1W8<�.�[	� X
�4tpKw���[�$/�[.<�$<=�[..�$
�[<K
�$J
�[<<w�$�[
M�$	�[���$�=><<JX
�,�!��-t�X�t�!t;L�JX��X��#�dXsKc?�<JXJXX�f�X
�&X�X
n<
o�<
oXX�?��Y[X�t=I=X��s��[t
.K
1	��$J<X	<�;<�mX	��;<�m�p�ym�M
�X
J<��}K
d�
X
JtO���}<����u��X �}J���/��z	XoX$	twJ	X�z�].A" f�XLx.=KKL��X .Jl�Z���f�}�
f, �% f�L.Nu
�
<	J!� �	!�<� �.Y
	$��	<��	 ��� � �m    X
 t K 
  w	  �+ ��	 f�	 	Y 
�	KJ�
	�
��sut	�~��u��Dt	�
��u�v���X��XW����tX����XZq�X
.b�v
&d�& �&�h o�u~�
tn.x$�$�$�$�
X
�t
�M�
�Ms
�M�
�Ms
�M�
�Ms�x�W
M�X
�x�U��t�x<
w�<
�xXU
w9��x
�
�t
�6(
�6s��`J��Ki�CyX
�}t�tv�}�<2z�y1DJ�}�X1�uw�y<��}J�<�t�}K��
XXb�w$fsbt�$\<������������z*u*t��z*�*���z*�*��f��| m ytg ��iqhtt�@f��	��vXO/ts.	Y�xX
tK
w	�)��f�tvv	H!	�!	�!	�!�E	Xt�	Kt;[�%:iX�P�ZJ�	�
 � z z< ^ � �	 ! � � X �1���)uh'�	�~��!�~�� �	!�z<	����rX�zuu���X
t�h�X
�z6�
�6s
�6�
�6s
�6%
�6s��X�x��u��<
o.oX�t2 �
�2I
���|JttmyJ5�!��;u��;��9G��9G��%G��9G��9G��%G��
	�*	g*	f�	;J�g!��� ,�T$�K$N,u�k��kJ
JK
w	��Jv,��k��kJ
JK
1	��J� f�J.�{���
<	6�!��V��M����X/�
 	m�y�	!u	��
J	0��##"uf�y���z�w��t�XX�&'�Y&UL1�!xJK!K!PIl[9�t�tK
t�
W����KP
2��	u�[�	Mg(�7�.	Bf�		�!Xt�"�Z"T�"Y2�YX M
	��oX<<
K
Kw	
�w	H��	=�o�JBB#KKBHA�BKA;#<L��~�� �- I�- �X �- V�z.(� �{�.f�
��f	�=I	g�{./�9�.<���"u�z�	 ��-U	M*� �� XȬ�!<t	���(./).6w�(XY)X�j�k!t�X�X�k.h��'!c�!�'K'W�'L'e�'K'$�'�L$v%p��X#�o}	{J� J\	�tg(0<.	�*	g* �"v�l?K�� Y3 s�]K
�\ZfJ{ X H O  fr� � H O  f	o�?�Jg�X�X�"X �H   j  �      /home/computerfido/Desktop/freetypetest2/freetype/src/type1 /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  t1afm.c   t1driver.c   t1load.c   t1objs.c   t1gload.c   ftcalc.h   t1parse.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   t1objs.h   tttables.h   ftmm.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   fterrors.h   t1driver.h   t1parse.h   t1load.h   svmm.h   svgldict.h   svpostnm.h   svpsinfo.h   svprop.h   svkern.h   ftstream.h   ftmemory.h   string.h   <built-in>    ftoutln.h   stdlib.h     	@�A     � Y-J=t?>�@�u(�.&�k��+�XuZ"K0,>+=	 �  *  �	 Y + � <	 Y/ + � X X J xXnfX�<$K-$=J<<h �f"u
��	J>	> X < <Zi9?@#t>
  X <	Z:	u-	KXXX.yXz.ZxXX.�wf!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��|�kKv]t9�Z
	Z	g%���~J�K]u�s��"tR�z�JX.�
	�>!	s�#Z#r	�	�O8N8~v�<�% � Jv�I��YI�Z�LVZJ?)'�K)'�K)'�Jt  ....	@tp�0tf=<tw
�  ��Y_LJ
�	Y:J	t�QX�.sJ3ww<$�J�	.wJ	<�"c�"r.�u����h�v��
X J	gH E <
�Jh�...	Jw.	<nt��$JJt�	.�"q�"�u������	z<tzJZ�
	K~fX$.Yf	 �  t I[�~�lpu���
.J �IY <.J	Et( �D ��D��D%	�=	� 	� us	u 	v �=  �! s ==  u! s u= ! J	 p_f�Z!��=" ��X<f��XX<�
JM(�3�
�M�	 K@ 5 � �\�t.tX�yu<X�LVO	t X <
QuX�=��YJ��
LsJt=ZJJPX 2.  ) N � =  � ) �' ; u I J zJ
fW=r�I=Z�~�^uX X��LLV�
�D��oYJY�	�	Z�	g	KW	KL��	��t	
J�	yJ �  ( L � =  � ( �& J J	 y t&X�f3�"X="�Kg<�S�  XuX(w<vX�U[L���?UYJZX.K�Gw���ZgK;KM
t�
�
&�.�>t	 L  2  K! L t2 � M G	 =2  J	 L!  K W	 = ! J J < < t t!]X�f3���Kf�x��JX�rvX�dvXX 	��A     �.�w�z=AE=<X�	 �  t I\���X��X�	  	 � 	 �  � F`�$��	 Y  � �	 z   � X �  J z	X��a.���X��X�	�	�	����ArL<=	=	�
J<��
J � �H W	�#���~f�
	�u��LQu
\ct
�	Z���Xs� X�-u�u
J	�	K�J  ....u�J YK ;	L#�~���X J..y�J �N ;	�# �~f? '�?s	�<�<	 �  % ) A < �v<	�f	t�t	�	�<Z� u ;=M%<�J�	0�t<	�J! J JZ! �� Xu�	�X JJ	�~�IWhAx� �H>/ Xy�"��DL!;=K<��2�$@2�@$"�L�#-�3.�Jh�& X�&� �!�!���Ku./%��w"�KY� Y8 s
�i���dB!vt�4:��"y<"{y<"�y<	<wJ	<�"c<"t�fw�u"pJx<� o�������yX~���K��[>
kE=�
	�ʀ	�	�.	��i?A� IL&	
J	� X�"	��) .���}J
XK
1	�N"�Jh�}
XK
1	�"�J	jʰ YIK	J5 .w ���}
JK
w	�"�Jg�}
JK
w	�"�Jf	�+%X�G	K%X?L%EX	L��J� J��~JL��	� <~	wZ�	�%[Wd%Ld	L%�V	�� �)�2�Z8J<���� o�X�~.�fB.�Jy� 	t �}   5 �<
 �}J K 
  w	  � �J u �}   
 J K 
  w	  � �J q Qʀ�) ��}�z�	XwJytuZ<X���x��X��X��X��X��X��X��X��X��X��X��Y���X��X��X��X��X��Xp�Y
���X ��~�!fF&�z.&P. H X>
�	KF2  �I/  W/� z �yJP=yX7Kv><�d�;� � � . � ��'	� JYJE<
t�~<Z
J J � . � � � X�JX��~f J � f � �	�tK(	�J�f	ZuJ�f�$ J JE � �	�1W	=1�t���w$ J JE ��J$ � J	�	L;	=/J	�&.<	h"< Y)xffW>�J�=� g9 ��9��v��Z�<G-��v�t�J	XX�xy�wt�K� $�M��(�<�wXY-Xh7>
d>
:	3t	+tw.X�-XA.
	Z	u.3Z-W�!.Z-WYwXY-XsX
	Z	u.mX
	�	u.�w�z4z.=vXX
<JL
tlMX ..	x �JK��	.wX	�w<M��L��	��K�FuwXY
	Z�
� M  . � t Y  J `h
<	Yv%u
fe0XK����AO=zJY	tw<Z=�X.'<Ok �_�+tUtYtYt)XS�� fv=
�
J X �	�J	� J�u
<�
�
k	�	�7���	�.x�WJ.u�	<�t	K	� �&X J&<	[ uG e �G �  	`&� �2 ;��JJ�!KY��=;Yv�LX	nJtI�� �wUw<
>f�Y*��M
�"M
��K
�XXL
��M
�"
 �  �f.J�~�<	K	M
J��	�J ��	�X�K�J�}�$XJ$�<.L
M$<L
P$<.K
 ��G ;
���M
�"M
�X$M
�$M
�$M
�&M
��M
��
�|XDoK9[??93 f�JK�,J<+ Y <C .H IX
�L
fu��� t�<� XN�$X$�<.K

� <
J	.�	��J	�!KYst=;	Y	vd	LXJ
	_�[w<L 
J �C ��vv�>5t
��u
�v <
J gD �	Muy
t	Z�	;Y
�$
�	�J���ff.�~JKu
<6 f	Z��ff. XKff.	� ���	M�	K�}�L	u�Mu<Jh^ZV<t
f�MxIYytu]Eu\puX]�u"X n<'�rvY�KY�YY�YY�YY)�w)&�<[Jh(
Jt�(J
X �
X�s ��	
Jt< tf
J,=K^,yJ;NK>ID
w<(<��XX 	��A     �}�u��.		�J<) w <v*f�
i
JZ�	Y)u<<tI/J...	xtA"H�hJXJ�~�.hV.Lvt���u�U�
	/2tx�
	/1tx�
	/0txX
	!/t�.X+�<Y
�	!JxX+�zX+�zX+�zX+b�
	/2txX
	/2tnX
	�/A .AX �o�
	!2t�
	/1fn�
	!2t��
	/DtxX
	/Ct	[Xt�.X\�/		Z$*�<=���,X��� .�}�
	/#fp�
;  	�6t.t	YW<K���*r
	/,%fq�
	�(.�<	=".oX
	�/t.x�
	/#fx�
	/1f�xX z.
	!$t`�
	���u.�<�~�
	!$t��
	�/t�|X
	���u��
	!2to�
	!2tu�%
t	�/A .AX �#�
	!2tK�
	/1fr�
	/34�%
t	�/H .HX ��
	!2tu�%
t	�/A .AX ��%
t	�/B .BX ���
	!2tr�
	/1fo�%
t	�/A .AX �v�
	�2t4�%
t	��B .BX ������}�uTuTuXu]uTu�~�J=.t.<JZ� qu�Y�}J7..OE@!:L<	XJoZ<<"t�J=�>
`
	[JmX�	�}�KI	=	L��|J
�J
��	�#1�?JLJ$=1<><g#1�?JMJ$K1J>JIL#1�?JMJ$K1J>JIL#1�?JMJ%K3J@JIMj�"u"��
�"/J<<g"/�<JJK"/�<JJ��gv�t<<<\� �  � IL�X !  t I\I/  �lJX.�X�v�t<<<��� K  � X IZ�f /  t I\I/f..kJX.�}J!uwXXK3J� O�
�<JO%IL��,ZUKZ# /IQ zXI=K N pO9F;K=;M
[
J	K� q�X-%<tJN�.ktJ	K�J	K�N8\	 �  X X t � X I t��s.oX�N�<v�
X0�<<<s+[�<	0-	�kg<	��~
K	hJ<J�X
	v!	Y!XeJ�f!�Y�'X?<u�J�y�KK
X	�\J	�	�t�	�	N	^J	 � 3 n JX	 `  X J J N5JYMJ�y�<Y<	<	g�1J��t	8HJ�X�t<Y�P��t� �� Y   IM�fJ�~�= @tYMK.  ��J. 	�B     �{'�uJZ,�!<Y>Z. 2Xt ><[ c?ZY6J3 <.Y� �<�2Z?Ys�
	K'�XY�JbP<Y
	Y6	Jh%� ta�z�y<l�f"��HX>�
X�0�v0�Jr���>Ko�Z<Z�
 
J<� J�KX<f
 �� �) INs�qKrLMEK�.O
JL
J b: N ��	Qtb"tT	Ya("XG	�	=W	K 	J@
JJL;H;�Hv;KGv;JL0;��0;��8C�Ju8C�Jv
	�	Y7	u[c�:;	��~JsJ�YJ�J<�<YJ���<>�J�J�=<<��
�<
X�j	<w<�ztBYLJ>
r>
J�XZ�LXY;/��	[G�s.KxX��K�$�� ��~X�� JȻ� t��	�Ys	Kf��z
^z.
�XJX .jJ!P � �M�L�Z:�XNX .��yc.�ot�.�oX�.�wT5utV�X5wt�P�<<*�o�<�o��<w��n�J�n�0Av��������XK�
� ��Gf�N��~~�X�ȑȑȑȓ���p�����o��i��K��m� K
�
��JK��
��X�3�to�H��N�o���
�X
��6;��!��/�o�HYY/���L��oz����� f��=J	f	Kn�	uW\����!#H<Z�	֟	�pX	�YI[fggh.��:�u�Y7X<7<<�#�,:�,X.;#�9�
��Z
		f	�	�	�	�
�
J�;�Y%�"�%X�;�Y%�"�%X	�%J;	Y	�#[	�#<�	��=�K�K�L!/��Y/IY��K��L�p� �J eK\.�B5g&<K�t�	K	�J � X

t���v0{y�u�����wt��s��u��!��uB!�B�!<u/ft�*��Y�w<	�*Z�xX	�.	�.	�	��Y.� X �>K�6w�6�Y4�3E���X��oL
V����ngX�	
�Z:	��u�	�	K	�X
	�����X�o�2]27K���
����t�� X"�"�"J�
	�	[�Jt��t�o
�B��\	�<	�s�	�	KL�X��	�pJvXX	� XW*�	��~<s�Xq�vtXXVs<t�v�t�z<w���ffu�K
�oO
	/�
	�
�u�K
	�	u�L<���tJJ�


��
t	/�
	ZJ �2 ;�<upu�<KIK1rL1u<s1KwpK<Jw
#0<Fu*/9v
u<	4yu<�		[� �!�
	�	Kr�	M	Z	�9 J	Mc	�	�W�WY	Y�.<�t	�~�tYM	��Q�
PP�JKJ�JJ���~J�f < .	���� �W�WY��~J�f fJ�</�%J.��$P�zX�.� W�WYk�-�IY �Y   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/cff /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  cffcmap.c   cffdrivr.c   cffload.c   cffobjs.c   cffparse.c   ftcalc.h   cffgload.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   svpscmap.h   pshints.h   fthash.h   t1types.h   cfftypes.h   tttables.h   ftmm.h   tttypes.h   cffotypes.h   cffcmap.h   cffparse.h   fterrors.h   ftstream.h   sfnt.h   psaux.h   svcid.h   svpsinfo.h   svpostnm.h   svttcmap.h   svcfftl.h   cffdrivr.h   svmm.h   svmetric.h   svgldict.h   svprop.h   ftmemory.h   string.h   <built-in>    ftoutln.h     	�B     %zB���1�fM�12h�		�	K	Pt	J�xJ/4f=?suy�v1�X�X�=wt< 	� B     =wt< 	� B     �wu�xX	JfZ<;.��<��tw>Z
	�<.�	vz4Z
�
V4
^f
.	Yt	.J�&�t< 	�!B     t< 	�!B     t< 	�!B     t< 	�!B     t< 	�!B     t< 	 "B     t. 	"B     t< 	 "B     �z � .���J[1�C>.Rf#
X		�)EO}	=f	K[WKJ�L�=J>
J	>X�W
.K	�	K h+#;K+=#=��t< 	0#B     
wYK�v�!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��w�":A�X�u ���JZt	 � . e	 = �  �[�G�Zf	 g , e	 K �  �[��XX�z�gK�]t9�Z
	Z	g%���}�>�>*#tK Y  � IM*#tK �  � IM+$tK �  � IM1*tK �%  � IM��� � �*#tu �  � IM+$tu �  � IM�!����<W[
QUM
	/tZ�0X <��:Jx� %<XuJuO<%zJY�
 X <	YzJl z �iJ.  [�<gu(�ufrf�,�Y �
 X <	YF@ . 	 (B     �|v
Yv;t<	.DXq�
	L
	M]=e/;=
Z	��gJ
	L
	M�tp<�X <�~�X	<�� J-KJ�W)< �� ��� <�<LJ�=
	��ifZ!�!hZ�g�<KI�<�	2K��q�	LM	�=e/;	=	��kJ	�� J-KJC�zfq�	LM	�=e/;	=	\�$J.iJ	�f�
J	Kz�B��� ��� �f	BX#<�X��IYI=X
h
�
x�<
m
		�<	�.<T�=IYI=TX<XX=<1<	� �tX�	�	�	�<X<	oX'<=;	�X�k<w	�ut��X<�J�	�/�f�J�~
[
�(tJJht<L
	w<<`�+J��
 X J�<�X	`� `J f  `J. 	0-B     ��z<�z�fXD�H^
�X�P=I u" ' J1 I Ji=jr�
�X<
.X�� 	<wX9 .X9t X9v.GO.J<J7W
X�~��I�
Jv<Z% J �L�X�~J�
j<8Jw
�
u�W	X<=
JX�O+M�.�1J<=

�
J	>	g 3   �J t>
	Z	�� �Jt� <LHL�KWKK�.tXii	�	�%<J$ Y1 I \(  <( < J( K�X\-J	    �uJ   �
 < K 
  w	  � J . �	tZ�/�X.�
6��w h	<uX�I�vmX� JJ t A� � M
 X J
 X8 -KU8���JX<..hXl<NA�WX�1�	��*�LZ���L=IY	   f& < J J	Z-J	�	��*&qJJ*J�		f<X�
	Y=
	��t�X���	J�X�w<K
X�
t�$�X
JdX�
-K
A<9�u9I0d\~N9�u9I2�KL	�Y-(JJ/	e\�X��� <J^N\X)<f���J��<X>X	��;(JKf	����	I
��s(JK�	��}�=
_

X�f.v<	J
a.[X.f
p	Jm.	�
[#tJ <'.<
.W�	&J
Z.[+J5XJ.J�
["fJ&<J.����t\fyfmfv.t
.�{fu).tM. 	`6B     ��wZ
f
	Zt	[M
	Zt	[R
	Z	�V0.X�\$Xc<.����}��u� X �X"�a�t�<
JM ��L Z�L Z�L Z�L XL&�&�(�(�Jf�u� X �>Xx���t�X<
JM0�>[
	Z�>[IC�`!Xv�<{#�#t�H\�X!\#.= /ut�|�$xTu�Z,�!<Y>h. ��L<Z��Qy�uvuxt	 /�K�	 | J n	h7�	K_J.	��~t.�w%yX<wz�
	Zv	ft �	 � XHh..,�f��y
C<ht
�	�����Qy�uvuxtt	�/�K�	 | J n	h7�	K_J.	I/.J	Q�/�X �~J ?;� [�K	wuX
�X�gt��L
Mt�� J	h!t	LH�X	�z�&�w	�<�1O<	�'XJJ;J=t.��/� � < <�o=
	�.	K�.J Q S    >^ �
J	�j
X	Z<<	>J�'�tX<K3J7I	X	uJ|X<J.�J	�&9M9?�J	MJ	/J	� C � �   =  Z f*J � �3 iX7 e=�w	�J[��KM�JL
XZZW*t� jt.�Xf�X$� 	y �|�4zJvK:�yX�<\bLZ
X�>	tX9JX ..	T�	�'��X JB�
X�LwZ
��
<^=/X*>:%LFK5:>5:LX
J��
�
�JL
	[�J�X ..	vX�O�}���ZDJ<<3u�X z.(ttXX {xR�Z?HL8<9K<�w��tX�|� ��Kv �: s\
	Z���z�f�
�|�idֻJc�X�ZXXou	�
 � K4 x��� ���~t�X!�YWY.;$kf�.nJ<tJ�/-=-Kp<tp�frXg<�
	��"���
�X=
	��	�� Z
�
t	�"	�!�	Y�OsYOI;�Os��x�8�SY��\&_&yt�&�&�n
<	�*	w*Wd	K*�e	K*�	�*	K*�~�.t�t
<	K<>'�u�~�X�FMI�XZ
	����	u"V	v��t��xJ	D�(*��?u��(?��=K��=K��.K��=K��=K��.K�NK8Lh.g.-
ft�2)Z)VL �A/�t2+.�Z	�z�.VvG[8�	� '�p/sY�[�)�eK)K)J		1	� ��/t	TY't[v�
fj!�!�	'	LX	�#	� X	#�	it) .��Z�|J"�X
�|XK
1	�\"�Jh�|
JK
1	�"�J	jXX��\ K 	�5� ���|
JK
w	�"�Jg�|
JK
w	�"�Jf	�Z+^%zX�%G<	K%��:G	Lg:9�	� �7�F�$.".3�ty� 	J �|   5 �<
 �|J K 
  w	  � �J u �|   
 J K 
  w	  � �J q �2)�K)� �<g�J� �X) F�pt>�H�$.".�	�t�6D<$�v$���~�6�+�/-c..g. �#?�-�/-j�~�[\[
�v�
.r�?�
Xf�#�
4Gw�J
�	�- ZJ V		�	�� � )  � �    �	 q �� 2�r�<
fv<>RxJJ^t�zJhK
	J�.J	RJ- `XJ  X	�	�� � )  � �    �	 q!X��Oo�Y���X��X��X�X �x�z�	�w
 suY?w
	��
pKYtYJYt\	M�}��J�����x��xJ���z�t���sJq�r���X��s�����Z�|�t��q�����q�u��X��X��X��X��Xr�Z����	�u�
��	�uX��wYf�|�  fX�z�8@\xR�?
X'y
_�'�	ft�f	��Xr
�'�t.wK'Jx�
J�~<�X��~�����~X��~�����~X��~�����~X���
.�}�
9?
PJx KK/H=7;/9/C<9	J_�z�;eJJ���t XsJXLHKL5	�	��	?����<�}LO�tt	��	�	=		�\VZttXA :	 J��X�}��+��~�+;XJ	J0 ����x.�� �	� J�<�x���!K� <g��+	X0��X`K�X<<f�~J��,7|L��J"MJ=h�J�=!�J%K�%Y�$K.�}JmXSO�YIYZ<�K;g�<J�t�X+�� =�!=X� vJ
XJ�}t<�u-Xw�Kuv .=�t��<t�<�	wt��t���ug�
JV
Z �qX @ Q � m    ]
  . t� `
 \ yX K
  t< � Y   
  X
 J X�K[�
X
 K �D - �X�z�����q��t .. V�
 v J V h�q����qJ��^�/�#91Z���
Zg!,#�w�"K X t^wU5��h2 k<X <�"K^��v.� �sX �~�.vK'J%�wJ	J%<Ys�%[q�	X�		.�.G'[JfVX JJlJm<J[G?
T	n8�	u8)J<	v	K	LX�4zX0K'Jf.tfJtJ	J<Y
^��
^�.  .�j X � K w� 	� t
	��v
��O�
�g��xq?�EK3IK3M7Uw�
sY.t< �:vv�5	J7yoEKZHv�;JfJ<J	X;JXAXJ;XX;;K;�(t	JwfP�=t.�f/t.�f/t�/t�<iJf��|&X�.'J��|��.���TuyS]�
�O=u4\T=s4<�4<	#,F	g0&<�4c	J��|&X�}<4zX�K'Jx�
J<D�w�nHt�����	M��%�X/	KZ�t yJ	��J��
	�	�,J�t�YX�� #Qy<Y�������.� �..
J�.f*�+y�%�@f�!2<.<� jJ	�	K	[/�	�	hZ+J�!2<.<JX	a	�Z&.	�	�	�	�	�	�3X J..�~ �� %<.<Jy�%<.<J���F��F��F��JqXqXXX=XJ .uXZY]�HX=g -f 	`dB     �yKuf�	wO)ZY܂..P<+uXJY�
X'dJXJ..Yf<	Y&ZJ&�  .Z.. 	 eB     ��q.�J
�q�X�
 v�t7x�J<sf`yvt�
�q<<�Z}��p<=�Y
zXY
7Y
t.
�X
JX�Y[�<:�h<>��LL:{0::kX�:l<������v���<��t��\� \�of�xX�����p���<J.�<
� K <5 ;�J[N<�Jg�J�
�	�	u� �  . W ��
�t�
���~�.�~t�.�~<�<�=
�.<�t���	�	b.	�,<	u �  ! e ? ��s�u�wrX<MrX<Z�<X"�X"["[Z�vX
SX
X���u�

�<u
	��	u�J� Jfu
	��ydfT��f��{�
<�JW;� Jy�YX
�[��stu�yQKIy<_�Y9�ZZ
]w�Z=
z<KKKM
X
tti�
%���
��
f
tt�+v:�+)X\)8u/M/Uw
�t
�j
$t
t4�vHvi�
X	�J�ft/x.|�
 
tt�rf�Jt�rX�tYsuj([�vtK��Y� ���X1��
�t
ti
�su
k
t�u
�$2	��Je.	��JX		ts.�XX	�
�rX�<�r.
X
tt&f#�1u���
X�?
�(,<�	't�z�Z
.4�Z��q�
�	E�	v}J	�X���Zt�q{
�
J&Y*Xp�uWuv(��*	?�' zt w1 N'z�	t�<u���
	�. � �	tzt	u �	�	<I	�wt��.�xb. f( Xg���#;X	Y �	�	    �	 g  X �	�.	=����eg"t ���ZY�YY�YY�YY�YY�Y<�~
	�fv
]�KX<	���	�Ȃ�u
		��A!t	y@Ft@vXsJ	K5@r;JuJ	L5@f	�5!�w@}L0�?<y<	v?9	�F'K;.2vtF;	=;04zt0BJ1�xt	�1J	�	
<		�>O"M<�'&��{� �{Z�	�	��		<.	Pp28�T@\��f K0 ; J	6,JYJ K? ;L	>zt<P
	�,Jo	��J?�v�.�?�J> vt	 < J  	y��yX	�	�Zd	>9 .	�	�	��rW���!���X�
�Zt
�qyf{
��
�|�<����
�t�
�%X

X�
�
tt&f
Jt
tf
J@X
�
�t
thN$uNsiN�uNsiN�uNsn
		���u
	�,	J� �}�<Z:v�Y;u�Y;u�Y;u�Y;u�Y;uX	�~	�	�X�� ��!��X�~!���|��J�|�"��%IKwXJKKXf"" <Mg�|+�.K
�	��@	�XMf	+?/	\	[XhY�;Zs<
Xt	�5�A��{�"�X	"�dKX�!��X  j�/���z����{X��{J>��|$�;=$Z�>k	L+-;+u;�4<f<	t�r	
X"	\"2</+<h�\7+K	� X	��+�|J��
�	Q��	v� 	�~�	��Z�
�qy��
������vX�X�wtZt
�px
�v�Xy�
�t
tg�3Wu3sk?[c[
X0
J	h	�X�
vrL[qwj�J�!w�s��JM�stY�� �v	#	�t	�XX�t	j(/�� X�	��
�
�	s�y���y��	f��G���	��.�
�	Z�Zr	vf
t�x�tL�Z � tJ	t�(�
J � �	�y�"�	�� t�	zX�{�t�	z	�z�t��~"&[9[&<w
Xt
tg/��/��?' �y��<���tj��<2?�t�X�;1-�w;,X*w�8<<J%nJ$X�����
�	�X�ti	����<j��&<�0�ƞ�#>#dZ#vXttiL0vJ[9M+�w9*J%ut<<J�X	� �-u"lXX	�z	�t	�XX�t	j'��%[9[%Jw
Xt
tg.��
��
tjZ�����<2vd5X�<3&t&J<Z<\s/ <>I9J =In�X�<.XX<� �Y��XY�zt����
v
	�t� �sX�	X	ft	�XX�t	j�X���	�tttX2 < �XJI�[ 	� ��f�XX� �
X�
Xg�0��
��
X�X�<	0X�<,d<��X
��
tg�:��:�h:��
��
ti��X<	8M�w�	Mt�J�7O7LX��g)��)�h�)W��JHLHK r	��.xXXI��XX�|j�uX֞�<)XX
X�
ti�	"%.�	M%�[J	�<�.rfJ	X�	���J1	 Zf1�<.�f��<,jX<�     A  �      /home/computerfido/Desktop/freetypetest2/freetype/src/cid /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  cidload.c   cidobjs.c   cidriver.c   cidgload.c   ftcalc.h   cidparse.c   ftsystem.h   stddef.h   stdio.h   ftconfig.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   tttables.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   cidparse.h   cidload.h   cidobjs.h   fterrors.h   cidriver.h   svpostnm.h   svpsinfo.h   svcid.h   svprop.h   ftmemory.h   ftoutln.h   ftstream.h   string.h   stdlib.h   <built-in>      	p�B     �t  J#�zJP-#,�v-<+<u+w<W�~�!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��|�w Y��.%�fYt>Yt>Yf0^Y>�Y0��kKv]t9�Z
	Z	g%��ZJ=KRqu�KtZ#tO�<J�L
�3's�V�"JIK9^`t>
�	�<�
�0-tu/K��.yz�gA	.wXJv0:�A�y.A{y<uuk
<�
	�X�
 	��~t�<(.�<J-%  <��I��YI�Z�L��<<M)'�K)'�K)'�t	�	���<�5�Kt..J�~�<	�X�0��#ZX#V	�(JX	Q�9N�9dv*�<��~�	'6/I=�	YYI	=�:Xt5<�X�6Fx<6Tut
 t
Jh�D��#3Y#sK��."JIK9^?'�t�"JIK9^� =�JIK9� X��� �
t2 �
	�<W
X0�� <
�J�
(��� �
t	\	��7	� <�X?.�X.pf�K^#Jc��u	JdiJX,�$y.J,Cl<v
"v<�,	w<� 	<wJ	<�"1" ����{JT���Kv�L�[J>���	ʀ�	�-�@#�B�
O#zfL#L
	/!�
�' .	���}J
XK
1	�N �J	h�}
XK
1	� �JjX	��	KM3	#y��Jy� 	� �}   3 �<
 �}J K 
  w	  � �J u �}   
 J K 
  w	  � �J q	_�}
JK
w	� �J	g�}
JK
w	� �Jf�)#X�GK#X
�:GL
f�~�<J?�	~w	Z��	#Z	��#W�#�#J� ��� JXJ `� t	�J	� JX' B��}�y�
�tJqw]	h	�JZ�K;uX�J x������X��X��X��X��X���X��X��X����X��X�XXf��y8.H.�t  ��yvf�<<0
W[X<�
_
%m� JQ%YJ� <uZwSu\Kwx.uu	k�)�r	vY�	KY�	YY�	YY�	Y	Y+)�u7u�<=XX-�w�X ..kf
)M�	 # "  f t z
X��XX 	 �B     �'�uJZ,�!<Y>Z. 3X @<Z�Y4J3<W� �<�2Z=1N1p�xX=
	K(�XX�JbP<Y
	Y7	Jh&� t��ufvrJf�
�� J�����|X.0�X�zt�<t�~t�|�=�fY�~��z.J.0:�
[[
X�
�
y<<.�Y�����}�}�<��X�{���u�K
�~N
	/�"v�L
	�	u�L<���tJt
��
	/�
t	ZJ�2;=u p� �=KIK2rL2=f�2�=�Jv
�%9<F�0/9�$2p$@p�X�}YX7h�T�A	>%J	�c>	u�	�	Z~	Z	<X'w�	J�g�FeN%��!J
Y;g
X
�9�$��s<�2:YY2��u�
;Yu�YZXX�
J�JJ���XX�
��B
DfZ�DWM	 .X&����|� � �<oJY�w		Y�X�	y$�	JZu�GeO�$xR	x���<
�J�zXM
<
Xt�f�&
s	[�
�X
��
�~t���~�
��=�d#�\J$<<	w�<.
	�<<C�
�JD<�
�
�Z<�<	�<��|CI�%��	�J	�0XJ	(t]Y���� ��~A;����M��}JKJ�JJ����
�~w�$M�.���\��Mt	�}	f�t� �'�f� ��	M��X:�+J	�!�J�0Kh:L�-ttn]�&Jb=�Y:�zut�sX��}XJ���7>S�>�kw&�M.�X�
t�~��	X�	=
J	P��F	=<	l��X	��&�;=<t�� +yt"�t	�
<wq��w
t�f�
	�
t<L`L0.IfJW�a�
J�.�
	�t
t�
��|�'����l�fJ�X�|XX�	�
	KX J=z����{���#����{X	 ��#�	� t	uX�Wt�{tX�t�/L<34J.L<34<?:
��|

t
wv�K[
X
���-�	</g
z�

<vJ
J
t	L<	?	�#�<�
��J��.�K	��|f�JvJIK9^1�=eM�	J	�t�`.f
�	�>�Z
<�<
�g6��6;j
��<�!�	b3�JXJz
t
�t/�ffX�}�KXuSuXJ�X�{<t� &���}���5���t	� <tXY�	0�X���s��t��|�
� JJ�WYWK�<	z��X����� f �0   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/pfr /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  pfrcmap.c   pfrdrivr.c   pfrobjs.c   pfrload.c   pfrgload.c   ftcalc.h   pfrsbit.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   pfrtypes.h   pfrcmap.h   pfrobjs.h   fterrors.h   ftstream.h   svpfr.h   pfrdrivr.h   pfrload.h   ftoutln.h   ftmemory.h   <built-in>      	 �B     >%gs=O	Z<	� f H Xq�y`��u&?@Z/I#<.u
Ji
v�#X.u
Ji
z..zX/t 	2F
4	KJ�4zJO;4	L=I'<<	uJ	f	pt'X.	gJ	fp.:X
>	ZL2=Jt=X yPKs.<=<�/=` =Htv]M>Z
	�)J	�.��y�u�K>f�?'qX� .��ff6up<J<2	�" XV<�fo;/'Jf.q.��zJ<
X �A �	�	K"TW	K'G@='E@F	K	g.0J><X�JNM0.��.J2MsJZ/.>�[t<		.tY.J	2LJY�@'J�tXJ�t.<%Xt.
��T�.fJ�>=<JL>X<�
�tXX<JM-#IK-�J =  f I�~ RxJ�=���Kc? �J��vKv=v=vJ�*�. JJX  � � : @  v  � � � < @  � � � . @  �( kJ J J � : l<�>J W � =:2 � J H @  v  � � � < @  � t � < @  �( jJ J H l<�
�.JpY�.M�9M�
�O�~#�~��~�wq?<X	w����Xq����Xn.Lr�~<�J?�~"u�X���
zzX�
?T�
<�J��JK'�9KJ= 'K)sB)z<N��Y�]�
.	�I<=>:�>	Z<<�JL:<.>X"su"="u(!Jff..zt�IY...��6t�J	f�<	h=L<.<�~��S�.�
wfX*z<B
<<X�N��X<��
P7�Y<X� � <�
t��
< W	J�<
JM�=�KX ..�`J.Kf..hJ�{tXX 	пB     A�@wY#f0Y"f0Z)J1f<)�Jc?1<�YLYL . ...n�WZ.�ZsX -<KY (JJjL(J=sJ=?
�	,J2�L=tt	�KI	Y�M=����O[*ffL
J]
JXt 	zXOt 	u<\FN
� .VwX�pJM/�tXrf��<��z
�zJ
4z<�
^X<� J .
 �� �0 ;NKJLt X� ��{��M���K=<IKJ��)��SJ
*./	X�<f<XD>,LkJ�>
	Z�<?
	m�JfX��~J��M�~
#�� f)���|
�
n�	<JYtt��?M.@<TN0�|�LLJ�J<��<<�f<��#JJ<.�JX�
�X
���J�VLh�	��	=	@ <�	��	=	@=?
	�J�<�
	�� ��*�� JX���?q1
	hJ�1<��
	Z�1��@�j�	�}�[
�r<���	� �J��J)�
���X	�	=,	L	[	�K�I	K<	1f, �� w�{J �� � �{   0 �<
 �{J K 
  w	  �= �J � �{   
 J K 
  w	  �= �J � X Je�	��� t��|XJ�)<LJh�~�>��J<��<<�f<.���~��<��~f�XZ	�	K>J:	>JX� XYfXN")X�XN.��X�yXYz^��� ���<K")X��<�.�	�X� <?Y	�� ��XWXoX�(Y;Y(�Y�o.�(�Y��XWX� X K�}J���}���X
X�}U[*�[�K�X�<�t����&J&<JK����&J&<JK	���<K�	���<<	=���<<	=��}M�?[�X
t��)����Kt �  = 0 G J �J6<XXX��|� ��}�M1b=1IJK=��X>L�9�}�X��}X!�
�<X�|=�X��X�|�2�MX�W�)Z��|X�Kh �_��0Ju��w���|tG[��Z���|J�tX<�|�tJ#=�
 X	��uo��K
	K�
	��"K"M��
	�!p	x � �~   5 �<
 �~J K 
  w	  � �J u �~   
 J K 
  w	  � �J	 q_�}<
<K
K<M	� �J	g�}
w	� �Jf��t�/)X/Y)W>HK)Z)H<K��� f� �su�J	2zJ	�gBWvZX.twX1X.%J?9?g=]<#t?q]J&X
X�D��}��X�}.%�<VJJ*X�}X�<%<VJ*X�}Ky.PK;K=-K=v!
�,J%��}J!H�L
	Xr<$t	<��$o<	<�9Y�@���X	+{�h=;/<>?
G	YJ�@
Z	/<f	�	�+.f�� ��X�	�|
fX�t����X��
�
Y,tsK
	u��%TN�p\t
��K;��2�}J
�L<��K=&<;KIKYt<�^�-� �t<�<K��	.;X.;XJAJ,<t�	'9h1C:U?F:3*;,O:8'F?s:A1KH?19'yJ2f1w<K
<1v<'yJ1m,KqX	�,HK,I*L,�	�*#M*q	M2	h�?��Y�=��~f$�f��|$*ug$>�>%<=%-<=�J�~J��.<�{<;nVX<	)	=	Y@cfJ.Zt<�
�
	K>
J
.<	0	=gHX	� .(�.JJ�~��K;/;<=	X��WY�=X=wX�KYX��YXY	X��I�;=�tYwX���KX�4X�J$<<�`���<.uyX�JX<X�X�<�SJXX�~JY	>x�X#X�	�<���|	�X�|@wfk=<mXy-DZ	.	/	K,dqf<L
X	KJL
	g>=
J
.<	0	/hIO�t��z<<��z.x<;
f*XR<	*�	=	Y:VfJ.Lt<L
J
[
<
.<	0	=hI	nX<j�[JJ=K=;K	jXX<f!.��~��xR{�t�ztM���<X��X��X��Xz��'�)�)�X���X����Xyt��	�	=�8^!��zJ!�<���zX�XXt	�0�.�~�JXJ�~X�t>�N3f�~3��!;j�~�,����~�
 J
�+�
�	<!�J(J9e�<9;��~�<���
��~��t
XJ
�+��X�
�J
�$�
�$��
KfX
qlX
J�%��KL����\*hv
	�Y	�g>
	�If�<�
	Z(L&J(eJ&�$:	jg#�?
	Z$>&��$/":k
J	0�}�><2�<�%f<J�	���g�
	Z� >J<�9�X�~X&�JX�x�J�}P���zJ
�f!:�z��t
z7hv�K
�J
�#��MLEv�$g$u$u$�$�$�$�$�"9ihJ�$J���h<d@*���Jm	Zt<<	hJ	��	K#�J	�I	K	��XtXL�� �t���uJ�xM�.eK.V:<�	Kt��J3 s	 <P�!�

f	YZO
iyf$
	K^&tK
�D
t8U o8zq �L2%kz<�.x=<7K=9uD,�D9/DI=0-/I�
�
	�&�:#rIvXo#vXvIfIsX&Xu&f&t.	�	�\
	�	^�	g	w�.�*�	J^&�	Zw��	�<	u �*  = +4 J L K2  ; K2  ; K  K 	 zJ`"�	X��J�f/�KrX��{XZX.X���+L+�>!�v�
��
t	�$�I���%��%�(8�'t\'F&sO)u>
	u>��=�>=t>J�
�X
t�
�t�DvX		<	L�J�:	@���. g<<J	�ZXW�/@zX	2�s��z�Z otX<>Z�ZX	�Vv>H'J	JX%fJ'.\<Y��MX�zXt�<�z���Xt��J	 �   !  �      /home/computerfido/Desktop/freetypetest2/freetype/src/type42 /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  t42drivr.c   t42objs.c   t42parse.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftdrv.h   t42drivr.h   t1tables.h   pshints.h   ftserv.h   fthash.h   ftglyph.h   ftrender.h   ftincrem.h   svpscmap.h   t1types.h   t42types.h   t42objs.h   fterrors.h   svgldict.h   svpostnm.h   svpsinfo.h   tttables.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   t42parse.h   ftmemory.h   ftsizes.h   ftstream.h   string.h   stdlib.h   ftlist.h   <built-in>      	��B     � u�.&�k��+��X,�t>=JZ�K(t*  ._.t>=JZ�K(t*  .� .tc�KxJq<J��XwXtzt.��x ��YW/LZt ��y�
XtJwtY[���X��X��X��X��X��X��X��X��X��X��X��X��X	w�	�X� ��X �� AJ�^<L/ zt^ �|.!f~	�w.&Pw� EZM
* X& �	Kk�.tI/f.;/�X�b<��J�><> �' t�g<�
JW�Xbf <�>[<4��<	Z	�	��	:	>K	" >�	L��
	�
�

� Z :>	& � J� X��~��
J	�J	=X�k�wf�b�&�Xt�&/X&�J#� JJ�<� ��/#Xt&�J#� JJ�<X�1!X&xJ%RK!x<�tm1EX!X<&0,K&!<fv��XJXt��1!X&_JJ%!XK!_<!!�:t ��X/ 
(2 ! J < � p�f./5 Y= e X�X?��fJ  ��- f  Jg<	���K	�9CX9<CfI<	�<l	#�X<	MY;	=	KXS� <�	��J	=��~X����{�LwtMw<	Jh^ZV<�
f
�ZxIzXuu\KouuX`XuX p���KY�YY�YY�YY)��XX 	 �B     �~J=.t.<JZ�  �  �fqKz<K><�
��
uIu
�
�7)<<).A<
J	Z(t
�"��<� t�"��<� t�"��<� t��� X/�����X
Mu
<�
�
J�\�
v=
\
J K# IYuv#�� �LVvn
�
��
��?
�Xt�
�t�
��
�t�
Mt�
Mt�
�~�$X�XK��~Ju
�u>w�t	Pu	�st<	Z<K<�u=	� X'�J	�	K.<	K<[	�	�� �&J	� uG e KG � � �	`v�	v>:	Z	K<	�.Z.r	h	�	�&t �&t	��L�J	�	K.<	/<J�z.ArL<=	=	�
J<��
J � �H W	�#���~��
	�utX@
�u
\bt
�	Z���Xs� X�-u�u
J �: '�:s	�<�<	 �    ) A < �v<	�f��	�<Z� u ;=M%<�J�	-�t<	�J! J JZ! �>�ufJ YK ;	L#	�~�	��X J..y�J YN ;	L#	��X J.	�~�	K�J  J..	�~fIWfr<CK
� �H>/ Xy�"��DL!;=K<��2">2�>" �L�!+�01H�k�' X�'��� �!�!���K/.�*=.t.� 8OJ�1;.�X\p@T�'JYf'JY<���"]J�!_t��������y�t^�x��1 JK1 JL'g�g��vK+fg+fh-fg-tv-usuwf....��y"'y<CJttYZ�� �|�w
<vt�XoJXoJXXUXvt�v���w��~�	.
�v�v�u�	=�v
�
Xt� ��ȑȑȑȓ�w���X/���xGu�K�pN/�yt	<w�QL�u
��<Q��tJ�<LJKJJT�f�}�� ��X�� T�0
mX����
�.��qf�~N��J�4
t	YN	wtuxX������
	�uV	����t�tq�(Ys�%vqKu%tu%tv.tu.zz�v�/�gZg[
	�	Kr�	�	�	�9 J	�c	�	�YH��	Y�< pXYH��t�JJ��
d�;�
*���zXPf
.�
��6I��!�~����/?�~��7��v�2�$�J	�	L;	�/t	�&.�	h"J'����
��JY?;	� �YtJ�f�y<�~��r��~N��YH��kX/H��f	�Y�	��t��v�Z#XJY�;e	JZ�#��	�=t�vL���f"�f`
.<.X)v<�[�9�Z9��~J<�X�~
��/� 5�J>X� �J� <�t>�kx"� w�v��h0��st�u��!��uB!�B�!<u/ft�*��Yw�	�*Z�xJ	�.	�.	�	��YJ��>Y�6w�6�Y4�.X� t�X�� �"��"�"�" &2O27A7���
��X��/X�x��tbX�uX/ �   #  �      /home/computerfido/Desktop/freetypetest2/freetype/src/winfonts /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  winfnt.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftwinfnt.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   winfnt.h   fterrors.h   svwinfnt.h   ftmemory.h   string.h   <built-in>      	�C     ��J=,EJ�B=2[>B19?UQK
	Z<2/kt-./�.�+w�~X'y.�=%vZ'0J*u0IK!5/�'3Jvt .X�=��
vXB ���@g!X�)vB/ f J <��Xw��L&�:nx�)w
frJ=973nw<�w = K K �3L[fjF�u+�Ku
# / f fC ; �J� X���f�J� ��t/B>)dv� � 
�k�	�%f	? � + ; K> ;5 t	 < X)J	X��x�.1w[x�|/t��d�X���XX 	�C     �~y<=J J %  , J L�q�
XXxX�.�o(J/�
JvX�z�x
�<<X0JX  Jt
 Q@ �O#JX|#J h nh��n
�
KO
E� 
�e �YJ'X  ��.t.Xt<�tf�|t�t�|J��Mu
�|.�?�|
<X����u��t
�
MEL�
�
	gZ
	�[
't
t�%MvJ	�xX\wX	K?9L?:O9G:	L�yJ	L	M	�,
vJ:
Jv<:
Jv<	
J	�	�	�	�	�h�	�X	xP1J
JR1916H�
t�����~v����t�~��t�
�{.C�s��fM�u	6��P
&�Fvu�Xv
	�	����|
�E�W�
� ���
<�
�
J���� �K�3SAoA<
Xt
t��&�
:�KH�
f	��	�{+w-Y`3w<.	<XJ�>�	�		��Z�'<<�X	m	�o</X	Zb����X	��	�|�K�	�
N"	%�	vfX4;uX	<�Xf�t\���X�}�"KXt�.tIZ	6y	�x<�	Z		�t	�	>	�	��	�J�H�	�*=�X*u ;=<	�*=XJ	x 8=<	�	hZ�JX� v�	��HW	���	Z"�$��;X	.���DW�X��7��9[XJ�J��$<&��=J.���FW�X��7����L��1J@,&;(��?<.���HWO��XKL�OX%�>��J<hXfXJ�� �����~X"M(K�K7F�(�?(vXK�JJ��S`xRvZ��uX X �   b  �      /home/computerfido/Desktop/freetypetest2/freetype/src/pcf /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  pcfdrivr.c   pcfutil.c   pcfread.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   ftbdf.h   pcf.h   pcfdrivr.h   fterrors.h   svbdf.h   svprop.h   ftmemory.h   string.h   ftgzip.h   ftlzw.h   <built-in>      	  C     � >usKLy���K	L.	u1ZJ=!�
^
t�J=!�
^
w.<zX.	uf 'J	=z 
	<	�J
�**		 yJK	**u	>ZJ=!�
^
t�J=!�
^
w.<XZ%JX%r *<= 'J@�DvX_<).I	et J'eJ	=` 
	<	�J�<t=t>�)�%���|�)�?<Z4�K5�K2Bt�t Bmz<=J J %  , J L�/q�
XXX<xJ` f;N.<Z4�K5�K2Bt�'I/  m�(J/�
JXcJX �=�V�v.�v0TKZWMvqw9yXC>:v7h�07<><�s�.4<�2HNz<;j79|"H-C:D="LL7==zt">RsuJu>"ytK"HL\tj-th:L��
�
 �2 �
��2t.[	
��|t�J�=+zJP=G>K=<u��� .��f� �I 7X ...A<07<><��07<><�� �� � Xtj<�{t?&O/..6.f<//.<6<f<//.<6<>0<w�	��{t�<�=+zJP=<y�X.���PI)
P�
t  e JTXu	k�%JJ^	�X~	
�KW	=J	>Jd.Xu��XX 	@'C     �{	w	�v�X��Xq�]<tJ	�	�Z�e�/�����s�X��������Xq��XX�Y�XXP<+���xJD�
�JH
X/<.	y�<M [..;/�� @p@f<X=dXZ
	�	gJ2 	l�	 ?*	g �}���<�X XdXXX
XM3EXg3EXu3EXu3EXu3EXu qfX�tz4z<�tt�P� JX �J
�M	�d<tyX0
	J
��;�u
��=�uZrJM�Zr�M�
���usu�kXr�M
�Zr�� �
�vt.�	Y�v
XtJ�Qf3�s�

t7;N�+s\Jk&-J��w
.���#tN#F<�
f� Js��K�u���y#uXP�
J
JX���!��
�
�J�4<�
X
X<[<f�JJ�A
yX	vC�#X�\y<�<��J�K��x�Y
�K
t �JX��K
�xX<��zzJuXP�
J
JX���t	�
�	����!
<	��
��
�v
<X
J���L�
�
&�XXA-	M#	u#	g#	u#	u#	v,jJX��j�{y#uXP��K��:Y�X\��	J�
�J�.X�	wXN!yJ�
e	wX��|�� ��
	��� X�G��K�v.Hv!��A>	>*�'J<*J<'J.tJZI<K�>dt�	M8�K;�rX
'cXXJ6�L
J$�5e�M
J$�5e�'w	<'wJ<XJ�<gJ���v��X�!
<	q�X<	yX�X� XXX
�}X
��
���[�X� <�+���
��
�X
X<��K�
��cvh?
7<�<	�	C XJ�		XJ�?
�C
 X
J�(X>
J	�f��v��
�	�[
�uJ..#�~i
J,X	_-�J!v�JX��J�K��|tu#YXP��K��8Z�Y;YY;KY;YY;YXt��L�x%
?%/
0%V0-
?0V;=-�
9
?.X
X���KO�X
	\h'<PzJJ'<=L*mJ	�;wX.�J�K��
�pN
	/h�~��sX�v�zX�YXg'J<=��13>1V3>�]�Xg'JGeMY��Xg
JH;
LH;L��tg
JH;
�H;�H�^�
	ZX	�&zXJf
�<Z�X�
�J
J�	>	[	�	\�<	L�@	
X<dJf
?J� 
J�g
 X	� �	�4we4rJL
XJ
t	�J	qft ��ti	�	g�J���		�_ ��			��J���	m	��� .^J�V�JM	�	Y�J�	
�� JvX
fK	��J			/ V= ���X�} �Y<H�� �K
(�}�XJ��XZ
�
JX�uv��H�Xt	�}XX� Y;YY;KY;YY;YX��|
�J	�	���!�}��
XJJ>�(��xXX�?�t"�f	?�X���w	Y	;=
X�Ȑ	�Z JKE.�֐	�u	�X��X� JK� $.�� �xX�XX!<Xth��X�	�x	�X�#��|L>�
�v<�v
JYL�&� ��		�	�
"�u�vY
�.
� .	�uu
	"f �- s�-s�K�f K> IL�*eN< KA ; f	x�	YQ�~��~XJ�X J	d�	Y	�.X	��	�
� ��~X��HZ 	�~ &�f	Y��
 �2   I  �      /home/computerfido/Desktop/freetypetest2/freetype/src/bdf /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  bdflib.c   bdfdrivr.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fthash.h   bdf.h   fterrors.h   ftbdf.h   svbdf.h   bdfdrivr.h   ftmemory.h   string.h   ftstream.h   stdlib.h   <built-in>      	`DC     � � = -�	=�
�X.Xv
	YJ+qMG�X�kJ.zf��q�JeJ/  � = -N	=�X.XZ
	g"+qM<9�X�kt.zf]�q�JeJ�W�j�z�=(usKM*K%���K	L.	u1ZJ=!�
`
r�J=!�
`
u.<X.	uf	�x 
<	�J
�-)		 yJK	-+w	>ZJ=!�
`
r�J=!�
`
u.<XZ%JX%r *<=.fv.Dx
.I	etnJIff^ 
<	iJ�<t=t>�~�,�<wZ6�K8�K-4Jvt 0�/=�9l�!t'fJ�!J�XJJLOag<gZ�tWuuw";9M
JtJ=j":v)?j"=:K"d7�:"9K"9K"cK9"<P6>�;��� .�t_�uj�t�u�u�{� f.\G�Z4fY
X�?J��
tMJ�vXX_�MT&f<X� J��
^zX
&pu
��
��Ov�LMxX ..�XX 	 KC     �}

��.�
	Y+9MJq[G.�z &��.�
	g+9M+<q[9.l^ Z�y<=J J %  , J Lx�t-q�
XXx �.�n(J/�
JvX��u�vfXq�Z������)�J��
J	g)q	MX��?9XXG��#r-JLX��X�m<XJ?rJLX��X�mx8X���t[,r6JLX��X���t9�[�t&.#�+JI��
e�
	/��w��X �oX�`xRv�t��o���X��Xs�X�������X J� �w
fI�Z<u����q. � J �  > V�O	AvX�	3J,.)<L
XgcJ	.0<4.pf��X<���	Y/J<N
�4tJ!�L
�
XA�L�
���!����	k�<LX��_X�J�I%<s	<�<��0IJ	JRX�	j�	��
4��MxF2Jnt_! _XY$��[�<���	w 	ftZ/#X</Ju/K/W/ �s��t-�:f�s��<Z"�XY 	`tI	g	K3 Y 	o�L		g!	=3 	e�L		g 	=3 �Y��yfytuz<�X]<
J���J�.��(t�=	�t�
�qg�tJL<=<K>:L�
�-
Qy�{
/	�.����	
t�|-X��"�
	�.���uI
JK<�t<�
�	�t
<�|-X��KnJN
of�K
�0
u
�<
J�%
�	�	���	K� JX ..���}
yfu�
X XJ�K
��	�� t��|t
2�u	L9JK�	
\�K
<���Odq�:LXK����� X	Y�	��
p�x�i
tr.��L
XJ�Jt
���q����q��#�
X<J��p�
�J��K\
�rt�XY�pJ��u
�r��v
�r�~<s���J�pX��r
s.Y�
�<t�]:@yX�y�Ku�	�	�	=
�		���YY��<��4�t�JL���
	g�4J+J
J	h�
J'�	�XX<.1<XZ / eK	�h!eK!	�&XheK	�'Xh#!/dK#!/#�K	J<1<XZ!j�
t	��Jt	�
2J �r��/��	�I!�/�])MFK4��JkT=
���
��pK����.X�:<X	�:<��	wtY�<	 �
"X�^�.�Jo�pt�.X�o���J�pK
��xJ| J�u������p
 X	����p
 � J	�����~�u0�����nX��t�nX��t�nX��t�nXy���n��n.f�
	ZX	�&zXJf
�<Z�X�
t�<	�	M	�	\�<	L�@	
fdJf
?J� 
J�: Lu:qJL
�	��)J��	*Jt�	7�.�p�	Z�.	�p�6Jt��	��	�p�*Jt��	�tX	�p^'Jt��	�tX	�q�J	w�� <^vd�t	i�X	�q�	MX	�Z XYX	b	K.	�	�	J'�z�6 � . u J	 ��+%>#H=�#��}<KY<H<t	��=&�>r>d>Z��}HI�<
�H;���?�A�� SI I)�g	��~GI'�g�Y1>1V>�<HI�<
�H;�u<GI'�Ge�Yt��	�q�"	�q��	�q�;�����[9M�1ztz��)M�Gt	
�� XvX
fY�<	�!���~���J�ktJZXJ�#eX$.����p+;J?X*.�	?�B�&f n���� �X�X5  �'�5I���J<s� t  �1 s �1s�K� KB �L.�N� KE �P%#x��%�Xf�xX
� XY� #�#�.�}t.XvJ[=.;=XZwJJ	�JIX�
J	Y�JwX�L=n .G�J[m�Z�yt���tt
pX
�pX
Jp<
�.  t��J�t
�{J��<��
�{��v*�JZ�
�
 �"
Y	KfY�/
 t� (	nJ-	Y-�	K-	=u	3�.	��,	Y,W	K,	=�		M
J���
�{�y�X�yJ����	I<M��~�/t�
���~f
t-Mqg��g?Xf��
�v:>Y��/	QXJ<�y<M	�Y;I�J:Y;I����y�?�~�1/t���?M@=
IKJ�	H<+��	�
�JTX�lX[�~�zfX�~<���~f�x�fxJ�Yx
XX<. ��(J	�L	Q�	/���~�J�f tr
t����
J�rL#txfu	�X.	K�f)u1J	I�M�L�
 ��
�Ȟ.K
�&t&J�uJ���
$rvHL
	�	��
 ��
�Ȟ.K
�0t�uJ�
.�uJX��
IY�u;X�<�
Z�Y�Z;?;+[ZZ�
 ��t��.K
���
�J�Ldv
��x�wJ�J'����wJ�z�J�z<��v�z��z<X�>	XL�������Z�~�KJ��
 ��
�Ȟ.K
�2t�tJ�.�tJX��IK�t-X��IK�t-X�
�M
	f�Z�
  ��

�*Y*�K�JL
� K+���L
��zXv��	�$����	
"	L	�iY�Q�
��1JK
�&JJ=�=�xX��		�g��K�.�wX	L	u_	uS	u	X���y�u
.iX
Xi<J
Nt.�w
 � � <J� ��fK
�$�{����"�tM
�	�$J	K
�
	�J	��
 ��
	�	� �f��|�L	K
��K�.��.�|�
 ��W�L��x�	�<	��<��	�|�
	KJ� �( ��
 ��
	�	�#�
� �����J
X	��Y�yX�.K���|��		�X
fX
JX � X�
	�	���|�Z��x��(I���x��k� �vrX���K
���
�X
�X
J�>
��}JZ��~
 "�
�
gsK
i'�x�X�<�Y�y�.���}��K
�(t�N
�
l
�
	ZJ�W��	J��
�-�-I<K=7�M		��dL��XK(:JL<	h=;	/.� l J/	}u;	/.	� ,<= I<f	/XB	 Y
 �3 eZ3I	w	��Y�
 ��
M
gsK
i'�x�X�<�Z
��� ���
 ��
MfK
�0t�xJ��<�IY�x��<�Y�IY=X[7=2SYb\�YL/LHLYWK��KZ
	�]
J��	�}�J	���� J3	wgW	K� Y
0�'�<	>.�
�� X
 ��
	�0 �'X,>6V<<fLK!	{Z
fX
Ji��x�.�	�}�� 	/�
	��X�	J	
f;(��	KK)J�T.	=&�L�vX�	nX	�X�}XXtk	� 	�X�~tBtXXtk"��	� X7)���x���	�<.�	��VZ2J����}��J" K�   Q  �      /home/computerfido/Desktop/freetypetest2/freetype/src/sfnt /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  sfdriver.c   sfobjs.c   ttcmap.c   ttkern.c   ttsbit.c   ttload.c   ttbdf.c   ttmtx.c   ttpost.c   stdio.h   stddef.h   setjmp.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   tttables.h   ftmm.h   tttypes.h   sfnt.h   sfdriver.h   fterrors.h   ftbdf.h   svbdf.h   ftvalid.h   svttcmap.h   ttcmap.h   svgldict.h   svpostnm.h   svsfnt.h   svmm.h   svpscmap.h   svmetric.h   ftbitmap.h   ftmemory.h   string.h   ftgzip.h   <built-in>    stdlib.h     	 �C     � ��u'5p0. �h�u uw�7 �x�u#5 ��.�f-[/.'.X/<<'t!./� � <��Xgh�
.�( v < JZ
 f	v	ifg(u.<J�.� W u w� t��~;=W
�2�}�K� �3# �& J3 <K�=�0K
Jq<�<=�M�%�h��1�
)Ku
<	3.	=tp<	�.	>^�"Xt	?[-t&zJBX=3Z	wJK�?>f<.A=Jf<.
A�zJ	�	Y<	�</vt+
..<Jf.�*=KK��
	Z	�<0�'
	�<Dt�� J>	uJJJ�
4X
�I��
�x	Jt9X<wof.jX	Jh��tJ�<0-.=-y�	<.f1+XM�%�h� �L.����HK�rXfr<$.o<.. 
�<V�0<Y�:��:��:��
.Y	i T# @  ��u	0.�. 
 v.	 K  6 wJ	 = tY	vf0' X0 < < .	Y	�y.�<z�	<<<��.t|� <�
XM��K
EL	OZ1$f.@dJ�<qJJ�<02.=L$K6$J K5��Z,LW�=Jz�N=��<4<b�;<?JL"K"m K�1 ^J�'.
.��r.�KqfqXX�hJuf.hh�fKtsYX..X�Z�gW��KX>
	L�
�ZV�HL%_y<%QV%>V	u.�� ���0JL X	<��=�
� r� � �� .w�X� � .�	DJ	iZ$1$919J?��KJh0<K��\;��X.l�.	p���\�� .�/ f��%..#�t.�K0tiut.��J�aX	Xt	�u<ZX/&<Y�;hHK�L
zX:X�.�
	Z	=�
�	�	�K	D��~>i�
.	2���~�<-�t
X.
X	Q	�X�	?��~�.�~X�sY+tUf	+�<YKIWh:LV	K�<	NJ�K�% � �Z	z�Yy	�.�	�~�t^�"XZJ>$< \�4�Y�:L�xJ4XYL�BYJ�;h:K�;>H=�XLJh��X4��,JY�=Hh�9Kh:K�uK;Y�t		�$X<[�~��.�t=<h0X<=���X<��0L0V<> f0�;�L;VL��~X[�>�	o�J��X)X�v��H\X �0tYu=Z:v�<>��<fx�H�HZ:>,/u:=J8<C=/pJ�;>H0:=ZHLJltt��~�t� �<Xc�<X/ � �%..�~Xz<�)�XJ���XvJt�����L,K�sg[�Y'�M�%�h� �KJ<�I>1f<+1@L	.Y�@�Y-u�PX�KtQ	gJZZJJ�
J4
y�J�
<4
�t<Xm."./hf.qf</] ..�M�%�h��Kft/	�
wJZ�Y/
tJ.4x .	.&1&+1XK
/��>vn�.�&<u��gY<>
	[4&.<4<&J<	[X0�=q
	[4&.f	[M.0<[X9.,/	s�b��p.9.,/�E 9./�M�<.Z� �KoM	0XL.Y�@�K
btO.)=[>[	gJ>ZJJ�
J1
�J�
<1
[w<X.=i�.ay<
<=s Z�M�<.Z� �L>dh� �J�u.HLs(JJt&<t��=./X>N
	[&t	[1�0�=q
	[	�Zf�=q
7 u� J J.�-K�	q�	l
w.	J.v.	K	L�
.v.!LKu�	<�nd	<�	�uJZJ/"fZ�>
zX:XU+.L
	Z	=\;KKh	�flJ�
iJ	f4<<&J	J�Lq<KKKh
	��<JK-KXY!�M�<.Z� �L>dh?�J�(JHLt�7  J JZ�.0hM	v
.X XhKKLPK�
.v.!LKu�	<�nd	<�	�uJZJ/"fZ�>
zX:XZ&.L
	Z	=\;KKh	�flJ�
iJ	fZLq<KKKh
	��<�K-KXY!�M�<.Z��L=�0�K� �g�V�>�	@<foZ J=#�YKMz
Bz� J/#tYgI=
zJ<X/s.B#<	YJZ
�	@cZJ=!JY#.1
�J/!<Y#f?
E<X/r 
Ah	KJ	�JX
f	@cZ!J=%�Y��
A�!J/%fY<<?
E<X/ttJA	KJ�u-/�JJY[�>R]�. pt
 2 .I �OX|�x.2qJ<j..*�Y-/!JJYW[�>Nw	X^J tJ
 CD � 4D z. 4D z. ^ sX
 2 . �I V J��=xD�t�f 	��C     ?t< 	��C     ?t< 	��C     ��Y?�b�1uxp
 zf?�J"�Xqct,<
[J%f�axX�<DJ>w
�KLc�<
t	Y-�Jk<���L[1���M1 � J v �"�:</	� J�<� � JJ��@Z%J=%f=J0]t�%J/%<.=J0]t.<X��!)<h�J�!.a<�J��� <  ��=J�zJPK����L
J[XY� JZ
,K	=tt,�[,K	=��KEKY j� .( �@ J	J(TJ �JJ"<)<t<�g&J<JJfK<��A<� 	yJ �0  J g 	 G(�	4<KA2<AJ5...* s < JU.� .�� � X] 7�tf	1� �, * J6 K ; /6  06 : . =  K 	 )(X	RJJK7(.7J&<7J3@>+z<<	@3f	hZ6=XJ* f < J f	Q9	1�`J	]3X3<.	Z�G� X	Q<� �t�Ks<EKnXK( �@ J	J(TJ �XJ<%J+<f<�	 _&!J<qX&;J.<q;!$JX3Wx<�efK	tf/!<l.!J3.J3-23TNtJn�
	����	`�:23FJ	>@�	 �  J K I	 /  > : .	 L  t	�
<	Z�Z<uJJ/w93<</W=<>( J X JJf� .`�.Xg;3./;Y�	� � XT�KXtt=;Jl<J.X� XX 	`�C     �wv
.v<
�vX
��=�\b�
�<�r"G>J���
J�KIKI=W/L
t�Zf<"./'.]� � � & � <�?G?
��WY�L
�hw
J2
 �( I\X�!f<<
�	Y/<tZB
	�J	L!f	<Lu<�g<� ? K 	 v J.<��<".� �ggx�� J$p@tY�� �~.C=��tJ>!�J\
	ZJX6
	Y>J<�Xz�huh.��#}k=�u�XIsXXJ;Ke�"1T=?
�t�?
^<.<twX� f�..JXJ<��
	�2	�./ YA �*[s*gWXA;�*	JOe�w.�yL� X�tvV� ��XY�1W
�1��!t�w =�gI== :L/
> JJ.I�.IxXJ"&;"KxsEuEu�	�zRxJ<�BX	>vX
X�ff��zh � �Yl�t* � X* � X, W�W�Y��Y�.	uXuX�XYJX .qJ�
	L6 tfE\  .w.��wfy�LurX�<f/MY;KXMt ..r urX��x.fqt#RyztutstXu;@LZ_<tB
	��	=J�/-Y\Z��
		X<Y	�JY �  �  �X<...	o�JY	�J�	[�I<	=J�	��tJ g*  �* W	�<YI/WJ	=J�o�	t�fJ g*  �* W�*�*Wf�JX�Jg��~�
	JwX
	 wX	QFK
<��LJL
�SJL
JM
<�v<X>X<nJ.  
t�M�
	XwX
	 wX(_FK
<(V	<L
�����>
��J��>
[
fwv<XL��nJ...
tf��g=�
J/�w<>dLtX<��M��udn�*�=IK^
dL
XMX�#��1 �	  	 /  I	 =  X tX
h�<mJ.JZ<
XXMX<Zy	�
<XM	YztJ �  � Y �hJ.u . .x���-2�JJZ�f=V0�J;
�w<	<�
=�J�� �~�~�=IK^� 
�
�t<
X�YHKz<[YKai9uW/-g/>	<X�K<J[K�<KI�/f	<X� ?  . �[���JW�=�~�� 
	K� �Jf� <��f� �J� .�	��f� �J<� ��-��� 4  .	 s � <M��W/f =  . e�y�Jv�\t
	]J	=X�!�K<<�~�
�y<�KK
JX�Xy�Q<J	<J wZtY1
 F 3 �H �	�t
�sJ�	fqX
��Jo�5Hǂ�t�<[� �KK
<XMYwtJ    �   tOhJ�u . .x��p�	.wX�LXfK+JXX�
M�;uZ:v[��eJX  .hX�
%
 �= ;�v v   � ; K   X L  X�u�l�u�	uv�		t=x.9;; �   / G< J�
" f	v&  X��K;��� X XX(K<�DL
��JMX$J=5��~.�.Kf.M�F�=�u!<(f
X
�h(K<����'X	'�G	w�<XJJ K? ���-�-K�?;�X	��z.��yt{
�	�uX	i��	0�	v� � - s = � 	 ���	-�	��	-��<�xpKZ%tJ?	 � # s	 K X �����Z(!�JM	 u # s	 K X �������f.���	J�u[
�	Y1
�	Y]�r<��s���s�����X���X-�ytw�yt���n�-�wY�������� w��X��X��  .�r<
	��v��J����Xs���u� @J�v�� ��Mu X JSP<X� .��":A�X�u �f�tt<
.JuX
Xv<�
�
��
XJ
 �0 �J%VL%<<��
	ZtNvJJ< rJ JXZ��.]�k7X0rY�X�w$�
�v��
JX
JX�
�J
 �0 JdL�A
X	NZ<J7 tJ JXL��JJ`t�/��gX�v<�m�ym[�|t��|tJ>X�X	�|fJ!zXJ\
X��� X <
X
t<v�>o�K
Xt:
<X 	��C     �}@t�K
e\D�	� �w�	-<s�	t�X< K �: ; �,� 	�~�6t�	Z,J	K,=J	L,V2>t	K2Jf		J	Z��	"��	J1"IQ_"t<6H/48p	�[�	MX	N�?�~�yf
m'<t�J�21=2I1=";K"�02�;K2V�"Ȭ	� �;	=	ZD	xJZ	�	YE	Z0�	LZtc	L+%t=.7t.��	M\�	O[�	MX	N��4"=4�"�K"��XX 	��C     �~w.u<�uX���U�g�
���X
	����X �~��f	4��	��;	=Y;	=	Z:	>Z		�,J		t		X�Y+1J	L<	�#��	uX	� vf�~�Y
	M�	r<Y
NY
	��	Xf	�r	�.</	�C � Zw	�	
�h.�JY1+�1J	� f� f��\Wut	�W���
LY
	KY
	KZ
��	�	r��	u��X����b b.<b< bXtgRX �sJ
|� 
X 	 �C     �{1.O<"KvX�K� JX<J��y�
	t�>
XJ
J/(tfY�X	X(�
"
 �> ��su�	�XfJ	2X	\1*t<	�" YH ;		t	
�b�J.�<t"<Mwz<w[��<
� �7 � K7 ��
" �F �	�tw		<*#tJ	��?3,t<�+ Y$ JJ ;x!%vf	Jf�) "�! X�"X= �K �j�.��i i.<i< iXtgJX u�\J
t� 
u X 	��C     �{]#.]X#X]X#�f/2Jt<��%t
�.M't�0'v���v0
�	J
	�%�
	�'lX'.N.�z�a$ \.��<0Uw/
J
�M��fm�u
Mt��/�w�.�J�mJJg�K<.t
>MxJJhJ�IKf<.
>	�-�~1�=J����YWYL�w<	t=
J[Ju�/.0
���f...frJX X.rtX� J	�	[L�	JZ�	M1�7�9	1	��w�s�.U<.M+.?��J<�?�* 	 J .KJ	�G	[3 � <9 f b@ 2F I	���JJ<.?}��? �* t	 J �f<	<=
J��gWY�=X>
� ��}�����}	<���~<8;y�J
J�
�>�����~��X�~J<WY#.�J	�	�v�Z<��2M12U?	�	K<�XX�X	W��	�\f
�
�fW.p�$Jvf;K3(;9=<?1<@0K<Y�e��<3>=�H=�=	 J	%<X�}X5K�XyX� t_�t	'�zlvJ
J;K.>=tvJ%�+;K+=g
JM�[��M	��{�K=gw.-;K3/3e=w.-;K3=3e=w.-;K3=3e=XX��t.0JDX��tXtK�<-t�J6f������ �ZK�z�zz�^z<=_
JJ$euKVY$K$�$�$�6&JK;K&D\���uusY>
^xXK � ��
#�*LJ ��� �7��J  � ��ZV'%Y�u6.v
.0 f t0 . �	�7(X	Y1(�	K(	�	X .�	Xh�YXJZ'�M Z VtvXP"t	J./t�t� XZ�X���O*�j.ufvs�;%<X�=(�E	Z<%�cX
 �<yk � t��-JO	<,�
��eJ@bJ=eJDxJt� ftY �          � e J          = � J          
< � t� J    .  	�. w� R   ' f�
	�<�
�
�Q=v=:>��x
7 X	��
	�M
	�M
	�O
	��u�
��utJ>!J�
	���!zJ�
	�t�
	u�uXJ�
J	��	*+%�*[�	K*$�*\�	K*	�*	�	 �+�	�9	#����*���?��?	�"�"	� f5�"x�	�H�#0H�#�	�	��|��J
	� .�
N 
	�J���
	�'f<�$J�
�t�#J#J�
	�<J�~X�
 �w  �� �wt        J > �!�J\
	�!z�JX<t!J\
	���	�w�!z�J�
 	!z�J\
��		�	#o�#�A �D ;�1=��X� �x
xXQ
	f�	��J	�%�zf�M�vX�	X�v��J�0
	L.<�<�	A�fJ	 tf�		v�u�� � � f�+ �= � J5�.5�t<5�<5J���w<*M�K<F#	X;X<wXtC8�Y+t,L;:;i,u$,Xf[[ g(,X(X,J� kJ�"�"#Hv#"I�#��yX�};  ��	��	�<Jt5XX��z<Y[Z; J��� 
 	�}<�
�<gXX � �	�}<�<��#o�#�	� �J��<����5��-�-,-0��X�|XX<tk�x�v
.vJ
 J� J(��
M<t
tXtwZJ�F@
1 X	K�r�.)�J�Jl�Xf�H=
<a=RyJ�x
�vX	� tt. <  .� X�r
f	h<	Y2 t% J <u	�JJ" _ J5�fJ...m ,X=aXX�ZJ�<0,.=gX�Xy�XJX�X<!����w	.wJ	 J� \F�8@<Z
J� J?�H>f[
���J[!ZW���=!?
�K
 YC ;	��)t�=IY�JZ#	�Y�
f ��6'tY.6'�	hJ<XZ<�#	j>9<?�* u6 .* � t? ;Z�.<	 �   �X = b �	>ZYJ�YY9M+=�;�	KuW	K��f�� $�<8 X��X]��* �5 .* J t= ;�<�C�fJ���<<t =�ZJ�<0..>YxȺtWXy�J�n�� ��= T� < J	��K��H>f[
	K�atX<8��<J�QBCW!s�/�Cs	w�XX�K
��	W� J<���JJ�i hE��dL7 X S( AN<O�J	Z	KJ<�=Y�XJo�w�X<�ty5yt#'J�%-tX71)7�SK1�7t � �e,� �t	J��=	���	�J�@F2: K> �Z�XL>�n4..4<<f,XX.xJ<v+19?4X,<XKJL�	� �%BJf�� �Je�tbX'  �.�<�04..4<<f,XXKy<�X��X.����JJ�$N,�8/<>6�J6;Z�XOXJ..��J	0	KJ<�=t�kX<��z�zJ�J�$k}0,0:L6��J<6IZ ς		�XY	�JL2F2: K> eLX��	 % i M 9	h��	=	=�XXJJ�Q�X<��z�zJ�J�$k}0,0:L6��J<6IZ ς		�XY	�JLX	 j% n M 9	h��	/	/Y�X�%q�J	[q9fJ�VfX<�tz4zJ#�zJ^�$[,�cY;Y6�J�6�Z 
Ȃ	"	�	"��M	��S	!�	X	[	#u	�	��Y JJ�-5�c>?GM � �^�t+t [  J( t Jh�iJ��Y�J(t
JZtf	JX�]EYJ�1C�9�UC19MCJ � ��� ��:L uJ J7 t �* r J��׹./u�XZ��<��� �*p�JXp�X��� tgX�z�te�Xz�tR��it�t\K
W[!.J&t<=&J=&J�uX�
�
.wj
	`�q�.ef	�Y	=K<<  ��3 f .fn Rx(Y
z.	hI	=<	.�.3 f .fn Rx(Y
z.	hI	=<	.�r.$8@p$TxgRX S
XK�X 	�zXw.tX	�w�=JlX
�"}X>w
X<N
�c�#ww��~

v�K
XXX	X� f��
�X
X��7s�-	��I� ]�	\	Y�Ih�vJX� 
XJ
X����~J�X�~<��w+�1e�	f�JJ�<7	��X_�	cX��	�J�4C4y<[<�X��
	w�K
X��3/J,J3T�
&J
K5�
u5s	.	�1	Mt	�1X<MZ����~�����X	���t��
�X
Xjft� ����X� �wX�fXX�%J<M! N	8XXX���tl�u�<.XLv
�
��I/  ..W<
�
t	Z5t<	Mw3t.i
	��-JI/  ..nt
�
t	�XQI/  ..	\ 	��#FJ:XJ	s�	��t[t�?X�<�}�z�J
Z��	�t���}
M
�	H y<yX.mf>��	�gJ[t�X��d 	��}	��[uetX.X<�}J��� �	�J�}f�X�h<�K
Z�Z
��JXX
 �~t> WJX���
�v
�M
J
 �2 I	�X�/	���+ n J��;=Y;KY;=\!
JZ-<(X	�	�J V`	'+<'J<J+<���~
Xp<
Jp<L
XJ�,l�<�k.=� ��.,�<�
X�!X
J]-X�	_	
 L
	Z		���2�	�	�e��	��<	]� n��� �� ��:<>�3��J�~X/� �fK_.<! _<!tgJX vJvJ
v� 
x X 	@D     t 	PD     ut 	`D     �5	�� .�X� X�X� �f//Jt<T�	v
�.M"Z"v�����v1
�M
	��	M�rJ� <r.�m.�}f'h

tttLK��wf��~�J� Xp�Y�?
��>
X<J���
J��}
,T�K�
��XxX�CW�JC��-J�CI��?gC�!��
�JB��z<�<���/�xu�[���t
M
t�� �X�C�{�!�
	f8IJ�u��	-19O%V<0NFJ����Y
	JvXK
	wXK
x<J
y<
Qx.=
��
� �<J
�3�
�3I�
X�
tJiXX��b<XXJJb��;KY;YY;YY;YXZ

J	Z��Z	������J/K
 � X�=
�u<�J�"0�T��&� U� �
.�#?� ���M�?U
ntt
�J��K�Mk�vM
�C J�)X
K�;X� ��
< K; ;L;;�
	�f�pNK��~�>.�f���q��<<J��|��
�J � J� 6� �@ � K@ ;��;!�	�!6X	
X6v�	
<6v.	Y	KfrJJ� �   1 I : L 	  <�3�Z3:<	Z	t	w�� 	� * wX	 J��NXJ�X��~<
��
$�
��.	�!'t!<'�%XI��J� K<�..��{.��CIYC;�C�YC;��CWuCIh�CW�C;�C�C;hCe�C-�Ce�CW��f�
7v"�J"X7�"L;7�xue,e>,;7:	z!e<!ftW�f� ���~X���}��\{[U(<J(YJLG�Zhw
J�$JAW(�Ae�$JA����`*KFM0=;=<kZ?
gAI(ZAeZA�-ZAf�� ������X�<X��|�Z
Y<�t�[#J>
	X<w��,.
	��f�
�
�<kbN����z<����������������
��0��X&X
�	��	[X	M	���	�	YGJ+HXX+JJ�  .Y!MH�qK�vX	I�����X�XJ�|�3E�J� hH�(f�<L	Yt�	Z	KKY�XJn��z.X<���&�~)t>���t<@��D;@
� 
��.-��;=Z:>Z�g6e�6s/6;�
��
��K-����w
X	h	�;	KYV�tY@<D����X��XX�X	�wz�^0)q)�
@t)8
NX.�sxX_Yu�YwoZqYvVZ2,t�/�
J�	Z%J#.Y%X#.Y#J\
&�F<JH�	��8�tg�wU?[��/
	KX���x<`Z7��XU��	�	\T	K	Mq	K	�Y+��z��t$X`X�6 .4�
f YNXJ�7H7�:�v�e�}q�vv� fl
�2��EHvEX-K.>�
e	J	��	��J<	��f	=>V	L<�fX�.KF<	P<	L���9V9�r���HL
���e=	>�}."[X	�	�	=X�}X���}J0	JK1M<��"	<"J�=;<=Q�XK	JJI�\
?GMML	.Jf<L
XixX\ KJ	�X	uX�ft	K<	KX�ft	K<	KX�ft	K	=Jf�<�/i%J7</JX�<<��z�CAC)OC)<> t<�W��
g
Jot=
f
=of0
p=
q<.s<9v
s<g0
st=

<�t<v
g>=
/�V.�X�<J�~<<f	Q�</�=	JIq�
#t�)�	Z�	�<�
X	�	>:X	ZX�{	
.X	/	g	=g	?#X	Z#X<	0"X<	0X	/	g	=g	?"X	Z"X<	0"X<	0X	/	g	=g	1"X	Z"X<	0"X<	0J	/	g	=g.//=>==0/=�~�.0�~�/.gg�//gic=wv��~<>0��~J=gX0��~\.��~</��~.g<J=gt>�
��{X02H0-P�
k�{JP	��{<J�JMv	L�.K;<�	XJ!�J.�{.K�	6#X<.vXu	Q#X<��	c<<<#�(	�	�E.��  \
�
�	�9H9�:��4
	Ze	['u'��?wX	y�X�	;l
	�l
	�;V;�r�X�{eeW� P�   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/autofit /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  afangles.c   afcjk.c   ftcalc.h   afhints.c   afdummy.c   afindic.c   aflatin.c   afmodule.c   afwarp.c   afglobal.c   afloader.c   afshaper.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftoutln.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   autohint.h   ftserv.h   ftincrem.h   afblue.h   aftypes.h   afhints.h   afglobal.h   afblue.c   afmodule.h   afscript.h   afstyles.h   aflatin.h   afcjk.h   fterrors.h   afwarp.h   afdummy.h   afindic.h   afloader.h   ftdriver.h   svprop.h   afranges.c   ftmemory.h   ftadvanc.h   stdlib.h   <built-in>      	�3D     �x
�x.`�&�	@	 [  I	 �  J	 �  J J yt XHXByJ5/ � � :ZfJ
t	
X�y� 	X  =  t	 G�	�Z;gj���
	g.X<. G^u	 `�    </ x<	 
< ���JY0t>Y0t=�.,0rOo0H+1LGK�w%�JJQ�wX�XQyXY�w��w<
.K
1	��J0
��h�V.��=[	�f	�y0V>yLuI=;=;=;KI��ZJj��v
<g
w	��J=�<J X0�
	YJ$HJ:���z�*�zJ;u
�z<K&J�ztf�K���JgAi� (JuWb<6i*gnXg<#���h	=�K
[
9< vJXJL_
Jyr Jv
J�t�*;uf�z����&�X 	�8D     �
Y0t>Y0t=�.,0r�:0K2,J�=K&<���MtO�r=<E�6�J�
Xm�8  J	ZG	[)�(X<>\&N.bXi�9Y&J..�?hKM�K�
L
	Zh�J6 wJ JX...� 	wJM�qu*
�<z<K&J�qtf�K���JgAg>
XE f�@ (Jtg?g+he<g>Y	<Etv�Y	<�o��s�M�w����	�|�z �  f I[	EL;E	JK�tJ@LK�/>#-t�nftb<J<���?	!�X,`
� XK
w	�	� 	:��� J	�J,;>g,	 �,  t � I � X w X�<1 y� . J z	Z	KM\ = JH= K JsX/v t<�BHQztF�YK@oY!z<u!u!�!��
�!,X=!1�
�="
	J.9"ztB.�
XZ0u0�VKKKZ�LG��O&,J&uJ	JKvJ5M,	ttJM:,	JG,[wJ	t"x<1<	y�..	[9X�<W=���#J#KI.?�J."> �<YLKK<�9 Z@ JG J	 J�KL$=IK�z
<�JK�z
<Kw	�"�J?< <JK�z
w	�"�J?< <JL.�=IKL��X�

<�J
t�>�:<ZX
��!xXR,=!1�

<�J
t�>.�>:>X
�M	� �	K3JJI=	=X�J�~�"XJ"<<�!+W=!�Y�	`�	K3JI=	= z� . | 1 H8 J L J �( 	 XJ� X��	Z4fX=L��
uKWJ.Xv<f$
<�"<<u�
%uX%/W<.Xv<f$
<�"<<X<<?oJX
�i+��K�Z�LJf=J>:>H>$<<$<J$<"�J^&f�Kv�|f�
d�f�X�t�KJ�}<� �  K 9 G J]L(?(9<�Kv.�J �	 J� �q�-<J9 b	 J�<[�&IN&GIKIN+IK&zX? X? S& J X [  X( >],>9b<JL,<�K	at� ��i,XXJ9 W�	 J�JMN�|�
	`	=f
x�<>fX�`(9Q(yXKIKIK9(S-PWS�:2Z-,2g:-X2<.�	�.f�Kv��~<<.X	�~us	K!,X=!1	n�	�	y�us	K��.[rJ�<u��Qy��5Pz�Pz��w��<�w!. i����	 v # V L	 K  � X��t��!��rX�X"��IYJ
��	S&<gX-1s�xDq�84
fq�;X��x�fpXXrX	��	
t K8 s6�	7�J�}	�v�	^	8JJ�}	KtL<NK[<>[f@hvx.Xt�A X  J�6IKB <Y6Bf <].�# gE ev L!
7xf$:Y� 7�.$;Y7Z!h� <!�<�i���r�X��
J'�2<2J<J?�	�wt	 zJG�!JsJ!XKtJ�N�!s�;CgtX
�r�)J�
�XY
�X	��
J	��XX��M2[<GM2JJM��)�<@!sf;n<	�r�Ys	K$J2<J2J<M��~�.5 geY��'XK'Z'XX&X!�!+j;�qJsfZ ,Y!h<!fX <Y!e<lf% Z)u<�~�X�A�XB0X%zXK�z��0t% �G e�'jC+�YC+�Y�2"TK"Y2":Z' KI ev$L;(,Y%;zX(-Y;[!w%_!yX%�S!:%�!zf%�WXLt'
�s�X�� 
�q�YfX-�����1+JJJ?
�Y7@<;;M�Y4?<;;J@ l J	Z	K	K	K	MJJXY4@<;;MJJY6?<;;@]JJX\�rȂXXX�	�.	%�2<GM2JJM�� �~2 X	x�K�L�XH	 � # V L	 K  ��t��7��J
<'�<�L �
 f^
��I4tZJ X
 f XX�=X ..." t�
T�&J�<�
�X<Y
X<�X
�		XX�ZX&.���	^us	KXwX.XXf\.X	�Xa.�	��N*2px8\K-'J�yfY�/t�I(K�<5��	MX	�	��IY		Y	�Y����uJ' � J �\�Y���v�	�v<.
<K
w	��	J<	Y	NJ7 � J �� fJo��JKp�IYt JK
�;.ZJ=�YL�J=JJYLT:XZ@�YJ/�6�-��(sKfXX�z y
�
.z.KE���tQytuvKM��, � J J��|<��|J
<K
w	���|JF�<y.
�|<J;�.
�|<�JKK�|
w	��J=<<KK�|
1�	�|��J
f	�M9J	MAX	Kf	1�{
<K
1	��J	>-mJ	K)
J)vJ<	Ld�	�{��|<
<K
<M	��J	0��# M� ȞJmX	KJ<�%)��YI� X 	�VD     �z. 	�VD     �/-=4�q2�Iv<XqtY2�rJ<,ttr�Y=* � Q  "  < X ^X" "XD�q���X�p��q�X
�K�
�p<1	��J0�X?�� dXxJ��J3 T J�
� Y3 WZ3Wl
 u; I ] �	�<J	=	�- X � J vX�y		\	$X%X	K	KJ	=X	=�p
g
w	�J�	K	KJ3DJ�3 � � JZ
���J z	Z<X	=	�X	' J	Y 	� 3`JJ�:�#N#8JK2J	Z	K �   K  L2wXJ	�yJ-D	�$rJJ:K+ �: J s g ?  ��K<�Z. J'<<=*�HL$X<=�XL�KJJ	�X�$tJ<:K�XvK:t	4��	J tu2 �� J � .� ��~�	' J	K 	� ���1 W�J.%� �}    
J v< Q* q < X ��x�yfl<
�2KE����<�{f	L�	�$f. � < J� �L�$K$ R t . � �& - ,& > J w �w   
 < K 
  w	  � �J . K  L   xX�w��w�
tK
1	��J;
�����}t�	�x�L�xJ��
�x<K
1	.���xJ=�Js	=	K4ffZ4VE		X<	L
��5KL$K$# ���tf9 ��;h�O7O7K+x �J	��w<��wJ�<
�w<K
<Kw	�
=;KM	H���w.=�J
�w<�<x<	K
�w�JyJ	K�w	��J?<<	K	K	��w	���tJ� � J	�	>t	 MZ<Z[. ��g.R��~�$d> �   J < < � G^�w��x.<��x<
<K
<M	�J���<<uv��%).�&<=.&<K.&<>YI� X 	�`D     �yk
<�Jo�
	Y<X�Jr�
	Y�u�tr�
	Y��tr�
	Y��   J tY��Jq�Y���u
�}JWi#�	�XZ6"s$@�YXZ�� sJ�h ,XJXX 	�bD     �p�	 
X^X��
	Z.t3�J
�
	��<� <?��.=iX+�%ft<.Z	�Xl<%X<<Xr<>	3WfJJX
<�X	�	g�N�Jf+gJ<��t
.JJ��JJ����KJ� �x3SRf.�
- �	�X$JK�-<=X@/J'�/s'=;'=<=Kz<g<���h
j  <$<��;?;;=>=>�<v
t
<<
Jf�y�
�X�ZK	JX ..J	�Xtx
6	Z[*VX*f\�<O_KMX ..J�<.�x
��<J�{�&<�=	�!z<(J/JJZJ=JL
<L����2��n
 v. �=[�Y
�J	h�
	�'w'9	Z�	L		��#6EJtM��"JJ� ?[M<t��'XfZ	�W'fJJ��~l
+�
�<� �'ft<.Z	sX�JJ��J�� �i�M9Kf<L�XjJ<��?9=�y�Jp��8(�#6EJtMZ�'�X%.J<>g<U'X%.J�<�<X^� J|xX&-IKqMf�?<<X&%<L.�i�z�<z<PYNX q��LX �	f�|J��|�<��|X�u2=Y2z�,<�<hz<KK8=0	Z	K<>,	L		K	h<,	AYX3mJX��|3u��tX2uKP,ytQN,uJ[rC<�6�J�
X	�.�J�*XM<j%#vkJ<+��-YF;1YhKKM#+J�-YF;1YhKKt8[J6�J�8>�J	�	KX4fAX,X	iJ:Xt.	JZ&J�KX.fw'�J+X]'�<�;vJZMZ��	���	Ptu�2�J�.� �3�|t� �L
	ZhH�JX-JgJ6uJJX��}2�q]7Y2F<,ytFYK,J�*��yfX
<K
1�	�y��J�.
�<V�S�J<�<l�	L	i<J.	=�:	L�OZK-=
�gXJtXMZXXtJ<X1 
	�' J	K 	� J3�XJX� �#��YKA2�J	Z	KXgKL2wXJ	�G;@	f$zJP,XhJiZ. J'<<=�HL�hXLZKJJ	E�[$FN,XLZK��x��	�~	�	�t#X	K	KJ	=X	=�x
g
w	�J�	K	K.�~��*4�!XX<�\J�&����t<JJ<CKK=;=>��	BuJuJ	Z	LZ�	NuJuJ!XX<J.of<<X��uX.��
	BuJJ	Z	LZY<v�u�
�u.
<K
w	��
J<<f.�IKG'L/L'HJ=K�	 � 7 H L	 K  _�=K	:�-�J� X�	 � 7 I K I[�� 	 � 7 H L	 K  X�=K		�J�	�<	[xJ	XX� 	 � 7 I K I�~<<� J Y6 I � <J	\�J�[J�	xJY
	��~'<	���~J&��-�J*�	��~���	��
	��~MJ�IK<I"[J�"IK<I�X-�J��<X� <�x<.n<�vTLX>.�=KK��|��|J�
<K
w	�J�<c�< �h-?�lT.,.<b�K==J`<N
<J
�X
�<<	�	=	�	�x.=C$=I�e=WXtP"J<�<<������	*�1c	�	[J	#x.YCx<$	<I�e=WX�^�|
<K
w	��J<<�"<�L�?<U��[
�x,Y;`x<D"�X;"=J�X
�}Xv.

 v�

JX��J JuJ.�c�.�~J(�t)=@(uqL(K(�(�(�(�(�(��~YJf��[��'fuX�J��
_
m	;\�rL/1�JKwXhKI���>JoJI	;X�	;��ZrL/1�JEwXh"tE�Z��ZV>JoJI	;�JM�� ��
"J.	gfJzf�!�J	0<�KXEX1�)"���}.�J�/J� J�~�Z&<� �~�<t<=�{�Ȃ��{><���}ruh�9K�o�Z�*JLX_'�='�(<5�~J�t���u�}����
� �<�0�?�K��~0;?�J��\J�
�r>
fLd�X=�4(�u�� �k�}.�J��}J.�.K�}
K
=w	��Ju�}
JK
w	��Jw
�
���YY�KKKYIYI�.:J�.K."=$M.T">$MWK
O.v�K$�K
gMI	��}J.��
�}�K
1	��J	3	�|J#�JM#�
�}JK#�
�}Jw�	�}�#�J2�i�|���|<���Z �~�
� 0��vXJ�MGwU[X
�� [V
L�= 
J	��V	Lh$J�>�XX�~� f8s6g4g��}ttX�z�Y1&z1zXM1�Z)J&Y�t=;Y^��Z�f?;?��	�EX�	�*	�$LX	U7<J
.K
1	�HJ�(�*Y(Vu*(;*KM*U(s�	�*	�	U$f	\X?J[7.
zK
1	�[J�*�,Y	X*iXu,*;,K	J,k<X	t*j<�	"W�'Y����\~�W���
X�@
	KJ	t��~J���
�~��J���~
�<
�~�M	��J3/
@}�
k 
J	��
	�#	�"��%�	�IxJ^xJLgO��KIKI��)��,��+;=�uf
J�~�	��5f�{�XX=
	�"��	v�	���y<��_	�I�	�)L:	�);	u)t<	��� ���u;KI���}GW� ��S�x-RtYXiX r.XY
	L"�X	vo�X��Mv�
�.X
�f
�f
	�<
�f

�f
�f�Y0��M�Z� X��f�
	KX�� X��J08X�X3X0�nf�
	KXh�J/uuuuuuv��}t	�wX	JwX	X.�L
+J)}� J �	�? Ji"=t
	tL
J� *X�
�~�J
JtM
	�XfP J>��.�~�
W�t�/
	�$��
!t�

 KX#J	zJ	X .	K-X	#X
K
Y
�Z-[�
v�9
X
xJZ_'�-�M = K = K = K = >�
tM
	J%#X�	�t	�Z��� ����	� t	�%	�~td"�^XJKMNKYJ XKxJKKIY=?�K�I1M.>.<yJX�I<<
�K
J
Yw	�
<J
	-&J	[J�<	&J @y<=H	-$> NFK#NFGLM xz<KM#z<PLx<L=LLL�K�NKO
&
f�&
J�$(J�Yv$(J�Yt^�..�	�F@Z fu#�
	�$<O�Y9O9K�~	��~f
<g
w	�	�~�	��~<	�J>X�R.f�
�	�sJ<�<=�KM�~	�W�~X
<XK
1	
�\
F	�J��~
1	�	�J���JJ	fXJt	M	��o"KIK
>���6x<�x�XK�
t	��j"�
XLX��
'X	OHYH;	��{	�X�{�K,&<J&jX�K�	��|JKe	KX	
�t2OJ	�J	M	K	L\!XJ	_Ks	K�~��J]�%�~f��f��
	JJ)UX�
M �w�w��|X;�<�XqX�<���~��	b��}���}JH�]%J��}JL	�X0RJ�
XjK
�
Y0I.�

��
f
�
� f.XKY0�~��JY�~�<X��0�@�#�0�Z��/
J[
J	Z�|,�J,�|<�J�|J�J�|<	�J0wJX0�J�
�J	geJY	�eJ\
	Z�|,�J�	�X�	���|,JJJ�'�	��{	�X�{�K,&<J&jX�K����M
J	 �	�Jw�;KD[pJ<_;K?^J	f0�JX	��e���$J	f�Jw�;KD[JpJ<_;K�� �,�z��J�zJ%�=	��t8�X
�tJK
w	�2�JsX�<�	��~�,&<�K�<	�~t���}��
J�}XH�]%J�%�}J<L	�
�� � �	��~X�~0@�#���~X��
�	R	�twKsu�L
�_�	Q�;	u�Jt� 	��~�^%<<YJ�}<<��(;8M:0L/,.%��!�%I�!J%J	0"J/<tKI	=Y	MZXu	w	Y	x�Z�	w	Y�p X 	��D     �y��y<t�XK�
t�&�x�<�
XLl��M
XFuYFW�'	M,�{IJuX	�<�{�&J;Y&�=&g� X���� �
X�K
	�
�
>	� X�"t� J		�	LGt�JX<.0�~J����.��	��m!2,J�=	�	K	[	K	KKIK�	xJKLX5oJX	��f���JEX�wX�X�w<Y��
V*JQ��wX���wfYL3��wX3���wtZ��
N$2J
J	��w+su%V�r�
�<�nX<��nX
.K	/��J<&r��n��VZ J	�<	Q3E	L	u��(J=�L�n
<K
<M	��J="�8<,�%i�.K�L�m
<K
<M	��J/�K&@�'�	��{t	�<�{�<,Y&XJ;Y!&_<�=p2v;<��'�v$M�;�<			KX	J;K;	K@�	{t2�J	�J	MuJ	J	��	_JKI	K�X�{3��wX3�t�wJZ��
�	�| !	O*� �1:J*L<<�
Jv�L�,g,>ffL,=<fL+>:L+t!<+=;!=;u!L�	�~X	�	�	�	�	Rx�	LX�~�	Ke	K�G�\�+K>A+y<;KK<<L�g=<<L7�K��}� <#��.��V��	,�	�J�+JK�	M��|Jt�			vXG�4JX<
f	��	� �m!2,J�=�	�	K	[	K	KKIK�	xJKLX5oJ.����J<J��J�#�"'J��J			vF�!lJ�t�GZ�U�tY<;eJ\Y<<�JXJ(J7J>J%IJ��}WX/f=JL,g,>ffL,=<fLv+!�"=;K"�F���	� �m2IK,�=��
	�X	K	uwKsu�L
	�"J"J/<�	=	Kt�	M�Xu	w	KJ�
����};�<	 �J�'-(	�	�t��y
	Z	KYJ$�J�	�h,�q	�J�q�%X�=	��t8�X
�tJK
w	�2�Js�	���	w	KX��m!2,J�=X�W�l��zPt�ltX 	@�D     	.zz&<�I<M<J f  �   t � f�JJs<M��	wJ	� . r�  � � f  J f 
< 
f 
J 
� 
J 
t �   t J J t �  � .  < f < 
� 
� 
J 
f 
XjJ<�gF� . rJ  J �   <�{�u�.�{tJ�t2�{�tX� X�2�{���<=4�{�J� <X�{v
<��X>�|t<	��I		XY�	=	2�L	�{X���|�
 � t�><u��v��{�������{Y
�?	0U	�	Z		��W	Y�	>.X	q�.<�sM X* �!�	J�:	W�:u.�	;Z�N�^X���|	 �   * ,�*�	M.'=.s'�.r*�.i	uv*,J*�	M.'=t.g<'�.r	Y�*c��t.e#JJ.=��.&f.J8tp. =�t�}��XX�}>��>�}t�0u�i�t�gf�<<J�I<		J		�/W	=	2�>	�}	^	�	��tx.vt	tX�*
�A<M��<t�<' J t1 ; < J J8 o < < X�<' J t1 ; < J J8f<<X9f	��t�~<��
>�1�~J<��7<E�.�~ K?� ���' J t < I
 �' J t < I ��}&xtDzf	><	[	KJy<XJ�XJ�xtDzf	><	[	KJy<XJ�X��JM�	��t
t	Z�Z!<)X�)�<�w
�WB��tX
ZHh
	�'fXW	$�	f�'JK's.	��X��x819	��<[%Xh�wX��X>i�Z
/W=
1� KLX��
[
X	ZXk�s./Xz�*=X ...r<.f!xp=w!V><XQ� <.y<���{�!yo>w
!V>
<XK�� <.u��	Ju�.�{tJ�t2�{�tX� X�2�{���<=4�{�J� <X�{v
<��X>�|t<	��I		XY�	=	2�L	�{X���|�
 � t�><u��v��{�������{Y
�?	0U	�	Z		��W	Y�	>.X	q�.<�sM X* �!�	J�:	W�:u.�	;Z�N�aX���|	 �   * ,�*�	M.'=.s'�.r*�.i	uv*,J*�	M.'=t.g<'�.r	Y�*c��t.e#JJ.=��.&f.J� tr.oX�=qXq<X�Z�<tX�}��.�}�Z�XL�}t<D�u7-:AJ��I	n�r	>	P[���$ N	 J��v�~^!v,t�.m<8m�t-h�s B[<' �_twJJh�L �zJJXJ<X: S J < X' "t_t wJ Jh�L ȺX�� .����J$�|�JX	�|�J	���"�t�|J 
�<�<
� �1�{fX.���}J��	 +  < ��zXJJf��z<v<	@Z	@	[	KJ<j	�<j	L\	LXmJ��$�}�#<��� t
JvX
�v<Y#Cm.<�Xi.�<�g><JJf���.X@XXJXXX�֐X�Xk<�<�g>�J><J���<J2XtZt1@X1X@J[@�<?q[J.i& Y( /& �? .B ; ��"I�z�z^��t �~� <�t+"tX�XX�XX.JXXXX�|!.t�})xtDzf	><	[z�	KJy<XJ�X+xtDzf	><	[	KJy<XJ�X��JM+	��t
�	Z.Mf[!<)X<t)J<�w+[+M9M+uvi
	K�
	K
	�DX
ZHv
	�)f�	
�)KI	u).�����~.v�t@$<���[/~B]X'JY<'<Y�'Xd��*Jf�Xg��5wf/�J<M<�����2<��.=J�I< X�J�X�J	RJh	NZ<J c	�<	f<	>Jj<.X#�~J�X��v��8@J��g.
X��@JJC.��J,Xg!<SX�J��=�!v!V><XQ�t y�HfvX� <Y���|���|��t}��|��|XX��|�>�<h
/W=
1�|KLX��
[
X	Zfk�s./f�|��*s�<�|X �>YyQX.<_Yv�  s;   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/pshinter /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype  pshalgo.c   pshglob.c   ftcalc.h   pshmod.c   pshrec.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   pshglob.h   pshrec.h   pshalgo.h   fterrors.h   ftmemory.h   string.h     	��D     � <#U.�
J
<[zJr<  EA�\�<=�C<<	� 	>�.>Y>;� XKY*.tL�)p�J�<.tu}_�t
<K
w	��~J=IK�K�.	L� �~<
�<K
w	��~J	/�	L	�(rJ	KJ�qX��Y�A& ��u<,v[& ��u�vY�|t!����~J<
<K
w	��J�~�
;=
;M	��J	Y<1wXz$-K�	h�}'�J
�~JK
w	��JA<	u�}
JK
w	�N�J
�~<A�J	u�}
K;KM	��}
w	��J	w�}��J@xȐ i<Z�t��}�� 8�}.�<owt	�p?u�f	*Z"<f/�}���}<
.K
w	���}<�Jy�"f/�}���}<
.K
w	��JX,w	J*yXJ�jT�.<	�	wt	=u�X&*nJJK&JK&JK&JKj�|<u�u�u���}uv�}#u#u#t��}#u#u#t�)��}uv�}#u#u#t��}#u#u#t��w�K��z�>M��YJ�z�����z��������wv��������wv�J<X�qu�X��r��X �J�=Mt!�%� t�JX�uut� ����fJX�~t�K%MqX�s�#Bw.�vf.
�^
	Z	wJh�Y $f�SJZ
	L	KXK*�AX	v	K>&.dZJMY	xXX���.e y��v֐�m<�'�X[
-�	[�	��&�JZ
<[zXP
	`t��=*<M?#X <Zg&`JJ=_�XL��=*<M?#X <�zJ	!X��L�?f(Y9e[Kfe�=$*<$J:<Mi#X <�zJ	Xf���=$*<$J:<Mi#X <ZgI=�"eK=��v�eK=�u.q
Xq.
Xq<
.q<
Xq<
<qX
Jq<
J 6JX
K�6$
�6�
K6Ij&�/{&x<LrKF��	>(,0JL	=<	=<8
X�9ML�<	/�ty5y<5X
ZP
M$uJZ
	L	YWJ\
	K$wfJ		<X>uX'� J�`J
�J	� &e	KWXKX.e��9ML�.! z�/<
H>Q%fY,gu1KX J[ft]�E��q.t
J	KL�f��w
	JfX=X �}��<	A�}eL�t!J�X	�	M�}e<L�t!J�	�JX ��y�*37%7*\0*�O)K_�g<;<ft�J
J	K"<?$Jt3	J ./%. W.=
;K%.
.1  t��JY
M�JzZ:l�YxK!M?$ �, < J	L Jf�|KQ#JJ[��
M
	Y<f...Jf.	�{
HL_ A EJY	�	/	KN�|KL#��|J!Y�
�f...Kt
Wl�{�]�1=�=<W�t
J	��	�;i���	k	.kX	X��A
J'uJXX<.	yX	YX<.� <YI���}��X .%����� 	 > 	 Y   U �	 |%  t I\�}<��k<�t�{�=Z=(u(�*�*�*�*���~�fz�(�f� X&�} �X�HJ�~<�L�	��~z�K�
J�
J[	AK	zJ	XM(� f� .5 H < J X :	M�.� �tn<@�
J�\&tK=
&yXJL	C	�H	KJ<>u	FX
u�.f�
	M)�	Ix	8GX	[\	�@�Jf<t<��~��� ������}[/&< -/= ;=&J�0�J		�� .��=Jp�y�}J<�=�}�~L�tX�%J<X�
	L�}�~<L�t�%J�<  �}.��  .�x�y{/x(=�Xo�
<	�>Jj.@	>	�'aJ<	0X�	J.��;[=>
	YAJ�.� �/=  	K�>H	>vfA	mXKL	1<dXAQKz�fK><�EA�u
t�<<+wZ�K?X�X	M	=J	uJ�h<g	  	 =,  X s XJv
�gY	w,;	K,<	uJ�	 m,  ;	 K,  < s Xcf		 X   � � < a< �	h[@>���:54yJ<Cr<ZKh�N(=?(F=(Mr<X>:	L�9<�# X.��=t� f<���S�XX
<J�*xt	N*�	�s	u "  > I I = 	 _+	t1w
<X1v	�+	Ys	u 0  > I I = 	 _2F AI2F\ Ht �zJ �E$	&�~Xf.�80.�)<J	X	��~X�h80.�)<J	X	��~XXJh80.�)<J	X	��~XXJh80.�)<J	X	�J	�'#��!�!)>���!��J=X .�}�<z�.xR<z<t^�}<��~<
tK
<M	��J<�J�}J
K
w	��J>
 � �& �MCw�� ��MZ��}B�.fB:.f@B9�}J
<KB�<J
�}<w�	�}��J(=<<<<��<��~0�08[�L
	hX�
	�	gdy���~�X�~JKWKI2=;=?
<
<J
J<<���;K
	�I	K�J	v�K<<�JL!<KmX<.8 �~��&��MCw	
�� J�	��� J�Z�.�
f[&
��pY
[&
t%z�J`
��=JJ�Z�=;=
<[)
fȺ�g
[)
f%z�J
[.��	�)W	K)	u�d�Mz	s<	[:	L9	K�X ..	]����JJ�~�Mz+<� 	e�)X	u�	K� �_-Y-Iuw�XK	Lt��&I&gX	���K&J�Ff�=W���X)P)zfPz<K<K<�utXXX	�~XJJwXJ�.�x.�.
�x<�<%�x��<#X�x
��X�xJX>
�X
�xXX.%9X�
JJ��v������X�
�xt?�
K?��YN}�wa	"f	K<b.X	L<	=	L!JK;	=0#/#I*J��Z#JKK<E_	M	K<b.X#KA.�<	
�J<<KI<=s	g�~;=IK;=;=;=��,|�,	LJ<=I	=	>�~=;KI����,��G	M�h,t5<J	�0�0)�I=;KI	K0	KJ��~��U	M[�9W0
�~�JJ[)��U	M[
�~�JfJ�)�W��~����~�J>-z<&JLu�		KJyJX�~�� �,�XJ�
�j>�		K	[	�L:LȂtt<	K[�	L:	ZZ0t<X�	v�f	<K�JgL:hZ	0Lt<<	<.	fgX8A\J�X�"V"�H�O�"V"�H���$��qX��qt�t�qt�<
�qX�JY�p
1	��J=L
J	"m�<	>	��y�
�!Gfu��!f�!�|��X�!<��|�	��w���K�	
�-zP	K&yQyJZtu�
	_-uJ	K&tJtJX�X�<
8�,BJJ� X<ZtK
<�*XJX	��u�tK%�K�W�	�
�{&
X&vXJK=4Z4VKx� \XJ��J��YX�	�/pL:	�	�Z@b=,JM�%�X�}�z�		=�J>		�K�(J	JZh	X	=r��KLSKL��
�z��)J	Jz�=��f	�t<Y(dJX	��pf �(J	Jf&`J�M
	Zt[]&<v�"���s�*-�s<
<K
<M	��J:;��<J�<	#f�|#�y�/(tJKx�
Jg4cJ^n��W�u
<4�JZ
i<X	Z(JJ	�J	iE7J_=4pJJp>Xt.	^J.X	\4t�J�
J�
<	JK.t+�	<X�!<J�f!XJ�-H.XJ�!�����	���~���w�r� �"zJ=JKX9/	whw/z<JX
��w<	Y� X6�JX	��w�o�XKM.	�@
	K�J*gJ<�
X	[L
	K.�	�Kl$X�	�=;=?��$�q�.�[�q(��q<
<K
w	�(�J<DLLgXv[�q
<K
w	��J<?LLX	>�sf�q
<J��
f<��	F/�rJ�
�rJK
<M	�"�J.	>�Y�r
JK
w	��J=.1r	J.��gf����wYLZ ��s
<K
<M	�,�J*<�� �r��r.<
<K
w	��J'-J	+J�D����{X�0�*W�	�}<`zfK�
)X	���~��.f	���.��
�J
<�� Z�r��r<<
<K
1	��J*-J�$J���<2�{�J�
tKCsO
i	pMv	�!t?q	i��	G!J<	?	[!�Y6�%tZ LHK1sJXt=!JJZ	�qM9	?f�	�J	?	�$�Y5�%tZ LHK1sJ��|W���~Xr�U	M��~��U	M��$� KfW ,��� <<8.! t� f� 	��D     �u��i
Jp�<`4�=;Y:4gKH4=;\�	zJ4X	JXX�~�&KI=]+�{�4X.4f+<f+<4<f4J<+�4<<4f<+t���{.M
���{�[/���{�[/��(�	X$X$�XY
O��
N_��X<X.�~�Q_Z�	���~X�
�z��XJ�|K���zJ���}�J��|���t�|<���}YJ��|����u��zX�itqJe<LJJ�!J�<X	JX<J.o�}[=�#JJ[!M6+=<S@+6;>I-=\	�	>Vf<.	y+	00K	[.0KlX<.�X ....�}t�Y��X ....��vx.nKN!
JJJ.�a�<fnXJf�
Mv
J=  ..��vx.n=N!
JXJ�a�<�n<J.<fZ
Mh
J=  ..  &   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/raster /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftraster.c   ftrend1.c   stdio.h   stddef.h   ftconfig.h   ftimage.h   ftraster.h   ftsystem.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fterrors.h   ftrend1.h   ftmemory.h   ftoutln.h   ftcalc.h     	�E     �'�u��K��vXsJ�Wgw/e�
	K<o�t/]�ux�uu /tJvt50oJK
	ZKkHvL�LK<�mv/x�uZ�u>�KI=<M9?<".J<<" J XY-J�
kK#<<;=#+m�j.��<?< 	   q	 1   	x�	u� KIK!=';�K'<x'F<K<<vH>!L=EL'�K'<�K<<�N�!L;H!M9K%WWJ==:KY\yJK=?GKX:KFL!GK%!W>W%;L;I?UKW=<KX:KK��v�u<.uJ	
�K	IW	JK
#<<
<.X>w��.t<Kw�X<"��f	�J	K<<J��= X_Xv
L
	X0u<JLJ	>>X�i;K-KX��t=;
X=
@	�	j�<	P>H	>"t$<h$:<$J"�vJ<f�KWu,X f.�.Kt� X�KKKKYL<:�<fZ X�!tLK  .� �yo�IKruLru;u�
&	�#�@t
	_
	t Z  : h @ J K+ ��ւ	���N�K,LX<	NtY	./f	g Z  /��IY <%��o�IKz`ruLruuuu�
�f
�
&	�4f	i �  J � � J K+ ��ւ	���NX�.
	tY'�ZK,LX 	U��	� �  : h < ���IY  ��=�"J<=�W�E	X
L�	�	K	LXlJZ
	
�	=J	K9	L?lJXJ���.u<JJuY/f5<J�	�
LiX
<.>
H�> � c ?( <: I� � ���
	Y<>?#X:>#/.U#M8K
"=+0
u9+0<
H0
<	L<	A��J=�	]�[
<h*�	b<X	�_!f	�;=	=� tX> X JZ6?<U&M6�&.2��
<!S	�(���<iX<	
<.Z.&�J�	 B 	 Z   ! � J �6 @ F N J6 t <6 <> s!��<	� X!�<3 `X��!<J; 4 I�<h!<J;9f�u 	�J<<<Zt
.=
>X	h�.	>/ X f <Z(&s.$W&K=IK$LvY0JJ>.	�i�	�;=	=� tX>+ X �Z#s!-K!e#K=I=�
	Y/<J>@��
<!S	����<iX<	
<.Z8Xf<�	 B   o" 0 ,	 >  "  M" 9 M J	 u Y+f1<J	>$ �* e$z�.$f<*C!��<	6�!�<3 `���!<J;4 �Jh!<J;� �����g�ufJ .J>`>J'JJ< 	�E     �fX 	�E     �ow	.w<	.>u�t� l
�
.=;g<
<1��-=
�
	�*X�*I.��	=
..����
fKt�����=X
JY
	X	=W=��JL
=
<	0	=>uXYI/���
Wg
;=
?�
�	h	��\X<<f
�Y
�K=0��#]J#X  .J.hJ/
YVgX
JY
	���1�
JX�}��< <Zt�!tL
�PK,LX .	]�$J$.X�#�EJ;X  .A�
J	�/&f$ 
f ID W Jf�
�d<
J	Z$<$.��$ �	n $t;<.�t$ t ���f��@.!�xJH|�<;�Ju!�x�F;���xJ�v��J~LJL�xuK���B\�~t<���~J�J��~JL�muHt><?G=I==H===:==;=>�<<?<<t?<Y�>?�M
X	�!=.;=;KI=;	=.@KMKL��JKL<�K�u;=;==�<<��p9�� �J>��KFK==Hu==9===;=>�<<><<�uI=;=<>�<<�Xk�J��� �
�	��K�u;=;	=	>�<<	�t�&Z,:&�,J?,9�X�	c��K9KZ=s=;=<>t=<<��fX�	�	�xt	�J=su>+	/ .	v 	(0	u%9?0:	�9	vXt4�I/��wf�	�(X�	�vtI<<f�	� X<�� +t[M/�?
<#Xg	�t0Y2�[�
J,�	�wJ
��
t	YJf!Z�)��v�v�f.0W	.��0�	�JXd.	M+u+	�Jm4=4;/�ut	���
�	#�t��}�{�u�{f���{���{�<<Y�{t��<<Z\"K	GL"..>
fh
�u�z�
�
hKE`K<�qX��r��
�	&����}���<xZ���	G`J�.&JJ/Ih
�{t���	Zf�	�I	K0�zZZ
�
�BwJX�<��zY�
�
ZKEXK<�<���*J3J&<3J%JK$��f	N	Y	Z3h=LXfCMc=U/W<=;@�&�<�f�KTJ	2�	�fv		Y�	�W	K/�zZZ
.BwJZ
^	F	=<�`	Y�	�W	K/�zZZ
�BwJZ
^	F	=���zY�
 
�KE`K���Y�u�/YZ�
	v	x�KpJ��=8M u��z	F	=�ZX���fu�y.XKs�XK�X�X�X�X�~Xf����zJ^ <..t�wXX�� ��V��l���K��X+ �! J�J( � J�ewJ7
XI�Wd�<� � <MyJM	Z#�#��J	Z#�# � <Y�/.Jf/�G9tK[~����U���~�m�u
�KKJ�L��<4nXBz�Cy�x8}�8;8��zt�Y}�ZXN��1w��;�z���;8��;�X�tQ .�~.��m<u�.�uX
�JL=N4?f  �h����t<X 	�+E     
Lr�Ru<���/B
� �t��K�t.HtU_��M
&�"	r&wv"U&=qL";KI=>Z=NQ�3�H�4XY�?qMh��k�� �XtW�XȞXXtW��J4zf2Yt<Zt<Y�t[ e   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/smooth /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftgrays.c   ftsmooth.c   stddef.h   stdio.h   setjmp.h   ftconfig.h   ftimage.h   ftgrays.h   ftsystem.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fterrors.h   ftsmooth.h   ftoutln.h   ftmemory.h   <built-in>    string.h     	0.E     ���p�ufJ .J>`>J'JJ< 	�.E     �fX 	�.E     �z>8J>K?�?UZ	�wt	<.ZrL~YUg<Yf��X@D�@<D<<���.K.K.K.K.K.K4j�<X<X	�fX�v����t<X 	 0E     � < J9? .K=
X[
1wJK
 X	Jtj,J,Jt�/<=>H>>	oJ<=ptm.� 	�0E     �	XZ�
XJ�Km��K
	u�K�==;&O*K&?z<KLi�J�-KXj%�8�Xh�FL�4�4GK	�tr�:MSK3Tf?YTL�	�.	l;	KL<�[�	b	gZ�7	�	K	L	ZL�|J�$<$JXKX*		�%f	=f.	i"uJu<	Z.XK.t
	YJ,iJ .X�K Q� .X��=Ws�J�J+ �! J�J ��7f;e� �La<<�h
J���<[J) �" X �< W)�"X�KMz<K$KHK$HYY[�KH-<uuu9KHKKL#�XX�t� .�f�� X@�
\
<t�t� .��- %� <M
J[
<	M$*<<�v�LJ
� �YJJJJ\ved�u.u�
=[
9? Jw�9U=>9& X X > X9 � � > X �w�X��o]7^IK	<MX �5 e��u	[8=	>?z<KPW	z<=	:ZN	8=	t>
>
��"<=�"JJ= X = �.  < tJ F. � tX T f < <v�	����.�\;@J�zXvVK.K;�	׬�<tXt�u	[8	?:I	KZ	9=	J=	t><� 	<ZH	J>/;	+[K	�(@<w�����A
S��<	 F    M = ~ �  � �   V	 ? � X? �[Z2zJKWK.J=h:geY�? �[Z\J~,�@9�)K.K;�h? .�.ZwJ:9�.J=h:<Y��f<JWX�y�	U>Y;�<<	 �    K  > = 9 M U u   V	 i �Uf�.J=t<j�y=L9�L)<<)JJZ�,�  .���uX
�JL=?f  �q��rux
Js<�Ktf��u<;
�.P[Kt..��~<Z�n<;
�.L�s�Mg��~<��[
�
J���dLYW;38;A9r=/,@Z=N<�G:tF�:XJ� �
9�$��O�X�~<a<;�.�~��XtW�� �mu�wXrKfK.L�Z
=�K
.����  �XYVZVv
��K
�Jt+z�
vXyq�
=sK
i�Y�v
�sK
�JJS.J;YL�>HvZ
KeK
l�
��
<�J..�g�=�<	a	� �!  J /!  X J K!  X � J	 F^!w�		JXwXX����JWYVZVv<�K
�!�/eg��� 	 BE     � 	0BE     � 	@BE     �.KrJ.KpJJu��uzt�YW$	�y<_w<YzJYYY[Y,s$�.�Z,sZ,sZ,s.�=;=>���
�9N;9N=<�?J
>\�<=JJ
>&f-J%ff
<Yf-J%fJ8;\�<Z
��f���!=K!Dv<==
<t<KFKH=ByJ>;!
<wJ:Kw<KDuJK=Dw<KI=Cx<=;KBzJBy<KPz<A=IEA7L>� <�JK8K;<KI=� <�f=;K<;K�J� V�it,s�,s�uu:. K;=�J<<Y�~�
.I�u�.o< oJ�$x9qYKYYY[Y,sL,s$�.;Z,IL,s�
<	J
wf=I
�t�hK9f^<+���\	;�!K� <�.K'=?>J'�JKI=;=<Kf:K!xK'I8'@FL'=s=;K'<K<�J	:��Jg�.�ptYJ\�uu#t��J=�f<Y�v.4zf2Yt<Zt<Y�t[ N(   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/gzip /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  inftrees.c   infblock.c   infcodes.c   inflate.c   adler32.c   ftgzip.c   infutil.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   fterrors.h   ftzconf.h   unistd.h   zlib.h   errno.h   zutil.h   inftrees.h   infblock.h   infutil.h   infcodes.h   inffixed.h   ftmemory.h   ftstream.h   <built-in>      	�HE     � e .`<�a�G`�� !� 	  J �YX	�.K�f� Iw0
Xgt I <1y.j<�Np	<:�n��qKfI?j�.J#.J" � .[.f�N	:�	<�=JJ	IX�<K
J<JJKY_=�y<x��7<
��� �� tmfDJ<.J�3�� J���#J =X8Y=;=I==I:>YNJ\�	�<
z.	K..e�i	`JJ	��IJ	�
�Xf�<Z � .<� J<.L@*X
X	cJA � XZ.h
WW=
�f	�
.J=s</�	 �
 ! ;
 / J �NJ	 � ' - .L	1g;J=.�	�=
:	=J.8.��XB�Xu-g	� �X�	��CXXJf� �)��X
.f�N�	<���YJ=.<YJJYY�2��~GguJKH�Y�J0KX c  X JW.Or.�,�.
-�.I</'u
/yX_� X J- X) JW[MJY��Y��0���}g%�
I/ yX_J</KH0:hY��	uX�-	=	g�tg�I���<��<ft�< �ffffff��	t	��W�	�s&�YIKI=s�X � 3   J J = 	 = ��n X���uKM[�~M[���~f����uv�u��X"�v..��� .�|�X 	�RE     kX 	�RE     q%.-KOXY�c%..hJOXY4�
%)
�XJ� JX
 A<$ WP' �uu|XJ�	�J	M�!	�J	��[�.
J � �% I  #��~tzCMFK( X K2 ; = Y   J <[/s=JYJX.JM�;Y?fK8MX J.Pt�
IK<\=Y�"J�=
GM���JM�;Yn�Mw<	<Xu��s 
s����WJ���|<�%btJ[%b��[�%f�GJ��J�=MTK:4uY	+_�
/ g�/u�$��vg��i���z��g�*X` .t � J �- �) <�#� f#�XL#:Y fX%X � )  u2 e � @ � *  u3 e  J K @ J *  u3 e  J K @ J *   t �  K  W g=X�<� f � *   t �
 	�	g	�	u�� yJ_�� � $ " t
 <	�	g	�	uw.;X �  " g ;" � ;- g( X - =-  .
 <	�	g	�	ueX7�gV�u8X�<� X � *  u3 e  J K @ � *  u3 e  J K ��<�=��� X � )  u2 e � 3��4��
J	h	g_<(<�JJ�J����<� <X��<XX
� ��2�� �JXX�6M
	�	��~	��~<���JJ��,#MJ:g<=q2ff�J�f<�f#J
<�JYI&	�vuBX<�JJ��<JJ�~
�
��'X,Y:.@<,<@<4.s	�	YXX�J�f<�(X�	K;	Y�0XI<0=W<4�;YX;�%<<	����J�<5<"X	u5;DX	=DI	g;X;X%<<�	><�5<5X"X:tsX[2�X?X@.�2�X3X�<�X���0h����/�

X8��<� JJ��<JXX�~��JP0�P<0<JfY<�X�/	�6
	�}X���}��X�}<��}X;"UK�J�}X�J��}XgK3	�Z="�~�X�~<�XXXtJ<Y�}� ?�t,� �JKX'*<f�J�f<�>:Z:Z
"�(<<	�)u�)
<�
XkJJ*:��X��B	;<A
�X�X�X�J��	Yu=	JYV=	<=	<=
Xy��f�JJ�
��~�='	���<Y
	�@�@[	`� J�Jt�f<���;=.�gY�YY�֐J�Jf�.XX��J�Jf�'	���;<
	�<	Y=�	Y�� 	YX�J�Jf�1/Z#�#;.�L.Z	=	I=Y	�;Z�	��Jt�f<��t=	I.	�	bd	h�X�<<X��<XXX�s<
	i	K
	K
L.XX
���
	�<	Y=�	YY:	YX �J�Jf�'/YdwZV?V;Y@�X�� 
3�Je1JJY
J	v	g�	?�
J	g	u��!'<
<	Z	g	�	up� �	yf 7�.	�J��<J�gqf-�JX<��J�<JXX�~� X�~ ��	�~��<�<f�� �cXXcJXZ�	�	�	�gJ�<�Xj��Y&�	Z��=�	W��u<	"J��<J�<�~<<X�<XXX[	0�J�� ��K����J�f<�hX:<�&<tj<<�	�3.t3J<.�!%JKK�	'<f	�~��J��<X!��sJ<JXX^.�J���B	;� ����~X,� .�4�}�Y;1� XJK�<gWL�3�!� Y�^X*<JNp9u�NNJJ<Xqf�X�%<�� X��/��	�u	K��X��<XXX�)�
	�vX!<	��X�	��<�� �zֺJ=�	Q�<<�<J<XCX
	L	Y!<	���<	��X��~<
=�		gM� XX�� <3�}��JJ�<�~J�Xt	9	u	�X� XJJJ=[�u�JJJJ<X�
���fXJ�	it	u	�X� t�zY
��t
Z`�	JtQ�/ p�	
q�tt���~g�7XXtf<�<JXXQ<<3�J� !8�JJJJ�	� tX<�<<g��.3pKs.t�uKvVt�
�.LK>	�
�Jk<�
	vF=�Xu
�
zJ��	-	�XX<.L�t1	&J	u�zJ4 <.
C�YXX0XMXf� �y'ytC��k��+&t�
	Y:�us<v
 <Jo<g=:Yu8:vY
P < .JUt�~t���3< f.]�>M<Y+t&tg
	Y=;uv�;uv
<i�
�<�MZsuK!�tuu)u��� JX 	PuE     z �n<JPXK�M�KI�XJ<��}Ku<=N�Z���Y
�l�
XyX��I�Z��Z
X6����"J�sK�	J:!MfM�u��XX�Y�<
�Mb=
M[:
J	�.J	J��}��K	�S�[:!c./X��	��}t��".�}[[	���}f����������X(���=��X	
J�fX"tytXtJ;_VZv<KZL��YM�/Z�

J[[�G?  V�*XXfzJ^  qXZ:>tcf*Xw� "   P  �      /home/computerfido/Desktop/freetypetest2/freetype/src/lzw /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftlzw.c   ftzopen.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   fterrors.h   ftzopen.h   ftstream.h   ftmemory.h   string.h   <built-in>      	`yE     � 
%)
yXJX
 v�$ OzF\  � � XU��zJ=f }. A�
	h<	=	�/ � �dA
�C�%�I\;Ks�=u���,>XH=/>NZJJ/s0:/KtJ/JJ1XVt
	�	u%Y	u.n�X  ^�<,�#t<c.Z((x<((<Zvt
JyJu
`
<	��XA�X
J�v/�	m��	�zJ.
�5X�K�uuuzs=J#uL�vrvK�c�K�uut� tz �	k<J	JXKMM�KI�
�JJ��u��X .�Yn<�}H	Js<KKLtuu�YQ	�cK	X�~��[�"�~�&zt�\JJwY��uut Y<X����f� �KKUP�~<JZ���~<u��~<��X"����-�:KK?[.f�X:KK>J<  J.	�t  ��u;9M	k	�J� gUthY*�LJy�<	J<Z(J�*,JY*,JL	M	g	M�~��X �D �	�&u�=;	=.f	�	[=,	u=y<A=�;	>�	@	Y	wY	>	�n��� _ �.  g��	.�	< . s	 = h i�l<��  �  J zJ�� � � ��~u�f
�
�
JJ�/L/VLrL\�X�f�<i � �  �	 � � � ��~Y�� r� tUpf�5x�gM�t�1t:<t:<<
<	Z=s	�bf�<t� &=
X	�=;Yuv2�X	�t���$![�'tK��u�U�uu	� ��� �5�0t=� t�<0?w=;uv<	��
��nth
[�
X+�=@7Yv�y<Ov�tJv/u ��   '  �      /home/computerfido/Desktop/freetypetest2/freetype/src/psaux /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  afmparse.c   psconv.c   psobjs.c   t1cmap.c   t1decode.c   pshints.c   ftcalc.h   psarrst.c   pserror.c   psft.c   cffdecode.c   psintrp.c   psblues.c   psread.c   psstack.c   psfont.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   tttables.h   ftmm.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   afmparse.h   fterrors.h   psauxmod.h   psobjs.h   t1decode.h   t1cmap.h   pstypes.h   psfixed.h   psarrst.h   psread.h   psglue.h   psfont.h   psblues.h   psft.h   psauxmod.c   svcfftl.h   pshints.h   svmm.h   psstack.h   <built-in>    ftmemory.h   string.h   stdlib.h     	P�E     �Y-J=t?>�@�{�>;E<[tll
fJ<LK
\X
<wJ<sX<.=�>Xp�~>K�Z�Ybf..=
���	�frJZJ< ��	v
 � J�
 X	iJ<ut�>J�  6xX�CyXYZX[XLX< r<ZMZZ
X_pJ. <�  ?Z �n
vJZ<	ZjX�
<XZ
FX
vJX=�=�2���QX<>
L
		J	\	J�K`�>X>g�Z<V A/  A E�<J	DJ	�JhJL8� �K=�J�<�
X[
�J
< N  U^
lJ.= x�<Xz��	�	�> m� � XL	QJ	�>z�� X�>X	p<	��~.�
<JL
F�	��J_Kl.>XU 8��IAX7YYT2�
<<������ 1%
y�� �A�� .D�
�; `�[I=X JV=KfUf
�
 ���PX�
J Xf
�	p���
�Wf�3�.<X��;t �
�z�uu�iJX=IY[<�K:�=Y
;=
	��^=X .��u�L
X	
J3�Z�F.u�L
XJ	<JHJ6<u=B8HXX=<ZXx<n�	
X	=���	� <lX X	x<YJMJ0JK (��iXZ tX .JbJWKY"JN%�WK%JZ		��	"Jt	���<�	>WKZf....l �.�z��� 	��E     �y��y�J��y<X�3>J�Z
�
M�x��y
MY'.@ k��x@<x���y��ffZ�i
[!	<u
[</
	ZJ	Km<Xm<<<�<Y<��AXY<+. �x�	<<x��y<>
  ��d X�x��y<� uKK=Kn�� �MY&�  K[�$ f, J$ J X @1  J��]�2`v6$I-J=;KI=Y
�\'t
<	P4J q� J	gJ� 		=I	=efg�.MY& M�-oJ<qJ-IJK	,Lc	=t�� �K[K$ f, J$ J \ F @ h6$I-J=;KI=Y
��'<
<	P4J[e F2 	�	�J��		=I	=� fMY&� �p��pJ[.wsX<<>"=;="J?.g<y&zX=yX�%X/X/Z1�l�u����  �=wgs=K���  �=wgs=K���   =2gg2s-=Py.=����91& K8 ;LfMl0H<'yJZJ.K
t�K
JA._1/vXD/y.,�#�KB=xD�t�f 	P�E     ?t< 	`�E     ?t< 	p�E     �
,
v.uw,�v<uuuuw� ��f<J�� <	<� �X<	� �%�K�K��%�	���J� <��f� <<X	��J	_\	f�0	?%X	*<f	
�J	gt�~�	/�	�� �	<� �X<� f�JJ�JK%-f<J�%-f5<<t�	5  �%�%����s�J ��?J* /. f7 Ih,]2Jֺ�t2 J J	�-M0X:vJJ	.�~��~J
XK
w	��J4Wt�~J
<K
w	�J�	.�~J�.�><<�JY�|�fl
X�|���7" . t�&?J
J.&J
<6�<+X
�}J��|f9�2�C
���
�	�m=
���h9X��
�~�j
N
J J]�| �.J
J�
�}J� �|f 9 ��
	��	��|��|J�J�|.
<K
w	��|�#��|.#�J-.	K#f�m�=4<J < > 
 ��./	t�(N"!��
	�('�(I'u
J	O�<t�	[X" Xj
�}J�.�|�9�X�Xy<";K3y_���tv�1�t<<��tJ1<;=9;�.NL
	�J�.t	��u
u
1	�J�
<�t
tu
1	�J<���;.� �
.	\ J�.t	X�t
u
1	�J�<�t
tu
1	�J�<��u� t	j. <JP%.t[Yf<	��<JP%.t	X�t
��u�+<yf�t
<�� �OfXu�����X���}f�J?�|Y&�t�t/��f�t� @tX� �~t":A�X�u ��.i@zX	J
�X
J<	J�yX��~(KH>H=�
<	Y#cJX�KeKXX�
�S
O7
OXX<JM#J=Mv=K��X ..�|�
37
]S
O7�K
.<�
JJJ��X .
 oJ1 ��WKKuu��(�X ��&
v�&
.v.Y/QG�&
<	Y	�J� 	�.Xgf� Xa�	JwtC
XJ
J	L	K
vX	Li	�JXgf� KtJ. <� ��Jf2K8KMYXX n�J
��
�M
�u.�w<-=-�JKY;��;Kfhu  ..�t��<Y
�tf<�j<��WZV>
�
g
e� XY�e� .J' X f��� X>����
О	V	�t<�qJh
��
	�X<���
\J
<��
.�~Xf�\�70e	$�4`<$<' 9Z
X�
<�>;�vX��X\�7+.�	�J�P&e?�Jm�	�< �	+	�	�"XL�J<X80�	�J@
<iuJ0�
	�ftXJW	�<�����<X��~<X,XP<e� .�t��.�;Z:�Y��
�W�
�u��
�
�"�	Y�-UM
	��
X]J_�Y
X� �N�
+�<XR	�	K�f.c���y�J�y<J��yfX��HX 	ШE     �|ufXuX�Yt�
[:WY
M
�d����2#�]X2"X�X�~:X-XA:S<K�f�Y���^z<Pz<YX<Jfk0-v  k� fJ#� >  U M  X =.  X � K.  t � K.  J � J xX�	�t���=�K�K�	L.�$JJ	t	�� 	af�YJX
	�JtY
� �XY	� �=	p�	��0[�	Xwt0KfD��KsY<ZȻ.J��L	>��	��/�/�N
�
�Y8�  I=�~���J<3$]KLx�=N$=$:LY
=Lj�
�	h	
�
go�	��X��~���J��y��8��$XXX<ZJ�'<�E=N4 ., < � X�"X4sJ+J�L?�=�]

J=N�.fWJ.�A	Km���T,X� <�y��z.�< �yJJX��z�<�zJY�=
��[
��u<�
�
�X"�7Y"I	u>
X	^L
t]JZ�
XX =��J�zf
+�<XR	�	K�f�c���y�J�y<JX�uIX 	 �E     �s=J%�g����LHLL K LnJLY�� �K�f ��� 
�t�v
.vJ
�y)Jt
t�NK�KKLX kX�}t���LXL�
h�
J(d<J
�	�~t
�
J�{�E�  �<Ov� i	�~J�	�~.X��,XL��>
�
�$�
	�m7B�iKHJ<KZ-!T� <�f� ��  .��X
	y�� �J� f7LKKM
l<<
K
<M	�J=��
	L� f7�� X=IKMZ-!V<	�~��	� f7��	T.7f7�XX
	Lf7�X	�f7�X��]J�]�g1*$Ju �  � IM*K$-u �  � IM+K%-u �   � IM1K+-u �&  � IM�����*u$-u �   IM+u%-u u    IMySg��vrv�<\g
	 �  &   X /  X /  Z 	 V��6�wX-.=$�h�~�!- =J)�f\"� ���������!�!�� f�X\0#tu%�#� � � � � � �#�!��'�'� �z�!K^�J
J	Y&4I&K4;�� q<K.  u� � 
J ltX �.%pK4J
J	Y&4I&K4;��  u� � L
Jy�K. �|��xo�KK>Z�?IKK�Z.J=�u
	Y/t�������XX� /W�wrKK>Z�f?IKK�Z��
	�	�Z"<u8"t�������XX�r�xy�/.u<
tv/JIJ<?f-LȂ H X>[
/ X�/�	LF2 X�oJXfo X��/-gJ;J�Xy���X
�wlKvqgN�gZ�v,ZX ...XkJX  ...�t�%4V*%�� : < X�
f��X$E	.Z �Y	ft.�|�
�
�wst�
��
�Y
�\�_�w@J	L	X	u i< �
 ��]�Xk	�	u$	u��
� <�<�� -[A	E�	
X	u uJ �
 ��	u�	u��	�w.�K
=
;	�X\
[vHL	X. �	 0 R<J:X�...	m��	0 W < JZ
=
;	�X	(J��	pf�	>uX�X�<��	� f � �	 0���[�$f,J$JX@1J��]�2`v6$I-J=;KI=Y
�\'t
<	P4qJ	gJ� 		=I	=efg
�o.u MJYK ��v�y�#tu2rg�pt-�tg�p
0W
� �j�vrvU/.  "Y��3.t@?
U�!>��!	�<\ <X�v.w�x<��x <��x<�t�x<�<�x �t<
�x<K
K�l	
�M	:���0V>:0�x
�K
K<Ml
	=��
�xtM�J	�x.��
FJ�
�x.�Jy�x
wl
	=��
�xtM��x �J	�x.��Jy�}���=u. X �{J ���z���T�+�z��z�� ֐�$�Cy<
<	i	K2 Xf J�
	iJ�"�zX�J g3 I / �zJ 3 ��" �y<	�<X.Kf��z
�	�wg�Jt ��!�f,�	XCy<<iK4 cf J	�hJ�"<�<O
: �-�:s>��z��z�~��<��{�N��~J��L�~
�	�%D�uf�s	K%_y�	M%	�	Z"tf<<	?"�="�5I�$YK$sK9:�	<�}J:��	<"$<"<$J	L�$�
	�:<J>JJ><<><XK,�&�X�~�����|�6�}� �6J��|J<[	�~J�����	?sK IK ;=
�	k"	M�}�h(IJXi<X��z���x�XM�xJ	���z��z<	�J�y�X	�G	��y�	�-��z��z�~��� �
X	L>JJ><J><JK,t&�Q
�J<$YK$W=$-K9:	3t"$<"<$J	ZY$�E�f�5
��otw)�]X>�~X<8xX>`��>�}Xf�8�~X�0�	Mf[B�%z<J�
$f�}'�	Z�[Br^ Jg.�K�}
�		�	K�}��f��z��zt��0YL6dIKL[9X��<I]o.2X-<���z�t�<�z��z�~����N< p t	��yf�j�yJi	�~J�	�~.X���,XL��y�����~�z�JsX�z<��\rfI�z<�Jf�z�����z<>�X9�}�<�~<:��%H>TZ%LXJ��|. J/.�
5KX�~.!�JPJ/(�}	��}�X�}
��<��f��.J�X.J��.J�X	X�}!�J	L�}X��}�~�	J<Xgf3�	�JXgf� v�-&<J&JJ^/IuK��-&<J&JJ^/IuK��Jl��0 J� F_�	�Jtg���J#� �P. J�� J�sJ	�~Jtg� ���~J#��O.Ju~	�~JXg
<�T^zP?tX���X �6� � U�J(<tJJ�
fg	 u�o�X
P�� ��
z<Y
X
�����XY\(KHOUME=Z
<	Y#cJXX<�X�� ��L;KJ)J>)dKKIKZK.f.
��<X� t�ZJ&X��K� X .f� f�~�#�~�J��w	Ji���~<�<[�1v<C-M_bL�-NXoX�Kf..J%`fg�
�<�{��s.pt�qt�|p.�t<JJJ! X\�~"KYYU/==9=;>KH=KG/===�w
K
K<wl
M	��.f� <'.��<� �	
T	��
�	j"=	s�
	$�F	�9	[h��X ..�t(��9�]##J��y+��XX�~��w�/	Cx<=;=;=
�w<K
J�l
M	���	.�<�wJ.�V�wX
<K
w	���wJJ�,L:>�w
<K
<M	�J�J<
YH��
YH��J
uH��J
uH��
&s
�L�� 	x���Jf� <�	
UF�	�
U	f|
�	��	2�
3  	��"=	s�
) �d��Xf
�{Xv#
��YJ<<
.�ZuIL$t1Xm..:u.s.KM�	�	w uf 	<v�
� -u v v 	t<%�	I�~���~���~t�<.�~1=AG1q�u1tv�u�
 �s.6 � �0Jt�! < X�~��E�N�v�		.�I�J�g�uX .p���
�s�.t�<t �� f�	�KIgh-;-3q:=>9YYt�du�u�`uu�. �� <& �8�tJn%#Is�Z u v+�zBz.Pz<�ff�_	��r.=;<�<�rJ�1�rX=;=�<>�r<<�>1�r<<�<9�rf�.a@IK0?zJ0H=>?0vxt:Y>y.Y��
lxtu�u����q���uuXt<Y�Z[ ztu vwk#=Iq%�J��s�y.u<
JU=x.J8YGK:.Jt N XX>
WY
	/<J��`���=:Xg;K�[
	_KI	K  J % � �   � �  �  K X   J	\�=I	KX

	x
LVL
	2JJ_ 	��
�SA
O	/���	�J�t 	��E      � ��\J!�NX .� XLX .+��oX
��Y
J  .	F�  *X 	��E     �=�t 	��E     8	EM�-cJ<cJ-IJK		=Ltt(X
v_�+JKR��4JJ�
X	Y&4I&K4;�t	���� XJ=X<.[�Yd�.�< VJX).
�oXYuXLj�t<`
�o
	���
�q��M$�t
�p�$<X
�p�$X
�p..w��J-cJuIK	KI	=LtJX
�p�6�
�pX�J-cJ<cJ-IJcJK		=L<JJX
�p�6�
�pX�J-cJ<cJ-IJcJK		=L<�
�p
X	�...� �} J�t 	`�E      �.�NX/� �KQ�[X0J-pJ<-oJJK	<	=LttJ$�	�rX�uY
J  .	p�  *X 	@�E     �p� �<� X� t#�g�f�t=<<�<� .T<`</K
� TJf<K-
w	�Q1XJO=-w<
?	�Bz.B
<Y�I?H*JW<M&<ZJ&J�f�?��[Xw-y;R(�<;(=<:�X�3<	�J^<
".K\
#<<M	�JZ
	�$J<�#�fN?cK[�x-KCxf(	<I�e=:WX�	$J$<<�L�11<	�	�	[	$x+=Cx<Rx<D&�J;&=J8�X��r%..s%fsJ<K?<!L�JHX>	fX�2�J
cJ. �bJ��v[Bz<�S�
RK  .o.1K <��K	s<u<	Z	�	�(Yt]�-?�Y#�?��.�K�u�<cY �
 � �9 Wv�f�Z�	�X�~
rJ��Yb
X��f	���rvX�vL�o�	c��	�X	[	�s��	�X	�	���~����J��}
��
X�Z��
��
JU	��
 �X� �	Q�	�X	�	�[�	�	�	�	�X	�	�	�	�	�a��}
��
X�	��f	���
�J�� �Y�~
X�L� ��,4f�X�i�f����}�L��f��~f���	")�	K�f�<�	�}
V	L	�Cy�JL�QU~	Z	�	�X	�	�	�	�	�	�X[�
��� �
��z��Bz���Z���Y��V/uJm=,�	@JX�	Y�	K�$,PX.y.u��]1xJ!xJAJ�<˯4seu�qt-�tg�q
0W
� �j"Vv"u"�  .�o�Zm0LUK6LHL`�CJ�<?Y,Jh�J�� Y,JfIX	�<X.Kf
� �u�Lj�t<`
�o
	J����X� M
�p
X	g1X<J� ..X 	��E     LJkh	�Jtg�� L:LtX	�Jtg��6.JJ�Jy<yv>v<4X��
�~���}4XcXs�
�J�}tL����{��Y
��}�|���g��|���������|���.�w���������|���������|���Z�yXF�#o�����w���t�yJ&�tTu&M�yJ�tw��{t�}t�~�������yu���yu���yu��v&��{��}��%vzt�%�z.�%v;%u,%vQ%y�7�%�
�}J%�X
�}X#��%�{.#�Xy�{
��}t�
��~�
�~�,�X � �{   � �   X t <M=XN
�
tJ�K� J��K�
�|m���
OE��|J��
���~.
���}<�s�}W
����~	�{
�	��
	Z u+ WN);	 ) �+ :	
." t/ f f .
t
�
Xl	�.<���kJ�	�{
�	��{�<	� � 	���	�x�J��q�w����X���h���X���h���X���h���X���hZ?������lf7 ��}���f�j����jJ��<�#A7.AX	�~�%�kJ#��.=0�� �l	�J�X<><<A;=Y;KYCx<=[�KZ��h�5�yJX��B%�kJ#��.=0�.f��>;=Y;=ZBx<KZ�LL��h���<><<�A�k#�<���lzJZHv[qw.wYJx<X��;�Y;�Y;KY;KYBy<KZ�L>�up�	W	�k#��- X	�V	�	��t	0�qt�Z��"	�l#��	�V	�	�	�Zd�	v�	���lJ#�� �lX0 �		�5	M���mU�t�mJ��~��?�t�l���u�~J��u����~�X����l���l�\XJ��q��3J.tfO&�t@� ��X!�
f�	�hJ	�	�X����	 �   >��n��X�mJ� ����n���m>���6�nJ �y�����n<[	�~����J�<
�'�f�'X�L�s �yJ#���y<.�?��ttt 2  �* t J < X t��Mt��Y�zJ#�.�J �  � : v+  @ [ q w  . w yX J �(�{J	�J��	�z#��- X	�V	�	�	�r.	vQ���z�		� . XS2��z�		� . X �* `  3�%�jJ#�� C y<Q=;KQfq<Z,u�=XK;KY-K	XwJLy.�XZu<uP�t�e�rfY-�XK;KY-K	�w<>����q	��yJ�	�~��	�~.X���,���y<�L�Z% � �Z.X@UY<
�~��
�~LV�g�!tfL�
t	�4<<�	���N�y#���y�<�0fY;�Y;�Y;KY;KY;KZ�L><�up.����m	���s%�x�t�t���l	�J�j.�
XX��<���g=�i �O��	�qu�y.�	�~��	�~.XgX.�,���	��x���- ���l"�<��j�<	 �@ 	 � �@ 	 ��t
�}LVvg�"t'/";JIL"JL�	VX	���k �|!�!X.!J=�Z&�E�iX�tX�����l��l	�JZ.0X�jg<��{fX����g=�i�JJJ<�/]73�
�o&!<J��X���s�0���\[�[���X�x�����i��<��iJJJ��<��i��J��i��<�&=<.lX&0.I=.�l]7X��ot�.X�t!��6 � J��f��m�J�s.�:v[qw.w[�{X��}#�}X�J#�}f�J#�}t�JM�}�=L>vwcM[?.f	u<JJ�~XJ.�
�~<K
1	�J�;�B�~�J#� �^t=t�J�ft�	�f<t�
/�>XX+K>;<	u&J��������n#���� -M <.0<X.��#�i	��m�.<[	��	�	��{�	� �m� # + ����dl�X0XuZ�vX=��
�q���`
�q8Z�8>���!-=�'
�q8Z�8>�������1��x�ւXX��
�u"��W=YW=\T>�xX�J#� ���<�x<�t�xf���xX�J#� ����x<�t�xt� � � ' ����uXv) �v< � X X X X����XY�{���X<�sJ�����*X;th�X/D�|�<X/ZO�|.�<f�|�0�|X4���VX�!X=!X=!X/!Zf..NfiZE ��@ts�\�X>E ��1WY1-uJ0�}X���XX�$X=$Z�.<Wt_�#X=#Z�r
.K
1	����&X/&Z...X`�$X/$Z..X\#[#Gw�Z2 �+ <B ;�$7X.$��X�X#�	�2$�Z>f#�r�$���< K @,f$�,b@ /#  � J �rX    . <D �
 �sJ K 
  1	  � J! � < I _ �s   �J #  � ��t=tJ �.�<<�0�~X4������tJX�
�� &8f<g&<���X�|�> � L* / <* u/ ; = - u/  � ��0�P�-�����X�|�2�<XJi��s��� X���s���r<0*�X�r����X�. t X=���Y�0WX2(��X�&7�h�X/@�}�<X/ZK�}.�<f�}X_�X=X/Zf.Xe��.�h�Z�$��z�+)�+X).+JK+)X+JZuZ�>���X�u��~	�&]v�L&�&X0#X=#X=#]#}MmX��9�?-t��'K 'S�= �Y �=l�tX� X[#/-	#w<h-#y<�#K#�-%X�X-� J%J�-,\%T-X,M%U?,I�,u,�5�X�"!��� J �  <3 W5 ; < . < ��z%�Zd0%X<. eXF s�9�?� X�������X
'�z���
�zJ�'>rv<JY8J<�J�5	X5w<K"I�JY"<6Lu"`"x�ZX?� J$`
'�zX��J
�z��'>rv J Y8J<��&4X[&94J�&4JX0����Z�o
.K
1	����Zf��X�� X�m.�7<= �7 . < .=-D�"X=\.X�z�w.tK"�"Z*..X     0 % : X	t"Y;="[*fWtL � Z*.X:�e0�0Z!tD�w<���uX�X>Y<X�w��hX�Z.�fX�Z16X.J��X <X�X0�o�J�~JJ#J���;[>��P<1�:	X2)n<)JJ<KulfZ
	Z	K:>J<M/
L	K..N.<.)	�~JXYfXX�X
�t�U� X�
tM�)yJu `Jypv�#�l<�X� Jm�Z�X#� t���%v
f��� 
�Lu
 J7 X	wL<utg�����=@agj�~� 
	L�}J(�X��)<�"tJ�4�~�zt�<��~�t��}xt��x
��~�uih
��~
v�*
���~Z=j#
@��
��!l\!w��!y�K�L
L	�w
$
��~t�
� ��h
�
t	�#	}�}f:��.�
� �t
� J��
'J<	���!�|�::�<j��tJ
u
WX�}����}e.t
�J�|X��w�|
��
�1qi���|
��|
4�t��|
�4��|
�4��|
�4��|
��|1f	.5.f5rt0/e	�		$.ej'R�J�	irv9.<	�
C	y<g+i
<4|
�	$.c	v.�
7Ct�KCt<�J� 
�L	�~֐��	g-.<	K.;	M:g	+;i
.4,
<�"h,9ifaJ(X�<J�
G1
	.flxfhlG�)?>��'/,qt	JX%IJJ� ft'�t���t	$�~%�+JM�Z
�	m�~%�wtJ	JwfX� �wt�
�t#���}t	�
�
\
�
�t��}�<M	�{�
�
��}tgft���~f	ZXi�:>��'/1t�	JX���LX�'%U.JJX�7�t
PD(�XX<
�XL
V�vH>>
	Y9t��� J�J�Lu� �t�<
�<�f�	�� <	n�}	���}f:�t�
	�vL�	�vJ<��v�~<
�%�t� z.���
� tJ�~X	t
�XX<�~	?	�+t.��b�	Ow	M	�	�J
�~��	��}fV��.	D�}:�	��.
TA�~�?Y�=��=��=��=��(&s�&^
"�&]f
#f#iJ
fn<#p
�u
w	�(TJ=��'Bet#b<h
K
1	�%`J:����	�{�
�g�	.X	,t�X
�}
 �
     �      /home/computerfido/Desktop/freetypetest2/freetype/src/psnames /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal/services  psmodule.c   pstables.h   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   svpscmap.h   psmodule.h   fterrors.h   string.h   stdlib.h   ftmemory.h     	�/F     �/-/-g\Jx
`03p�
0.t��	K>!:�<0#JL
.#qJ�
[
	KJjZ<#<JL
.PZ
M
	�JhX+\�L�'72%�/	�%	/.	L<t�.	�/o<	Z<%..=I	=<	^	hY<	LpX
N
>	L	Ky ;	=t=f<`XK=Y..XX��$g3�2.$��11�XX 	`1F     �u K	WA)J/+6\�	�v
g
]
s�)J/+6\�	�v
g
]
s..� X/�.J
`	�=
�	L
W9tJ
	Z)W. Xv(XX (t
HX	/Jp� �g�JvL	�<�	v�t	9<��	vf�%JX�t�_�< � J �V�	 ,  �HJ
J	�XX��`X[ �f I6XMF7<W	4J	KZ K[	M	 [  <- m J J . m <	.	Z���`. e
��	fMF	4J	KZ K�	P	 �  <- j J . jX	J	L�.1G|u�uXXuXJ<u.Xu<[/X
tJ
��	�	�X���
�Hf� �	�XY�% k < X��	J]gKH== wJf<L
	
�!t	�\�tJ.	�~���g� �<J� Z��Mt
JHf9=I=	J�4>IK<	�2Xo	,�!��� �   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftsystem.c   stdio.h   stddef.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   stdlib.h   fterrors.h     	�6F     � =JZ � � u � Xbmy
QLi�Y -�.<Xi�~�<X 	P7F     5<X 	`7F     e<<X 	p7F     � ��y RP yX� u � � �X=S`�#�K_� Ky.��X p �sJX  ZX&X<N�Zu����X  �   �  �      /home/computerfido/Desktop/freetypetest2/freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/freetypetest2/build /home/computerfido/Desktop/freetypetest2/freetype/include/freetype /home/computerfido/Desktop/freetypetest2/freetype/include/freetype/internal  ftbitmap.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftmemory.h   <built-in>    fterrors.h     	�8F     "Y/t���#�=0;=;KIK0L�$.a>yJ=.
XL�t4.<XL
�JYIK
	�(b	Y/<fJ	>� > � : X >  	 7 J
J�J.B�u
	YZ:.	[<�XJ
J ��J� X�.� X^��X	��(���OJ:�</��8KK3X	f=Y3f	t>#WXlf	<#H$?#+.$2!8M=A!wJ	>:LJ/	�.X�	�; � L	��,	�Z<Jf. >  w/  = ; K  Z   wJ ��K1f 0  J =  J <	 h < f;KX �~�J<	�:	��<��>�}lz.=X.Ygf2oKKHuu<r=<>q.J<..�LE�<=J<	pJ��:	��<Xf� �  	< I/ E + 1/  ? 9 K/  / ; = = : = ; K     u�<fJ=J<	[J�h:T	K	L � � >  J =  J	 7 J �A:	��<Xf �  < I/ wJ + 1/  C y< K/  ^ z< u/  X u/  X u/  X u/  / - = ; = ; K     q �J<.J=J<	VJ�; f �8<M �  0 I - g   �� <M Z  0 I ; u   �� �}J�X�}.�X�~�<�� �2<>�p. X� pX; se.	 ��z�J�zJ�<�z< �Y
Mgs�NX6[yX
J<JX�,w x�`u<�{�� ��H(ZJ �( J> I�n<.?j.
.m<
f[k.J
+K
L
h�t<� .Ztu% d J J �0XJ.	�	� u  f	 I �  z < 
X	 % �< J% . <� �uh/	���}�JX�}X�	��}��	Y	M�L��~J:�J�~J�.�~J�<�~X;/;=>��ci�~�%�gf��$I$�JM
	�7?dY7:M9	=��*.8<	<<hv=LY�.S%�ufX�J�~X��J�~�/;=�%�ufX���~J:�J�~J�.�~J�<�~X;/;=>IgKX��2y�~'�
<�J�f�*�
X�	*��	;Y�uyX
f�9M�J� 2�"	�D�� t+rt	�\	F��<,<Xf,<<<�</$J0<<" e�	 <�htMY X�tJJX\	�=<+<	J<�X<.J� �Xw�YJ��X	"�	;YJ�yX�
m �    '   �       src/gfx/sse2.asm      	@RF     !>==ALLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""�� �    �   �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include  syscall.c   types.h   stdint.h    g 	�UF     �� �   7  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../sysdeps/lemon/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../options/ansi/include/bits/ansi ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   lemon.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   pid_t.h   time_t.h   types.h   stdint.h   debug.hpp 	  type_traits   sysdeps.hpp 	  string.hpp   <built-in>     2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	;VF     

�(5>� �
�J
�	%tY
uY00
�Y$0
�'>K�2
�	'
u=:0
0	&�
�uY2&�,�!  # +�� # 6���?	KY1L  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�ZF     � �/  	�ZF     � 	 	[F     
�/K 	 	,[F     
�/K 	 	T[F     !�t��K  	�[F     � �  	�[F     � �  	�[F     -�1%  	�[F     ��2  	\F     ��0  	T\F     � �/  	z\F     �=/  	�\F     �/4  	�\F     0��  � .��gt��������y�	X  	�]F     �	/fY%* � � � .�%  	[^F     � �3  	�^F     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	O`F     �� J J . K  	x`F     &  � .��gt���J����� 8     �      ../options/internal/generic ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/include/mlibc  debug.cpp   type_traits   optional.hpp   string.hpp   logging.hpp   debug.hpp   <built-in>    formatting.hpp    1 	,aF     
��2L�� �	   {  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/mlibc  new   formatting.hpp   ensure.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   type_traits   string.hpp   debug.hpp   <built-in>     2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	maF     &�,�!  # +�� # 6���?&�+�!  # +�� # 6���  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�ZF     � �/  	�ZF     � 	 	[F     
�/K 	 	,[F     
�/K 	 	T[F     !�t��K  	�cF     � �/  	�cF     � 	 	�cF     
�/K 	 	�cF     
�/K 	 	dF     !�t��K  	�[F     � �  	�[F     � �  	�[F     -�1%  	�[F     ��2  	\F     ��0  	T\F     � �/  	:dF     -�1%  	ndF     ��2  	�dF     ��0  	�dF     � �/  	z\F     �=/  	�\F     �/4  	eF     �=/  	FeF     �/4  	�\F     0��  � .��gt��������y�	X  	�]F     �	/fY%* � � � .�%  	�eF     0��  � .��gt��������y�	X  	afF     �	/fY%* � � � .�%  	[^F     � �3  	�fF     � �3  	�^F     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	RgF     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	O`F     �� J J . K  	x`F     &  � .��gt���J�����  	�hF     &  � .��gt���J����� �   �   �      ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  essential.cpp   stddef.h    . 	�iF     �� � � � W	vKN0�� � � � � < -	vK90��� � � � � < -w �. �5 � � �5 � < -	wK0	�� � ! W	vK e    :   �      ../options/internal/x86_64  setjmp.S     	*kF     =KKKKLYKKLu%=KKKKL=K �/   �  �      ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  random.hpp   new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   stdlib-stubs.cpp   optional.hpp   strtofp.hpp   logging.hpp   utility.hpp   mutex.hpp   errno.h   types.h   stdint.h   stddef.h   locale_t.h 	  stdlib.h   string.hpp   type_traits   debug.hpp   charcode.hpp   mbstate.h   <built-in>      	�}F     �  	�}F     
�� � �# u( �+ <4 �9 �< <> �- < .H f �F � . � �"  	l~F     ���� t � �, t/ f1 � X Y �  � X0 .3 f& f J �k t � �, t/ f1 � X Y �& �! X6 .9 f, f J �k�,t.fXY!�X1.4f'f.	�����f=fX=fX=f
>= 2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	<�F     5//
�!  	r�F     �F  	ÀF     ��  	րF     �6J7tXK�  	�F     �Ju ! 	{kF     �X�/�Y/�Y%/�YE/�+t�D/�/K/$�0��M/2	tKt�X	LU0$ ��KtK	K[g f�#X\�	tKt J tK<$�X	xzX	.u� f t .J!S/0YX00��	w�<g��1g	u�<	�g�<g f  fgt  J t
K�gYvg f t X&=	f&/$f	 =�u�XKg�X�� J t X?�# f J4 f, J> f��u! r�<g]>	 g	�gtKu f � JuK]/0Y2-L<�Y0���=>�?X��4>��	u
g	v L)/�K
uu	�K3K ��	YY'/���Y���� ����/�	��
��
�<uA���gg	
g�%�i �	�Y/0v �*�&�	tK �+�'�
tK<X
N�� � �
 � g � � < / � co  ��>���#��"��	t=�	=K&/�2��-�#6�,�6�,K)�,�L�A;�#�&g�J KQu��AX�� �� �� �� ���t<	/Y&/�A�#=�//�3�)�3.L;v+�Jg
�2i#�Jg�J
�K	�.
g LX0=�"!�f��� ���Y5�?����!>!%�Z!�fK����	�K'0�'��!�fK��  +��	�K;0KJ
g��t
Yu7�".!
uw <�	�Y[v=�� f�}���<J  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/ 	 	.�F     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	ZY 	 	{�F     	�t�t J tKZt J! � <1 J6 �( <K�� K&�J� t � J K��X�!Y
�J�S6����<# J( � <8 J= �/ <K��YX"L)���S	s.<
z<'u�g	LY 	 	ǅF     	�t�t J tKZt J! � <1 J6 �( <K�Z K&�J� t � J K��X�!�
�f�S6����<# J( � <8 J= �/ <K��YX"L)����	s.<
z<'u�g	�= 
 	�cF     � �/ 
 	�cF     � 
	 	�cF     
�/K 
	 	dF     !�t��K 
	 	�F     
�/K  	�F     � v
�<g�ut�t!J�u �&�)J�  	��F     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	��F     ��Y  	��F     �
�t�  	܉F     �
=*t/ 
 	�F     �� X J . K  	�[F     � �  	�[F     � � 
 	:dF     -�1%  	ndF     ��2 
 	�dF     � �/  	7�F     ��2  	|�F     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	�F     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	��F     �Nu�u
/� ���g�u � .
�f�*�$t��	�gu	�g
0� � � .� � � .��g	hgu%u	�/
0_J #�  	eF     �=/  	��F     �=/S  	4�F     $�/�  	f�F     '��K�  	��F     ��=��'g !3�(�	<(g" � � � .�	jY  	V�F     ����uf	u.u
fy.�"k  	�F     7� � � .���  	b�F     ���  	x�F     �	���# f- �+ � < f t Y  	F     ���fK/[���fKg0#�fKg0t�X  	��F     ����uf	u.u
fy.�"k  	r�F     � ��uu���
0K  	ʙF     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�F     ���fK/[���fKg0#�fKg0t�X  	�F     1� � � .���  	N�F     � � � .�t�J/	PK 
 	�eF     0��  � .��gt��������y�	X  	�F     �	=fY&* � � � .�&  	��F     �  �u  	��F     � �(�K  	��F     � �)�K  	؝F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	9�F     � �/�K  	X�F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�F     �  �u  	��F     � � � � .��/1  	`�F     ����  	��F     � �(�K  	��F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	ݤF     � �)�K  	��F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	4�F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	��F     � �/�K  	��F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	@�F     �6h:J  	��F     � � � � .��/1  	�F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	F�F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	~�F     �3g71  	ɮF     � �4  	 �F     7��  	6�F     � �-�K  	T�F     � �uu�(<g  	��F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	I�F     <�*�=  	f�F     ���u�<L�0#  	��F     ���  	εF     ���  	�F     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	D�F     7��  	Z�F     ���u�<L�0#  	��F     � �-�K  	��F     � �uu�(<g  	�F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��F     <�*�=  	ҿF     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	(�F     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��F     � �uu�(<g  	�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	B�F     &
�Y  	Q�F     &
�Y  	`�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	 �F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��F     � �uu�(<g 
 	O`F     �� J J . K 
 	�hF     &  � .��gt���J����� g	   
  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/ansi/include ../options/internal/include/bits ../options/internal/include ../subprojects/cxxshim/stage2/include  formatting.hpp   charcode.hpp   charset.hpp   ctype-stubs.cpp   optional.hpp   string.hpp   logging.hpp   stddef.h   wctype.h   types.h   stdint.h   mbstate.h   type_traits   debug.hpp   <built-in>      	&YF     2&�*M  	ZF     1�  	��F     /KJ	=J J �K�)�&�)�(K%�(�K$0�JgZ �� �� Y - 	��F     !1u" f1 f? f1 � t 
Y  	��F     #���
g+u.J =0#���
g+u.J =0#���
g,u/J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g+u.J =0#���
g"u%� =0#���
gu� =4)��t
g+u.J =0)��t
g+u.J =0)��t
g,u/J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g+u.J =0)��t
g"u%� =!.!�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 J�6 Ju�/�5 T��	� Y 0��#���
g+Y K0#���
g+Y K4���  	6ZF     �<  	ZZF     7�  	�F     �h��K;0  	l�F     *��JYu � �gt�$J�K r
wY  	�cF     � �/  	�cF     � 	 	�cF     
�/K 	 	dF     !�t��K  	�[F     � �  	�[F     � �  	:dF     -�1%  	ndF     ��2  	�dF     � �/  	eF     �=/  	�eF     0��  � .��gt��������y�	X �)   O  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   environment.cpp   optional.hpp   string.hpp   logging.hpp   vector.hpp   utility   mutex.hpp   utility.hpp   errno.h   stdio.h   stddef.h   types.h   stdint.h   type_traits   debug.hpp   <built-in>      	r�F     �F  	ÀF     ��  	րF     �6J7tXK�  	�F     �Ju 2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	<�F     5//
�!  	(�F     ��#f 2 	��F     % �"�#JK� � �" �1  	 7: � ���K vf
�u4�CK �B JC X	8u0������ � � � � �v�
�w�
 Q0)� #�gu�J.[ ��J�=�
��/��� #�g t � .�   < t X J)��4��w
�� ��*
u!�"J!� t%�,�/� = 0�/�u�Y	5Y@v"����!�0 57��	�K� 2� ��Y	D Y ��Y	&Y  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�F     �h��K;0 	 	R�F     6" �  �gt�Y dxu 	 	�cF     � �/ 	 	�cF     � 		 	�cF     
�/K  	��F     
�u 	 	��F     &
�� 		 	��F     
�/K 		 	dF     !�t��K  	 �F     � = t � .�1t#  	l�F     *��JYu � �gt�$J�K r
wY 
 	r�F     �N.R$ 
 	��F     �� � � fvJ�� 
 	�F     � 
�� 
 	�F     � � � � fv� 
 	L�F     ���/��J<��
=K 
 	��F     ��2/���J<�u
=K 
 	J�F     � 
���= 
 	l�F     � 
����= 
	 	��F     � 
�� ! 	��F     0�u  	��F     ��
K�
u�u 
 	�F     ��="�!�t	�K  	�[F     � �  	�[F     � � 	 	:dF     -�1%  	ndF     ��2  	M�F     ��6 	 	�dF     � �/  	��F     �#f ! 	��F     0�u  	�F     � v
�<g�ut�t!J�u �&�)J�  	��F     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	��F     ��Y 
 	��F     ��	��� � �# g, �" � � � ew � � fvJ���t�   	eF     �=/  	��F     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	|�F     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�    	��F     �
�t� 	 	�eF     0��  � .��gt��������y�	X 	 	�hF     &  � .��gt���J�����  	��F     �=7  	4�F     $�/�  	f�F     '��K�  	��F     ��=��'g !3�(�	<(g" � � � .�	jY  	V�F     ����uf	u.u
fy.�"k  	�F     7� � � .���  	b�F     ���  	x�F     �	���# f- �+ � < f t Y  	F     ���fK/[���fKg0#�fKg0t�X  	�F     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	FeF     �/4  	��F     �  �u  	�F     1� � � .���  	��F     � �(�K  	��F     � �)�K  	؝F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	9�F     � �/�K  	X�F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�F     �  �u  	��F     � � � � .��/1  	`�F     ����  	��F     � �(�K  	��F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	ݤF     � �)�K  	��F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	��F     ����uf	u.u
fy.�"k  	r�F     � ��uu���
0K  	ʙF     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�F     ���fK/[���fKg0#�fKg0t�X  	N�F     � � � .�t�J/	PK  	afF     �	/fY%* � � � .�%  	 �F     7��  	6�F     � �-�K  	T�F     � �uu�(<g  	��F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	I�F     <�*�=  	f�F     ���u�<L�0#  	��F     ���  	εF     ���  	�F     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	D�F     7��  	��F     � �/�K  	Z�F     ���u�<L�0#  	��F     � �-�K  	4�F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	��F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	@�F     �6h:J  	��F     � � � � .��/1  	�F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	F�F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	~�F     �3g71  	�fF     � �3  	��F     � �uu�(<g  	�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	B�F     &
�Y  	Q�F     &
�Y  	��F     <�*�=  	��F     � �uu�(<g  	`�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	 �F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	�F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	ҿF     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	RgF     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��F     � �uu�(<g 
 	O`F     �� J J . K D    >   �      ../options/ansi/generic  errno-stubs.cpp    �5   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../options/ansi/generic ../options/ansi/include/mlibc ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/posix/include/bits/posix  new   formatting.hpp   rbtree.hpp   slab.hpp   allocator.hpp   file-io.cpp   optional.hpp   list.hpp   logging.hpp   utility.hpp   allocation.hpp   utility   intrusive.hpp   mutex.hpp   file-io.hpp   errno.h   stddef.h   types.h   stdint.h 	  ssize_t.h 
  stdio.h   off_t.h 
  type_traits   string.hpp   debug.hpp   <built-in>     2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	r�F     �F  	ÀF     ��  	րF     �6J7tXK�  	�F     �Ju  	$�F     /V�D��������!�/> K��Y�Y���Y��-��Yv<
����Z��"MB' ���XK!��0��g��tY�
�� J �Y�Y������ g� g�;�)g��tY���!$ ��/�-�fBJ� ��JY�	� YT>' ���XK!��� �1��g�� ��
���Y g� g�� J �Y�Y��� ��(�&�:�X:<wK�,Y�u�
tuM ���	t��<"��+Y�3��<'�0��7��<�����-��$�:��<��g�XKw	 Y#> ��
����<g5L� J�	�Y0������L���Y�g[�
gY	�Y00.���
g)Z#�;<3� <t	u Y30/�
g�&g �8<0�<6��<�/[ f f1��<g/^	� Y!>�t
K"v�f
gY �	�Y$>�t
K v�!<XKu �	�Y">��
g���
Y�tVZ��3<��g��� �� J���V�3�A��f&�$�J.g/Z ��gxf	XY >! 
g����/<�9��g��5�?���
Z	v Y0��
g�tY J� J���	�Y*0� ���[$�g�$B$/(/L	�u>!��Y�Y��<
g	YY0>�"	g
�u	�
�v >30��	�
��<	g
�u	�
�v�&X��ZJ>v�
gY	� YQ>v�
gY	� YC>g�
g	YY
<�L" 1 � / �g�Y� � �]&D� t � X K �0��&-<E�7�S�&<S�&<S�1U��"<��K
g���K
g�	v��6�7�?�K����	���K�	�K�	�
Ku��7�? K���v�X�	u
g5v'�TY X f Y&6E�7�S�&<S�&<S�(z�u�Y��5�'�TY X fY0� t � X K u � XKu��XKu	�=50/ t � X K �	ug	vY0� t � X L X	ug	� K&0� t � X K � X
K	uY/��C0h t � X K"g<
�g�"g<
ugv"g<
ug	�K	wY0� t � X K Y /$>� t � X K	 = = 0� t � X K ��{<�Kv.�*K3�*<	�3�	J3�=��Kv.�*K3�*<	�3�	J3�=��� ��{���X�X�X��&<J  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�G     � "�&f  	G     3�7�  	,G     �  � � .(�� � � .� � � .� � � .��Y���.K�f>�.Kg 	 	�cF     � �/ 	 	�cF     � 		 	�cF     
�/K 		 	dF     !�t��K  	�F     � v
�<g�ut�t!J�u �&�)J�  	��F     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	��F     ��Y  	�G     � � � � .�g  	*G     � � � .� � � .1�!.�,K.�JY  � .�� 0 � .�J�Nu � � .�J�� / � .#�. ��.? � � .�.u.�.
LK 	 	�ZF     � �/ 	 	�ZF     � 		 	[F     
�/K 		 	T[F     !�t��K 

 		G     �� X J . K 

 	�F     �� X J . K 		 	4G     
�/K  	��F     �
�t�  	\G     �(�%  	�G     ��K  	�G     ;�.=  	�G     ?��uK  	G     4�u 		 	 G     
/K  	JG     �v/�#  	�G     �K  	�[F     � �  	�[F     � �  	�G     
�K  	�G     $��� ! 	�G     0�u  	�G     1�� 	 	:dF     -�1%  	ndF     ��2 	 	�dF     � �/  	|�F     �� ���gu � .
�f� � � .�g��.fJ<��<t�t��\ � � .��� X � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY�p�R"�   	 	�[F     -�1%  	�[F     ��2 	 	T\F     � �/  	
G     ��0  	�F     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
  	NG     8�t� 	 	pG     ,� ��  	�G     ��4  	�G     �=� 
 	G     !��  	4G     ��  	eF     �=/  	4�F     $�/�  	f�F     '��K�  	��F     ��=��'g !3�(�	<(g" � � � .�	jY  	V�F     ����uf	u.u
fy.�"k  	�F     7� � � .���  	b�F     ���  	x�F     �	���# f- �+ � < f t Y  	F     ���fK/[���fKg0#�fKg0t�X  	z\F     �=/  	NG     �/4  	��F     ����uf	u.u
fy.�"k  	r�F     � ��uu���
0K  	ʙF     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�F     ���fK/[���fKg0#�fKg0t�X  	�F     1� � � .���  	N�F     � � � .�t�J/	PK  	�G     �K��/[4��K � � .�t)�#t� # � .'�J��� � � .�JtK � � t X J � 	.��u�gg� X, �6 � JY s�k�$  
 	�G     �K 	 	�eF     0��  � .��gt��������y�	X  	��F     �  �u  	��F     � �(�K  	��F     � �)�K  	؝F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	9�F     � �/�K  	X�F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�F     �  �u  	��F     � � � � .��/1  	`�F     ����  	��F     � �(�K  	��F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	ݤF     � �)�K  	��F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1 	 	�\F     0��  � .��gt��������y�	X  	�G     �	/fY%* � � � .�%  	4�F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	��F     � �/�K  	��F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	@�F     �6h:J  	��F     � � � � .��/1  	�F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	F�F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	~�F     �3g71  	 �F     7��  	6�F     � �-�K  	T�F     � �uu�(<g  	��F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	I�F     <�*�=  	f�F     ���u�<L�0#  	��F     ���  	εF     ���  	�F     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	D�F     7��  	Z�F     ���u�<L�0#  	��F     � �-�K  	~G     � �Fg	<Y3,3  	��F     � �uu�(<g  	�F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��F     <�*�=  	ҿF     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	��F     � �uu�(<g  	�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	B�F     &
�Y  	Q�F     &
�Y  	`�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	 �F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	RgF     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	G     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��F     � �uu�(<g 

 	O`F     �� J J . K 	 	�hF     &  � .��gt���J�����  	�G     � �!  	�G     � � �~   �  �      ../subprojects/frigg/include/frg ../options/internal/include/mlibc ../subprojects/cxxshim/stage2/include ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix ../options/internal/include/bits ../options/internal/include  rbtree.hpp   slab.hpp   allocator.hpp   new   formatting.hpp   stdio-stubs.cpp   optional.hpp   utility.hpp   logging.hpp   utility   mutex.hpp   string.hpp   errno.h   <built-in>    stdarg.h   stddef.h   ssize_t.h   stdio.h   types.h   stdint.h 	  type_traits   debug.hpp   list.hpp     	r�F     �F  	ÀF     ��  	րF     �6J7tXK�  	�F     �Ju 2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	<�F     5//
�!  	(�F     ��#f  	4VG     � �f  	ZVG     � 	���  	�VG     � 	*	�/  	WG     � 	=�g  	VWG     � �f  	|WG     � �
t�<g��  	�WG     � � � ! � t � < < /	 � �x  	 XG     � � � � � t � < < /	 � �x  	�XG     � )�-#  	�XG     � ���Yt�<g��  	YG     �� � !
 � �v  	`YG     �> � �
 � �v  	�YG     �&�*#  	�YG     ����)�"� �3t5�@�K �
��
t	�t�
�� J�  	�ZG     �	�
t�<g��  	4[G     �� � !
 � �v  	�[G     �= � �
 � �v " 	G     ��4���	�KvX	ug	vYV/Y�K��f�=?���J?Y-	&gI/Y-	&g00Y-	)gL.�-�0�0�0� 0� 0�0�2�"/�<Y\�Y-	*gJ/Y-	&g2�	�0�t�t	�Ov.YX�-&g[/>�02KA�tuJYt � fY0�tuJYt� � fYZl.= t � X J � �' f !@/��@/�7�"
u�'��5J)�f*<,<= K[�>�02JJ<=K`/=@�Y?�YL�<K�<�YJ�YW�tV�t-�Y,�Y9��8��ؼ�
u	u uP0= t���g�=i�
fu�=iw�[g�=`f"XY)0�g�t
K	u Y /�L0�/'t
K	uYC/�/!0��0��0K!0K!(0�g�t
K	u =/�0�g/��08�� X � X	 L ��'WLu	JYww�.�X
K	w Y0�=�. ��9����׺�J��׬ ��H�uuP0uuC0�3�� ���>�$t=0�$t= 0�= t t
K	"+:B� �	�K�	���
Y��2u<X��fK�
��=�=�E�O1�����F�g3�Y-	&gD0>��
2�JJ<=JuK2!�NX��>!�PX��>!�QX��)>��$>�$t=&0�$t="0
��t
K	uJ =Q0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��&�-�t�WM�Y��/t]s�
X&� mf
�vX0' � � X K �
��
��0WM�Y��/
t]s�
X
&� ��-�4�t�WM�Y��/t]s�
X&� mf
�v+0/�y�	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=�}.	� u"	< � t% � �/���3	�# J �K�K�K�$ ���<% J � J t	 XL�_�u	� K �Y�" LE /" � � �Y�! LC /! � � �Y�( J  �Lu �( J  � K, � � Y � 6u	u;�Ku�Zu�[u�[�Ku�Zu�[u�1u�1u�1u�1�- J# �Ku�0u�	$;$w�)- ��'�1<�u5g�!!g#�$* f!g+�5�!�$�1 f!g+�5�!�$�1 �!�+�5�!�xt )X fg'�1<�ue.<C"�K$[�!! fg�)<�u3�K$\�!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X�K[�!u% f � J t XK�+u�g!K fz�5"+��=[�!ugu ���+��g!E
.�u�Ku��v�K(��!��K(�� i!�' J��- J% �K-�#�5 f0 �' � t �+���y�
��u! f�$�t�L+��g!yJ1&'��$��!g�!g�$" fg#�-���) fg#�-���) fg#�-��xt X��1�+����~.<<<<.<	'  t�}fD�<�} ��=  	6ZF     �<  	ZZF     7�  	�[G     � 
��  	vZF     )���u�K&<f/ 
 	�F     �� X J . K  	�[G     #�'f  	\G     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	�bG     #�'f  	
cG     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X 
 		G     �� X J . K  	�iG     #�'f  	 jG     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	�F     � v
�<g�ut�t!J�u �&�)J�  	��F     � ���tK t# < �Y�tK �i>���.��O�5U<ZJJ��tK  	��F     �
�t� 	 	�cF     � �/ 	 	�cF     � 		 	�cF     
�/K 		 	��F     
�/K 		 	dF     !�t��K  	�pG     #�'f  	�pG     �0	!�K� J KW	0��[� � � .	��	 K  �[
��KK� � � .�
�KK� � � .
�KK�   � .
�KK�   � .
�KK�   � . m�X$ � � .� � � .	��K� � � .�0Zu� J �K��Y� � � . �3	i��� � � .
���� � � .�3	;u � � � .�� J �K��.=� � � . �36	u��� � � .
��Ku� � � .��	�Ku� � � . � ? �� 
m�� X  	�[F     � �  	�[F     � � 
! 	�wG     0�g  	�wG     =�  	xG     K  	.xG     "=�/  	|xG     <�/K  	�xG     $(=�K  	�xG     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	�|G     =�  	�|G     K  	(}G     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	 �G     =�  	2�G     K  	\�G     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	�F     �����= f � .�("J��	���K � � .� � � .�t X. � < � J t XK � .�t	�t���g.�	�v�K � � .� � � .�t X. � < � J t XK � .�t	�t"������/fJ<��� � � .�g� X- �7 � JYu��
�KJ(7ȟ!������.fJ<�(�/�v< �
 	 	:dF     -�1%  	ndF     ��2  	M�F     ��6 	 	�dF     � �/  	4�G     =�  	f�G     K  	��G     (5+�'Z+�'Z+�'Z �� �� �� �� �� f��t�Z ��	�.�J�[2���  	g�G     � �  J �*KJJ�	�' J � < KJ�*>�0./�	<' J �!KJ�)>� 1��� 
 	�G     �K  	d�G     � � � � .�K  	��G     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	z�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	T�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	*�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	ڔG     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	��G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��G     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	?�G     ��_/0 � .� 		 	 G     
/K  	��G     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	~�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	X�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	.�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	ިG     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	��G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��G     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	C�G     ��_/0 � .�  	��G     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	��G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	\�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	2�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	��G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��G     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	G�G     ��_/0 � .�  	4�F     $�/�  	f�F     '��K�  	x�F     �	���# f- �+ � < f t Y  	��F     ����uf	u.u
fy.�"k  	r�F     � ��uu���
0K  	�F     7� � � .���  	ʙF     ��t �!�	����0 � � .�J5P�! � �4 g= � t t K � �	�K  	�F     ���fK/[���fKg0#�fKg0t�X  	�F     1� � � .���  	F     ���fK/[���fKg0#�fKg0t�X  	N�F     � � � .�t�J/	PK  	eF     �=/  	��F     �'� � J	� f f+ fgJ
Y fgJ
YgY
 �J
Yg
ug
ug
ug
ugL/B i�  	��G     �%� � � .� � � .� � � .� � � .�0/1%Z � � .� � � .� � � .� f � .� f � .� t* � < Y �h0Z � � .� � � .��	t.u$��= f) . . X t XK.Z�K t � = �h" f � � �i" f � Y �h t � u �j f � .�	t.u3��= f) . . X t XK.Z�� t � � 'h" f � � �i" f � Y �h t � � 'l � . �*$   	��G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	`�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	6�G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	�G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p   	��G     �.t � t. � f t t X 	J 	w � t U w � x � J U w < �~   	��G     ��.t � t. � f f t X 	J 	w � t U w � x � J U w < �p  	��G     ��2 � � .� � � .�gJ	3gJ	3gJ0 f � .�-h-� J( � .- J t t X1�� J t X = � J X $[ � � .�	��K	g=U f � .	�;[ � � .� � � .��	g=U f � .	�;Z � � .� � � .��	g=	V;Z � � .� � � .� < � .�i� J t X =	rXi� J t X =	vXi� J t X 	=S f � .�� J t X <0 � . ��.�    	K�G     ��_/0 � .� 
 	��G     ��
=�
g�g 
! 	��G     0�u 
 	
�G     ��
=�
g�g  	T�G     � �4  	�F     �h��K;0 	 	��F     &
��  	��G     �h�K;0 	 	�G     &
��  	�G     � �Fu	Ju4,4  	��G     � �3  	�G     � �4  	�G     ��4  	c�G     � �4  	��G     � �Fu	Ju4,4  	Y�G     � �3  	��G     � �4  	�G     � �4  	\�G     � �Fu	Ju4,4  	��G     � �3  	P�G     � �4  	��F     �  �u  	��F     � �(�K  	ݤF     � �)�K  	4�F     �K��uJ�KuJ�L�<fK�K��2       t 
X J � .��u��	tKJ�h f � .�J�LuJ�>�����u����u/  	��F     � �/�K  	��F     �K���u��	tKJ�h f � .�J�LJ�=$�<�>J�KuJ�>J�KuJ�?��J<,K��(K��K��J<L�����u����//  	�F     �  �u  	@�F     �6h:J  	b�F     ���  	��F     � � � � .��/1  	`�F     ����  	��F     � �(�K  	�F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	��F     � �)�K  	F�F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	��F     � � � � .��/1  	��F     �K � � .� X � .�J�KJ�?�uJ�KJ�KJ�KJ�L//1  	��F     �K � � .� X � .�J�KJ�?�J�KJ�KJ�KuJ�L//1  	~�F     �3g71 	 	�eF     0��  � .��gt��������y�	X 	 	�hF     &  � .��gt���J�����  	��F     �=7  	��G     � �4  	��G     � �Fu	Ju4,4  	��G     � �3  	��G     � �4  	I�G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	8�G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	NG     �/4  	��G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	0�G     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	w�G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	�G     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	f�G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	D�F     7��  	��F     � �-�K  	��F     � �uu�(<g  	�F     � � � .����t� X � .�<#<f��� f � .��u�wL f � .� X � .�<"<fK�/ f � .��u�w�<% J < J t XK�<fK�u/Z�u�u]�g�t�<$ J < J t XK�0�u�v� � � .�/�u<�=<� f � .�<% J < J t XK�0�u�v� � � .�/�u<�=<���    	��F     <�*�=  	Z�F     ���u�<L�0#  	εF     ���  	��F     ���  	ҿF     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	 �F     7��  	9�F     � �/�K  	f�F     ���u�<L�0#  	6�F     � �-�K  	�F     ���u�u\�u�<f�� t < t X J � 	.� �( f  < J t XK�u�u<v/Y'�/ f' < J t	 XK�u�u<v/[�t�	�tK//��/�v�� f � .�	�tK//��/�v�S�/   	FeF     �/4  	�G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � $�v � � . �J��gfŖg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	^�G     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	��G     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	O`F     �� J J . K  	�G     �	/fY%* � � � .�%  	��F     � �uu�(<g  	`�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	 �F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	Q�F     &
�Y  	B�F     &
�Y  	I�F     <�*�=  	T�F     � �uu�(<g  	�F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	��F     �� t   t X J � 	.���uJ�=J�KJ�=J�KJ�>u��	tKJ�h f � .�J�M//  	afF     �	/fY%* � � � .�%  	~G     � �Fg	<Y3,3  	�fF     � �3  	RgF     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h  	G     � #�v � � . ����g��g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h �   �   �      ../options/ansi/generic ../options/ansi/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include  string-stubs.cpp   errno.h   stddef.h    6 	��G     ���	t K�<�-0	uKH/�	��t J ��<�/V
2��=V	2KA0��	YKS/=���	K�t J ��<�/V2	uK70� �8��8g�g�u� zt	|Y*/	���=�= fgv�u�uY/+0�/<0	���u�=�= fgv�u�uY/T/=1��� ���<2K �	wY$/	��	!#Y�U3"g	�Y1/	�
�� J �  X t XKgV 20/	��!�f#K�U	3Y%/�� ����*Y.� �	xY0/	�
��  J �  X t XKgV 22/� �YK �!� J �+ � �
MK+|#g u�	�YU/= ��u�t	YJ
��t J t  X t XKW3�t J t  X t XKW1tKu
J�ZJ	vKD/��'1	��	!#Y�U!3�@0�?��F��C�.I�.M�.S�.A��J�<�<7�<A��J�<.��/��7�<E�<7�<+��2��4��,��1��3��W�<<��� ��J)Y,� �	wY 0�.�.�v35�Y.�Y2�Y3�Y0�Y4�Y0�Y&�Y5�/9�/-�/D�/9�/7�/*�/1�/7�0�K33/	�h�t
K	uY80=*�uA0���� �   $  �      ../sysdeps/lemon/generic ../options/internal/include/bits ../options/internal/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/posix/include/bits/posix  filesystem.cpp   types.h   stdint.h   stddef.h   ssize_t.h   off_t.h    K 	~H     
h'�tg
v YE0j'<Yv
� YD0])�uv
� Y81
0&uv
� Y0
�(Y00�	L<K�u Y �   �  �      ../subprojects/cxxshim/stage2/include ../options/internal/include/mlibc ../options/internal/generic ../subprojects/frigg/include/frg /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include  new   allocator.hpp   allocator.cpp   eternal.hpp   utility   slab.hpp   rbtree.hpp   stddef.h   type_traits   types.h   stdint.h   mutex.hpp   <built-in>    sysdeps.hpp    2 	YF     	�K  	H     �� ! 	�H     (� � J=u � J<' �; J1 �< J��0B� ��K@>= ��  	.H     ��  	ZH     *�K  	hH     �K  	vH     '���  	�H     *�K  	�H     �K  	�H     '���  	2H     *�K  	@H     �t  	RH     ��  	xH     �/ G X  
  	�H     ��  	
H     ���  	$H     ����  	HH     ��( ! 	H     �  	�H     � ��  	�H     ����  	�H     � �� �   �  �      ../options/internal/include/mlibc ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../subprojects/frigg/include/frg ../subprojects/cxxshim/stage2/include  charcode.hpp   charcode.cpp   stddef.h   types.h   stdint.h   optional.hpp   string.hpp   logging.hpp   type_traits   mbstate.h   debug.hpp   hash.hpp   formatting.hpp   <built-in>      	�H     � S!W(  	�H     � J  	H     �'f  	$H     �#t  	6H     .�)t	<=f�JL��u�u��u�u��u�u� � ��x ��t$Xt.uf
�t�Y  	�H     ;=	tY f
�tYt�t�Y  	�H     +�X�*��5K � J
5uB0��Y)0
Lu  	<H     � E�I(  	tH     � �!  	�H     � �  	�H     � � ��/� � � t X�Xg�LJuKut�/tt�XKu Y  	H     � v ��/� � � t X�Xg�KJvKu�t/tt�XKu Y  	bH     �v ��/���XgZKJvKuv XKu Y  	vH     �v ��1 � � t X�tY<K�+��K�
hgZ ��t�Jx�y XJtYu Y  	�H     
�t�  	�H     
�t�  	H     
�t�  	.H     
�t�  	NH     
�t� �   �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/generic /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   charset.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   string.hpp   debug.hpp   charcode.hpp   charset.hpp   <built-in>     2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1� # 	nH     	�Y%>u# � � J t X!K �! �. �! �9 X! .9 X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y&0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X;K �! �. �; �H 	�; �S X; .S X/��-X�	�Y%0u# � � J t X)�z� �+ �7 �C �� � �* �6 �B �� � �� � �) �5 �A ��� � �* �6 �B � � � �) � �1 X) 	.1 	X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��)�3��	�Y%>u# � � J t XGK �  �- �: �G 
� �O XG .O X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y%0u# � � J t XK � � X . X/��-X�	�Y*0u# � � J t XK �����-X�	�g*0u# � � J t XK �����-X�	�g0
Lu  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�cF     � �/  	�cF     � 	 	�cF     
�/K 	 	dF     !�t��K 	 	�cF     
�/K  	�[F     � �  	�[F     � �  	:dF     -�1%  	ndF     ��2  	�dF     � �/  	�dF     ��0  	eF     �=/  	FeF     �/4  	�eF     0��  � .��gt��������y�	X  	afF     �	/fY%* � � � .�%  	�fF     � �3  	RgF     � #�v � � . ���g<ňg � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	O`F     �� J J . K  	�hF     &  � .��gt���J�����    �  �      ../subprojects/cxxshim/stage2/include ../subprojects/frigg/include/frg ../options/internal/gcc /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0//include ../options/internal/include/bits ../options/internal/include ../options/internal/include/mlibc  new   formatting.hpp   guard-abi.cpp   optional.hpp   logging.hpp   utility.hpp   stddef.h   types.h   stdint.h   type_traits   string.hpp   debug.hpp   <built-in>     2 	YF     	�K  	&YF     2&�*M  	�YF     1��  	ZF     1�  	<�F     5//
�!  	�'H     �"u!��N�+$0��uF<��)�3���R>���J8<XK
�vZS/��Ju�  	6ZF     �<  	ZZF     7�  	vZF     )���u�K&<f/  	�ZF     � �/  	�ZF     � 	 	[F     
�/K 	 	$)H     
�/K 	 	T[F     !�t��K  	�[F     � �  	�[F     � �  	�[F     -�1%  	�[F     ��2  	M)H     ��2  	T\F     � �/  	z\F     �=/  	�)H     �=/S  	�\F     0��  � .��gt��������y�	X  	*H     �	=fY&* � � � .�&  	�*H     � �4  	+H     � $�v � � . � ��gf�g � � .��w.�K/ t . � � hfK! t � Y �h< f g �h 
 	O`F     �� J J . K  	x`F     &  � .��gt���J�����         extensions FT_ENCODING_APPLE_ROMAN FT_Face_Internal FT_ENCODING_ADOBE_EXPERT xMin user /home/computerfido/Desktop/Lemon/Applications/Init FT_StreamRec_ 20bitmap_info_header_t fbInfo FT_Face_InternalRec_ closeButtonBuffer num_faces FT_Size_InternalRec_ _ZN8ListNodeIP8Window_sEC4Ev FT_SubGlyph FT_DriverRec_ senderPID FT_Glyph_Format_ _ZN4ListIP8Window_sE10get_lengthEv FT_ENCODING_MS_BIG5 _ZN4ListIP8Window_sEixEj windows __mlibc_uintptr n_contours FT_ENCODING_NONE FT_UShort FT_ENCODING_MS_GB2312 FBInfo lsb_delta __buffer_size lastKey platform_id FT_Generic 10win_info_t FT_ENCODING_UNICODE RemoveDestroyedWindows recieverPID renderPos horiBearingX horiBearingY FT_Bitmap descriptor FT_Vector_ main fb_info_t FT_Stream_IoFunc mouseDown remove_at _ZN4ListIP8Window_sEC4Ev main.cpp uint8_t FT_Generic_Finalizer _ZN4ListIP8Window_sE8add_backES1_ FT_ENCODING_JOHAB compression FT_LibraryRec_ mouseX mouseY FT_ListRec_ environ unsigned char FT_Stream ownerPID FT_Int linePadding FT_ListNodeRec_ vertAdvance FT_ListNode add_front _ZN4ListIP8Window_sE10replace_atEjS1_ y_ppem yMax num_subglyphs FT_BBox_ mouseData underline_position __dirty_begin __offset FT_SizeRec_ 20bitmap_file_header_t _ZN4ListIP8Window_sE6get_atEj windowInfo hdrSize rows _ZN4ListIP8Window_sED2Ev vector2i_t decltype(nullptr) FT_ENCODING_ADOBE_STANDARD FT_Vector __mlibc_uint16 replace_at __static_initialization_and_destruction_0 FT_ENCODING_PRC operator+ stdin windowFound stdout vres __io_offset Vector2i FT_ENCODING_MS_SYMBOL descender _Z13AddNewWindowsv keyMsg FT_StreamDesc_ ascender finalizer ListNode<Window_s*> __mlibc_int8 style_name FT_ListRec FT_CharMapRec_ AddNewWindows __mlibc_uint32 linearHoriAdvance __dirty_end RGBAColour FT_Encoding_ _ZN10win_info_tC2Ev optind closeButtonLength _ZplRK8Vector2iS1_ FT_Generic_ __priority available_sizes mouseDevice add_back FT_GLYPH_FORMAT_BITMAP FT_Size num_fixed_sizes operator[] rsb_delta FT_Size_Metrics this active uintptr_t FT_String FT_ENCODING_MS_WANSUNG FT_Library FT_ENCODING_SJIS _GLOBAL__sub_I_keymap_us colourNum closeButtonSurface pixel_mode List<Window_s*> __mlibc_uint64 __initialize_p FT_Face long long int __mlibc_uint8 FT_StreamDesc yMin num_glyphs mouseEventMessage underline_thickness FT_SubGlyphRec_ 13ipc_message_t FT_Fixed FT_FaceRec_ rgba_colour_t renderBuffer FT_Glyph_Format FT_GLYPH_FORMAT_OUTLINE GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions FT_Bitmap_ palette FT_Size_Metrics_ __io_mode importantColours FT_ENCODING_ADOBE_CUSTOM FT_Encoding FT_ENCODING_MS_JOHAB FT_UInt32 FT_Glyph_Metrics autohint FT_UInt FT_Bitmap_Size_ _ZN4ListIP8Window_sE9add_frontES1_ fbSurface FT_GLYPH_FORMAT_COMPOSITE __buffer_ptr FT_BBox __valid_limit FT_CharMap FT_Short x_ppem long double FILE data2 get_front _Z10DrawWindowP8Window_s FT_Size_Internal FT_Glyph_Metrics_ FT_MemoryRec_ FT_Pos mainFont optopt _Z22RemoveDestroyedWindowsv style_flags FT_ENCODING_BIG5 surface_t uint16_t palette_mode FT_Driver _ZN4ListIP8Window_sED4Ev DrawWindow FT_GLYPH_FORMAT_NONE FT_Outline_ opterr mousePos FT_ENCODING_GB2312 FT_GlyphSlot max_advance control_data FT_ENCODING_ADOBE_LATIN_1 FT_Stream_CloseFunc ~List num_grays xMax get_back encoding_id FT_ENCODING_WANSUNG get_at FT_Alloc_Func num_charmaps max_advance_width _ZN4ListIP8Window_sE5clearEv horiAdvance FT_Bitmap_Size _ZN4ListIP8Window_sEC2Ev _ZN10win_info_tC4Ev stderr handle_t short int uint64_t drag colourPlanes linearVertAdvance redrawWindowDecorations FT_GLYPH_FORMAT_PLOTTER _ZN4ListIP8Window_sE9remove_atEj backgroundColor FT_Long get_length _ZN8ListNodeIP8Window_sEC2Ev FT_Slot_Internal FT_Free_Func windowHandle FT_Slot_InternalRec_ vertBearingX vertBearingY face_flags __dso_handle uint32_t dragOffset optarg _ZN4ListIP8Window_sE8get_backEv _windowCount title short unsigned int magic closeInfoHeader control_len hres FT_ENCODING_OLD_LATIN_2 FT_Outline max_advance_height sizes_list __in_chrg units_per_EM _ZN4ListIP8Window_sE9get_frontEv bitmap_top tags __mlibc_int32 FT_ENCODING_MS_SJIS closeButtonFile FT_Memory __status_bits FT_GlyphSlotRec_ FT_Realloc_Func face_index bitmap_left autofit_module_class FT_SpanFunc done_slot FT_Span FT_Byte FT_Renderer FT_Err_Corrupted_Font_Glyphs FT_Err_Max FT_Init_FreeType property_value glyph_size FT_Parameter FT_Err_Too_Few_Arguments FT_Err_Locations_Missing FT_Err_No_Unicode_Glyph_Name bearing_x no_stem_darkening FT_Err_Syntax_Error FT_Err_Array_Too_Large FT_Err_Invalid_Stream_Skip FT_Module_Class FT_Matrix_ FT_IncrementalRec_ FT_SIZE_REQUEST_TYPE_SCALES glyph_copy FT_Glyph_CopyFunc service_POSTSCRIPT_FONT_NAME request_size FT_Raster_BitTest_Func FT_Err_Invalid_PPem slot_object_size FT_Renderer_Class winfnt_driver_class FT_Size_RequestRec_ FT_Err_Invalid_Driver_Handle FT_Err_Invalid_Reference FT_Module_Interface FT_Incremental_GetGlyphDataFunc FT_Err_Invalid_Vert_Metrics FT_RasterRec_ glyph_format FT_Face_GetAdvancesFunc glyph_hints FT_Err_Invalid_Frame_Operation transform_matrix FT_Err_DEF_In_Glyf_Bytecode alibrary FT_Raster_RenderFunc FT_Incremental_InterfaceRec psnames_module_class FT_Incremental FT_Err_Invalid_Opcode FT_GlyphLoaderRec_ FT_Raster_ResetFunc FT_Err_Invalid_File_Format size_object_size FT_Err_Missing_Startchar_Field FT_Err_Invalid_Horiz_Metrics incremental_interface FT_Err_Invalid_Glyph_Index extra_points FT_Size_SelectFunc FT_Raster_SetModeFunc clip_box get_glyph_metrics FT_Err_Missing_Font_Field FT_Err_Stack_Overflow FT_Glyph version_major FT_Err_Invalid_Composite FT_Incremental_InterfaceRec_ FT_Size_RequestFunc FT_Err_Invalid_CharMap_Handle FT_Glyph_PrepareFunc FT_Size_Request FT_Err_Missing_Fontboundingbox_Field FT_GlyphLoader FT_Err_Horiz_Header_Missing FT_Err_Unlisted_Object ft_smooth_lcdv_renderer_class FT_Glyph_Class FT_Raster_Funcs_ FT_SIZE_REQUEST_TYPE_CELL FT_Module FT_ServiceCacheRec FT_Face_GetKerningFunc init_slot FT_Err_Invalid_Offset FT_Err_Invalid_Pixel_Size FT_Err_Unknown_File_Format render_glyph psaux_module_class FT_New_Library FT_Err_Bbx_Too_Big FT_Err_Bad_Argument FT_Err_Raster_Overflow FT_DebugHook_Func getenv FT_Err_Stack_Underflow FT_Raster_Params_ bdf_driver_class glyph_transform FT_Incremental_FreeGlyphDataFunc FT_Err_Code_Overflow FT_Err_Cannot_Open_Resource FT_GlyphRec_ FT_Render_Mode bit_test FT_Err_Raster_Uninitialized max_contours FT_Slot_InitFunc version_patch FT_ServiceCacheRec_ FT_Err_Invalid_CharMap_Format FT_Slot_DoneFunc FT_Face_DoneFunc transform_glyph FT_Err_Ok FT_Err_Could_Not_Find_Context FT_Driver_ClassRec_ FT_RENDER_MODE_NORMAL FT_Err_Missing_Encoding_Field property_name ft_raster1_renderer_class FT_Err_Divide_By_Zero service_WINFNT horiResolution module_requires max_subglyphs FT_Err_Invalid_Frame_Read extra_points2 FT_Err_Invalid_CodeRange bit_set FT_RENDER_MODE_LCD FT_Incremental_MetricsRec_ FT_Err_Corrupted_Font_Header version_minor FT_Err_CMap_Table_Missing FT_Set_Default_Properties FT_Renderer_SetModeFunc FT_Raster_BitSet_Func FT_Raster_Params glyph_class FT_Err_Raster_Corrupted FT_Incremental_MetricsRec module_interface transform_delta glyph_delta FT_ModuleRec_ renderers FT_Add_Default_Modules num_modules FT_Err_Too_Many_Function_Defs GNU C89 8.2.0 -mtune=generic -march=x86-64 -g -O2 -ansi FT_Glyph_TransformFunc FT_Driver_ClassRec FT_Renderer_Class_ pfr_driver_class FT_Err_Missing_Size_Field FT_Matrix FT_Glyph_InitFunc FT_Incremental_FuncsRec done_size max_points target module_data FT_Err_Too_Many_Drivers FT_Err_Invalid_Character_Code FT_Err_Out_Of_Memory FT_Err_Post_Table_Missing autohint_mode FT_Err_Missing_Chars_Field ft_property_string_set FT_Raster FT_Err_Cannot_Open_Stream FT_Renderer_TransformFunc FT_Err_Invalid_Face_Handle FT_Raster_DoneFunc FT_Error FT_Err_Too_Many_Hints cff_driver_class cur_renderer FT_Size_Request_Type FT_Err_Nested_Frame_Access t1_driver_class FT_Err_Lower_Module_Version FT_Err_Hmtx_Table_Missing FT_GlyphLoadRec_ module_flags FT_Render_Mode_ FT_Glyph_Class_ FT_Char ft_default_raster FT_New_Memory FT_Slot_LoadFunc FT_Err_Debug_OpCode faces_list raster_class transform_flags glyph_matrix bearing_y FT_Glyph_GetBBoxFunc FT_Size_Request_Type_ FT_Err_Too_Many_Extensions ft_smooth_renderer_class FT_Add_Module FT_Data FT_Err_Invalid_Handle FT_ModuleRec FT_GlyphLoadRec FT_Done_FreeType t42_driver_class module_name ft_smooth_lcd_renderer_class FT_Int32 refcount FT_Face_InitFunc service_MULTI_MASTERS FT_Glyph_DoneFunc FT_Err_Missing_Bitmap FT_Raster_NewFunc FT_Err_Invalid_Stream_Seek FT_Err_Table_Missing FT_RENDER_MODE_LIGHT module_done service_GLYPH_DICT pshinter_module_class FT_Parameter_ get_glyph_cbox FT_Err_Invalid_Stream_Handle FT_Err_Execution_Too_Long black_spans FT_RENDER_MODE_MAX autohint_metrics FT_Bool attach_file FT_Module_Class_ FT_RENDER_MODE_LCD_V glyph_bbox FT_Incremental_FuncsRec_ FT_Renderer_RenderFunc /home/computerfido/Desktop/freetypetest2/build module_size FT_Err_Invalid_Slot_Handle FT_Err_Invalid_Outline FT_Err_Raster_Negative_Height module_version FT_Err_Missing_Startfont_Field FT_Err_Invalid_Library_Handle FT_Err_Invalid_Cache_Handle FT_Err_Glyph_Too_Big FT_Err_Invalid_Table FT_Err_Cannot_Render_Glyph FT_ULong FT_Err_Missing_Property FT_SIZE_REQUEST_TYPE_REAL_DIM service_PFR_METRICS init_size FT_Module_Constructor FT_Err_Invalid_Stream_Operation vertResolution FT_Err_Invalid_Size_Handle FT_Renderer_GetCBoxFunc use_extra FT_Err_Ignore FT_Module_Destructor FT_RENDER_MODE_MONO glyph_loader FT_Err_Invalid_Version FT_Err_Invalid_Stream_Read FT_Err_Missing_Module FT_Err_Name_Table_Missing FT_Err_Invalid_Post_Table_Format FT_RendererRec_ FT_Span_ module_init FT_Err_Too_Many_Instruction_Defs FT_Err_Nested_DEFS FT_Err_Invalid_Glyph_Format FT_SIZE_REQUEST_TYPE_NOMINAL FT_Err_Unimplemented_Feature auto_hinter FT_Size_InitFunc FT_Size_DoneFunc FT_Err_Invalid_Argument pcf_driver_class select_size advance_v FT_SIZE_REQUEST_TYPE_MAX debug_hooks FT_Err_Missing_Bbx_Field FT_Pointer /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftinit.c FT_SIZE_REQUEST_TYPE_BBOX FT_Err_Invalid_Post_Table FT_Module_Requester gray_spans FT_Driver_Class FT_Done_Memory FT_Err_ENDF_In_Exec_Stream glyph_prepare FT_Done_Library t1cid_driver_class face_object_size FT_Data_ FT_Err_Too_Many_Caches tt_driver_class sfnt_module_class FT_Raster_Funcs service_METRICS_VARIATIONS FT_Face_AttachFunc FT_Incremental_GetGlyphMetricsFunc glyph_transformed ft_default_modules FT_Property_Get version_number CheckSum_Adjust ft_raccess_sort_ref_by_id font_program_size FT_Frame_Op_ vertical vec1 vec2 glyph_locations FT_GlyphLoad FT_Set_Char_Size GX_BlendRec_ FT_Sfnt_Tag_ rdata_len isFixedPitch instructions maxInstructionDefs TT_SBit_Scale FT_UInt64 ft_glyphslot_alloc_bitmap FT_Properties_SetFunc usWeightClass p_index xMax_Extent xAvgCharWidth hash_str_compare block2 TT_MaxProfile FT_Properties_GetFunc TT_GaspRec result_offset error2 ft_frame_schar FT_Stream_ReadUOffset FT_New_Face FT_Done_Face panose debug_hook min_origin_SB reset_face TT_SbitTableType_ num_kern_tables FT_Service_TrueTypeEngine glyf_offset ft_service_list_lookup FT_Stream_ExtractFrame FT_AutoHinter_InterfaceRec_ hori errors FT_Outline_New_Internal ft_frame_short_le vfs_rfork_has_no_font hash_insert first_point FT_GlyphLoader_Add access_glyph_frame Mac_Read_sfnt_Resource strstr result_file_name short_metrics FT_SFNT_TableGetFunc doblend FT_Get_Sfnt_Table kern_order_bits kern_avail_bits FT_Get_Module_Interface FT_RFork_Rule_linux_cap render_mode FT_GlyphLoader_CheckPoints ft_frame_end driver_name max_profile FT_Outline_Get_CBox ft_frame_ushort_le FT_Get_Font_Format ft_hash_str_insert nouse padvance TT_Post_20Rec_ ft_corner_is_flat test_mac_fonts map_len raccess_guess_apple_generic _ft_face_scale_advances FT_Hash args2 kern_table_size ft_hash_num_init face_index_in_resource ft_hash_str_init FT_Outline_Transform var_postscript_prefix FT_SFNT_HEAD yshift FT_Get_Kerning FT_MulFix ulUnicodeRange3 FT_Face_GetVariantSelectors forget_glyph_frame advance_Height_Max FT_GlyphDict_GetNameFunc maxCompositePoints maxStorage subg xshift langID anoutline FT_RFork_Rule_darwin_ufs_export usWidthClass FT_TrueTypeEngineType maxPPEM FT_CMapRec_ original_name engine_type FT_RFork_Rule_ ft_glyphslot_done Line_Gap FT_New_Size aslot p_arg2 in_y FT_ServiceDescRec astream raccess_guess_linux_double stringOffset structure is_sfnt_cid sbit_num_strikes FT_Get_Postscript_Name FT_Get_Sfnt_Name_Count FT_List_Up FT_PIXEL_MODE_GRAY FT_CharMapRec FT_GlyphLoader_Done pfb_len left_bearing __builtin_memset languageID p_arg1 FT_Offset fsSelection Fail agindex FT_Vector_Unit min_advance_SB v_prev hash_bucket ySubscriptYSize entry_length maxMemType42 TT_Loader_StartGlyphFunc angle1 angle2 acmap FT_DriverRec load_flags FT_Stream_Read FT_Property_Set raccess_get_rule_type_from_rule_index ft_cmap_done_internal vcmap TT_GaspRangeRec_ FT_SFNT_OS2 pfb_lenpos TT_Postscript_ FT_Matrix_Invert service_id numPoints FT_Stream_New aminor raccess_guess_linux_cap FT_Vector_NormLen FT_Set_Charmap achVendID ulUnicodeRange1 ulUnicodeRange2 ulUnicodeRange4 head2 vert_resolution FT_Get_First_Char last_charmap horz_resolution get_track FT_RFork_Rule_darwin_hfsplus new_count FT_ServiceDesc hash_num_compare maxComponentDepth destroy_face minMemType42 FT_Outline_Done_Internal TT_TableRec_ FT_Angle_Diff ft_mem_dup Index_To_Loc_Format FT_CMap_New FT_Stream_EnterFrame FT_Vector_Polarize FT_Hashkey_ FT_Service_GlyphDictRec_ hash_init hdmx_record_count TT_SBIT_TABLE_TYPE_NONE FT_Stream_ReadUShortLE caret_slope_denominator FT_ValidationLevel_ usFirstCharIndex FT_AutoHinter_Interface /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftbase.c p_error is_cff ft_hash_num_insert FT_Set_Transform FT_SFNT_POST size_index buffer_max FT_PIXEL_MODE_GRAY2 FT_PIXEL_MODE_GRAY4 padvances ttface FT_Raccess_Guess is_owner d_hypot sfnt_data get_table TT_Header desc theta FT_Atan2 Modified FT_CMap_ClassRec_ FT_Stream_GetUOffset get_global_hints FT_Face_GetCharVariantIndex linear_def FT_Get_Charmap_Index raccess_guess_apple_single variantSelector char_height rfork_offset ft_mem_realloc TT_Header_ is_light_type1 TT_Post_NamesRec exec FT_Cos Load_Ok FT_MulFix_x86_64 ySubscriptXOffset FT_Set_Pixel_Sizes FT_Load_Glyph FT_List_Iterate num_locations FT_CMap_DoneFunc right_glyph variantchar_list FontNumber var_postscript_prefix_len external_stream number_Of_HMetrics stream2 FT_Frame_Field FT_Hashnode min_Right_Side_Bearing ft_validator_run FT_SFNT_TableInfoFunc maxContours FT_PIXEL_MODE_LCD TT_Face Mac_Read_POST_Resource usWinDescent TT_GlyphZoneRec TT_SBIT_TABLE_TYPE_SBIX glyph_indices ins_pos hook_index swap FT_Vector_Rotate ft_open_face_internal file_names FT_Service_Kerning language ft_raccess_rule_by_darwin_vfs FT_Stream_Seek TT_Name cmap_size memory_stream_close TT_NameTableRec_ allzeros usMaxContext ystrength ft_frame_skip jmp_buf FT_Get_CMap_Format FT_List_Finalize FT_Get_Track_Kerning TT_MaxProfile_ usBreakChar FT_ORIENTATION_NONE acbox strncpy degree char_width sTypoLineGap magic_from_stream cvt_program_size FT_Hypot pads CharacterComplement FT_Service_TTCMapsRec_ frame_accessed FT_Outline_ConicToFunc FT_GlyphLoader_New FT_Vector_Transform FT_Remove_Module new_max FT_Attach_Stream FT_Stream_Free Font_Direction after FT_Outline_EmboldenXY FT_CMap_CharVariantListFunc FT_PIXEL_MODE_MAX darken_params cur_size resource_cnt FT_Load_Sfnt_Table ulCodePageRange1 ulCodePageRange2 FT_CMap_CharVarIsDefaultFunc maxFunctionDefs rpos ft_glyphslot_init error1 FT_Service_PropertiesRec_ numLangTagRecords FT_SfntName_ FT_DivFix FT_CMap_Class FT_Vector_From_Polar maxPoints FT_Outline_MoveToFunc FT_TRUETYPE_ENGINE_TYPE_PATENTED advance_Width_Max Table_Version old_max FT_Stream_Open TT_LangTagRec_ pixel_width TT_Loader_EndGlyphFunc num_sbit_scales font_program FT_Get_Char_Index FT_Service_SFNT_Table ps_property_get n_base_points caret_slope_numerator TT_Interpreter langTags horizontal FT_GlyphLoader_CopyPoints x_left set_property FT_Request_Metrics FT_MulDiv_No_Round FT_Select_Charmap FT_PIXEL_MODE_LCD_V TT_Post_25Rec long_metrics missing_func FT_ValidatorRec_ num_tables numRanges v_middle v_start FT_SFNT_VHEA Destroy_Module FT_KERNING_DEFAULT nameID Calculate_Ppem FT_Get_Name_Index FT_RFork_Rule FT_ServiceDescRec_ metric_Data_Format FT_Stream_GetUShort sTypoDescender IsMacBinary FT_ORIENTATION_POSTSCRIPT ySuperscriptXSize FT_GlyphLoader_CreateExtra xtemp FT_FaceRec TT_VertHeader_ FT_Outline_Reverse FT_Open_Face FT_Service_GlyphDict cvt_program raccess_guess_apple_double ft_mem_strdup read_composite_glyph FT_Get_CMap_Language_ID d_in FT_RFork_Rule_linux_double xOffset numGlyphs platformID ps_property_set FT_PIXEL_MODE_NONE TT_SBit_LineMetricsRec FT_List_Insert d_out hdmx_record_size FT_Set_Renderer FT_CMap_CharVarIndexFunc FT_Select_Size FT_AutoHinter_GlobalDoneFunc longjmp FT_TRUETYPE_ENGINE_TYPE_UNPATENTED Magic_Number FT_CMap ft_mem_qalloc FT_SFNT_HHEA FT_Get_Renderer char_var_default TT_SBit_LineMetricsRec_ arctanptr FT_GlyphLoader_Adjust_Points FT_GlyphLoader_Prepare raccess_guess_linux_double_from_file_name TT_CMap_Info_GetFunc FT_GlyphDict_NameIndexFunc FT_Raccess_Get_HeaderInfo FT_AutoHinter_GlobalGetFunc hash_lookup number_Of_VMetrics FT_RFork_Rule_vfat sbit_strike_map TT_OS2_ FT_Set_Debug_Hook maxComponentElements x_shift top_bearing yMax_Extent FT_GlyphLoader_Rewind minMemType1 ft_recompute_scaled_metrics ft_lookup_PS_in_sfnt_stream serv_data variation_support FT_VALIDATE_DEFAULT ySubscriptYOffset maxMemType1 ySuperscriptXOffset y_ppem_substitute alangTag v_control PS_DriverRec_ ft_raccess_guess_rec FT_Get_TrueType_Engine_Type Lowest_Rec_PPEM FT_Raccess_Get_DataOffsets FT_Stream_GetChar TT_OS2 min_after_BL aname PS_Driver Created FT_ORIENTATION_TRUETYPE __builtin_memcpy FT_New_GlyphSlot FT_SFNT_MAXP level ft_synthesize_vertical_metrics result FT_Outline_New raccess_guess_darwin_ufs_export parameters strings_size encodingID Fail2 hdmx_table raccess_guess_linux_netatalk raccess_guess_darwin_hfsplus open_face read_glyph_header FT_Library_Version numNameRecords is_num StrokeWeight TT_Post_25_ FT_Stream_Pos vert_metrics_offset tag_internal sCapHeight filepathname FT_Face_Properties FT_Outline_Funcs_ vert_metrics_size FT_CMap_Done FT_Stream_ReadULong FT_Orientation_ TT_NameRec ft_frame_bytes x_ppem_substitute entry_offset raccess_guess_vfat num_params TT_BDFRec FT_CMap_CharNextFunc ptrdiff_t TTC_HeaderRec TT_ExecContext FT_GlyphLoader_CheckSubGlyphs FT_Outline_LineToFunc FT_CMap_CharIndexFunc sbit_table FT_RFork_Rule_apple_double max_before_BL ft_glyphslot_clear usLowerOpticalPointSize new_memory_stream stringLength FT_F26Dot6 FT_AutoHinter_GlobalResetFunc FT_Stream_GetULong maxStackElements caret_Offset ft_frame_uoff3_be FT_KERNING_UNSCALED FT_PtrDist FT_Get_Glyph_Name aface TT_HoriHeader FT_List_Add maxCompositeContours caret_Slope_Run FT_Get_Sfnt_Name SymbolSet TT_CMapInfo_ find_variant_selector_charmap sfnt_ps subcnt FT_Stream_ReadAt pbytes new_name FormatType ft_frame_off3_be TT_Loader_GotoTableFunc kern_table v_cur memory_base read_bytes akerning usWinAscent TT_PCLT_ FT_Service_KerningRec_ TT_SBIT_TABLE_TYPE_CBLC yStrikeoutSize destroy_size dlen FT_SfntLangTag ft_glyphslot_preset_bitmap FT_Outline_Get_Orientation is_cff2 FT_Load_Char FT_HashnodeRec_ FT_List_Destructor FT_Stream_ReleaseFrame FT_Service_Properties FT_Pixel_Mode_ ft_trig_arctan_table ft_glyphslot_grid_fit_metrics Mac_Style num_names FT_Sfnt_Tag l_anchor TT_CMapInfo TT_SbitTableType FT_Reference_Face map_pos yOffset ft_mem_alloc TypeFace apatch FT_RFork_Ref is_darwin_vfs ebdt_size ft_frame_byte FT_Vector_Length base_file_name FileName FT_Match_Size ySuperscriptYOffset hdmx_record_sizes TT_SizeRec_ name_table FT_Outline_Translate FT_Stream_ExitFrame yStrikeoutPosition FT_Outline_Embolden FT_SFNT_PCLT gaspFlag FT_Size_RequestRec FT_Sin FT_Tag FT_Tan Fail3 FT_TRUETYPE_ENGINE_TYPE_NONE y_shift FT_Face_GetCharVariantIsDefault num_properties ft_module_get_service TT_Postscript new_names newpath TT_Loader_ReadGlyphFunc FT_Open_Args_ kern_mode ft_trig_prenorm ft_lookup_glyph_renderer FT_Done_GlyphSlot FT_Frame_Field_ FT_Get_Advances memory_size FT_Outline_Decompose table_end TT_BDFRec_ FT_RFork_Rule_uknown p_transform pfb_pos horz_metrics_size FT_SFNT_MAX FT_Stream_GetUShortLE FT_Stream_ReadFields FT_Kerning_TrackGetFunc face_index_internal max_width sub_index ft_frame_ulong_be TT_Size slash FT_Hash_LookupFunc serv_id resource_fork_entry_id FT_PsName_GetFunc done_global_hints FT_MulDiv base_file_len _tmp_ strlen abitmap FT_Render_Glyph caret_Slope_Rise sxHeight insertion FT_Open_Args FT_Service_PsFontName ft_frame_long_be FT_ORIENTATION_FILL_RIGHT FT_Select_Metrics FT_Hashkey ySuperscriptYSize sFamilyClass ft_hash_str_free FT_GlyphLoader_Adjust_Subglyphs pstable_index data_offsets jump_buffer FT_Stream_ReadULongLE ft_frame_uoff3_le read_simple_glyph end0 hash_rehash FT_Get_SubGlyph_Info psaux CheckSum FT_FloorFix open_face_from_buffer FT_Stream_ReadUShort FT_Service_TTCMaps FT_Get_Sfnt_LangTag usUpperOpticalPointSize TT_Loader TT_HoriHeader_ FT_SFNT_TableLoadFunc maxZones Font_Revision FT_List_Remove ft_property_do raccess_make_file_name FT_RFork_Rule_linux_netatalk aloader TT_LangTag init_data FT_RFork_Rule_apple_single FT_RFork_Ref_ FT_AutoHinterRec_ value_is_string TT_Post_20Rec FT_Stream_TryRead scaled_h FT_Get_Module interpreter TTC_HeaderRec_ reads scaled_w FT_Int64 func_interface FT_ORIENTATION_FILL_LEFT sfnt FT_Matrix_Multiply_Scaled FT_SfntName ft_raccess_guess_func TT_FaceRec_ TT_LangTagRec underlineThickness strcat ft_remove_renderer FT_RFork_Rule_darwin_newvfs Do_Conic null_outline FT_HashRec_ open_face_PS_from_sfnt_stream cmap_table mod_name FT_TrueTypeEngineType_ orig_x orig_y before glyf_len load_mac_face qsort numTables in_x FT_List TT_GlyphZoneRec_ flag_offset FT_CMap_VariantCharListFunc find_unicode_charmap new_length TypeFamily TT_SBIT_TABLE_TYPE_MAX horz_metrics_offset composites fsType ft_validator_init resource_offset FT_Stream_ReadChar FT_ValidationLevel TT_PCLT usLastCharIndex pfb_data ebdt_start ft_glyphslot_set_bitmap left_glyph FT_Stream_Close FT_Sfnt_Table_Info ft_frame_off3_le FT_AutoHinter_GlyphLoadFunc FT_Outline_Funcs ft_corner_orientation FT_KERNING_UNFITTED FT_RFork_Rule_invalid postscript_names usDefaultChar FT_Get_Advance ft_frame_start ft_raccess_guess_table n_curr_contours TT_Gasp_ ft_raccess_guess_rec_ gloader ySubscriptXSize FT_Face_GetCharsOfVariant FT_Orientation offsets_internal FT_Reference_Library FT_New_Memory_Face IsMacResource n_subs TT_Table Success numContours FT_CMap_VariantListFunc FT_Get_Next_Char ucmap min_Top_Side_Bearing min_Bottom_Side_Bearing p_flags dir_tables sbit_table_type maxTwilightPoints FT_CeilFix ft_frame_ulong_le ft_add_renderer FT_Activate_Size ft_lcd_padding out_x out_y Units_Per_EM ft_glyphslot_free_bitmap ft_hash_num_lookup FT_Incremental_Interface FT_Pixel_Mode pixel_height base_name FT_Stream_OpenMemory ignore_width item_size gaspRanges FT_Service_PsFontNameRec_ italicAngle FT_Service_TrueTypeEngineRec_ ft_frame_short_be TT_NameTableRec asize FT_List_Iterator ft_trig_pseudo_polarize min_Left_Side_Bearing cur_count FT_Outline_Get_Bitmap FT_Service_SFNT_TableRec_ TT_GaspRange destroy_charmaps FT_Angle FT_CMap_InitFunc ft_set_current_renderer hdmx_table_size raccess_guess_darwin_newvfs type_list language_id hinting_engine WidthType FT_Request_Size SerifStyle sTypoAscender ft_frame_ushort_be external FT_Hash_CompareFunc TT_ExecContextRec_ num_contours ft_validator_error FT_Matrix_Multiply service_descriptors FT_Outline_Done sign_shift ft_trig_pseudo_rotate ft_mem_qrealloc amajor FT_PIXEL_MODE_BGRA TT_Post_NamesRec_ ft_frame_long_le FT_UInt16 n_of_entries sort_by_res_id FT_Stream_GetULongLE FT_RoundFix load_table FT_Outline_CubicToFunc ft_mem_free ft_trig_downscale ft_hash_str_lookup Exit2 FT_AutoHinter TT_SBit_ScaleRec_ FT_Face_GetVariantsOfChar strtol FT_PIXEL_MODE_MONO strrchr origin TT_LoaderRec_ xstrength FT_Done_Size FT_Vector_Transform_Scaled FT_VALIDATE_TIGHT num_points Glyph_Data_Format GX_Blend FT_Render_Glyph_Internal ft_mem_strcpyn cvt_size FT_VALIDATE_PARANOID FT_Outline_Render file_size FT_List_Find FT_Validator FT_Kerning_Mode_ TT_VertHeader sbit_table_size ttc_header Reserved FT_Attach_File FT_SfntLangTag_ new_size load_face_in_embedded_rfork allmatch FT_GlyphLoader_Reset rdata_pos underlinePosition storageOffset Destroy_Driver charvariant_list caret_offset TT_NameRec_ FT_Outline_Check format_tag TT_SBIT_TABLE_TYPE_EBLC FT_Outline_Copy FT_Stream_Skip v_last FT_Lookup_Renderer maxSizeOfInstructions FT_Get_X11_Font_Format /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftfntfmt.c FT_Library_SetLcdFilterWeights FT_LcdFilter_ FT_LCD_FILTER_LEGACY FT_LCD_FILTER_LEGACY1 FT_LCD_FILTER_DEFAULT /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftlcdfil.c FT_LcdFilter FT_LCD_FILTER_LIGHT FT_LCD_FILTER_NONE FT_Library_SetLcdFilter FT_LCD_FILTER_MAX filter TT_Err_Invalid_Table TT_Err_Invalid_CharMap_Format Ins_SHP TT_Err_Syntax_Error inline_delta tt_face_load_loca nIfs TT_Err_Invalid_Reference is_composite tt_size_reset dualVector GX_HVVarTableRec_ old_range sfnt_id out1 out2 FT_SizeRec TT_Err_Missing_Font_Field TT_Get_Name_ID_Func codeRangeTable TT_Err_Invalid_Stream_Operation TT_DotFix14_long_long SFNT_Interface_ TT_Err_Horiz_Header_Missing TT_Err_Raster_Overflow axisSize Update_Max TT_Err_Too_Many_Function_Defs tt_coderange_font FT_Service_MultiMastersRec_ GX_TC_RESERVED_TUPLE_FLAGS FT_Multi_Master_ GX_TI_RESERVED_TUPLE_FLAG strid avalue cur_range shortDeltaCount delta_cnt tt_prepare_zone innerIndex projVector TT_CallRec SFNT_Service dummy2 Ins_GETINFO TT_Err_Name_Table_Missing compensations TT_Project_Func tt_service_properties storage_size tt_size_run_fpgm TT_Err_Glyph_Too_Big TT_Err_Ignore codeSize Compute_Point_Displacement FT_F2Dot14 netAdjustment FT_Get_MM_Var_Func TT_CallRec_ all_design_coords Round_None Ins_S45ROUND TT_Err_Invalid_Horiz_Metrics Ins_ODD Ins_SFVTPV Caller_IP tt_size_init y_ratio namedstyle tt_loader_set_pp Ins_MPS Ins_JMPR aIdx1 aIdx2 next_coords_size GX_AVarCorrespondenceRec_ TT_CodeRange_ gv_glyphcnt GX_ItemVarStoreRec_ tt_face_load_prep iupx_called Ins_GPV start_contour GX_DeltaSetIdxMap tt_get_var_blend Compute_Round Ins_INSTCTRL incr_metrics F_dot_P localpoints tt_driver_done opcode rotated Ins_DEBUG Ins_PUSHB TT_Err_Hmtx_Table_Missing scalar ref2 TT_Process_Simple_Glyph Ins_DIV iupy_called discriminant TT_Err_Invalid_Face_Handle Ins_PUSHW instanceSize TT_Err_Invalid_Stream_Read Ins_SHC control_value_cutin TT_Err_Invalid_Pixel_Size Ins_SHZ psid refp GetShortIns func_write_cvt tt_check_trickyness_sfnt_ids Ins_NPUSHB TT_Err_Missing_Fontboundingbox_Field FT_Set_MM_Design_Func TT_Err_Locations_Missing Ins_CLEAR Ins_NPUSHW grayscale get_mm Ins_FLIPRGOFF GX_TI_INTERMEDIATE_TUPLE instruct_control GX_VarRegionRec_ Current_Ppem num_axis TT_Init_Glyph_Loading im_start_coords TT_Err_Invalid_Offset TT_Clear_CodeRange Ins_NROUND tt_face_vary_cvt Ins_RTHG TT_Load_Context Ins_DELTAC Ins_FLIPON tt_face_done_loca FT_HAdvance_Adjust_Func cont_limit __builtin_strcmp Exit1 tt_face_load_hdmx TT_Err_Invalid_Library_Handle Round_To_Double_Grid Move_CVT_Stretched incr get_psname Ins_UNKNOWN Ins_SCANCTRL Round_Super node2 scan_control dotproduct Ins_SFVTL TT_Err_Invalid_File_Format Ins_RTG cur1 cur2 FT_Get_MM_Blend_Func Round_Down_To_Grid ft_var_to_normalized Normalize TT_GraphicsState_ FT_Var_Axis_ TT_Err_Out_Of_Memory TT_RunIns TT_Err_Invalid_Glyph_Format load_eblc curs tt_face_free_hdmx Ins_SMD cur_dist vvar_table varData TT_Err_Invalid_Driver_Handle Ins_SANGW table_len GX_TI_PRIVATE_POINT_NUMBERS next_name FT_Service_PropertiesRec axisCoords glyphSize tt_service_gx_multi_masters delta2 TT_CodeRange_Tag_ IUP_Worker end_point Ins_LTEQ ttsize TT_CodeRangeTable hvar_error glyphoffsets FT_Set_MM_Blend_Func FT_Service_TrueTypeEngineRec current_outline header_only mapData Round_Up_To_Grid namedstyle_size new_top mvar_tag LErrorCodeOverflow_ loopcall_counter_max subglyph FT_VAdvance_Adjust_Func round_state ft_var_get_value_pointer TT_Err_Missing_Bitmap GX_DeltaSetIdxMapRec_ Ins_MDRP Ins_ENDF delta_x delta_y GX_TC_TUPLE_COUNT_MASK TT_Err_Ok Ins_NOT TT_Get_Metrics_Func TT_Face_GetKerningFunc num_axes stackSize subpixel_hinting_lean TT_Load_Any_Func TT_Err_DEF_In_Glyf_Bytecode Ins_EQ tt_size_ready_bytecode TT_Err_Raster_Uninitialized point_cnt tupleIndex tt_face_load_fpgm coderange TT_Err_Invalid_Version FT_Get_Var_Design_Func has_fpgm outerIndex rsb_adjust tt_get_kerning Ins_IP do_scale Direct_Move_X TT_Set_MM_Blend tt_coderange_cvt TT_Err_Table_Missing step_ins p_limit _pbuff temp2 vertical_lcd_lean TT_GlyphSlot Ins_ABS sharedpoints func_round tt_size_run_prep TT_Set_Var_Design TT_Err_Corrupted_Font_Glyphs Ins_EIF TT_Err_Missing_Encoding_Field tt_interpolate_deltas axisTag tt_size_select TT_Err_Invalid_CodeRange vvar_error Ins_SSW GX_FVar_Head Ins_MSIRP TT_DefRecord_ TT_Get_PS_Name_Func Ins_WCVTF TT_Err_Too_Many_Drivers reexecute Ins_ADD widthMap_offset TT_Err_Missing_Module TT_Err_Invalid_Stream_Skip TT_Load_Simple_Glyph TT_Err_Stack_Underflow regionCount points_out TT_Err_Execution_Too_Long Ins_GT flag_limit Round_To_Grid callStack instanceCount ttslot Ins_SUB Project_x axisCount TT_Err_CMap_Table_Missing innerBitCount in_points cvtEntry table_start TT_Err_Unimplemented_Feature tt_driver_init GX_AxisCoords GX_DeltaSetIdxMapRec default_GS func_project Ins_SZP0 Ins_SZP1 Ins_SZP2 TT_Access_Glyph_Frame FT_Service_MetricsVariationsRec _iup_worker_interpolate instruction_trap has_cvt TT_DefArray TT_Err_Lower_Module_Version LNo_Error_ free_psnames n_ins Ins_FLOOR tt_glyph_load glyphCount vec_limit tt_vadvance_adjust need_init opcode_length single_width_value Ins_AA tt_get_metrics_incr_overrides Ins_IUP TT_Load_Glyph TT_DefRecord max_function_defs num_function_defs tt_glyphzone_new Ins_SWAP Caller_Range phase TT_Err_Invalid_Post_Table Ins_EVEN TT_Err_Invalid_Slot_Handle round_mode Ins_IF numIDefs func_read_cvt tuplecoords TT_Err_Invalid_CharMap_Handle fvaraxis_fields correspondence GX_VarRegion prev_cont func_cur_ppem TT_Forget_Glyph_Frame tt_hvadvance_adjust TT_Err_Bbx_Too_Big Ins_IDEF Ins_CEILING touch Init_Context TT_Err_Missing_Bbx_Field first_delta TT_Err_ENDF_In_Exec_Stream tupleCount deltas_x num_coords FExit TT_Size_Metrics fvar_fields TT_Err_Bad_Argument ft_var_load_mvar tt_apply_mvar TT_Err_Corrupted_Font_Header ref1 neg_jump_counter_max SetSuperRound Ins_ISECT manageCvt nump tt_check_trickyness_family TT_Err_Invalid_Opcode TT_Err_Missing_Startfont_Field TT_Err_Stack_Overflow max_ins set_mm_design Fail_Memory tt_services GX_TC_TUPLES_SHARE_POINT_NUMBERS GX_GVar_Head first_touched cur_base regionIdxCount tt_property_get scale_valid dummy1 numFDefs TT_SBit_MetricsRec FT_VOrg_Adjust_Func TT_Free_Table_Func Ins_DEPTH TT_Goto_CodeRange sph_fdef_flags glyphIns endCoord free_eblc ft_var_apply_tuple tt_default_graphics_state Ins_WCVTP tt_sfnt_id_rec_ defaultValue tt_interface vvar_checked avar_segment neg_jump_counter tt_hadvance_adjust subpixel_hinting Ins_Goto_CodeRange Ins_SPVTL Compute_Funcs FT_Set_Instance_Func Ins_RTDG TT_Err_Max func_move_cvt TT_Round_Func Ins_AND period TT_Get_VMetrics inc_stream pedantic_hinting callSize Ins_JROF TT_Set_Named_Instance majorVersion Round_Super_45 TT_Err_Cannot_Render_Glyph TT_Err_Could_Not_Find_Context has_delta TT_Err_Too_Many_Hints TT_Done_Face_Func tt_get_advances tt_size_request TT_Get_Name_Func mcvt_retain interpreter_version TT_Size_Metrics_ TT_Load_Table_Func TT_Driver multiplier GX_TupleIndexFlags_ Ins_UTP glyph_data_loaded num_matched_ids tt_synth_sfnt_checksum func_dualproj TT_Err_Invalid_Vert_Metrics orgs Direct_Move minimum_distance Direct_Move_Y Ins_SROUND mapCount ft_var_load_gvar GX_MVarTableRec_ tt_face_get_location Direct_Move_Orig_Y axisList axisScalar itemStore maxFunc callrec gep0 gep1 offsetToCoord FT_Set_Var_Design_Func valueCount runcnt tt_face_init cvt_ready FT_StreamRec Ins_SZPS only_height mac_yscale TT_Err_Raster_Negative_Height varRegionList Ins_LT tt_service_metrics_variations sfntd Ins_MIN tt_sfnt_id_rec pairCount num_instances TT_GraphicsState Ins_MD vorg_adjust TT_LoaderRec Fail_Overflow Ins_FLIPOFF TT_Err_Cannot_Open_Stream bsb_adjust FT_UnitVector_ Ins_SRP0 Ins_SRP1 Ins_SRP2 pindex TT_Load_Strike_Metrics_Func Ins_SxyTCA max_instruction_defs tt_get_interface FT_Get_Var_Blend_Func Ins_NEQ old_stream mvar_table deltas_y deltaSet TT_Run_Context axis_size Ins_NEG mmvar ft_var_get_item_delta load_truetype_glyph Move_Zp2_Point cur_delta Ins_MPPEM normalized_stylecoords TT_Get_HMetrics tt_check_trickyness Ins_GETDATA Ins_MAX use_aw_2 Ins_OR in_twilight FT_Var_Named_Style tt_property_set GX_ItemVarStore opened_frame size_metrics tmp_o TT_Get_CVT_Func TT_Err_Missing_Chars_Field FT_UnitVector FT_MM_Axis_ cvt_dist Direct_Move_Orig_X TT_Err_Too_Many_Caches ft_var_readpackedpoints fvar_start TT_Err_Cannot_Open_Resource maxIns ft_var_load_hvvar spoint_count Ins_RCVT context Ins_CINDEX ft_var_readpackeddeltas axis_rec next_coords num_designs grayscale_cleartype lsb_adjust new_dist ft_var_load_avar tsb_adjust Ins_POP num_base_points worker hvar_table vvar_loaded TT_Load_Composite_Glyph tt_size_done_bytecode TT_CallStack single_width_cutin Ins_ROFF FT_MM_Var peak FT_Service_TTGlyfRec_ num_base_subgs FT_TSB_Adjust_Func /home/computerfido/Desktop/freetypetest2/freetype/src/truetype/truetype.c TT_Save_Context Ins_RS GX_ItemVarDataRec_ peakCoord innerIndexMask Ins_MIAP set_design_coords _iup_worker_shift SkipCode TT_Load_Metrics_Func Ins_SCFS compensation x_ratio Dual_Project Current_Ratio linear_vadvance toCoord TT_Err_Code_Overflow TT_Err_Invalid_Stream_Seek TT_Err_Debug_OpCode TT_Set_CodeRange pedantic tt_loader_done ftsize FT_Int16 ft_var_to_design FT_Metrics_Adjust_Func func_freeProj tt_slot_init TT_Set_CVT_Func Ins_FLIPRGON Ins_MDAP FT_Done_Blend_Func FT_Service_TTGlyfRec num_records FT_MM_Axis TT_Err_Invalid_Size_Handle fvar_axis_ TT_Err_Invalid_PPem pointSize tmp_r TT_Err_Invalid_Post_Table_Format GX_AVarSegment TT_Init_Face_Func GX_Value TT_Load_SBit_Image_Func Current_Ppem_Stretched named_style tt_delta_interpolate widthp hvar_loaded auto_flip normalizedcoords widthMap FT_Get_MM_Func im_end_coords aRange sbit_metrics minValue num_instruction_defs TT_Err_Missing_Startchar_Field TT_Get_Var_Design gep2 TT_Err_Invalid_Cache_Handle tuplecount TT_Process_Composite_Glyph temp1 FT_Service_MetricsVariationsRec_ out_points cur_touched GX_FVar_Head_ Ins_SFVFS TT_Load_Glyph_Header GX_AVarCorrespondence offsetToData Ins_SPVFS Ins_SSWCI Ins_WS GX_ItemVarData FT_MM_Var_ FT_Multi_Master startCoord mcvt_load avar_loaded SFNT_Interface Ins_FLIPPT Ins_ROLL TT_Set_SBit_Strike_Func func_move TT_Err_Unknown_File_Format Ins_GETVARIATION GX_HVVarTable new_loca_len curRange maximum Ins_MUL scaledDelta linear_hadvance Ins_SxVTL TT_SBit_MetricsRec_ Ins_CALL TT_CodeRange storeSize LSuiteLabel_ func_move_orig Direct_Move_Orig tt_size_reset_iterator Cur_Count Ins_ALIGNPTS Project_y TT_Get_MM_Var have_diff Read_CVT_Stretched IUP_WorkerRec_ cvtSize TT_Err_Raster_Corrupted region_offset tt_get_sfnt_checksum mac_xscale max_func Ins_SLOOP ft_var_load_item_variation_store GX_TI_TUPLE_INDEX_MASK GX_TupleCountFlags_ axis_flags points_org maxValue gvar_fields delta_base callTop TT_New_Context tt_check_single_notdef axis_flags_size GX_ItemVarStoreRec TT_Load_Face_Func fvar_head mmvar_size Ins_GTEQ Ins_RDTG gvar_head TT_Err_Invalid_Handle here Ins_MINDEX GX_AVarSegmentRec_ orus1 orus2 Ins_LOOPCALL tt_metrics regionIndex stretched Ins_SDPVTL minimum recurse_count tt_get_metrics Ins_SCANTYPE GX_MVarTable TT_Err_Invalid_Composite gvar_start TT_DriverRec_ TT_Err_Invalid_Character_Code delta1 has_prep TT_Err_Nested_Frame_Access ttdriver ins_counter TT_Err_Nested_DEFS trick_names regionIndices Ins_FDEF TT_Err_Invalid_Frame_Operation mcvt_modify tt_size_done tt_coderange_glyph tt_face_load_cvt Ins_MIRP ttmetrics Ins_SDB FT_BSB_Adjust_Func Ins_SHPIX Write_CVT TT_Get_MM_Blend TT_Err_Too_Many_Instruction_Defs tt_face_done Ins_SDS next_name_size fromCoord Round_To_Half_Grid Ins_GC Ins_JROT tt_size_init_bytecode ft_var_load_delta_set_index_mapping Ins_ELSE TT_Err_Invalid_Stream_Handle freeVector tt_done_blend tt_coderange_none TT_Err_Too_Many_Extensions orus_base itemCount orig_cvt maxFDefs tuple_coords bytecode_ready tupleDataSize tt_service_truetype_engine byte_count TT_Err_Post_Table_Missing usePsName Ins_DUP Ins_ALIGNRP tt_delta_shift TT_Err_Missing_Property TT_Err_Array_Too_Large Move_CVT Ins_ROUND Bad_Format have_scale FT_Var_Axis TT_Process_Composite_Component scan_type TT_Move_Func globalCoordCount org_dist GX_FVar_Axis glyf_table_only TT_Err_Divide_By_Zero GX_GVar_Head_ tt_face_get_device_metrics TT_Err_Unlisted_Object tt_loader_init TT_Glyf_GetLocationFunc Ins_RUTG gvar_size tt_glyphzone_done loop TT_Err_Too_Few_Arguments ft_list_get_node_at IUP_WorkerRec entrySize tt_service_truetype_glyf hvar_checked Ins_SCVTCI ft_var_done_item_variation_store TT_Err_Invalid_Frame_Read Fail1 GridPeriod TT_GlyphZone Ins_GFV TT_Err_Invalid_Glyph_Index mmvar_len xy_size TT_Vary_Apply_Glyph_Deltas backward_compatibility tt_set_mm_blend num_twilight_points TT_Err_Invalid_Argument FT_Service_MultiMastersRec Read_CVT GX_ValueRec_ TT_Cur_Ppem_Func dataCount maxIDefs pCrec org1 FT_Var_Named_Style_ org2 FT_LSB_Adjust_Func TT_Err_No_Unicode_Glyph_Name Write_CVT_Stretched loopcall_counter hinted_metrics GX_AxisCoordsRec_ TT_MulFix14_long_long Ins_DELTAP TT_Err_Invalid_Outline unmodified TT_Hint_Glyph Pop_Push_Count old_byte_len GX_TI_EMBEDDED_TUPLE_COORD TT_Err_Missing_Size_Field num_namedstyles FT_RSB_Adjust_Func LErrorLabel_ dataOffsetArray TT_Done_Context records_offset compute_glyph_metrics mm_axis_unmap header_string T1_Err_Invalid_File_Format CFF_SubFontRec_ t1_services num_other_blues axis_count T1_Err_Ignore PS_GetFontInfoFunc local_subrs_offset t1_cmap_classes cff_decoder_funcs PSH_Globals PS_BlendRec_ PS_DICT_RND_STEM_UP PS_DICT_FONT_NAME sids T1_Err_Invalid_Composite T1_Err_Invalid_Vert_Metrics T1_Token T1_GlyphSlot PS_DICT_BLUE_SHIFT t1glyph top_font CFF_Builder_Add_Contour_Func units_per_em t1_get_name_index PS_DICT_ENCODING_ENTRY num_blue_values T1_FIELD_TYPE_NONE PSH_Globals_Funcs T1_FIELD_LOCATION_FACE T1_ParseState parser CFF_VarRegion num_hints incremental get_glyph_callback design_pos t1_ps_get_font_extra global_subrs_index num_strings AFM_FontInfo PS_Private T1_Driver_Done T1_Load_Glyph max_elems point_tokens T1_Err_Cannot_Open_Resource PS_DICT_OTHER_BLUE T1_Err_Too_Many_Extensions paint_type ps_parser_funcs T1_FontRec adobe_expert_encoding AFM_Parser_FuncsRec_ italic_angle code_last CFF_Size T1_Err_Corrupted_Font_Header T1_Err_DEF_In_Glyf_Bytecode PS_FontExtraRec T1_TokenRec_ T1_Builder_Check_Points_Func PS_DICT_SUBR PS_Parser_FuncsRec_ parse_blend_design_positions T1_Loader T2_HintsRec_ pos_lf CFF_SizeRec_ CFF_PrivateRec_ CFF_Decoder_FuncsRec CFF_Decoder_ font_offset t1_get_ps_name cid_uid_base global_subrs T1_Parse_Start T1_Err_Divide_By_Zero width_table_length parse_weight_vector FT_CMapRec PS_FontInfoRec_ PS_DICT_NUM_FAMILY_BLUES PS_DICT_WEIGHT parse_private T1_Err_Invalid_Glyph_Index PS_DICT_BLUE_VALUE charset_offset axiscoords single_block blue_scale PSH_Globals_SetScaleFunc T1_Err_Invalid_Stream_Skip T1_Err_Invalid_Offset PS_UniMap nominal_width PS_TableRec T1_FIELD_LOCATION_LOADER T1_Get_Var_Design keywords_encountered T1_FIELD_TYPE_MM_BBOX PS_DICT_FAMILY_OTHER_BLUE read_width PS_ParserRec_ PS_FontExtraRec_ T1_FIELD_TYPE_FIXED T1_Err_Invalid_Post_Table_Format the_same PS_Builder_FuncsRec char_string standard_height T1_ParserRec t1_decrypt T1_EncodingRecRec_ CFF_AxisCoords test_cr PS_Dict_Keys cid_count cid_ordering t1_make_subfont path_begun font_dict_index T1_TokenType t1_get_glyph_name lengths PS_DICT_NUM_OTHER_BLUES usedBV pos_x pos_y PS_DICT_FAMILY_NAME PS_DICT_STD_HW CFF_Font array_size lcoords vstore_offset in_memory afm_data t1_decoder_funcs t1_font PS_DICT_BLUE_FUZZ CFF_Decoder_Get_Glyph_Callback PS_GetGlyphNameFunc T1_FIELD_TYPE_FIXED_1000 private_size T1_Set_MM_Blend PS_GetFontValueFunc T1_Driver_Init token2 t1_ps_get_font_private T1_Err_Table_Missing hints_globals T1_Err_Too_Many_Function_Defs PS_DICT_UNDERLINE_THICKNESS T1_Err_Too_Many_Caches PS_DICT_PASSWORD string_pool private_len CFF_Builder_Start_Point_Func len_buildchar CFF_EncodingRec notdef_glyph parse_subrs T1_Err_ENDF_In_Exec_Stream AFM_ParserRec T1_Err_Too_Many_Hints T1_FIELD_TYPE_STRING cid_font_version T1_FIELD_TYPE_BOOL encoding_table T2_Hints_MaskFunc private_offset encode start_binary charstrings_offset T1_Err_Invalid_CharMap_Handle t1size PS_DICT_FORCE_BOLD FT_Service_KerningRec t1_builder_funcs swap_table have_integer T1_Err_Raster_Uninitialized T1_Err_Cannot_Render_Glyph T1_FIELD_TYPE_BBOX PS_Decoder_ lenIV vstore PS_UnicodesRec_ T1_DecoderRec ndv_idx strncmp PS_DICT_CHAR_STRING T1_Err_Too_Few_Arguments CFF_IndexRec CFF_SubFontRec T1_EncodingType T1_Err_Bad_Argument CFF_Decoder_FuncsRec_ blue_fuzz T1_Field off_size Again locals_bias FontBBox local_subrs_index T1_TOKEN_TYPE_NONE PS_DICT_NUM_CHAR_STRINGS T1_Face_Done T1_Decoder_Callback CFF_FDSelectRec T1_Reset_MM_Blend AFM_Parser T1_ENCODING_TYPE_ISOLATIN1 cid_registry t1_get_index num_locals T1_Field_ParseFunc cid_fd_array_offset glyph_names_block temp_scale T1_Decoder_ZoneRec T1_LoaderRec T1_Finalize_Parser T1_Err_Invalid_Argument is_t1 PSHinter_Service hintmask T1_Err_Invalid_Handle T1_Parse_Have_Width T1_Err_Invalid_CodeRange design_tokens PS_DICT_NOTICE T1_FIELD_LOCATION_BLEND t1_done_loader afont_extra T2_Hints_OpenFunc AFM_Stream globals_bias T1_Err_Missing_Startchar_Field T1_Err_Invalid_Version t1_service_properties force_scaling T1_Hints_SetStem3Func CFF_FDSelectRec_ PS_Table_FuncsRec CFF_FontRecDictRec start_pos PSH_Globals_DestroyFunc builtBV T2_Hints_Funcs initial_random_seed T1_Encoding PS_DICT_NUM_SUBRS T1_Err_Invalid_Stream_Handle lastVsindex n_axis pshinter T1_Compute_Max_Advance T1_Err_Invalid_Library_Handle T1_FIELD_LOCATION_FONT_EXTRA PS_PrivateRec FT_Service_PsCMaps T1_Err_Missing_Fontboundingbox_Field check_type1_format parse_callback parse_state width_only num_flex_vectors T1_EncodingType_ T2_Hints_FuncsRec_ T1_Err_Post_Table_Missing T1_FieldRec embedded_postscript PS_Decoder_Zone CFF_FontRecDictRec_ T1_Err_Invalid_Stream_Operation FT_Service_PsCMapsRec_ unique_id T1_Size T1_Err_Bbx_Too_Big T1_FIELD_TYPE_MAX range_count PS_DICT_PAINT_TYPE FT_Service_PsInfoRec_ charmaprecs t1_service_kerning PS_DICT_IS_FIXED_PITCH T1_FaceRec CFF_CharsetRec_ read_binary_data data_offset PS_Table_FuncsRec_ T1_Hints_ResetFunc CFF_BlendRec_ T1_Builder_Close_Contour_Func T1_FIELD_LOCATION_PRIVATE T1_Decoder_FuncsRec_ T2_Hints max_objects T1_Err_Horiz_Header_Missing no_recurse array_max cache_first blue_shift t1_set_mm_blend t1_parse_font_matrix T1_Err_Syntax_Error notice T1_Err_Stack_Overflow T1_BuilderRec_ synthetic_base T1_Err_Invalid_Frame_Read PS_DICT_ENCODING_TYPE glyph2 ident T1_Get_Kerning PS_DICT_MIN_FEATURE ps_table_funcs T1_Builder_Add_Point_Func flex_state PS_DICT_NUM_BLUE_VALUES T1_Err_Stack_Underflow T1_Err_Invalid_Size_Handle password T1_Hints T1_Read_Metrics T1_Builder_FuncsRec_ cache_fd T1_Decoder_ZoneRec_ notdef_found psdecoder T2_Hints_CloseFunc PS_DICT_NUM_STEM_SNAP_H t1_face PS_DICT_NUM_STEM_SNAP_V T1_Err_Out_Of_Memory T1_ParserRec_ PS_DesignMap_ num_elems T1_Err_Invalid_PPem T1_Err_Invalid_Slot_Handle T1_Err_Missing_Startfont_Field max_ptsize T1_Builder_Start_Point_Func round_stem_up PS_GetFontExtraFunc CFF_Builder_Close_Contour_Func PS_HasGlyphNamesFunc PS_Unicodes_CharIndexFunc T1_FieldLocation_ T1_GlyphSlot_Done custom count_offset T1_FontRec_ full_name T1_Err_Raster_Corrupted T1_Err_Code_Overflow CFF_Decoder T1_Err_Missing_Module T1_Get_MM_Blend CFF_Builder_Check_Points_Func num_snap_heights T1_Size_Request PS_DICT_FONT_BBOX T1_Err_Missing_Font_Field T1_ENCODING_TYPE_EXPERT T1_Font code_table T1_Err_Invalid_Reference subrs_block ps_decoder_init T1_Err_No_Unicode_Glyph_Name blend_top design_points T1_Err_Hmtx_Table_Missing adobe_std_strings T1_FieldLocation index1 index2 encoding_offset PS_Blend pair2 final_blends PS_Builder_FuncsRec_ T1_Err_Invalid_Driver_Handle t1_service_glyph_dict language_group CFF_VarRegion_ min_feature T1_FieldType_ glyph1 T1_Get_Private_Dict old_cursor T1_Err_Cannot_Open_Stream PS_DICT_FS_TYPE T1_Hints_Funcs T1_Decoder_Funcs adobe_std_encoding T1_Decoder_Zone cid_font_type CFF_Builder_ T1_Err_Invalid_Glyph_Format PSHinter_Interface T1_Get_Track_Kerning TrackKerns CFF_VarData_ PS_Macintosh_NameFunc default_weight_vector T1_BuilderRec T1_Hints_OpenFunc T1_Size_Get_Globals_Funcs PS_DesignMap PS_DICT_STEM_SNAP_H point_token T2_Hints_StemsFunc CFF_EncodingRec_ only_immediates CFF_Builder_FuncsRec PS_DICT_STEM_SNAP_V T1_Builder_FuncsRec cff_random T1_Set_MM_Design T1_Err_Invalid_Outline T1_TOKEN_TYPE_ARRAY PS_DICT_FAMILY_BLUE PS_Decoder_Zone_ bboxes afont_private T1_Parse_Glyph_And_Get_Char_String num_family_other_blues notdef_index PS_Adobe_Std_StringsFunc T1_Loader_ AFM_TrackKern T1_Err_Lower_Module_Version num_chars base_offset font_infos t1_allocate_blend num_default_design_vector CFF_Builder_Add_Point_Func current_subfont weight T1_TOKEN_TYPE_KEY T1_Decoder cid_supplement NumTrackKern T1_Err_Corrupted_Font_Glyphs CFF_SubFont T1_Get_Advances user_data midi CFF_GlyphSlotRec_ T1_Face_Init IsCIDFont fontdata T1_HintsRec_ CFF_PrivateRec code_first dummy_object T1_Err_Invalid_Table AFM_KernPairRec_ charstrings_block T1_Get_Multi_Master CFF_VarData CFF_Builder PSH_GlobalsRec_ T1_GlyphSlot_Init T1_Builder_Add_Point1_Func base_dict AFM_StreamRec_ T1_DecoderRec_ cffload atag blend_alloc T1_FIELD_TYPE_INTEGER hdr_size oldcharmap T1_Open_Face PS_FontInfo T2_Hints_ApplyFunc T1_Private charstrings_len T1_Get_MM_Var T1_Err_Could_Not_Find_Context T1_FIELD_LOCATION_CID_INFO PS_Builder T1_Err_Nested_Frame_Access cid_font_revision T1_Err_Nested_DEFS min_kern font_dict stroke_width cid_font_name PSAux_Service T1_ENCODING_TYPE_STANDARD AFM_KernPair T1_Parse_Have_Path T1_New_Parser t1_interface CFF_GlyphSlot subrs_len CFF_CharsetRec PSHinter_Interface_ PS_Table PS_Unicodes_CharNextFunc subrs_hash value_len_ CFF_IndexRec_ PS_TableRec_ __builtin_memcmp axis_token max_kern CFF_VStoreRec_ top_dict_index T1_Err_Ok blend_points PS_FreeGlyphNameFunc default_width T1_Done_Blend full PS_Decoder T1_TOKEN_TYPE_MAX gname T1_Size_Init axismap FT_Service_PsFontNameRec T1_Err_Debug_OpCode PS_DICT_VERSION PSH_Globals_FuncsRec_ T1_Err_Raster_Negative_Height CFF_Decoder_Zone_ PS_BlendRec T1_Hints_ApplyFunc num_snap_widths T1_EncodingRec locals_hash T1_FIELD_LOCATION_MAX p_design parse_blend_axis_types fs_type PS_DICT_LEN_IV T1_Err_Unknown_File_Format num_globals pair1 PS_DICT_LANGUAGE_GROUP char_name CFF_FontRec_ FT_Service_GlyphDictRec T1_Err_Missing_Size_Field KernPairs T1_ParseState_ T1_Err_Invalid_Character_Code PS_FontInfoRec min_ptsize PS_Unicodes_InitFunc T1_ENCODING_TYPE_NONE max_cid T1_Parse_Glyph T1_Err_Invalid_Cache_Handle axis_names parse_buildchar T2_Hints_CounterFunc T1_FaceRec_ T1_Err_Name_Table_Missing AFM_Parser_FuncsRec charstrings_index T1_Err_Invalid_Pixel_Size the_blend T1_FIELD_LOCATION_BBOX FT_GlyphSlotRec T1_Err_Raster_Overflow T1_Err_Missing_Bitmap base_len T1_CMap_Classes hints_funcs blend_bitflags T1_TOKEN_TYPE_ANY copyright t1_keywords T1_Err_Too_Many_Drivers header_length T1_FIELD_TYPE_FIXED_ARRAY T1_Err_Missing_Bbx_Field T1_TOKEN_TYPE_STRING T1_Err_Too_Many_Instruction_Defs CFF_BlendRec read_pfb_tag PS_Unicode_ValueFunc PS_Dict_Keys_ T1_Err_Missing_Chars_Field private_index T1_Read_PFM T1_SizeRec_ lenBV T1_Err_Execution_Too_Long force_bold num_subfonts t1_load_keyword T1_Err_Max T1_FieldRec_ afont_info T1_Size_Done T1_Err_Locations_Missing num_maps mmaster PS_DesignMapRec in_pfb T1_FIELD_LOCATION_FONT_INFO T1_FieldType encoding_type T1_Err_Invalid_Horiz_Metrics CFF_Builder_FuncsRec_ T1_TokenRec T1_Parser min_char num_family_blues PS_DICT_UNDERLINE_POSITION NumKernPair lenNDV PS_Parser_FuncsRec standard_width T1_FIELD_TYPE_INTEGER_ARRAY PS_DICT_MAX cache_count afm_parser_funcs T1_FIELD_TYPE_CALLBACK max_char T1_Err_Invalid_Post_Table old_limit T1_Hints_FuncsRec_ PSH_Globals_NewFunc PS_DICT_NUM_FAMILY_OTHER_BLUES T1_Builder PS_ParserRec T1_Parse_Have_Moveto t1_service_ps_name is_fixed_pitch PS_DICT_CHAR_STRING_KEY must_finish_decoder T1_Done_Metrics cid_fd_select_offset T1_GlyphSlotRec_ /home/computerfido/Desktop/freetypetest2/freetype/src/type1/type1.c retval PS_Unicodes T1_Err_Invalid_Frame_Operation T1_TokenType_ glyph_width blend_used T1_Err_Glyph_Too_Big force_bold_threshold PS_UniMap_ T1_Err_Invalid_Opcode PS_Builder_ header_size T1_Hints_SetStemFunc T1_Builder_Add_Contour_Func reader PS_PrivateRec_ cf2_instance t1_ps_get_font_info blend_stack T1_Err_Unlisted_Object cdv_idx FT_Service_PsInfoRec AFM_ParserRec_ value_len t1_service_ps_info T1_Decoder_FuncsRec CFF_Decoder_Free_Glyph_Callback PS_DICT_STD_VW T1_Err_Invalid_CharMap_Format T1_Err_Missing_Encoding_Field T1_Err_Unimplemented_Feature privates free_glyph_callback T1_Err_Invalid_Face_Handle PS_DICT_BLUE_SCALE has_font_matrix T1_Err_Invalid_Stream_Read fd_select T1_Err_Invalid_Stream_Seek T1_Err_Missing_Property parse_blend_design_map PS_DICT_UNIQUE_ID top_dict_length PS_GetFontPrivateFunc PS_DICT_FONT_MATRIX data_size CFF_VStoreRec PS_DICT_ITALIC_ANGLE T1_Err_Array_Too_Large CFF_Builder_Add_Point1_Func CFF_AxisCoords_ AFM_FontInfoRec_ locals_len T1_Hints_CloseFunc string_pool_size mm_weights_unmap T1_FIELD_LOCATION_FONT_DICT num_subrs metrics_only dummy T1_Face PSAux_ServiceRec_ PS_DICT_FULL_NAME T1_CMap_ClassesRec_ t1_ps_has_glyph_names local_subrs notdef_name T1_ENCODING_TYPE_ARRAY lastNDV T1_Set_Var_Design standard axis_tokens t1_service_multi_masters AFM_TrackKernRec_ CFF_Decoder_Zone t1_init_loader PS_Parser t1face T1_FIELD_TYPE_KEY t1_ps_get_font_value T1_Err_CMap_Table_Missing PS_DICT_FONT_TYPE FT_CMap_ClassRec Populate cff_hadvance_adjust CFF_Err_Too_Many_Hints cff_parse_vsindex CFF_Err_Nested_DEFS start_def FT_CID_GetIsInternallyCIDKeyedFunc CFF_Err_Bad_Argument CFF_FDSelect CFF_Err_Invalid_Stream_Operation cff_parse_font_matrix CFF_Err_Invalid_Frame_Operation cff_get_kerning FT_Blend_Build_Vector_Func CFF_Parser CFF_Err_Invalid_Opcode exponent_sign have_overflow CFF_Err_Too_Many_Instruction_Defs start14 cff_parse_fixed cff_service_get_cmap_info num_ranges CFF_InternalRec_ pbyte_len cff_charset_cid_to_gindex cff_get_cid_from_glyph_index FT_CID_GetRegistryOrderingSupplementFunc numOperands CFF_Err_Missing_Property cff_make_private_dict cff_vstore_done CFF_Err_Invalid_CharMap_Handle CFF_Err_Invalid_Reference CFF_Load_FD_Select cff_get_var_design cff_cmap_unicode_class_rec qcount subFont cff_service_ps_info invert Store_Number cff_face_done csindex cff_get_glyph_data CFF_Err_No_Unicode_Glyph_Name cff_sid_to_glyph_name sub_upm sfnt_module CFF_Err_Invalid_Vert_Metrics CFF_Err_Invalid_CharMap_Format CFF_FontRec cff_field_handlers cff_service_cff_load cmaprec next_offset cff_kind_fixed_thousand CFF_Err_Invalid_Frame_Read cff_size_done cff_blend_build_vector FT_Service_TTCMapsRec glyph_sid CFF_Err_Too_Many_Function_Defs cff_set_mm_blend cff_kind_max end14 cff_parse_private_dict CFF_FontRecDict CFF_Err_Missing_Size_Field pchar_code CFF_Err_Missing_Bbx_Field CFF_Private CFF_Err_Invalid_Stream_Seek cff_encoding_done CFF_Err_Invalid_Size_Handle cff_load_private_dict CFF_Err_Invalid_Face_Handle cff_fd_select_get FT_Service_MultiMasters cff_font_done CFF_VStore CFF_Err_Missing_Font_Field power_ten_limits CFF_Charset cffslot CFF_Err_CMap_Table_Missing CFF_ParserRec cff_cmap_encoding_done cff_size_request cff_get_mm_var FT_Service_CFFLoadRec_ CFF_Err_Debug_OpCode CFF_Err_Name_Table_Missing org_bytes cff_charset_done cff_get_ps_name CFF_Err_Invalid_File_Format cff_parse_fixed_dynamic cff_cmap_encoding_class_rec cff_get_advances FT_FD_Select_Get_Func cff_service_multi_masters cff_index_get_pointers CFF_Field_Reader FT_Service_CIDRec CFF_Err_Invalid_Library_Handle CFF_ParserRec_ cff_blend_doBlend CFF_Err_Lower_Module_Version remove_style p_end CFF_Err_Hmtx_Table_Missing topfont poff cff_kind_fixed style_name_length cff_size_get_globals_funcs CFF_Err_Raster_Overflow power_ten CFF_Err_Table_Missing CFF_Err_Too_Few_Arguments cff_parser_run errorp min_scaling cff_service_ps_name cff_get_ros CFF_Err_Invalid_Composite cff_index_get_name CFF_Err_Invalid_Driver_Handle cff_size_init CFF_Err_Cannot_Open_Stream cff_header_fields cff_kind_bool cff_parse_real FT_Service_CFFLoadRec cff_cmap_encoding_init CFF_Err_Invalid_CodeRange CFF_Err_Cannot_Open_Resource cff_service_properties CFF_Err_Array_Too_Large FT_CID_GetCIDFromGlyphIndexFunc CFF_Err_Invalid_Handle sfnt_format new_bytes CFF_Field_Handler_ cff_cmap_unicode_init CFF_Err_Unlisted_Object peak14 cffface cff_parser_done CFF_Index cff_get_mm_blend cff_isoadobe_charset vsOffset cff_services CFF_Err_Missing_Encoding_Field CFF_Err_Missing_Startchar_Field CFF_Field_Handler fullp regionListOffset blend_top_old CFF_Err_Corrupted_Font_Glyphs numBlends family_name_length CFF_Err_Corrupted_Font_Header CFF_Err_Ok cff_slot_init cff_blend_clear cff_set_var_design Missing_Table CFF_Err_Invalid_Slot_Handle CFF_Err_Invalid_Outline cur_offset CFF_Err_Locations_Missing CFF_Err_Too_Many_Drivers CFF_Err_Invalid_Post_Table FT_Blend_Check_Vector_Func exponent_add blend_stack_old CFF_Blend cff_get_interface CFF_Err_Ignore cff_index_forget_element CFF_Err_Stack_Underflow cff_size_select CFF_Err_Execution_Too_Long CFF_Err_Invalid_Offset CFF_Err_Horiz_Header_Missing charstring_len CFF_Err_Post_Table_Missing cff_free_glyph_data half_divisor num_args subfont_index CFF_Err_Syntax_Error FT_Load_Private_Dict_Func region cff_get_is_cid max_scaling top_upm glyph_code integer_length cff_kind_num cff_expert_encoding CFF_Encoding cff_index_init string_index CFF_Err_Invalid_Table cff_parse_maxstack CFF_Done_FD_Select cff_get_cmap_info CFF_Err_Invalid_PPem FT_Get_Standard_Encoding_Func CFF_Face CFF_Err_Raster_Uninitialized cff_service_metrics_variations cff_ps_get_font_info cpriv cff_vstore_load CFF_Err_Missing_Bitmap Skip_Unicode CFF_Err_ENDF_In_Exec_Stream CFF_Err_Invalid_Stream_Read cff_cmap_encoding_char_index /home/computerfido/Desktop/freetypetest2/freetype/src/cff/cff.c varRegion cff_parse_blend cff_ps_has_glyph_names CFF_Err_Invalid_Pixel_Size cff_index_access_element cff_parse_multiple_master do_fixed cff_kind_string CFF_Err_Too_Many_Caches cff_index_done CFF_Err_Code_Overflow CFF_Err_Invalid_Horiz_Metrics CFF_Err_Invalid_Argument cff_get_name_index CFF_Err_Invalid_Cache_Handle continue_search CFF_Err_Raster_Negative_Height CFF_Err_Missing_Chars_Field dict_len cff_driver_done cff_slot_load CFF_Err_DEF_In_Glyf_Bytecode cff_get_var_blend CFF_Err_Invalid_Character_Code cff_get_standard_encoding gids cff_expertsubset_charset CFF_Err_Invalid_Glyph_Format CFF_Err_Out_Of_Memory cff_blend_check_vector CFF_Err_Bbx_Too_Big fdselect CFF_Err_Raster_Corrupted cff_expert_charset scalings CFF_Err_Invalid_Stream_Handle CFF_Err_Unimplemented_Feature cff_index_get_string cff_metrics_adjust cff_charset_free_cids cff_ps_get_font_extra CFF_Err_Could_Not_Find_Context CFF_Err_Invalid_Version Glyph_Build_Finished cff_parse_integer cff_subfont_load cff_cmap_encoding_char_next exponent cff_cmap_unicode_char_index remove_subset_prefix CFF_Decoder_Funcs pure_cff cff_glyph_load kind cff_done_blend cff_subfont_done CFF_Err_Stack_Overflow has_vertical_info cff_kind_callback CFF_Err_Invalid_Glyph_Index cff_get_glyph_name CFF_Err_Unknown_File_Format absolute_offset object_code cff_encoding_load CFF_Err_Invalid_Stream_Skip nleft cff_index_get_sid_string offsize CFF_Err_Invalid_Post_Table_Format cff_slot_done cff_face cff_kind_blend cff_parse_num CFF_Err_Glyph_Too_Big cff_cmap_unicode_done cffsize cff_parser_init fd_index CFF_Err_Divide_By_Zero cff_cmap_unicode_char_next cff_font_load cff_parse_fixed_scaled Load_Data CFF_Err_Missing_Fontboundingbox_Field cff_kind_delta start_fstype cff_index_load_offsets cff_parse_font_bbox cff_charset_compute_cids cff_standard_encoding CFF_Err_Max CFF_CMapStdRec_ new_fraction_length Fail_CID cff_service_cid_info cff_charset_load CFF_Err_Missing_Startfont_Field cff_set_instance CFF_Err_Nested_Frame_Access CFF_Err_Missing_Module cff_strcpy cff_driver_init FT_Service_CFFLoad cff_parse_cid_ros FT_Service_MetricsVariations power_tens CFF_Internal cff_index_read_offset FT_Service_CIDRec_ cff_face_init cff_service_glyph_dict CFF_CMapStd CFF_Err_Cannot_Render_Glyph CFF_Err_Too_Many_Extensions cff_kind_none fd_bytes max_offsets cid_face_open CID_Err_ENDF_In_Exec_Stream cid_get_offset gd_bytes CID_Parser CID_Err_Invalid_Frame_Operation CID_Err_Stack_Underflow CID_Err_Invalid_CharMap_Format CID_Err_Invalid_CodeRange CID_Err_Glyph_Too_Big CID_Err_Hmtx_Table_Missing CID_Err_Missing_Chars_Field num_dict CID_Err_Missing_Property cid_size_request CID_Err_Code_Overflow CID_FaceDictRec_ CID_FaceInfoRec_ CID_Err_Raster_Uninitialized upper_nibble CID_Err_Horiz_Header_Missing subrmap_offset CID_Parser_ cid_done_loader CID_Loader CID_FaceDictRec CID_Err_Invalid_Stream_Seek cid_slot_load_glyph CID_Err_Raster_Overflow CID_Err_Missing_Size_Field CID_Err_Invalid_Stream_Operation cid_service_cid_info cid_subrs CID_Err_Invalid_Pixel_Size CID_Err_Missing_Bbx_Field /home/computerfido/Desktop/freetypetest2/freetype/src/cid/type1cid.c CID_Err_Too_Many_Hints CID_Err_Missing_Fontboundingbox_Field CID_Err_Unknown_File_Format glyph_length CID_Err_Unlisted_Object CID_GlyphSlot CID_Err_Missing_Font_Field cid_driver_done cidface CID_Err_Unimplemented_Feature CID_Err_Table_Missing CID_Err_Invalid_Cache_Handle CID_Err_Invalid_Face_Handle CID_Face cidglyph cid_hex_to_binary CID_Err_Invalid_Outline cid_slot_done cid_version cid_face_done CID_Err_Invalid_Glyph_Format cid_services CID_Size CID_Err_Ignore cid_service_ps_name CID_Err_Invalid_Post_Table CID_Err_Corrupted_Font_Header cid_parse_font_matrix CID_Err_Too_Many_Extensions CID_Err_Could_Not_Find_Context CID_Err_DEF_In_Glyf_Bytecode newlimit cid_interface CID_Err_Post_Table_Missing dlimit CID_Err_Invalid_Handle cid_driver_init CID_Err_Raster_Negative_Height CID_Err_Divide_By_Zero CID_Err_No_Unicode_Glyph_Name CID_Err_Invalid_Stream_Handle font_dicts CID_Err_Invalid_Character_Code CID_Err_Lower_Module_Version binary_length CID_Err_Too_Many_Caches CID_Err_Invalid_Offset CID_Err_Max CID_Err_Ok CID_Err_Invalid_Library_Handle cid_get_interface CID_Err_Invalid_Reference CID_FaceInfo CID_Err_Too_Few_Arguments CID_Err_Too_Many_Drivers CID_SizeRec_ cid_get_ros CID_Err_Invalid_Opcode CID_Err_Stack_Overflow CID_FaceInfoRec CID_Err_Too_Many_Instruction_Defs forcebold_threshold CID_GlyphSlotRec_ CID_Err_Invalid_Composite CID_FaceDict CID_SubrsRec_ cid_ps_get_font_info cid_parser_done CID_Err_Name_Table_Missing CID_Err_Invalid_Version CID_Err_Bbx_Too_Big CID_Err_Missing_Module CID_Loader_ cid_ps_get_font_extra CID_Err_Out_Of_Memory cid_service_ps_info cid_load_glyph CID_Err_Debug_OpCode CID_Err_Raster_Corrupted CID_Err_Missing_Startfont_Field cid_load_keyword oldpos CID_Subrs CID_Err_Invalid_File_Format CID_Err_Nested_Frame_Access plimit cidsize CID_Err_Nested_DEFS cid_size_get_globals_funcs CID_Err_Bad_Argument cid_slot_init CID_Err_Invalid_Argument CID_Err_Missing_Encoding_Field cid_get_cid_from_glyph_index CID_Err_Invalid_Size_Handle read_len CID_Err_Cannot_Render_Glyph CID_Err_Invalid_Vert_Metrics CID_Err_Invalid_Horiz_Metrics sd_bytes num_dicts parse_expansion_factor cid_size_done cidmap_offset cid_get_postscript_name CID_Err_Invalid_Stream_Read CID_Err_Invalid_Glyph_Index CID_Err_Corrupted_Font_Glyphs CID_Err_Invalid_Stream_Skip CID_Err_Execution_Too_Long CID_Err_Invalid_Post_Table_Format CID_Err_Invalid_Table postscript_len CID_Err_Syntax_Error CID_Err_Invalid_CharMap_Handle cid_size_init ps_len CID_Err_Invalid_Slot_Handle parse_fd_array cid_field_records cid_get_is_cid CID_Err_Invalid_PPem CID_Err_Invalid_Frame_Read cid_stream stream_len CID_Err_Missing_Bitmap CID_Err_Too_Many_Function_Defs CID_Err_Invalid_Driver_Handle CID_Err_Array_Too_Large CID_Err_Cannot_Open_Resource CID_FaceRec_ CID_Err_Missing_Startchar_Field entry_len cid_service_properties CID_Err_Cannot_Open_Stream CID_Err_Locations_Missing cid_parse_dict cid_init_loader num_xuid CID_Err_CMap_Table_Missing cid_read_subrs cid_face_init cid_parser_new log_font bct_offset PFR_Err_Out_Of_Memory PFR_Err_Cannot_Render_Glyph PFR_Err_Missing_Startchar_Field base_adj num_items PFR_HeaderRec size1 pfr_cmap_done stroke_flags Found_Strike PFR_Err_Raster_Corrupted Failure PFR_Err_Name_Table_Missing phy_font_max_size phy_font_section_offset phys_offset acount PFR_Err_Missing_Property PFR_Err_Missing_Startfont_Field PFR_Err_Invalid_Driver_Handle max_subs pfr_phy_font_load PFR_Err_Invalid_Horiz_Metrics local gps_section_offset kern_items pfr_face_done aformat PFR_Err_Unimplemented_Feature FT_PFR_GetMetricsFunc PFR_LogFontRec num_vert num_log_fonts PFR_ExtraItem_ParseFunc char1 char2 pair_count bct_max_size PFR_Err_Missing_Chars_Field PFR_Err_Too_Few_Arguments prev_code twobytes PFR_Err_Unlisted_Object pdata axsize pfr_get_kerning log_font_section_size PFR_Err_Divide_By_Zero PFR_Err_Ok item_list pfr_metrics_service_rec PFR_Err_Invalid_Cache_Handle item_data pfr_cmap_char_next PFR_Err_Invalid_Reference pfr_extra_item_load_bitmap_info PFR_Err_Invalid_CharMap_Format PFR_Err_Invalid_File_Format log_font_max_size PFR_Err_Horiz_Header_Missing PFR_Err_Invalid_Face_Handle pfr_glyph_curve_to pfr_glyph_end PFR_Err_Max PFR_BitWriter_ PFR_Err_Too_Many_Function_Defs max_horz_stem_snap found_offset chars_offset PFR_SubGlyphRec_ PFR_Err_Invalid_Stream_Skip twobyte_adj stroke_thickness phys PFR_ExtraItem y_count pfr_glyph_load_simple pfr_glyph_close_contour old_points pfr_face_init PFR_DimensionRec_ ametrics_y_scale anadvance PFR_Err_CMap_Table_Missing font_ref_number PFR_Err_Too_Many_Caches log_dir_offset color_flags PFR_DimensionRec item_type PFR_Err_DEF_In_Glyf_Bytecode num_bitmaps PFR_Err_Corrupted_Font_Glyphs pair_size y_ppm PFR_Err_Missing_Fontboundingbox_Field Line1 pfr_extra_items_parse pfr_cmap_init PFR_Err_Missing_Encoding_Field PFR_BitWriter PFR_Err_Hmtx_Table_Missing pfr_get_metrics em_metrics max_xy_control PFR_Glyph FT_Service_PfrMetricsRec pfr_bitwriter_init anoutline_resolution PFR_BitmapCharRec_ pfr_extra_item_load_stem_snaps pfr_glyph_start writer PFR_Err_Invalid_Version phy_font Test_Error PFR_SubGlyphRec y_delta phy_bct_set_max_size PFR_CMapRec_ pfrsize max_y_orus PFR_Err_Lower_Module_Version PFR_Err_Cannot_Open_Stream PFR_Err_Invalid_Table bct_size probe FT_PFR_GetKerningFunc PFR_Err_Invalid_Slot_Handle PFR_BitWriterRec PFR_Err_Unknown_File_Format PFR_Err_Invalid_Stream_Read PFR_Err_Too_Many_Hints PFR_SubGlyph max_vert_stem_snap PFR_ExtraItemRec PFR_Err_Stack_Underflow kern_items_tail pfr_phy_font_done PFR_Err_Debug_OpCode standard_advance PFR_Header em_outline pfrface num_kern_pairs PFR_LogFont PFR_Char pfr_header_load pfr_face_get_kerning phy_font_max_size_high PFR_Err_Missing_Size_Field pfr_header_check pfr_cmap_class_rec Too_Short PFR_PhyFontRec_ pfr_glyph_move_to format_low pfr_glyph_load decreasing PFR_Err_Execution_Too_Long PFR_Err_Invalid_Composite PFR_Err_Invalid_Size_Handle gps_max_size char_len PFR_Err_Table_Missing num_aux FoundPair gps_offset pfr_glyph_done PFR_Err_Raster_Overflow PFR_Err_Invalid_Frame_Operation PFR_Err_Missing_Bbx_Field PFR_Err_Nested_DEFS pfr_get_service PFR_Err_Invalid_Vert_Metrics signature2 PFR_Err_Invalid_PPem PFR_Size PFR_Err_Code_Overflow PFR_Err_Invalid_Post_Table x_ppm PFR_StrikeRec ametrics_x_scale pfr_services miter_limit found_size pfr_phy_font_extra_items avector PFR_Err_Invalid_Post_Table_Format control1 control2 PFR_KernItem PFR_Err_Ignore PFR_KernItemRec_ PFR_Err_Invalid_Offset PFR_Err_Raster_Negative_Height Restart power PFR_Err_Invalid_Stream_Operation PFR_Face PFR_Err_No_Unicode_Glyph_Name PFR_SizeRec_ PFR_Err_Invalid_CodeRange PFR_StrikeRec_ PFR_Err_Stack_Overflow pfrslot PFR_Err_Bad_Argument size_increment PFR_Err_Glyph_Too_Big pfr_cmap_char_index PFR_Err_Nested_Frame_Access PFR_Err_Invalid_Outline pfr_extra_items_skip PFR_Strike PFR_Err_Missing_Bitmap PFR_Err_Invalid_Handle PFR_Err_Array_Too_Large flags0 PFR_Err_Too_Many_Extensions PFR_LogFontRec_ FT_PFR_GetAdvanceFunc org_count PFR_ExtraItemRec_ PFR_Err_Corrupted_Font_Header PFR_Err_Syntax_Error Found_It log_font_section_offset PFR_Err_Invalid_Frame_Read scaled_advance pfr_get_advance PFR_Err_Invalid_Opcode PFR_SlotRec_ PFR_Err_Invalid_Glyph_Format pfr_slot_done PFR_BitmapChar ametrics_resolution PFR_Err_Invalid_Glyph_Index PFR_Err_Too_Many_Instruction_Defs pfr_extra_item_load_kerning_pairs axpos PFR_Err_Bbx_Too_Big num_phy_fonts pfr_lookup_bitmap_data PFR_GlyphRec_ aadvance PFR_HeaderRec_ args_format phy_font_section_size astring PFR_CMap PFR_Err_Missing_Module max_x_orus max_blue_values gchar y_pos PFR_Err_Missing_Font_Field PFR_Slot PFR_Err_Locations_Missing PFR_Err_Invalid_Argument phys_size num_stem_snaps gps_section_size cpair pfr_log_font_count PFR_Err_ENDF_In_Exec_Stream signature pfr_bitwriter_decode_bytes pfr_glyph_line_to num_horz PFR_GlyphRec pfr_load_bitmap_metrics PFR_Err_Invalid_Stream_Seek pfr_slot_load max_strikes counts pfr_log_font_load pfr_slot_load_bitmap PFR_Err_Invalid_Character_Code PFR_FaceRec_ pfr_bitwriter_decode_rle2 PFR_Err_Post_Table_Missing pfr_header_fields aypos pfr_slot_init old_count PFR_Err_Cannot_Open_Resource FT_Service_PfrMetricsRec_ PFR_Err_Invalid_CharMap_Handle PFR_Err_Invalid_Pixel_Size PFR_PhyFont PFR_Err_Invalid_Stream_Handle PFR_PhyFontRec pfr_glyph_load_rec pfr_aux_name_load num_subs pfr_glyph_init PFR_Err_Raster_Uninitialized PFR_Err_Could_Not_Find_Context pfr_glyph_load_compound PFR_Err_Invalid_Library_Handle pfr_bitwriter_decode_rle1 character pfr_load_bitmap_bits gps_size bold_thickness aysize log_dir_size /home/computerfido/Desktop/freetypetest2/freetype/src/pfr/pfr.c PFR_CharRec_ x_control max_chars PFR_Err_Too_Many_Drivers pfr_extra_item_load_font_id t42_get_ps_font_name T42_GlyphSlot real_size T42_Err_DEF_In_Glyf_Bytecode t42_ps_has_glyph_names t42_services T42_Driver_Init T42_Size_Select T42_Err_Nested_DEFS T1_FontInfo T42_Err_Unknown_File_Format T42_Err_Post_Table_Missing T42_Err_Missing_Startchar_Field t42_ps_get_font_private t42_loader_done T42_Err_Invalid_Cache_Handle T42_Err_Unimplemented_Feature T42_Face_Init t42_parse_font_matrix T42_Err_Invalid_Frame_Read T42_Err_Invalid_Glyph_Format T42_Err_Lower_Module_Version T42_Err_Nested_Frame_Access T42_Open_Face T42_Err_Missing_Size_Field T42_Err_Invalid_Version t42_interface T42_Err_Out_Of_Memory t42_service_ps_font_name T42_Err_Cannot_Render_Glyph T42_Err_Missing_Property ttclazz T42_Parser T42_Err_Invalid_Frame_Operation T42_ParserRec t42_service_ps_info T42_Size_Init T42_Load_Status_ T42_Err_Invalid_Stream_Handle T42_Err_Invalid_Handle T42_Err_Name_Table_Missing t42_parse_dict T42_GlyphSlotRec_ ttf_size T42_Err_Invalid_Stream_Skip T42_Err_Missing_Fontboundingbox_Field t42_get_glyph_name status T42_Loader BEFORE_START T42_Size T42_Err_Divide_By_Zero T42_Err_CMap_Table_Missing T42_Err_Hmtx_Table_Missing T42_Err_Ignore T42_Err_Invalid_Vert_Metrics /home/computerfido/Desktop/freetypetest2/freetype/src/type42/type42.c T42_Err_Invalid_CharMap_Handle T42_LoaderRec T42_Err_Invalid_Table unicode_map t42size t42_service_glyph_dict T42_Err_Invalid_Glyph_Index T42_Err_Stack_Underflow ttf_face T42_Err_Raster_Overflow T42_Err_Missing_Module t42_loader_init T42_Loader_ T42_Get_Interface T42_Err_Invalid_Stream_Seek T42_DriverRec_ t42_parse_sfnts T42_Err_Could_Not_Find_Context T42_Err_Invalid_Face_Handle T42_Err_Array_Too_Large T42_Err_No_Unicode_Glyph_Name T42_Err_Unlisted_Object T42_Err_Invalid_Offset T42_Err_Invalid_Post_Table_Format T42_Err_Raster_Negative_Height T42_GlyphSlot_Init T42_Err_Invalid_Reference T42_Err_Invalid_File_Format T42_Err_Execution_Too_Long T42_Err_Table_Missing T42_Err_Invalid_Character_Code T42_Err_Invalid_Horiz_Metrics T42_Err_Invalid_Outline have_literal T42_Err_Debug_OpCode t42face OTHER_TABLES PS_UnicodesRec T42_Err_Missing_Startfont_Field t42_parser_done T42_Err_Invalid_Library_Handle T42_Err_Bbx_Too_Big T42_Err_Invalid_Post_Table T42_Driver t42_ps_get_font_info T42_Err_Missing_Bbx_Field T42_Load_Status T42_Err_Cannot_Open_Resource T42_FaceRec_ T42_GlyphSlot_Done T42_Err_Glyph_Too_Big T42_Err_Too_Many_Drivers T42_Err_Invalid_Stream_Operation T42_Err_Invalid_Pixel_Size T42_Err_Syntax_Error T42_Err_Code_Overflow T42_SizeRec_ t42_load_keyword string_buf t42slot T42_Err_Corrupted_Font_Header t42_is_space T42_Err_Invalid_PPem ttf_data T42_Err_Bad_Argument T42_Err_Invalid_Driver_Handle T42_Err_Too_Many_Caches t42_get_name_index T42_Err_Invalid_Slot_Handle T42_Err_ENDF_In_Exec_Stream ttmodule T42_Err_Raster_Corrupted T42_Err_Ok T42_ParserRec_ T42_Err_Cannot_Open_Stream T42_Err_Invalid_Opcode T42_Err_Too_Few_Arguments T42_Err_Missing_Bitmap t42_parser_init t42_ps_get_font_extra T42_Err_Raster_Uninitialized T42_Err_Corrupted_Font_Glyphs t42_parse_charstrings T42_Err_Invalid_Argument T42_Err_Horiz_Header_Missing T42_Err_Invalid_CodeRange T42_Err_Invalid_Composite T42_Err_Max T42_Err_Too_Many_Extensions n_keywords t42_parse_encoding T42_Face T42_Err_Missing_Encoding_Field T42_Size_Done T42_Driver_Done T42_Err_Locations_Missing T42_Err_Invalid_Stream_Read t42_keywords T42_Face_Done BEFORE_TABLE_DIR T42_Size_Request t42_glyphslot_clear old_string_size T42_GlyphSlot_Load T42_Err_Too_Many_Hints T42_Err_Missing_Chars_Field T42_Err_Stack_Overflow T42_Err_Invalid_CharMap_Format T42_Err_Too_Many_Function_Defs T42_Err_Too_Many_Instruction_Defs T42_Err_Invalid_Size_Handle T42_Err_Missing_Font_Field WinPE_RsrcDirEntryRec WinNE_HeaderRec_ winpe_rsrc_dir_entry_fields fntface /home/computerfido/Desktop/freetypetest2/freetype/src/winfonts/winfnt.c bits_offset dir_entry2 dir_entry3 WinMZ_HeaderRec_ WinPE_RsrcDirEntryRec_ root_dir FNT_Face_Done ne_header first_char A_space type_id aheader FNT_Size_Select pitch_and_family size_shift pe32_header WinMZ_HeaderRec bytes_per_row rsrc_virtual_address last_char winne_header_fields WinPE32_HeaderRec_ column new_format FT_Service_WinFntRec FNT_Face_Init winpe32_header_fields WinPE32_SectionRec FT_WinFNT_HeaderRec nominal_point_size face_instance_index fnt_font_done italic B_space fnt_font_load FNT_CMap magic32 winpe32_section_fields winmz_header_fields FT_WinFnt_GetHeaderFunc strike_out fnt_cmap_char_next Found_rsrc_section charmap_handle x_res lang_dir_offset root_dir_offset characteristics WinPE32_SectionRec_ rname_tab_offset winpe_rsrc_dir_fields WinPE_RsrcDirRec number_of_named_entries winpe_rsrc_data_entry_fields FT_Service_WinFntRec_ time_date_stamp rsrc_size C_space FT_WinFNT_HeaderRec_ name_dir color_table_offset WinPE32_HeaderRec FNT_Size_Request default_char winfnt_service_rec resource_tab_offset number_of_id_entries avg_width fnt_frame WinPE_RsrcDirRec_ WinPE_RsrcDataEntryRec internal_leading size_of_optional_header FNT_FontRec_ code_page horizontal_resolution pe32_section dir_entry1 winfnt_services device_offset offset_to_data FNT_CMapRec_ mz_header name_dir_offset WinNE_HeaderRec fnt_cmap_init WinPE_RsrcDataEntryRec_ FNT_FaceRec_ file_type major_version fnt_cmap_char_index winfnt_get_service external_leading fnt_face_get_dll_font bits_pointer fnt_cmap_class_rec res_offset family_size minor_version winfnt_header_fields fnt_cmap_class pointer_to_raw_data reserved1 fnt_size size_of_raw_data number_of_sections FNT_Load_Glyph data_entry break_char winfnt_get_header FT_WinFNT_Header vertical_resolution lfanew FNT_Font FNT_Face machine underline lang_dir y_res face_name_offset PCF_Err_Horiz_Header_Missing drawDirection pcfcmap FT_Stream_OpenLZW PCF_Err_Invalid_Stream_Read PCF_ParseProperty pcf_table_header PCF_ParsePropertyRec num_encodings BDF_PropertyRec_ PCF_Err_Glyph_Too_Big fontDescent pcf_read_TOC PCF_Err_Invalid_Library_Handle PCF_Face_Done orig_nprops PCF_Err_Unimplemented_Feature PCF_Err_Invalid_Stream_Operation pcf_load_font pcf_service_bdf PCF_Err_Code_Overflow pcf_cmap_char_index PCF_Err_Missing_Chars_Field PCF_Err_Invalid_CharMap_Format PCF_Err_Invalid_Reference acharset_registry ink_maxbounds PCF_Err_Invalid_Frame_Operation pcfface PCF_Encoding PCF_Err_Missing_Fontboundingbox_Field PCF_Toc pcf_seek_to_table_type ntables PCF_Err_Invalid_Character_Code PCF_TableRec_ PCF_Err_Ok PCF_Err_Stack_Overflow PCF_CMap pcf_driver_done constantWidth nbytes /home/computerfido/Desktop/freetypetest2/freetype/src/pcf/pcf.c PCF_Err_Invalid_Slot_Handle PCF_Err_Out_Of_Memory BDF_PROPERTY_TYPE_ATOM PCF_ParsePropertyRec_ PCF_Err_Invalid_Stream_Skip pcf_metric_header TwoByteSwap FourByteSwap PCF_Err_CMap_Table_Missing pcf_cmap_init PCF_Err_Divide_By_Zero PCF_Err_Invalid_Vert_Metrics hasBDFAccelerators PCF_Err_Invalid_Frame_Read sizebitmaps inkInside PCF_Err_Post_Table_Missing PCF_Err_ENDF_In_Exec_Stream isString PCF_Err_Invalid_Version PCF_Err_Invalid_CodeRange PCF_Err_Too_Many_Caches pcf_get_metrics PCF_Size_Request PCF_Err_Invalid_Size_Handle PCF_Err_Syntax_Error PCF_Err_Cannot_Open_Resource PCF_Size_Select pcf_property_msb_header pcf_property_header PCF_Err_Bad_Argument PCF_Err_Invalid_Table pcf_driver_requester PCF_Err_Too_Many_Function_Defs pcf_service_properties pcf_driver_init terminalFont PCF_TocRec_ PCF_Err_Stack_Underflow PCF_Err_Debug_OpCode pcf_find_property PCF_Err_Unlisted_Object PCF_Err_Invalid_Driver_Handle PCF_Err_Missing_Size_Field defaultChar PCF_AccelRec_ PCF_Err_Locations_Missing pcf_cmap_done firstCol PCF_Compressed_MetricRec PCF_Err_Invalid_Outline nencodings Bail PCF_Err_Name_Table_Missing PCF_Err_DEF_In_Glyf_Bytecode PCF_Err_Too_Many_Instruction_Defs PCF_Err_Nested_Frame_Access PCF_Err_Too_Few_Arguments PCF_Err_Cannot_Open_Stream PCF_Err_Invalid_Pixel_Size PCF_Err_Missing_Startfont_Field PCF_Face fontAscent PCF_TocRec PCF_Err_Raster_Overflow inkMetrics resolution_y PCF_FaceRec_ error3 pcf_accel_header PCF_TableRec PCF_Err_No_Unicode_Glyph_Name PCF_Err_Ignore PCF_Err_Missing_Font_Field PCF_Err_Bbx_Too_Big PCF_Err_Raster_Corrupted PCF_Err_Execution_Too_Long PCF_Err_Invalid_Glyph_Index FT_BDF_GetPropertyFunc bitmapSizes PCF_Err_Raster_Negative_Height PCF_Property BitOrderInvert pcf_get_properties acharset_encoding PCF_Err_Table_Missing pcf_toc_header PCF_Err_Missing_Property ink_minbounds PCF_Err_Invalid_Glyph_Format PCF_Face_Init PCF_Err_Array_Too_Large pcf_get_encodings pcf_get_accel pcf_compressed_metric_header PCF_MetricRec_ PCF_Err_Missing_Encoding_Field PCF_CMapRec_ PCF_Err_Corrupted_Font_Glyphs PCF_Err_Invalid_Face_Handle PCF_Err_Invalid_Post_Table_Format PCF_Err_Invalid_Stream_Seek BDF_PROPERTY_TYPE_CARDINAL acharcode rightSideBearing PCF_Err_Invalid_PPem prop_name bitmapsFormat PCF_Err_Lower_Module_Version PCF_Err_Missing_Bbx_Field nencoding PCF_Err_Corrupted_Font_Header have_change aproperty BDF_PropertyType PCF_Compressed_MetricRec_ BDF_PropertyRec pcf_interpret_style PCF_Err_Hmtx_Table_Missing BDF_PropertyType_ pcf_get_metric characterWidth BDF_PROPERTY_TYPE_NONE PCF_Err_Invalid_Offset leftSideBearing pcf_cmap_char_next cardinal orig_nmetrics PCF_Glyph_Load FT_BDF_GetCharsetIdFunc PCF_Err_Invalid_Horiz_Metrics resolution_x PCF_Err_Cannot_Render_Glyph attributes pcf_has_table_type pcf_services PCF_Accel lastCol PCF_Err_Invalid_Handle BDF_PROPERTY_TYPE_INTEGER PCF_Err_Max comp_source pcf_get_bitmaps PCF_Err_Invalid_Composite FT_Stream_OpenGzip maxOverlap lastRow PCF_Err_Nested_DEFS PCF_Err_Invalid_Opcode PCF_EncodingRec_ FT_Service_BDFRec_ PCF_Err_Too_Many_Extensions pcf_metric_msb_header PCF_Err_Raster_Uninitialized pcf_accel_msb_header PCF_Err_Invalid_Argument PCF_Table encodingOffset PCF_Err_Invalid_CharMap_Handle PCF_PropertyRec_ PCF_AccelRec PCF_Err_Missing_Startchar_Field pcf_get_charset_id PCF_Err_Unknown_File_Format PCF_Err_Too_Many_Hints PCF_Err_Missing_Bitmap firstRow PCF_Err_Could_Not_Find_Context pcf_get_bdf_property PCF_Metric comp_stream PCF_Err_Invalid_Stream_Handle PCF_Err_Missing_Module constantMetrics pcf_cmap_class noOverlap PCF_Err_Invalid_File_Format PCF_MetricRec PCF_Err_Too_Many_Drivers FT_Service_BDFRec PCF_Err_Invalid_Post_Table PCF_Err_Invalid_Cache_Handle pcf_property_set pcf_property_get orig_nbitmaps compr BDF_Err_Missing_Fontboundingbox_Field _bdf_readstream bdf_property_t bdf_driver_requester _bdf_list_shift BDF_Err_Table_Missing BDF_Err_Too_Many_Instruction_Defs bdf_options_t_ BDF_CMap _bdf_atol BDF_Err_Missing_Encoding_Field _bdf_atos bdf_free_font BDF_Err_Raster_Uninitialized buf_size bdf_load_font BDF_Err_Invalid_Driver_Handle BDF_Err_Raster_Overflow keep_comments client_data BDF_Err_Raster_Negative_Height BDF_Err_Corrupted_Font_Header bdf_bbx_t_ _bdf_parse_glyphs BDF_Err_Bad_Argument glyphs_size maxas BDF_Err_Horiz_Header_Missing BDF_Err_No_Unicode_Glyph_Name BDF_Err_Invalid_Face_Handle BDF_Err_Invalid_Post_Table bdf_get_property BDF_Err_Invalid_Stream_Operation vlen BDF_Err_Locations_Missing props_used BDF_Err_Invalid_Outline BDF_Err_Invalid_Table BDF_Err_Too_Many_Drivers nibble_mask _bdf_list_split bdf_cmap_init BDF_Err_Invalid_Stream_Skip separators nuser_props extmemory x_offset BDF_Err_Invalid_Stream_Read bdf_glyph_t_ BDF_Err_Invalid_CharMap_Format _bdf_set_default_spacing BDF_Glyph_Load BDF_Err_Nested_DEFS BDF_encoding_el _bdf_add_comment _num_bdf_properties call_data alen BDF_Err_Array_Too_Large BDF_Err_Invalid_Handle maxds nbuf BDF_Err_Invalid_Version BDF_Err_Invalid_Post_Table_Format BDF_Err_Invalid_CodeRange correct_metrics BDF_Err_Divide_By_Zero BDF_Size_Request bdf_cmap_char_next _bdf_opts oldsize _bdf_atous bigsize BDF_Err_Ok BDF_Err_Nested_Frame_Access nmod _bdf_list_t_ bdf_glyphlist_t_ BDF_Err_Corrupted_Font_Glyphs bdf_cmap_class default_glyph bdf_service_bdf _bdf_parse_start Missing_Encoding monowidth BDF_Err_Max BDF_Err_Could_Not_Find_Context BDF_Err_Missing_Chars_Field BDF_Err_Unlisted_Object bdf_font_t keep_unencoded BDF_Err_Invalid_PPem BDF_Err_Bbx_Too_Big BDF_Err_Glyph_Too_Big BDF_Err_Too_Many_Extensions BDF_FaceRec_ BDF_Err_Cannot_Open_Resource ddigits bdf_property_t_ nibbles comments_len _bdf_is_atom BDF_Err_Invalid_File_Format propid /home/computerfido/Desktop/freetypetest2/freetype/src/bdf/bdf.c BDF_Err_Unknown_File_Format font_ascent BDF_Err_Invalid_Frame_Read bdf_get_charset_id BDF_Err_Invalid_Vert_Metrics bdf_glyph_t BDF_Err_Invalid_Cache_Handle BDF_Err_Invalid_Composite BDF_Err_Invalid_Argument BDF_Err_Invalid_Size_Handle BDF_Err_CMap_Table_Missing props_size proptbl minlb font_descent _bdf_list_ensure _bdf_list_done BDF_Err_Hmtx_Table_Missing linelen BDF_Size_Select BDF_CMapRec_ BDF_Err_Too_Many_Function_Defs BDF_Err_Missing_Bbx_Field BDF_Err_Missing_Size_Field lineno _bdf_add_property BDF_Face_Init seps BDF_Err_Code_Overflow _bdf_list_t BDF_Err_Invalid_Offset bdf_interpret_style BDF_Err_Invalid_Character_Code BDF_Err_Invalid_Stream_Handle BDF_Err_Name_Table_Missing hdigits BDF_Err_Cannot_Open_Stream BDF_Err_DEF_In_Glyf_Bytecode BDF_Err_Stack_Overflow BDF_Err_Invalid_Pixel_Size BDF_Face_Done BDF_Err_Invalid_CharMap_Handle by_encoding BDF_Err_Stack_Underflow BDF_Err_Too_Many_Hints BDF_Face _bdf_parse_properties BDF_Err_Invalid_Frame_Operation maxrb BDF_Err_Missing_Font_Field _bdf_atoul BDF_Err_Invalid_Library_Handle final_empty BDF_Err_Invalid_Opcode BDF_Err_Invalid_Glyph_Index _bdf_parse_t BDF_Err_Invalid_Slot_Handle have BDF_Err_Missing_Module BDF_Err_ENDF_In_Exec_Stream BDF_Err_Too_Few_Arguments BDF_Err_Too_Many_Caches bdf_services BDF_Err_Out_Of_Memory BDF_Err_Raster_Corrupted BDF_Err_Missing_Bitmap bdf_get_bdf_property bdf_options_t swidth BDF_Err_Unimplemented_Feature BDF_Err_Invalid_Glyph_Format bdf_bbx_t BDF_Err_Missing_Property bdfface BDF_Err_Post_Table_Missing builtin bdf_create_property FT_HashRec BDF_Err_Invalid_Horiz_Metrics unencoded_used _bdf_list_join BDF_Err_Debug_OpCode BDF_Err_Invalid_Stream_Seek en_table bdf_glyphlist_t BDF_Err_Execution_Too_Long bdf_font_t_ BDF_Err_Missing_Startfont_Field mask_index glyph_enc BDF_Err_Syntax_Error umod BDF_Err_Lower_Module_Version glyphs_used dwidth font_spacing bitmap_size unencoded_size bdfcmap BDF_Err_Missing_Startchar_Field to_skip _bdf_line_func_t bdf_cmap_char_index BDF_Err_Ignore maxlb _bdf_parse_t_ BDF_Err_Cannot_Render_Glyph BDF_encoding_el_ bdffont BDF_Err_Invalid_Reference bdf_get_font_property avail bdf_cmap_done newsize rbearing _bdf_list_init /home/computerfido/Desktop/freetypetest2/freetype/src/sfnt/sfnt.c SFNT_Err_Invalid_Library_Handle lastVarSel tt_face_load_kern FT_Bitmap_Done tt_cmap14_char_var_index tt_cmap6_class_rec sfnt_get_name_id sfnt_interface NoBitmap table1 table2 sfnt_header woff_offset tt_cmap4_next min_after_bl SFNT_Err_Invalid_Argument cur_gindex char_type SFNT_Err_Invalid_Slot_Handle TT_SBitDecoderRec_ strike_idx TT_CMap tt_cmap12_validate instance_offset char_lo TT_CMapRec_ SFNT_Err_Invalid_Reference tt_cmap8_validate numVar last_end keys count2 SFNT_Err_Bbx_Too_Big SFNT_Err_Too_Many_Function_Defs SFNT_Err_Unimplemented_Feature num_segs metaLength SFNT_Err_Invalid_Handle tt_face_load_head num_pairs has_head tt_cmap8_char_next tt_cmap0_class_rec max_before_bl SFNT_Err_Invalid_CharMap_Handle old_pair TT_Name_ConvertFunc post_len tt_get_cmap_info tt_cmap14_class_rec tt_cmap10_get_info tt_face_free_name wval SFNT_Err_Invalid_Post_Table load_post_names maxProfile tt_cmap2_get_info tt_cmap14_get_nondef_chars cur_group sfnt_find_encoding p_delta bitmap_allocated num_components variantCode SFNT_Err_Nested_DEFS tt_face_load_sbit TT_CMap_ClassRec_ tt_face_load_strike_metrics tt_cmap14_char_index SFNT_Err_Missing_Startchar_Field SFNT_Err_Invalid_Stream_Read tt_get_glyph_name entrySelector TT_CMap_ClassRec SFNT_Err_Glyph_Too_Big originOffsetX originOffsetY subfamily_name tt_face_load_hmtx SFNT_Err_Invalid_Outline SFNT_Err_Ok TT_CMap4 SFNT_Err_Stack_Overflow found_unicode tt_cmap14_init SFNT_Err_Post_Table_Missing SFNT_Err_Code_Overflow woff_header_fields TT_CMap12 max_gid recurse_depth tt_face_get_kerning ignore_typographic_family post_limit SFNT_Err_Missing_Chars_Field sfnt_get_var_ps_name privOffset TT_CMapRec SFNT_Err_Corrupted_Font_Header image_format sfnt_service_sfnt_table TT_CMap13 TT_CMap14 TT_CMap4Rec_ sfnt_is_postscript PSname tt_cmap10_char_next tt_cmap12_init sfnt_is_alphanumeric pwrite report_invalid_characters tt_cmap12_next glyph_id graphicType charCode tt_face_load_font_dir num_groups tt_name_ascii_from_utf16 sfnt_stream_close get_sfnt_table tt_cmap14_def_char_count SFNT_Err_Stack_Underflow rangeShift totalSfntSize storage_start SFNT_Err_Corrupted_Font_Glyphs FT_Bitmap_Init sfnt_table_info TEncoding_ SFNT_Err_Missing_Module psnames_error sfnt_init_face NoData TT_CMap13Rec_ SFNT_Err_Invalid_Table tt_face_load_gasp tt_cmap_unicode_char_next load_format_25 TT_SBitDecoder_LoadFunc found_win SFNT_Err_Invalid_Frame_Operation tt_sbit_decoder_done duplicate tt_cmap14_validate tt_sbit_decoder_load_bitmap SFNT_Err_Cannot_Open_Resource prev_end sfnt_services get_win_string varSel default_values TT_SBitDecoderRec tt_cmap14_variants WOFF_HeaderRec_ image_size FoundStrike aprop NextTable tt_cmap14_char_map_nondef_binary SFNT_Err_Invalid_Stream_Seek eblc_base tt_face_free_ps_names tt_cmap2_class_rec check_table_dir tt_sbit_decoder_init SFNT_Err_CMap_Table_Missing SFNT_Err_Invalid_Offset tt_face_get_metrics new_map tt_cmap4_validate Next_Segment byte_size instance_values starts SFNT_Err_Invalid_Stream_Skip default_value_offset glyph_ids property_len fixed2float tt_cmap0_validate last_start FT_Gzip_Uncompress tt_cmap0_get_info tt_cmap13_char_index tt_cmap4_char_map_binary SFNT_Err_Invalid_Driver_Handle offset1 offset2 cur_end SFNT_Err_Raster_Negative_Height range_index found_apple_roman sfnt_ps_map tt_cmap13_char_map_binary valid_entries SFNT_Err_Raster_Corrupted tt_cmap13_validate metaOffset tt_face_load_sbix_image WOFF_HeaderRec TEncoding sfnt_offset SFNT_Err_Invalid_Character_Code nblocks bit_depth tt_cmap14_char_next post_fields SFNT_Err_Nested_Frame_Access tt_cmap4_class_rec image_offset ptable_offset SFNT_Err_ENDF_In_Exec_Stream tt_face_load_hhea SFNT_Err_Missing_Encoding_Field privLength has_unicode tt_face_get_ps_name tt_cmap2_char_index tt_cmap14_variant_chars tt_face_load_cmap cur_start tt_face_goto_table p_next SFNT_Err_Horiz_Header_Missing nuni cur_charcode tt_cmap13_class_rec SFNT_Err_Missing_Fontboundingbox_Field SFNT_Err_Cannot_Render_Glyph ptable_size SFNT_Err_Table_Missing avgwidth first_code tt_cmap10_char_index tt_cmap12_get_info tt_face_load_maxp sfnt_open_font tt_cmap14_char_map_def_binary cmap4 ttcmap numMappings maxp_fields metrics_loaded SFNT_HeaderRec convert validator tt_sbit_decoder_alloc_bitmap tt_cmap2_char_next tt_module tt_cmap_unicode_char_index TT_Validator instance_size ignore_typographic_subfamily TT_NameTable woff tt_cmap12_class_rec is_apple_sbit char_type_func is_apple_sbix tt_cmap6_char_next tt_cmap12_char_next TT_TableRec SFNT_Err_Ignore SFNT_Err_Array_Too_Large tt_encodings ppem_ tt_face_load_any tt_cmap6_char_index tt_face_load_bhed SFNT_Err_Locations_Missing tt_cmap0_char_next tt_cmap4_get_info tt_cmap_unicode_init load_format_20 tt_sbit_decoder_load_compound tt_cmap14_get_def_chars found_apple_english sfnt_get_ps_name FoundRange tt_cmap_unicode_done BadTable TT_CMap_ValidateFunc SFNT_Err_Invalid_Glyph_Index SFNT_Err_Invalid_Stream_Operation tt_cmap4_set_range woff_open_font tt_cmap12_char_index tt_name_ascii_from_other SFNT_Header ordered bit_height get_apple_string SFNT_Err_Bad_Argument SFNT_Err_Invalid_Glyph_Format tt_cmap4_char_next is_english SFNT_Err_Invalid_Opcode start_id SFNT_Err_Invalid_CodeRange sfnt_get_interface name_table_fields pclazz bsize_idx SFNT_Err_Execution_Too_Long Next_SubHeader sfnt_load_face key0 tt_sbit_decoder_load_metrics duni offset_table_fields SFNT_Err_Invalid_Cache_Handle upem sfnt_service_bdf old_tag tt_cmap4_char_map_linear retry SFNT_Err_Divide_By_Zero tt_cmap8_char_index strike_index_array pcharcode has_outline murmur_hash_3_128 entry_selector searchRange SFNT_Err_Too_Few_Arguments tt_cmap13_get_info SFNT_Err_Too_Many_Instruction_Defs nbits tt_cmap12_char_map_binary tt_face_load_bdf_props flavor minorVersion sfnt_get_glyph_name pclt_fields SFNT_Err_Invalid_Face_Handle maxp_fields_extra tt_cmap14_ensure tt_cmap4_init WOFF_TableRec_ nondefOff SFNT_Err_Raster_Uninitialized tt_cmap10_class_rec SFNT_Err_Debug_OpCode tt_cmap6_validate tt_sbit_decoder_load_image table_pos SFNT_Err_Invalid_Size_Handle rval SFNT_Err_Missing_Size_Field hexdigits tt_cmap14_char_variants SFNT_Err_Out_Of_Memory bit_width lastUni ttc_header_fields tt_sbit_decoder_load_bit_aligned tt_cmap0_char_index tt_face_build_cmaps search_range found_apple frac_part tt_face_load_generic_header SFNT_Err_DEF_In_Glyf_Bytecode tt_cmap8_get_info bit_size FT_Bitmap_Convert SFNT_Err_Invalid_Pixel_Size range_shift SFNT_Err_Missing_Font_Field strike_offset SFNT_Err_Syntax_Error tt_cmap14_char_var_isdefault num_segs2 SFNT_Err_Max storage_limit next_end tt_cmap8_class_rec tt_cmap_unicode_class_rec SFNT_Err_Invalid_Stream_Handle lastBase abearing langTag_record_fields SFNT_Err_Invalid_File_Format SFNT_Err_Unknown_File_Format check_length TT_Post_Names WOFF_Table SFNT_Err_Name_Table_Missing image_start tt_face_load_name os2_fields_extra5 line_bits os2_fields image_end SFNT_HeaderRec_ gaspranges TT_SBit_Metrics name_record_fields compare_offsets name_strings SFNT_Err_Raster_Overflow SFNT_Err_Could_Not_Find_Context SFNT_Err_Too_Many_Caches SFNT_Err_Invalid_PPem has_meta tt_face_lookup_table SFNT_Err_Invalid_Composite cur_values code_count sfnt_get_name_index astrike_index SFNT_Err_Too_Many_Drivers tt_cmap14_get_info next_start tt_face_done_kern tt_cmap6_get_info metaOrigLength metrics_header_fields TT_ValidatorRec tt_face_free_sbit SFNT_Err_Hmtx_Table_Missing tt_sbit_decoder_load_byte_aligned cur_pair SFNT_Err_Missing_Property max_results os2_fields_extra1 os2_fields_extra2 SFNT_Err_No_Unicode_Glyph_Name tt_cmap_classes tt_face_set_sbit_strike tt_service_get_cmap_info table_dir_entry_fields SFNT_Err_Missing_Startfont_Field SFNT_Err_Unlisted_Object output_len sfnt_service_ps_name array_start is32 SFNT_Err_Cannot_Open_Stream tt_face_get_name CompLength TT_Post_20 TT_Post_25 TT_CMap14Rec_ cmap12 cmap13 cmap14 dcnt tt_cmap14_find_variant FT_Service_SFNT_TableRec tt_cmap2_validate SFNT_Err_Too_Many_Extensions TT_ValidatorRec_ strike_index_count tt_face_find_bdf_prop sfnt_get_charset_id SFNT_Err_Invalid_Version sfnt_service_glyph_dict setjmp offset_table index_format SFNT_Err_Invalid_Frame_Read tt_cmap2_get_subheader SFNT_Err_Lower_Module_Version sfnt_done_face tt_face_load_pclt nameid SFNT_Err_Missing_Bbx_Field construct_instance_name OrigOffset fvar_len TT_CMap12Rec_ int_part SFNT_Err_Invalid_Post_Table_Format tt_cmap14_done old_p fmix32 tt_face_free_bdf_props defp tt_face_load_os2 tt_face_load_sbit_image num_selectors eblc_limit p_start FT_ValidatorRec tt_cmap_init tt_cmap13_char_next tt_cmap10_validate SFNT_Err_Invalid_Horiz_Metrics SFNT_Err_Too_Many_Hints char_hi tt_cmap13_next tt_face_load_post SFNT_Err_Missing_Bitmap TT_CMap_Class tt_cmap13_init has_sing tt_cmap4_char_index TT_BDF num_cmaps num_results TT_SBitDecoder SFNT_Err_Invalid_CharMap_Format SFNT_Err_Invalid_Vert_Metrics af_warper_compute af_latn_titl_style_class AF_BLUE_STRING_LATIN_SUBS_SMALL_DESCENDER af_telu_dflt_style_class AF_COVERAGE_ORDINALS style_metrics_size AF_BLUE_STRING_MYANMAR_TOP shaper_buf AF_CJKMetrics af_iup_shift AF_BLUE_STRING_TAI_VIET_BOTTOM AF_BLUE_STRING_MAX AF_AxisHintsRec_ AF_ScriptClass axhints af_lao_script_class height_threshold af_latn_c2cp_style_class AF_BLUE_STRINGSET_TFNG p_last AF_Err_Raster_Corrupted af_none_script_class AF_STYLE_LATB_DFLT af_grek_sups_style_class pp1x_uh af_face_globals_new AF_BLUE_STRING_GEORGIAN_MKHEDRULI_ASCENDER AF_Err_Raster_Uninitialized has_last_stem af_cjk_writing_system_class AF_BLUE_STRING_ETHIOPIC_TOP is_top_right_blue AF_Err_Ok af_osge_dflt_style_class AF_BLUE_STRING_TAMIL_BOTTOM AF_SCRIPT_KALI AF_STYLE_LATN_C2CP af_kali_uniranges AF_Err_Corrupted_Font_Glyphs AF_BLUE_STRING_LAO_BOTTOM AF_WritingSystemClassRec_ af_limb_script_class af_gujr_dflt_style_class AF_SCRIPT_SAUR AF_Err_Invalid_Reference af_dsrt_uniranges af_cari_uniranges AF_STYLE_VAII_DFLT AF_Err_Missing_Fontboundingbox_Field af_thai_uniranges AF_BLUE_STRING_GLAGOLITIC_SMALL_BOTTOM af_nkoo_script_class AF_BLUE_STRING_MYANMAR_DESCENDER prev_min_pos AF_Err_Unknown_File_Format AF_Err_Raster_Negative_Height af_axis_hints_new_segment AF_BLUE_STRING_GURMUKHI_BASE AF_BLUE_STRING_ARABIC_TOP af_cjk_hints_detect_features AF_BLUE_STRING_LAO_TOP AF_BLUE_STRING_SINHALA_BOTTOM af_nkoo_dflt_style_class AF_STYLE_SUND_DFLT AF_COVERAGE_PETITE_CAPITALS_FROM_CAPITALS AF_BLUE_STRING_ADLAM_SMALL_BOTTOM AF_BLUE_STRING_GUJARATI_BOTTOM AF_WRITING_SYSTEM_LATIN Is_Weak_Point points_limit prev_min_coord AF_AxisHints af_goth_script_class af_gujr_uniranges last_touched af_guru_nonbase_uniranges AF_BLUE_STRING_KHMER_SYMBOLS_WANING_BOTTOM AF_BLUE_STRINGSET_SUND AF_BLUE_STRING_LATIN_SUBS_CAPITAL_BOTTOM af_cjk_hints_link_segments af_avst_dflt_style_class org_len AF_Warper af_sund_dflt_style_class af_cjk_hints_init af_bamu_uniranges af_cjk_metrics_scale_dim seg_delta AF_BLUE_STRING_OLD_TURKIC_TOP AF_BLUE_STRINGSET_NONE AF_COVERAGE_SMALL_CAPITALS_FROM_CAPITALS AF_Err_Invalid_Character_Code AF_Err_Invalid_Size_Handle af_ethi_uniranges AF_BLUE_STRINGSET_THAI AF_STYLE_ETHI_DFLT AF_BLUE_STRINGSET_ARMN AF_COVERAGE_PETITE_CAPITALS AF_STYLE_ORKH_DFLT AF_SCRIPT_OSMA AF_BLUE_STRINGSET_OLCK AF_Err_Raster_Overflow style_metrics_scale style_metrics dist_score FT_Prop_GlyphToScriptMap AF_BLUE_STRING_SHAVIAN_SMALL_TOP af_loader_init af_latn_sups_style_class inverse af_avst_nonbase_uniranges af_geok_uniranges af_deva_dflt_style_class segment_dir af_beng_nonbase_uniranges script_uni_nonbase_ranges af_cyrl_pcap_style_class af_blue_stringsets AF_Err_Bbx_Too_Big af_cans_dflt_style_class AF_SCRIPT_BENG AF_StyleMetricsRec af_osge_nonbase_uniranges AF_STYLE_CYRL_SUBS AF_BLUE_STRINGSET_BUHD af_glyph_hints_done AF_CJKAxisRec_ AF_SCRIPT_ETHI af_tfng_dflt_style_class AF_BLUE_STRING_GEORGIAN_NUSKHURI_DESCENDER af_shaw_uniranges best_distort AF_STYLE_LATN_SUBS AF_Dimension_ af_orkh_nonbase_uniranges AF_BLUE_STRING_DEVANAGARI_HEAD AF_Err_Invalid_Post_Table_Format xx1max AF_BLUE_STRINGSET_ETHI AF_WRITING_SYSTEM_INDIC AF_Err_Invalid_Driver_Handle AF_Err_Invalid_CodeRange AF_Err_Invalid_Composite af_mymr_uniranges af_latn_script_class af_grek_c2sc_style_class AF_Module fpos is_round AF_BLUE_STRING_DEVANAGARI_BASE AF_BLUE_STRING_KAYAH_LI_TOP AF_SCRIPT_GURU AF_COVERAGE_SCIENTIFIC_INFERIORS AF_STYLE_CHER_DFLT AF_Err_Nested_Frame_Access AF_BLUE_STRING_LATIN_SUPS_CAPITAL_BOTTOM AF_STYLE_CYRL_SINF prev_max_coord af_warper_compute_line_best d_off1 darken_by_font_units_x AF_LatinAxisRec AF_BLUE_STRING_COPTIC_SMALL_TOP AF_STYLE_LATN_SINF old_rsb best_round af_saur_nonbase_uniranges af_cyrl_script_class AF_StyleClassRec AF_Err_Invalid_Table AF_BLUE_STRING_GEORGIAN_MKHEDRULI_TOP AF_WRITING_SYSTEM_DUMMY AF_SCRIPT_KNDA scale_down_matrix AF_SCRIPT_CAKM AF_BLUE_STRING_OSAGE_CAPITAL_DESCENDER num_segments af_avst_uniranges style_metrics_done edge_distance_threshold warper af_cari_nonbase_uniranges af_orkh_script_class best_score trans_delta AF_WritingSystem_ x2max idx_max AF_CJKMetricsRec AF_BLUE_STRING_CYPRIOT_TOP af_cjk_hints_compute_segments AF_ModuleRec_ AF_BLUE_STRING_TAI_VIET_TOP af_limb_nonbase_uniranges AF_ScriptClassRec_ af_orkh_dflt_style_class AF_BLUE_STRING_NKO_SMALL_TOP af_hint_normal_stem AF_Err_Too_Many_Extensions AF_LatinMetricsRec_ AF_Err_Missing_Startchar_Field AF_STYLE_NKOO_DFLT AF_DIR_DOWN prev_min_on_coord AF_BLUE_STRING_GURMUKHI_DIGIT_TOP af_tfng_nonbase_uniranges AF_LatinMetricsRec af_glag_uniranges af_buhd_script_class oldmap af_style_classes af_cans_script_class scaler af_grek_sinf_style_class reference stdHW AF_BLUE_STRING_ARMENIAN_SMALL_ASCENDER af_glyph_hints_rescale af_none_dflt_style_class AF_BLUE_STRINGSET_GLAG max_segments AF_BLUE_STRING_KANNADA_BOTTOM af_knda_uniranges AF_SCRIPT_CANS AF_STYLE_SAUR_DFLT AF_Style AF_COVERAGE_DEFAULT AF_SCRIPT_SYLO af_blue_strings AF_STYLE_GEOK_DFLT AF_Err_Invalid_Frame_Operation af_armn_dflt_style_class AF_BLUE_STRING_MALAYALAM_BOTTOM AF_BLUE_STRINGSET_COPT AF_Err_Invalid_Version AF_Err_Missing_Font_Field AF_BLUE_STRINGSET_GUJR curr af_face_globals_is_digit /home/computerfido/Desktop/freetypetest2/freetype/src/autofit/autofit.c AF_Err_Corrupted_Font_Header best_contour_last next_u af_geor_nonbase_uniranges AF_BLUE_STRING_MALAYALAM_TOP AF_STYLE_MAX AF_BLUE_STRING_CHEROKEE_SMALL_DESCENDER AF_Err_Invalid_Outline AF_LatinBlueRec AF_STYLE_CAKM_DFLT extra_light af_vaii_nonbase_uniranges af_bamu_dflt_style_class AF_Err_Missing_Property AF_Err_Too_Many_Drivers af_dsrt_script_class af_cjk_metrics_init_blues af_indic_get_standard_widths af_property_get FT_Prop_GlyphToScriptMap_ best_x af_latn_subs_style_class af_cher_uniranges af_osge_script_class AF_BLUE_STRINGSET_KALI AF_LoaderRec af_cjk_get_standard_widths AF_LatinAxis AF_BLUE_STRING_LAO_DESCENDER AF_STYLE_GREK_C2CP AF_BLUE_STRING_LATIN_SUPS_SMALL best_on_point_last af_geok_nonbase_uniranges AF_BLUE_STRINGSET_SAUR Try_x3 Try_x4 AF_STYLE_GURU_DFLT is_serif AF_Width AF_Script_UniRange AF_WarpScore AF_LatinBlueRec_ blue_stringset AF_BLUE_STRING_GEORGIAN_ASOMTAVRULI_TOP prev_max_pos AF_BLUE_STRING_GUJARATI_TOP af_deva_nonbase_uniranges AF_BLUE_STRING_SINHALA_TOP FT_Prop_IncreaseXHeight af_autofitter_init AF_SCRIPT_LAO AF_BLUE_STRING_VAI_BOTTOM prev_segment af_lisu_dflt_style_class AF_BLUE_STRING_LATIN_SUBS_SMALL af_lisu_script_class neutral2 AF_SCRIPT_CARI AF_BLUE_STRING_GURMUKHI_HEAD AF_SCRIPT_MLYM af_loader_load_glyph af_cans_nonbase_uniranges near_limit2 AF_AxisHintsRec af_hani_dflt_style_class AF_Err_Invalid_Frame_Read latin af_hani_nonbase_uniranges AF_CJKBlueRec_ AF_Err_Too_Many_Instruction_Defs AF_STYLE_TAML_DFLT AF_BLUE_STRING_GEORGIAN_ASOMTAVRULI_BOTTOM AF_BLUE_STRING_LATIN_SMALL_BOTTOM AF_COVERAGE_SUBSCRIPT org_delta AF_BLUE_STRING_ARMENIAN_SMALL_DESCENDER af_cyrl_sups_style_class af_mymr_dflt_style_class AF_BLUE_STRING_DESERET_SMALL_TOP AF_SCRIPT_VAII AF_STYLE_GUJR_DFLT af_latp_script_class af_shaper_get_elem AF_BLUE_STRING_KAYAH_LI_DESCENDER af_hebr_script_class AF_WritingSystem_DoneMetricsFunc AF_BLUE_STRING_KAYAH_LI_LARGE_DESCENDER AF_BLUE_STRING_GUJARATI_ASCENDER af_sinh_uniranges AF_BLUE_STRING_CARIAN_BOTTOM AF_Err_Divide_By_Zero af_sund_uniranges AF_Err_Stack_Underflow AF_Direction_ AF_LatinAxisRec_ x2min af_latb_nonbase_uniranges idx_min af_grek_dflt_style_class prev_v AF_SCRIPT_LIMB AF_STYLE_TELU_DFLT AF_BLUE_STRING_ETHIOPIC_BOTTOM af_latn_sinf_style_class AF_CJKAxis scaler_flags af_vaii_script_class first_v near_limit blue_sorted af_latn_smcp_style_class AF_STYLE_CYRL_C2CP AF_BLUE_STRING_KHMER_TOP af_latin_snap_width AF_STYLE_SYLO_DFLT af_cjk_hints_compute_edges af_hebr_uniranges af_tibt_nonbase_uniranges AF_STYLE_TIBT_DFLT af_tavt_script_class AF_ScalerRec AF_Err_Invalid_Stream_Read af_buhd_nonbase_uniranges af_face_globals_free AF_BLUE_STRING_SHAVIAN_BOTTOM AF_BLUE_STRING_GREEK_SMALL_DESCENDER AF_Err_Missing_Size_Field af_blue_1_2 AF_BLUE_STRINGSET_BENG AF_BLUE_STRING_SUNDANESE_BOTTOM AF_DIMENSION_VERT script_uni_ranges af_osma_dflt_style_class best_dist0 af_buhd_uniranges af_none_nonbase_uniranges AF_BLUE_STRING_BENGALI_TOP af_latin_hint_edges AF_BLUE_STRINGSET_CAKM AF_SCRIPT_GLAG org_scale AF_STYLE_GREK_SUBS AF_SCRIPT_MYMR warping af_latin_hints_compute_blue_edges af_arab_uniranges af_indic_writing_system_class touch_flag AF_STYLE_CYRL_SUPS stem_flags af_limb_uniranges af_dsrt_dflt_style_class af_sund_script_class AF_Point af_glyph_hints_init AF_BLUE_STRING_KAYAH_LI_ASCENDER AF_SCRIPT_TELU best_blue dist_threshold AF_BLUE_STRING_THAI_TOP AF_STYLE_CYRL_SMCP asegment AF_BLUE_STRING_BUHID_SMALL AF_BLUE_STRING_MYANMAR_ASCENDER AF_BLUE_STRING_GURMUKHI_TOP AF_STYLE_CARI_DFLT AF_BLUE_STRING_BENGALI_HEAD stem_width_per_1000 cur_pos1 cur_pos2 AF_STYLE_LATN_SMCP skipped af_latin_sort_blue increase_x_height edge1 edge2 ft_module AF_SCRIPT_MAX AF_STYLE_MLYM_DFLT edge3 af_armn_uniranges FT_AutoHinter_InterfaceRec AF_STYLE_GREK_SINF AF_Err_Invalid_Face_Handle af_autofitter_load_glyph af_cher_nonbase_uniranges AF_BLUE_STRINGSET_KNDA AF_BLUE_STRING_BENGALI_BASE AF_BLUE_STRING_CYPRIOT_SMALL af_glyph_hints_reload prev_max_on_coord AF_BLUE_STRING_AVESTAN_BOTTOM best_scale stdVW AF_BLUE_STRING_GEORGIAN_NUSKHURI_BOTTOM AF_BLUE_STRING_HEBREW_DESCENDER AF_SCRIPT_AVST AF_Err_Lower_Module_Version AF_STYLE_GREK_SUPS AF_BLUE_STRING_BUHID_TOP AF_BLUE_STRINGSET_LAO wmin AF_Err_CMap_Table_Missing af_cyrl_ordn_style_class af_mlym_script_class Hint_Metrics af_loader_compute_darkening AF_Err_Invalid_Stream_Operation AF_LoaderRec_ af_latin_align_linked_edge AF_BLUE_STRING_LAO_LARGE_ASCENDER af_saur_script_class af_guru_uniranges AF_SCRIPT_TAML af_dummy_writing_system_class af_saur_uniranges AF_SCRIPT_SHAW af_khms_uniranges af_cans_uniranges AF_BLUE_STRING_KHMER_DESCENDER old_advance AF_STYLE_GREK_PCAP AF_Err_Name_Table_Missing AF_STYLE_OSMA_DFLT AF_BLUE_STRING_MYANMAR_BOTTOM best_delta style_metrics_init af_tfng_script_class af_vaii_dflt_style_class af_indic_hints_apply af_lao_nonbase_uniranges AF_STYLE_GREK_SMCP AF_STYLE_GREK_ORDN af_property_set AF_STYLE_COPT_DFLT af_taml_uniranges AF_BLUE_STRING_TELUGU_TOP AF_BLUE_STRINGSET_BAMU em_ratio af_cjk_metrics_check_digits AF_FaceGlobalsRec_ AF_SCRIPT_LISU af_goth_uniranges af_cher_script_class best_on_point_first AF_BLUE_STRING_GEORGIAN_NUSKHURI_ASCENDER AF_Err_Too_Many_Hints AF_BLUE_STRING_COPTIC_CAPITAL_TOP af_lisu_nonbase_uniranges size_internal af_grek_ordn_style_class AF_BLUE_STRING_KAYAH_LI_BOTTOM Use_y4 af_cjk_align_serif_edge AF_Err_Invalid_Vert_Metrics AF_BLUE_STRING_CYRILLIC_CAPITAL_BOTTOM af_blue_2_1 af_blue_2_2 AF_BLUE_STRINGSET_CANS af_ethi_script_class AF_BLUE_STRING_SHAVIAN_TOP AF_ScalerRec_ FT_Prop_IncreaseXHeight_ AF_Err_Invalid_Argument af_nkoo_nonbase_uniranges AF_WarperRec_ af_latb_script_class xx1min af_shaper_buf_destroy AF_COVERAGE_TITLING af_thai_dflt_style_class af_osma_nonbase_uniranges AF_BLUE_STRING_OSAGE_SMALL_ASCENDER AF_STYLE_ORYA_DFLT AF_BLUE_STRING_ARMENIAN_CAPITAL_BOTTOM best_segment_last dist2 af_sinh_nonbase_uniranges d_off af_beng_script_class AF_BLUE_STRING_CANADIAN_SYLLABICS_SUPS_TOP contour_limit style_hints_init AF_STYLE_LATN_SUPS new_scale AF_SegmentRec AF_BLUE_STRINGSET_GURU AF_StyleClassRec_ af_cyrl_smcp_style_class af_olck_uniranges af_cakm_dflt_style_class is_under_ref AF_Err_Nested_DEFS AF_STYLE_CPRT_DFLT AF_BLUE_STRING_CHEROKEE_SMALL_ASCENDER af_thai_script_class AF_WritingSystem_ApplyHintsFunc af_grek_subs_style_class AF_CJKMetricsRec_ AF_Err_Invalid_CharMap_Handle af_axis_hints_new_edge AF_BLUE_STRING_LATIN_SMALL_F_TOP AF_BLUE_STRING_OLD_TURKIC_BOTTOM af_tavt_uniranges AF_BLUE_STRING_CANADIAN_SYLLABICS_SMALL_TOP AF_Err_Hmtx_Table_Missing anedge num_rounds af_cjk_hint_edges AF_BLUE_STRINGSET_DEVA af_deva_uniranges segment_limit base_delta ydelta af_khms_nonbase_uniranges AF_BLUE_STRING_ARMENIAN_SMALL_TOP AF_BLUE_STRING_OL_CHIKI AF_STYLE_SHAW_DFLT af_latin_writing_system_class AF_Blue_String_ AF_Blue_StringRec_ af_goth_nonbase_uniranges af_telu_script_class AF_STYLE_MYMR_DFLT opos af_get_interface AF_BLUE_STRINGSET_CPRT is_straight link af_latn_c2sc_style_class AF_BLUE_STRING_SUNDANESE_DESCENDER AF_BLUE_STRINGSET_MAX af_cyrl_nonbase_uniranges other_flags xdelta has_serifs old_best_point AF_BLUE_STRINGSET_CARI AF_Err_Invalid_File_Format AF_BLUE_STRINGSET_MLYM af_cyrl_sinf_style_class AF_STYLE_AVST_DFLT af_geok_dflt_style_class AF_COVERAGE_SUPERSCRIPT af_cher_dflt_style_class stem_darkening_for_ppem af_shaper_buf_create AF_BLUE_STRING_CHAKMA_TOP AF_SCRIPT_NKOO AF_CJKBlue AF_STYLE_OSGE_DFLT AF_Coverage AF_Err_Invalid_CharMap_Format AF_SCRIPT_DSRT AF_SCRIPT_ADLM a_delta control_overshoot AF_BLUE_STRINGSET_VAII af_arab_dflt_style_class big_max af_telu_uniranges AF_Err_Ignore AF_BLUE_STRING_ARMENIAN_SMALL_BOTTOM af_limb_dflt_style_class AF_STYLE_HANI_DFLT AF_STYLE_GREK_C2SC AF_STYLE_ADLM_DFLT af_glag_dflt_style_class af_latin_hints_detect_features af_lao_uniranges AF_DIR_UP af_khmr_uniranges AF_GlyphHintsRec AF_BLUE_STRING_HEBREW_BOTTOM af_glyph_hints_align_edge_points scaled_stem AF_BLUE_STRING_BAMUM_TOP EndContour num_flats AF_BLUE_STRING_NKO_BOTTOM af_latin_hints_init AF_Err_Unimplemented_Feature u_off1 u_off2 AF_Err_Too_Many_Function_Defs AF_STYLE_LAO_DFLT AF_Err_Locations_Missing AF_Err_Code_Overflow af_latin_hints_compute_segments scores AF_BLUE_STRING_COPTIC_CAPITAL_BOTTOM AF_STYLE_DEVA_DFLT passed AF_BLUE_STRING_KANNADA_TOP style_options AF_BLUE_STRING_KHMER_BOTTOM AF_BLUE_STRING_LATIN_SMALL_TOP AF_BLUE_STRING_THAI_LARGE_ASCENDER edge_next AF_WritingSystem_InitMetricsFunc new_lsb left2right AF_BLUE_STRING_CHAKMA_BOTTOM AF_SCRIPT_TAVT AF_SCRIPT_GEOK buf_ AF_BLUE_STRING_LATIN_CAPITAL_TOP AF_SCRIPT_GEOR AF_Err_Invalid_Offset AF_BLUE_STRING_CHAKMA_DESCENDER len_score out_dir best_contour_first af_taml_script_class AF_DIMENSION_HORZ af_mlym_nonbase_uniranges gstyles AF_STYLE_GOTH_DFLT AF_BLUE_STRINGSET_MYMR af_sort_pos idx0 u_off AF_BLUE_STRING_GUJARATI_DIGIT_TOP af_cprt_nonbase_uniranges af_geok_script_class embedded af_nkoo_uniranges AF_Err_Syntax_Error last_v AF_SCRIPT_BUHD AF_BLUE_STRING_OSAGE_SMALL_DESCENDER af_loader_done af_beng_dflt_style_class af_ethi_nonbase_uniranges AF_BLUE_STRING_ADLAM_SMALL_TOP standard_vertical_width AF_BLUE_STRING_LATIN_CAPITAL_BOTTOM af_latn_nonbase_uniranges af_sund_nonbase_uniranges af_buhd_dflt_style_class blue_ref af_grek_script_class AF_STYLE_LATP_DFLT AF_BLUE_STRING_KHMER_LARGE_DESCENDER AF_BLUE_STRING_LISU_BOTTOM af_lisu_uniranges AF_BLUE_STRINGSET_AVST AF_STYLE_GLAG_DFLT af_grek_pcap_style_class af_loader_embolden_glyph_in_slot AF_BLUE_STRING_OSAGE_CAPITAL_TOP AF_WritingSystem_ScaleMetricsFunc af_adlm_nonbase_uniranges af_cjk_metrics_init af_bamu_script_class AF_BLUE_STRING_OSAGE_SMALL_BOTTOM AF_FaceGlobals AF_STYLE_BAMU_DFLT AF_Err_Out_Of_Memory AF_SCRIPT_GOTH AF_SCRIPT_ORKH af_telu_nonbase_uniranges AF_STYLE_CYRL_DFLT margin af_dummy_hints_apply af_glyph_hints_align_weak_points prev_min_flags AF_Err_Array_Too_Large AF_SCRIPT_CYRL AF_BLUE_STRING_OSMANYA_TOP AF_Err_Invalid_Slot_Handle AF_SCRIPT_COPT fitted_width AF_BLUE_STRING_HEBREW_TOP af_loader_reset AF_STYLE_LATN_DFLT af_armn_nonbase_uniranges AF_Err_Horiz_Header_Missing AF_EdgeRec AF_SCRIPT_TFNG af_copt_uniranges af_taml_dflt_style_class AF_BLUE_STRINGSET_TAML AF_BLUE_STRING_SAURASHTRA_TOP af_indic_metrics_scale AF_BLUE_STRINGSET_SHAW AF_BLUE_STRING_CYPRIOT_BOTTOM af_lao_dflt_style_class AF_GlyphHintsRec_ AF_Segment AF_Err_Invalid_Glyph_Index AF_CJKAxisRec AF_Err_Invalid_PPem af_knda_script_class af_autofitter_done af_latp_dflt_style_class AF_Err_Unlisted_Object cur_idx AF_SCRIPT_HANI af_hebr_dflt_style_class af_orkh_uniranges best_pos AF_SCRIPT_OSGE af_ethi_dflt_style_class AF_BLUE_STRINGSET_LISU af_kali_script_class AF_Err_Invalid_Stream_Skip org_pos AF_BLUE_STRING_GUJARATI_DESCENDER af_latin_metrics_init_blues AF_STYLE_KHMS_DFLT af_geor_dflt_style_class af_saur_dflt_style_class af_mymr_script_class AF_Style_ AF_BLUE_STRING_LATIN_SUPS_SMALL_F_TOP af_tibt_dflt_style_class seg0 top_to_bottom_hinting seg2 AF_SCRIPT_GREK AF_BLUE_STRING_LISU_TOP af_sylo_script_class af_hebr_nonbase_uniranges AF_PointRec_ af_sylo_dflt_style_class af_latin_get_standard_widths AF_Err_Too_Few_Arguments AF_STYLE_KHMR_DFLT AF_SCRIPT_LATB best_blue_is_neutral af_cakm_nonbase_uniranges new_delta AF_SCRIPT_LATN AF_SCRIPT_LATP AF_COVERAGE_SMALL_CAPITALS AF_BLUE_STRING_GEORGIAN_MKHEDRULI_DESCENDER darken_amount AF_BLUE_STRING_NKO_TOP AF_Err_Missing_Startfont_Field AF_STYLE_KALI_DFLT af_blue_1_1_1 af_blue_1_1_2 len_threshold af_property_get_face_globals AF_EdgeRec_ AF_BLUE_STRING_OSAGE_SMALL_TOP AF_BLUE_STRING_AVESTAN_TOP AF_SCRIPT_DEVA AF_STYLE_CANS_DFLT af_grek_titl_style_class af_cyrl_c2sc_style_class af_khms_script_class AF_Blue_Stringset_ glyph_styles af_cjk_align_edge_points af_cprt_script_class best_y_extremum AF_SCRIPT_ARAB af_grek_c2cp_style_class blue_count AF_BLUE_STRING_OSAGE_CAPITAL_BOTTOM AF_Err_Execution_Too_Long af_latin_metrics_init_widths af_knda_nonbase_uniranges AF_BLUE_STRING_TAMIL_TOP AF_Err_Invalid_Library_Handle af_latin_metrics_scale_dim AF_STYLE_TFNG_DFLT trans_matrix AF_BLUE_STRING_KHMER_SYMBOLS_WAXING_TOP endpoint num_edges AF_Blue_StringRec AF_Coverage_ af_orya_script_class af_latp_nonbase_uniranges AF_BLUE_STRING_ARABIC_BOTTOM AF_DIMENSION_MAX AF_CJKBlueRec size_changed AF_STYLE_KNDA_DFLT AF_BLUE_STRING_THAI_BOTTOM af_warper_weights AF_BLUE_STRING_SINHALA_DESCENDER AF_Err_Invalid_Handle AF_WritingSystem_GetStdWidthsFunc af_sylo_uniranges af_autofitter_interface AF_SCRIPT_SINH AF_BLUE_STRING_LAO_ASCENDER max_edges af_latin_hints_compute_edges af_cjk_align_linked_edge scale_down_factor AF_BLUE_STRINGSET_TAVT AF_BLUE_STRING_GOTHIC_TOP AF_BLUE_STRING_LATIN_SUPS_CAPITAL_TOP af_script_classes AF_Script_UniRangeRec AF_SCRIPT_BAMU AF_BLUE_STRING_CANADIAN_SYLLABICS_BOTTOM AF_BLUE_STRINGSET_NKOO AF_STYLE_LIMB_DFLT AF_BLUE_STRINGSET_DSRT AF_Err_Table_Missing wmax AF_BLUE_STRINGSET_ADLM af_hani_uniranges AF_BLUE_STRING_NKO_SMALL_BOTTOM af_khmr_dflt_style_class af_sylo_nonbase_uniranges af_armn_script_class af_glyph_hints_scale_dim af_osge_uniranges segment_width_threshold AF_Script_UniRangeRec_ AF_BLUE_STRING_GLAGOLITIC_SMALL_TOP af_cyrl_c2cp_style_class AF_SCRIPT_CPRT AF_BLUE_STRING_ADLAM_CAPITAL_BOTTOM AF_STYLE_CYRL_TITL AF_SCRIPT_KHMR AF_SCRIPT_KHMS p_first AF_WritingSystemClassRec AF_BLUE_STRING_COPTIC_SMALL_BOTTOM AF_STYLE_SINH_DFLT darken_x darken_y AF_Err_Missing_Bbx_Field AF_Err_Invalid_Post_Table AF_STYLE_LATN_TITL AF_STYLE_BUHD_DFLT base_edge AF_Scaler AF_BLUE_STRING_CYRILLIC_CAPITAL_TOP writing_system AF_SCRIPT_CHER AF_COVERAGE_RUBY AF_BLUE_STRING_LATIN_SMALL_DESCENDER AF_STYLE_LATN_C2SC best_y bdelta pp2x_uh af_guru_dflt_style_class link1 af_knda_dflt_style_class AF_BLUE_STRING_VAI_TOP af_face_globals_get_metrics af_tavt_nonbase_uniranges af_copt_script_class AF_BLUE_STRINGSET_GEOK AF_BLUE_STRING_CHEROKEE_CAPITAL AF_BLUE_STRINGSET_GEOR af_khmr_nonbase_uniranges AF_BLUE_STRING_GURMUKHI_BOTTOM af_latn_ordn_style_class AF_BLUE_STRING_TIFINAGH AF_WRITING_SYSTEM_MAX segment_length_threshold af_latn_uniranges style_metrics_getstdw AF_STYLE_ARAB_DFLT ametrics AF_BLUE_STRING_GLAGOLITIC_CAPITAL_BOTTOM af_cjk_hints_apply seg1 af_cakm_script_class af_latin_hints_apply AF_BLUE_STRING_THAI_DIGIT_TOP AF_BLUE_STRING_BUHID_BOTTOM AF_BLUE_STRING_ARMENIAN_CAPITAL_TOP AF_STYLE_LISU_DFLT af_glag_script_class AF_ScriptClassRec AF_BLUE_STRING_SHAVIAN_DESCENDER AF_BLUE_STRING_LATIN_SUPS_SMALL_DESCENDER af_orya_nonbase_uniranges old_charmap AF_BLUE_STRING_DESERET_CAPITAL_TOP AF_STYLE_HEBR_DFLT af_grek_uniranges af_geor_uniranges af_latin_align_serif_edge AF_BLUE_STRING_CJK_BOTTOM AF_Err_Invalid_Stream_Handle AF_StyleMetrics af_cjk_hints_compute_blue_edges standard_horizontal_width af_dummy_hints_init AF_LatinBlue AF_Err_Invalid_Pixel_Size AF_Direction af_indic_hints_init num_idx af_goth_dflt_style_class af_mlym_dflt_style_class af_taml_nonbase_uniranges AF_Err_Post_Table_Missing af_cjk_metrics_scale af_tibt_uniranges is_neutral_blue AF_DIR_LEFT xmax_delta AF_BLUE_STRINGSET_GOTH in_dir AF_BLUE_STRINGSET_ORKH AF_BLUE_STRING_CARIAN_TOP af_khmr_script_class af_olck_script_class AF_BLUE_STRING_GEORGIAN_MKHEDRULI_BOTTOM old_lsb NextContour af_shaw_nonbase_uniranges af_service_properties AF_BLUE_STRINGSET_CYRL AF_Err_Missing_Encoding_Field AF_SCRIPT_HEBR AF_WidthRec_ af_face_globals_compute_style_coverage af_osma_script_class AF_WarperRec af_mlym_uniranges af_arab_script_class AF_Err_Debug_OpCode AF_STYLE_GREK_DFLT AF_BLUE_STRING_KHMER_SUBSCRIPT_TOP AF_SCRIPT_ORYA af_olck_dflt_style_class af_gujr_nonbase_uniranges af_copt_nonbase_uniranges af_shaw_script_class AF_Err_Invalid_Opcode edge_limit AF_Err_Stack_Overflow AF_BLUE_STRINGSET_HEBR af_adlm_dflt_style_class AF_Script af_direction_compute fallback_script d_off2 AF_BLUE_STRING_GREEK_SMALL_BETA_TOP AF_STYLE_CYRL_C2SC AF_BLUE_STRING_GOTHIC_BOTTOM af_kali_nonbase_uniranges default_script af_cyrl_dflt_style_class style_hints_apply dflt AF_BLUE_STRINGSET_HANI width_count AF_STYLE_TAVT_DFLT AF_BLUE_STRINGSET_OSGE AF_Err_Cannot_Render_Glyph laxis num_widths af_avst_script_class is_top_blue AF_STYLE_OLCK_DFLT stem_edge AF_Err_Glyph_Too_Big af_shaper_get_cluster AF_BLUE_STRING_THAI_DESCENDER af_shaw_dflt_style_class af_latb_dflt_style_class af_cyrl_subs_style_class AF_BLUE_STRING_DEVANAGARI_BOTTOM af_guru_script_class blue_edge AF_Err_DEF_In_Glyf_Bytecode point_limit AF_BLUE_STRINGSET_GREK AF_STYLE_DSRT_DFLT segments_end Done_Width AF_BLUE_STRING_LATIN_SUBS_CAPITAL_TOP AF_BLUE_STRING_SAURASHTRA_BOTTOM af_latp_uniranges AF_BLUE_STRING_GREEK_SMALL AF_Err_Too_Many_Caches AF_SCRIPT_SUND AF_BLUE_STRINGSET_LATB af_tavt_dflt_style_class AF_DIR_NONE AF_BLUE_STRINGSET_LATN AF_BLUE_STRINGSET_LATP AF_BLUE_STRING_DESERET_SMALL_BOTTOM is_major_dir af_cprt_dflt_style_class AF_SCRIPT_NONE AF_BLUE_STRING_GREEK_CAPITAL_BOTTOM af_cjk_compute_stem_width fitted af_vaii_uniranges dist1 AF_WritingSystemClass darken_by_font_units_y af_cari_script_class AF_SCRIPT_THAI af_latb_uniranges AF_Edge AF_SCRIPT_ARMN AF_BLUE_STRING_OSMANYA_BOTTOM AF_StyleMetricsRec_ AF_Script_ AF_Err_No_Unicode_Glyph_Name dist_demerit AF_SCRIPT_OLCK AF_BLUE_STRING_GREEK_CAPITAL_TOP AF_Blue_Stringset best_dist pp2x af_tibt_script_class AF_Err_Invalid_Horiz_Metrics af_dsrt_nonbase_uniranges AF_BLUE_STRING_CHEROKEE_SMALL AF_BLUE_STRINGSET_ARAB AF_Dimension AF_BLUE_STRING_CANADIAN_SYLLABICS_SUPS_BOTTOM AF_BLUE_STRING_BAMUM_BOTTOM AF_BLUE_STRING_CANADIAN_SYLLABICS_SMALL_BOTTOM AF_BLUE_STRING_SUNDANESE_TOP AF_BLUE_STRING_DESERET_CAPITAL_BOTTOM af_hani_script_class af_sinh_script_class af_sinh_dflt_style_class AF_Err_Missing_Module AF_STYLE_NONE_DFLT AF_STYLE_ARMN_DFLT AF_Err_Invalid_Cache_Handle af_latin_hints_link_segments Store_Point af_glyph_hints_align_strong_points on_edge af_services AF_BLUE_STRING_THAI_LARGE_DESCENDER xmin_delta AF_STYLE_CYRL_PCAP AF_Err_Max af_tfng_uniranges AF_Blue_String AF_BLUE_STRINGSET_SINH AF_Err_Missing_Chars_Field AF_BLUE_STRING_ARABIC_JOIN AF_StyleClass aglobals AF_STYLE_LATN_PCAP AF_BLUE_STRING_SHAVIAN_SMALL_BOTTOM fallback_style AF_Err_Missing_Bitmap af_bamu_nonbase_uniranges AF_GlyphHints af_indic_metrics_init AF_WritingSystem cur_len best_segment_first AF_BLUE_STRING_LATIN_SUBS_SMALL_F_TOP AF_DIR_RIGHT af_latn_pcap_style_class AF_Err_Cannot_Open_Stream base_distort AF_STYLE_CYRL_ORDN log_base_2 standard_charstring AF_STYLE_THAI_DFLT af_cjk_metrics_init_widths n_edges AF_BLUE_STRINGSET_OSMA af_cari_dflt_style_class digits_have_same_width AF_STYLE_LATN_ORDN edge_delta af_glag_nonbase_uniranges AF_BLUE_STRING_BUHID_LARGE af_cyrl_uniranges AF_SegmentRec_ AF_WRITING_SYSTEM_CJK AF_BLUE_STRING_THAI_ASCENDER af_cprt_uniranges AF_BLUE_STRINGSET_KHMR AF_BLUE_STRINGSET_KHMS AF_BLUE_STRING_CYRILLIC_SMALL af_none_uniranges pp1x AF_Loader slot_internal af_glyph_hints_save AF_WritingSystem_InitHintsFunc AF_STYLE_BENG_DFLT AF_STYLE_GREK_TITL AF_BLUE_STRING_TELUGU_BOTTOM af_latin_metrics_scale started AF_BLUE_STRINGSET_CHER af_blue_1_1 af_deva_script_class AF_LatinMetrics af_kali_dflt_style_class AF_BLUE_STRING_CANADIAN_SYLLABICS_TOP AF_BLUE_STRING_CJK_TOP af_latin_metrics_init af_orya_dflt_style_class af_gujr_script_class af_adlm_uniranges blue_shoot af_grek_smcp_style_class AF_Err_Invalid_Glyph_Format last_stem_pos af_blue_2_1_1 af_blue_2_1_2 AF_PointRec AF_BLUE_STRING_GLAGOLITIC_CAPITAL_TOP AF_Err_Cannot_Open_Resource cur_val af_mymr_nonbase_uniranges AF_BLUE_STRING_DEVANAGARI_TOP AF_BLUE_STRING_ADLAM_CAPITAL_TOP af_orya_uniranges af_latin_compute_stem_width AF_Err_Invalid_Stream_Seek a_scale af_sort_and_quantize_widths AF_BLUE_STRINGSET_TELU flat_threshold AF_Err_Bad_Argument af_latin_metrics_check_digits af_cakm_uniranges link2 AF_BLUE_STRING_CYRILLIC_SMALL_DESCENDER af_cyrl_titl_style_class over_ref contour_index af_shaper_get_coverage af_khms_dflt_style_class AF_SCRIPT_TIBT af_beng_uniranges AF_BLUE_STRING_GEORGIAN_NUSKHURI_TOP af_copt_dflt_style_class base_flags AF_STYLE_GEOR_DFLT af_osma_uniranges prev_max_flags AF_Err_ENDF_In_Exec_Stream af_arab_nonbase_uniranges vvector af_grek_nonbase_uniranges af_latn_dflt_style_class af_geor_script_class af_writing_system_classes af_adlm_script_class af_olck_nonbase_uniranges glyph_count AF_Err_Could_Not_Find_Context num_fills af_cjk_snap_width af_iup_interp AF_SCRIPT_GUJR af_thai_nonbase_uniranges AF_WidthRec cur_ab t2_hints_stems PS_Mask_TableRec_ align_top PSH_Err_Code_Overflow PSH_Err_Stack_Underflow psh_hint_snap_stem_side_delta PS_DimensionRec PSH_Err_Invalid_Stream_Skip PSH_Err_Invalid_PPem alignment strongs_0 pshinter_interface glyphrec PSH_ZoneRec PSH_Err_Missing_Property PSH_DIR_UP PSH_Err_Invalid_Composite cur_top PSH_Hint_TableRec_ ps_dimension_done PSH_AlignmentRec_ PSH_Err_Missing_Chars_Field PS_Mask_TableRec org_ab ps_hint_table_ensure PS_Hint_Table ps_hints_init direction psh_globals_scale_widths psh_glyph_find_strong_points ps_dimension_add_counter PSH_Err_Invalid_Character_Code ps_hints_t1reset psh_glyph_interpolate_other_points PS_HINT_TYPE_1 PSH_Alignment PSH_Err_Raster_Uninitialized hint_tables ps_dimension_init T1_Hints_FuncsRec old_y_scale PSH_Blue_ZoneRec PSH_Err_Raster_Overflow PSH_Err_Invalid_CharMap_Handle psh_globals_new PS_HintsRec psh_glyph_find_blue_points PSH_Err_Table_Missing bit_pos PSH_Err_Cannot_Render_Glyph cur_height fit_count dimension PSH_Hint_TableRec PSH_Err_Too_Many_Hints PSH_Blue_TableRec_ PSH_Glyph finished PSH_Err_Invalid_Argument ps_dimension_add_t1stem PSH_Err_Bad_Argument PSH_DIR_LEFT PSH_Width PSH_Err_Too_Many_Caches PSH_Err_Nested_DEFS scale_ab scale_delta PSH_Err_Too_Many_Extensions org_bottom PSH_Err_Invalid_Outline psh_glyph_compute_extrema cur_max PSH_Err_Nested_Frame_Access ps_hints_stem PSH_Err_Invalid_Cache_Handle PSH_Err_Missing_Encoding_Field PS_Hint_Type read_count PSH_Contour t1_hints_stem PS_HintRec_ PSH_Blue_TableRec PSH_Err_Array_Too_Large max_bits PS_Hinter_Module dir_in psh_glyph_compute_inflections PSH_Err_Corrupted_Font_Glyphs par_cur_center cur_pos PSH_Err_Syntax_Error num_zones dim_x dim_y PSH_Err_Unlisted_Object psh_hint_table_record_mask PSH_Err_Invalid_Version scale_mult fit_len PSH_ContourRec_ do_horz_hints bit_count PS_Hinter_Module_Rec_ PSH_Err_Horiz_Header_Missing ps_hints no_overshoots PSH_Err_Too_Many_Function_Defs PSH_Err_Too_Few_Arguments PSH_Err_Corrupted_Font_Header PS_Dimension normal PSH_DimensionRec sort_global do_horz_snapping no_shoots PSH_Err_Invalid_CharMap_Format n_prev is_others ps_mask_set_bit psh_hint_table_find_strong_points psh_blues_set_zones PSH_Hint_Table PS_Hints PSH_GlyphRec PSH_Err_DEF_In_Glyf_Bytecode PSH_Err_Invalid_Frame_Read min_flag max_masks PSH_Err_No_Unicode_Glyph_Name PSH_Err_Stack_Overflow psh_dimension_quantize_len PSH_Dimension PS_Hint ahint psh_blues_set_zones_0 wmask left_nearest ps_hints_apply t1_hints_funcs_init psh_globals_destroy mask1 align_bot PSH_Err_Invalid_Handle PSH_Err_Lower_Module_Version PSH_Blue_Zone num_masks /home/computerfido/Desktop/freetypetest2/freetype/src/pshinter/pshinter.c rmask PSH_Widths PSH_Err_Invalid_Opcode PSH_BluesRec right_disp orient_prev PS_Mask PS_DimensionRec_ PSH_Err_Raster_Corrupted blue_threshold PSH_Err_Invalid_Glyph_Format PSH_Err_Out_Of_Memory ps_mask_table_merge pshinter_get_globals_funcs psh_globals_set_scale PSH_Err_Invalid_Reference org_ac cur_a PSH_Err_Invalid_Glyph_Index cur_c PSH_HintRec_ ps_mask_table_ensure PSH_Err_Invalid_Face_Handle PSH_Err_Invalid_Slot_Handle cur_u PSH_Hint old_x_scale t2_hints_funcs_init PSH_DimensionRec_ PSH_Err_Missing_Size_Field hint2 ps_mask_table_done ps_mask_test_bit PSH_Err_Invalid_Vert_Metrics ps_hints_close PS_HINT_TYPE_2 PSH_Err_Missing_Module org_top psh_calc_max_height PSH_Err_Unknown_File_Format do_vert_snapping PSH_Err_Invalid_CodeRange PSH_ZoneRec_ PSH_Err_Too_Many_Instruction_Defs ps_hints_t2mask psh_blues_snap_stem count_top stem_bot T2_Hints_FuncsRec hint_masks PSH_Err_Execution_Too_Long ps_hinter_done PSH_Err_Invalid_Stream_Handle ps_dimension_set_mask_bits ps_hints_open psh_hint_table_activate_mask psh_glyph_load_points count1 PSH_Err_ENDF_In_Exec_Stream max_hints ps_hint_table_alloc zone2 count_bot point_dir psh_compute_dir pshinter_get_t2_funcs PSH_Globals_FuncsRec left_disp ps_mask_table_alloc psh_glyph_interpolate_strong_points n_next PSH_Err_Invalid_Stream_Seek stand PSH_Err_Glyph_Too_Big psh_hint_table_align_hints PSH_Err_CMap_Table_Missing PSH_Err_Name_Table_Missing PSH_WidthsRec ps_dimension_end_mask normal_top PSH_Err_Invalid_Table Next_Contour family_top max_scale PSH_Err_Cannot_Open_Stream PSH_DIR_NONE ps_mask_table_merge_all PSH_Err_Invalid_Pixel_Size counter_masks org_v hint1 hint3 flags2 PSH_Err_Cannot_Open_Resource PSH_Err_Invalid_Size_Handle points_end family_bottom cur_bottom PSH_GlyphRec_ PSH_Err_Max PSH_Err_Missing_Startfont_Field ps_hints_t2counter aindex PSH_Err_Hmtx_Table_Missing PSH_Err_Missing_Font_Field PSH_Err_Ignore psh_blues_scale_zones PSH_Err_Invalid_Frame_Operation psh_hint_align PSH_Err_Unimplemented_Feature PSH_WidthRec_ ps_hinter_init cur_org_center source_bits psh_hint_table_record PSH_Err_Raster_Negative_Height orient_cur psh_glyph_interpolate_normal_points counters PSH_WidthsRec_ PS_Hint_TableRec psh_hint_overlap cur_ref delta0 par_org_center PSH_Blues Extremum org_ref right_nearest PSH_Err_Too_Many_Drivers PSH_Zone PSH_Err_Post_Table_Missing psh_hint_table_done psh_hint_table_init PS_Hint_Type_ PSH_PointRec_ PSH_Blue_Table PSH_Err_Invalid_Stream_Operation PS_Hint_TableRec_ PS_MaskRec_ ps_mask_table_set_bits mask2 PSH_DIR_RIGHT stem_top PS_Mask_Table t2_hints_open normal_bottom PSH_Err_Could_Not_Find_Context PSH_Err_Invalid_Library_Handle psh_glyph_done PS_MaskRec source_pos pshinter_get_t1_funcs PSH_Err_Divide_By_Zero ps_mask_table_test_intersect t1_hints_open PS_HintsRec_ do_stem_adjust org_c PSH_Err_Invalid_Stream_Read PSH_AlignmentRec PSH_Err_Invalid_Post_Table_Format minor_dir ps_mask_clear_bit psh_glyph_save_points PSH_Err_Bbx_Too_Big PSH_DIR_DOWN org_a PSH_Err_Invalid_Post_Table num_bits num_strongs do_vert_hints org_u PSH_WidthRec dir_out ps_mask_table_last PSH_Err_Invalid_File_Format PSH_Err_Missing_Bbx_Field PSH_Err_Invalid_Horiz_Metrics PSH_Err_Debug_OpCode hint_mask ps_mask_done PSH_BluesRec_ PSH_Err_Missing_Bitmap psh_globals_funcs_init ps_hints_done hint_type ps_dimension_end do_snapping top_table ps_hint_table_done max_flag PSH_Err_Locations_Missing ps_dimension_reset_mask zone1 psh_hint_table_deactivate ps_hints_t1stem3 PSH_Err_Missing_Startchar_Field amask PSH_Err_Invalid_Offset ps_mask_ensure PSH_Err_Ok count_others psh_glyph_init PSH_Point PSH_Blue_ZoneRec_ bot_table PSH_Err_Missing_Fontboundingbox_Field PSH_Err_Invalid_Driver_Handle Line_Up Raster_Err_Missing_Chars_Field Raster_Err_Nested_DEFS High max_Y Raster_Err_Out_Of_Memory Raster_Err_Could_Not_Find_Context Raster_Err_Unlisted_Object y_turns Decompose_Curve ft_raster1_init lastY Cubic_To joint Raster_Err_Missing_Startfont_Field min_Y Raster_Err_Invalid_File_Format ymin2 Raster_Err_Locations_Missing TStates Raster_Err_Stack_Underflow TProfileList Horizontal_Sweep_Init Raster_Err_Invalid_CharMap_Format black_TBand_ start_arc Raster_Err_Missing_Fontboundingbox_Field Bezier_Down band_stack Raster_Err_Ok precision Sort Bezier_Up ft_raster1_set_mode Raster_Err_Invalid_Table Raster_Err_Invalid_Size_Handle Raster_Err_Invalid_CodeRange P_Right Function_Sweep_Span Raster_Err_Too_Many_Function_Defs draw_left Raster_Err_Invalid_Driver_Handle Raster_Err_CMap_Table_Missing Raster_Err_Raster_Overflow New_Profile target_map ymax1 black_PRaster Raster_Err_Unimplemented_Feature Proc_Sweep_Span Skip_To_Next Raster_Err_Invalid_Character_Code Raster_Err_Raster_Uninitialized InsNew araster Vertical_Sweep_Span y_min Raster_Err_Too_Many_Caches Raster_Err_ENDF_In_Exec_Stream Raster_Err_Invalid_Outline End_Profile ft_black_done Next_Line Raster_Err_Invalid_Post_Table_Format Raster_Err_Divide_By_Zero Raster_Err_Table_Missing Raster_Err_Invalid_Slot_Handle Raster_Err_Too_Many_Extensions Proc_Sweep_Drop Flat_State pool_base Raster_Err_Array_Too_Large Conic_To Raster_Err_Invalid_Reference TPoint Raster_Err_Invalid_Glyph_Index countL precision_bits y_change ymin Unknown_State Horizontal_Sweep_Step ft_black_render PProfileList cProfile band_top Raster_Err_Debug_OpCode Raster_Err_Invalid_Frame_Operation traceOfs Raster_Err_Missing_Size_Field Raster_Err_Corrupted_Font_Glyphs bTarget ft_standard_raster Line_Down Raster_Err_Missing_Encoding_Field Raster_Err_Invalid_Stream_Seek Raster_Err_DEF_In_Glyf_Bytecode ft_black_init P_Left Raster_Err_Cannot_Open_Stream Raster_Err_Invalid_Pixel_Size Raster_Err_Missing_Bbx_Field precision_half Scan_DropOuts ft_raster1_render ft_raster1_get_cbox precision_shift Raster_Err_Missing_Font_Field Raster_Err_Too_Many_Drivers gProfile numTurns Raster_Err_Invalid_PPem arcs num_Profs traceIncr Raster_Err_Horiz_Header_Missing Raster_Err_Invalid_Argument Raster_Err_Invalid_Cache_Handle Convert_Glyph flipped ft_black_reset Raster_Err_Max Raster_Err_Cannot_Open_Resource TProfile Raster_Err_Too_Many_Hints Horizontal_Sweep_Drop Raster_Err_Nested_Frame_Access Raster_Err_Invalid_Stream_Operation scale_shift mode_tag Raster_Err_Invalid_Composite Raster_Err_Cannot_Render_Glyph Raster_Err_Invalid_Vert_Metrics Raster_Err_Code_Overflow black_TBand black_TWorker Raster_Err_Post_Table_Missing Vertical_Sweep_Drop bWidth TSplitter Raster_Err_Too_Few_Arguments sizeBuff maxBuff Raster_Err_Name_Table_Missing dropouts oldProfile lastProfile precision_step Horizontal_Sweep_Span fProfile maxY Raster_Err_Invalid_Stream_Handle Raster_Err_Invalid_CharMap_Handle Raster_Err_Missing_Startchar_Field maxy ft_black_set_mode Raster_Err_Execution_Too_Long Raster_Err_Ignore traceG splitter Raster_Err_Glyph_Too_Big /home/computerfido/Desktop/freetypetest2/freetype/src/raster/raster.c Ascending_State aState dropOutControl black_TWorker_ ft_black_new precision_jitter ymax ymax2 fresh Raster_Err_Hmtx_Table_Missing Vertical_Sweep_Init Raster_Err_Invalid_Offset Raster_Err_Raster_Corrupted Insert_Y_Turn DelOld black_TRaster_ second_pass PByte state_bez Raster_Err_Stack_Overflow PLong Raster_Err_Invalid_Stream_Skip TPoint_ Proc_Sweep_Init Descending_State Raster_Err_Corrupted_Font_Header Render_Single_Pass Raster_Err_Invalid_Handle Raster_Err_Invalid_Stream_Read Split_Conic black_PWorker Raster_Err_Invalid_Opcode Raster_Err_Missing_Property Split_Cubic Function_Sweep_Init Finalize_Profile_Table Raster_Err_No_Unicode_Glyph_Name Init_Linked ft_raster1_transform Vertical_Sweep_Step Raster_Err_Invalid_Frame_Read lastX waiting Raster_Err_Lower_Module_Version Raster_Err_Invalid_Horiz_Metrics Raster_Err_Bbx_Too_Big Set_High_Precision Raster_Err_Missing_Bitmap Raster_Err_Invalid_Glyph_Format Raster_Err_Missing_Module Raster_Err_Too_Many_Instruction_Defs TStates_ Raster_Err_Raster_Negative_Height Line_To minY Draw_Sweep Raster_Err_Invalid_Library_Handle Function_Sweep_Step Raster_Err_Bad_Argument miny Raster_Err_Invalid_Post_Table Proc_Sweep_Step Raster_Err_Invalid_Face_Handle Raster_Err_Syntax_Error Raster_Err_Invalid_Version gTarget TProfile_ PProfile draw_right ymin1 Raster_Err_Unknown_File_Format Smooth_Err_Missing_Startchar_Field Smooth_Err_Hmtx_Table_Missing Smooth_Err_Too_Many_Extensions Smooth_Err_Glyph_Too_Big ft_smooth_render Smooth_Err_Too_Many_Instruction_Defs ft_smooth_set_mode gray_render_conic Smooth_Err_Invalid_File_Format bands gray_raster_reset gray_raster_render gray_move_to Smooth_Err_Invalid_Offset Smooth_Err_Invalid_Horiz_Metrics gray_sweep ft_smooth_render_lcd_v gray_render_line Smooth_Err_Missing_Chars_Field Smooth_Err_Stack_Overflow Smooth_Err_Cannot_Open_Resource Smooth_Err_Missing_Font_Field Smooth_Err_Missing_Fontboundingbox_Field dx_r Smooth_Err_Invalid_Handle TPixmap_ Smooth_Err_Raster_Overflow Smooth_Err_Missing_Size_Field gray_split_conic Smooth_Err_Too_Few_Arguments Smooth_Err_Invalid_Opcode PCell Smooth_Err_Invalid_Outline Smooth_Err_Invalid_Post_Table ft_smooth_render_generic TArea Smooth_Err_Invalid_CodeRange gray_PRaster gray_hline Smooth_Err_Bad_Argument Smooth_Err_Missing_Encoding_Field Smooth_Err_Array_Too_Large gray_raster_new Smooth_Err_Invalid_Table prod pcell Smooth_Err_Invalid_Slot_Handle Smooth_Err_Raster_Negative_Height Smooth_Err_Too_Many_Drivers ft_smooth_transform Smooth_Err_Missing_Bitmap TCell gray_convert_glyph Smooth_Err_Invalid_Glyph_Format Smooth_Err_Locations_Missing Smooth_Err_Unimplemented_Feature gray_raster_done Smooth_Err_Invalid_Size_Handle Smooth_Err_Bbx_Too_Big Smooth_Err_Invalid_Stream_Seek Smooth_Err_Max Smooth_Err_Invalid_Driver_Handle Smooth_Err_Code_Overflow cover Smooth_Err_Lower_Module_Version Smooth_Err_ENDF_In_Exec_Stream Smooth_Err_Missing_Startfont_Field TPixmap Smooth_Err_Invalid_Frame_Operation min_ex gray_PWorker ycells gray_convert_glyph_inner to_x to_y Smooth_Err_Invalid_Stream_Handle ft_smooth_render_lcd Smooth_Err_Invalid_CharMap_Handle max_cells Smooth_Err_Nested_DEFS Split Smooth_Err_Table_Missing /home/computerfido/Desktop/freetypetest2/freetype/src/smooth/smooth.c Smooth_Err_Invalid_Frame_Read gray_set_cell Smooth_Err_Could_Not_Find_Context Smooth_Err_Invalid_Library_Handle __int128 unsigned num_cells min_ey gray_raster_set_mode Smooth_Err_Divide_By_Zero Smooth_Err_DEF_In_Glyf_Bytecode Smooth_Err_Syntax_Error Smooth_Err_Ignore Smooth_Err_Invalid_CharMap_Format Smooth_Err_Invalid_Glyph_Index gray_conic_to gray_TRaster_ Smooth_Err_Missing_Bbx_Field TCoord gray_render_cubic render_span_data bez_stack gray_cubic_to Smooth_Err_Debug_OpCode Smooth_Err_Invalid_Stream_Operation Smooth_Err_No_Unicode_Glyph_Name Smooth_Err_Too_Many_Function_Defs gray_TWorker Smooth_Err_CMap_Table_Missing Smooth_Err_Name_Table_Missing Smooth_Err_Raster_Corrupted Smooth_Err_Cannot_Open_Stream ft_smooth_init required_mode Smooth_Err_Stack_Underflow Smooth_Err_Invalid_Pixel_Size Smooth_Err_Invalid_Face_Handle hmul gray_TWorker_ Smooth_Err_Invalid_Stream_Skip Smooth_Err_Raster_Uninitialized clip gray_record_cell Smooth_Err_Invalid_Stream_Read draw TCell_ Smooth_Err_Invalid_Composite ft_grays_raster Smooth_Err_Invalid_Argument Smooth_Err_Invalid_PPem Smooth_Err_Nested_Frame_Access Smooth_Err_Unlisted_Object Smooth_Err_Invalid_Character_Code ft_smooth_get_cbox vmul Smooth_Err_Invalid_Vert_Metrics gray_split_cubic Smooth_Err_Invalid_Cache_Handle Smooth_Err_Out_Of_Memory TPos Smooth_Err_Too_Many_Caches max_ex max_ey Smooth_Err_Post_Table_Missing Smooth_Err_Horiz_Header_Missing Smooth_Err_Cannot_Render_Glyph Smooth_Err_Invalid_Post_Table_Format band Smooth_Err_Too_Many_Hints gray_line_to Smooth_Err_Invalid_Reference Smooth_Err_Corrupted_Font_Glyphs Smooth_Err_Missing_Property Smooth_Err_Missing_Module Smooth_Err_Ok Smooth_Err_Execution_Too_Long dy_r render_span Smooth_Err_Invalid_Version Smooth_Err_Corrupted_Font_Header Smooth_Err_Unknown_File_Format WASH ft_gzip_file_skip_output ft_gzip_alloc voidpf Gzip_Err_Invalid_Vert_Metrics nowrap Gzip_Err_Post_Table_Missing inflate_codes_new Gzip_Err_Invalid_Table CHECK1 Gzip_Err_Invalid_Cache_Handle total_in Gzip_Err_Missing_Size_Field Gzip_Err_Ok window Gzip_Err_Invalid_Slot_Handle zalloc fixed_bd Gzip_Err_Array_Too_Large fixed_bl Gzip_Err_Missing_Fontboundingbox_Field Gzip_Err_Execution_Too_Long Gzip_Err_Invalid_Offset zstream Gzip_Err_Max z_stream CODES inflate_block_mode /home/computerfido/Desktop/freetypetest2/freetype/src/gzip/ftgzip.c Gzip_Err_Invalid_Horiz_Metrics Gzip_Err_Stack_Overflow ft_gzip_file_fill_output Gzip_Err_Hmtx_Table_Missing inflate_codes_free check_func inflate_mask inflate total_out cpdext Gzip_Err_Invalid_Size_Handle __mlibc_errno checkfn Gzip_Err_Invalid_Opcode Gzip_Err_Corrupted_Font_Glyphs Gzip_Err_Code_Overflow uLong Gzip_Err_Missing_Property Gzip_Err_DEF_In_Glyf_Bytecode adler DICT1 DICT2 DICT3 DICT4 inflate_codes_state inflateReset FT_GZipFileRec_ Bytef Gzip_Err_Ignore TABLE marker trees BLOCKS inflateEnd inflate_trees_bits Gzip_Err_Missing_Bitmap Gzip_Err_Invalid_Stream_Operation DISTEXT Gzip_Err_Debug_OpCode inflate_huft_s zip_buff Gzip_Err_Too_Many_Drivers DTREE Gzip_Err_Invalid_PPem Gzip_Err_Table_Missing next_out Gzip_Err_Nested_Frame_Access Gzip_Err_Missing_Bbx_Field INFLATE_DONE inflate_blocks_reset decode Gzip_Err_Invalid_Argument BADCODE inflate_flush Gzip_Err_Missing_Encoding_Field avail_out lbits Gzip_Err_Invalid_Post_Table Gzip_Err_Invalid_Glyph_Index program_invocation_name method Gzip_Err_Raster_Negative_Height Gzip_Err_Too_Many_Function_Defs Gzip_Err_No_Unicode_Glyph_Name CHECK2 CHECK3 CHECK4 zcalloc Gzip_Err_Unimplemented_Feature inflate_blocks_free ft_gzip_file_reset Gzip_Err_Syntax_Error Bits inflate_blocks_statef inflateInit2_ inflate_codes need Gzip_Err_Missing_Chars_Field inflate_huft dtree ft_gzip_file_done Gzip_Err_ENDF_In_Exec_Stream Gzip_Err_Invalid_Composite inflate_trees_fixed COPY z_stream_s ft_gzip_get_uncompressed_size Gzip_Err_Invalid_Stream_Seek FT_GZipFile alloc_func free_func Gzip_Err_Stack_Underflow avail_in Gzip_Err_Glyph_Too_Big Gzip_Err_Raster_Corrupted uLongf z_streamp bitb Gzip_Err_Invalid_Post_Table_Format bitk inflate_blocks_state Gzip_Err_Invalid_Reference BTREE Gzip_Err_Divide_By_Zero dbits zcfree Gzip_Err_Out_Of_Memory Gzip_Err_Raster_Uninitialized Gzip_Err_Lower_Module_Version Gzip_Err_Unlisted_Object Gzip_Err_Raster_Overflow ft_gzip_file_init ft_gzip_stream_close Gzip_Err_Could_Not_Find_Context opaque Gzip_Err_Cannot_Render_Glyph uIntf Gzip_Err_Invalid_Face_Handle ft_gzip_file_io inflate_trees_dynamic fixed_td fixed_tl Gzip_Err_Locations_Missing Gzip_Err_Too_Many_Caches Gzip_Err_Invalid_CharMap_Format Gzip_Err_Corrupted_Font_Header Gzip_Err_Invalid_Frame_Read what Gzip_Err_Invalid_Outline inflate_mode Gzip_Err_Too_Many_Instruction_Defs next_in program_invocation_short_name METHOD adler32 INFLATE_BAD Gzip_Err_Unknown_File_Format Gzip_Err_Bad_Argument Gzip_Err_Too_Few_Arguments Gzip_Err_Too_Many_Extensions LENEXT ltree inflate_blocks_new input_len Gzip_Err_Missing_Startchar_Field Gzip_Err_Invalid_Version Gzip_Err_Nested_DEFS ft_gzip_free Exop Gzip_Err_Invalid_File_Format Gzip_Err_Missing_Startfont_Field cpdist ft_gzip_stream_io Gzip_Err_Invalid_Frame_Operation Gzip_Err_Invalid_Handle Gzip_Err_Invalid_Driver_Handle inflate_blocks ft_gzip_check_header old_pos Gzip_Err_CMap_Table_Missing ft_gzip_file_fill_input Gzip_Err_Invalid_Stream_Skip Gzip_Err_Invalid_Glyph_Format Gzip_Err_Name_Table_Missing zfree data_type uInt Gzip_Err_Invalid_Stream_Read Gzip_Err_Horiz_Header_Missing Gzip_Err_Cannot_Open_Stream Gzip_Err_Invalid_Pixel_Size zip_size huft_build cplens DIST STORED Gzip_Err_Invalid_Character_Code Gzip_Err_Too_Many_Hints Gzip_Err_Missing_Font_Field Gzip_Err_Invalid_Stream_Handle stream_size Gzip_Err_Invalid_CharMap_Handle Gzip_Err_Invalid_CodeRange inflate_codes_mode Gzip_Err_Missing_Module internal_state border LENS blens Gzip_Err_Invalid_Library_Handle cplext inflate_codes_statef Gzip_Err_Cannot_Open_Resource hufts Gzip_Err_Bbx_Too_Big DICT0 wbits ft_lzw_file_done LZW_Err_Invalid_Glyph_Index LZW_Err_Missing_Size_Field LZW_Err_Out_Of_Memory LZW_Err_Could_Not_Find_Context LZW_Err_Invalid_Library_Handle stack_top LZW_Err_Invalid_Frame_Read LZW_Err_Invalid_CharMap_Format LZW_Err_Stack_Overflow LZW_Err_Missing_Bbx_Field NextCode LZW_Err_Invalid_Horiz_Metrics LZW_Err_Invalid_Face_Handle ft_lzw_stream_close LZW_Err_Invalid_Opcode LZW_Err_Locations_Missing LZW_Err_Syntax_Error LZW_Err_Invalid_Stream_Skip LZW_Err_Cannot_Open_Resource LZW_Err_Too_Few_Arguments LZW_Err_Invalid_Stream_Read ft_lzw_file_reset LZW_Err_Missing_Bitmap LZW_Err_Invalid_Vert_Metrics LZW_Err_Nested_DEFS LZW_Err_Debug_OpCode LZW_Err_Missing_Module ft_lzwstate_refill old_char LZW_Err_Max LZW_Err_Horiz_Header_Missing ft_lzw_stream_io LZW_Err_Invalid_Composite LZW_Err_Invalid_Stream_Operation FT_LzwStateRec LZW_Err_Invalid_Post_Table_Format prefix_size LZW_Err_Array_Too_Large buf_total LZW_Err_Invalid_Stream_Handle FT_LZW_PHASE_START ft_lzw_check_header LZW_Err_Cannot_Render_Glyph LZW_Err_Invalid_Argument LZW_Err_Post_Table_Missing FT_LZW_PHASE_CODE free_bits out_size ft_lzw_file_fill_output LZW_Err_Invalid_CharMap_Handle LZW_Err_Ignore old_size LZW_Err_Invalid_Offset LZW_Err_Invalid_PPem ft_lzw_file_skip_output buf_clear ft_lzw_file_io LZW_Err_Invalid_Reference LZW_Err_DEF_In_Glyf_Bytecode LZW_Err_Too_Many_Instruction_Defs LZW_Err_Missing_Chars_Field LZW_Err_Invalid_Driver_Handle buf_tab LZW_Err_Bbx_Too_Big LZW_Err_No_Unicode_Glyph_Name ft_lzwstate_get_code LZW_Err_Unimplemented_Feature LZW_Err_Too_Many_Hints FT_LzwStateRec_ LZW_Err_Invalid_Table LZW_Err_Invalid_File_Format LZW_Err_CMap_Table_Missing LZW_Err_Name_Table_Missing LZW_Err_Too_Many_Function_Defs LZW_Err_Cannot_Open_Stream LZW_Err_Invalid_Pixel_Size LZW_Err_Lower_Module_Version FT_LZWFile FT_LZW_PHASE_STACK LZW_Err_Invalid_Handle LZW_Err_Raster_Corrupted LZW_Err_Missing_Font_Field FT_LzwPhase_ ft_lzwstate_reset LZW_Err_Invalid_Glyph_Format stack_0 LZW_Err_Missing_Property FT_LzwState LZW_Err_Raster_Negative_Height LZW_Err_Divide_By_Zero LZW_Err_Too_Many_Extensions LZW_Err_Code_Overflow suffix FT_LZW_PHASE_EOF LZW_Err_Missing_Fontboundingbox_Field ft_lzwstate_prefix_grow LZW_Err_Corrupted_Font_Glyphs LZW_Err_Glyph_Too_Big FT_LZWFileRec_ LZW_Err_Execution_Too_Long LZW_Err_Invalid_CodeRange LZW_Err_Invalid_Slot_Handle LZW_Err_Table_Missing LZW_Err_Corrupted_Font_Header LZW_Err_Stack_Underflow ft_lzwstate_done LZW_Err_Missing_Encoding_Field LZW_Err_Hmtx_Table_Missing ft_lzw_file_init old_code ft_lzwstate_stack_grow LZW_Err_ENDF_In_Exec_Stream LZW_Err_Bad_Argument LZW_Err_Ok LZW_Err_Invalid_Size_Handle LZW_Err_Raster_Overflow LZW_Err_Raster_Uninitialized numread LZW_Err_Invalid_Stream_Seek LZW_Err_Invalid_Character_Code LZW_Err_Missing_Startchar_Field LZW_Err_Missing_Startfont_Field LZW_Err_Too_Many_Caches LZW_Err_Invalid_Frame_Operation LZW_Err_Invalid_Outline ft_lzwstate_init LZW_Err_Too_Many_Drivers FT_LzwPhase /home/computerfido/Desktop/freetypetest2/freetype/src/lzw/ftlzw.c LZW_Err_Unknown_File_Format LZW_Err_Nested_Frame_Access ft_lzwstate_io LZW_Err_Invalid_Cache_Handle LZW_Err_Unlisted_Object LZW_Err_Invalid_Version LZW_Err_Invalid_Post_Table buf_offset free_ent in_eof max_free in_code cf2_builder_lineTo FieldArray CF2_Err_Missing_Startchar_Field bitCount PSaux_Err_Syntax_Error moveUp op_endchar cf2_hint_isPair AFM_VALUE_TYPE_STRING haveWidth ps_table_new needWinding PSaux_Err_Missing_Startchar_Field aint CF2_Matrix_ cf2_cmdRLINETO cf2_stack_pushFixed vStemHintArray max_tokens summand1 cf2_escRANDOM AFM_TOKEN_CAPHEIGHT CF2_Err_Too_Many_Instruction_Defs AFM_TOKEN_XHEIGHT cf2_hintmask_setCounts charstring_base PSaux_Err_Invalid_Post_Table_Format cff_builder_start_point PSaux_Err_Table_Missing in_offset darkenX darkenY afm_key_table T1_CMapStd t1_cmap_custom_init PSaux_Err_Invalid_Glyph_Index currentCS PSaux_Err_Unknown_File_Format PSaux_Err_Bad_Argument cf2_cmdCALLGSUBR cf2_arrstack_init CF2_PathOpQuadTo topHintEdge initialHintMap csFlatEdge CF2_Err_Invalid_Version CF2_BluesRec charstringIndex AFM_TOKEN_STARTKERNDATA otherBlues PSaux_Err_Name_Table_Missing PSaux_Err_Invalid_PPem CF2_StackNumber_ ps_builder_done cf2_hint_isPairTop op_hlineto flatFamilyEdge CF2_MAX_HINTS curp familyBlues cff_decoder cff_builder_funcs ps_tobool captured currentDS ps_table_release PSaux_Err_Invalid_Reference cf2_escGET CF2_Err_Corrupted_Font_Glyphs PSaux_Err_Corrupted_Font_Header cf2_buf_isEnd PSaux_Err_Too_Many_Instruction_Defs logBase2 AFM_TOKEN_VVECTOR t1_builder_add_contour CF2_Err_Corrupted_Font_Header CF2_BufferRec AFM_TOKEN_W1X CF2_Err_Invalid_CharMap_Format normalizedV t1_cmap_expert_init emBoxTop emBoxBottomEdge psaux_get_glyph_name cf2_cmdRESERVED_17 PSaux_Err_Missing_Chars_Field renderingFlags upMoveDown CF2_Err_Too_Many_Extensions PSaux_Err_Missing_Bitmap cf2_escFLEX1 PSaux_Err_Raster_Corrupted cf2_cmdBLEND afm_stream_read_one intersection cf2_glyphpath_computeIntersection hintOffset t1_cmap_std_init PSaux_Err_Missing_Module CF2_HintRec PSaux_Err_Cannot_Open_Resource CF2_Err_Invalid_Handle cf2_cmdCNTRMASK emRatio FT_Fast op_hsbw cf2_stack_popInt dsCoord AFM_VALUE_TYPE_INTEGER PSAux_Interface sizeItem t1_lookup_glyph_by_stdcharcode_ps AFM_TOKEN_STARTCOMPOSITES AFM_TOKEN_W0X AFM_TOKEN_W0Y AFM_TOKEN_AXISTYPE CF2_Outline factor2 cf2_getNominalWidthX AFM_VALUE_TYPE_FIXED PSaux_Err_Invalid_Slot_Handle CF2_Err_Bbx_Too_Big blueFuzz cf2_cmdHMOVETO cf2_getT1SeacComponent CF2_Err_Debug_OpCode cf2_cmdVSINDEX PSaux_Err_ENDF_In_Exec_Stream AFM_TOKEN_STARTKERNPAIRS1 cf2_stack_clear PSaux_Err_Lower_Module_Version op_vhcurveto CF2_Err_Invalid_Face_Handle cf2_hint_isValid flatEdge CF2_Err_Invalid_Stream_Read get_callback cf2_getOtherBlues AFM_TOKEN_CC AFM_TOKEN_CH ps_parser_skip_spaces cf2_hintmask_init CF2_StackNumber cf2_glyphpath_curveTo PSaux_Err_Glyph_Too_Big AFM_Token cf2_hintmap_dump CF2_Err_Code_Overflow cf2_cmdVSTEMHM t1_cmap_std_char_index have_underflow hStemHintArray cf2_hintmap_build ps_table_add CF2_Err_Glyph_Too_Big PSaux_Err_Invalid_Argument chunk PSaux_Err_Missing_Bbx_Field PSaux_Err_Cannot_Render_Glyph AFM_TOKEN_FONTNAME pflags cff_builder_add_point known_othersubr_result_cnt op_hstem cf2_escDUP AFM_TOKEN_NOTICE scaleX scaleY snapThreshold cf2_escMUL cf2_escNOT darkenAmount CF2_GhostTop fracUp PSaux_Err_Execution_Too_Long pathIsClosing glyphWidth ps_builder_add_contour afm_parse_kern_pairs bottomHintEdge doConditionalLastRead cf2_escPUT ps_parser_load_field_table end_section CF2_NumberType_ CF2_Err_Missing_Chars_Field emBoxBottom CF2_Err_Missing_Module skip_procedure CF2_PairBottom CF2_Err_Missing_Font_Field cf2_hint_lock curX curY skip_literal_string op_div CF2_Callback_Type t1_cmap_standard_init cf2_getScaleAndHintFlag afm_stream_read_string CF2_NumberFrac cf2_cmdVHCURVETO ps_parser_to_fixed_array ps_parser_to_int lsb_x lsb_y subtrahend CF2_Err_Invalid_Opcode CF2_Err_Cannot_Open_Resource doEmBoxHints instructionLimit afm_parse_kern_data CF2_HintMaskRec_ dsMove ps_table_done CF2_HintMove cf2_builder_cubeTo cf2_getBlueValues cf2_arrstack_finalize CF2_HintMoveRec PSaux_Err_Invalid_Stream_Seek CF2_NumberInt op_rrcurveto PSaux_Err_Raster_Overflow cf2_cmdHHCURVETO CF2_Err_Missing_Startfont_Field AFM_TOKEN_ITALICANGLE AFM_TOKEN_C CF2_Err_Post_Table_Missing CF2_Blues AFM_TOKEN_L cond2 AFM_TOKEN_N PSaux_Err_Invalid_Post_Table PSaux_Err_Stack_Underflow arrstack AFM_TOKEN_STARTAXIS cf2_arrstack_push t1_cmap_unicode_char_index PSaux_Err_Debug_OpCode AFM_TOKEN_ENDCOMPOSITES AFM_TOKEN_METRICSSETS cf2_glyphpath_closeOpenPath cf2_escRESERVED_8 CF2_HintMask shared_vals cf2_free_instance dummyWidth cf2_escSETCURRENTPT prevP0 cff_decoder_init xOffset1 xOffset3 ps_parser_to_fixed afm_parser_read_int elemIsQueued Unexpected_OtherSubr cf2_outline_init PSaux_Err_Missing_Fontboundingbox_Field AFM_TOKEN_ENDAXIS ps_builder_funcs PS_Conv_EexecDecode CF2_Err_Stack_Underflow PSaux_Err_DEF_In_Glyf_Bytecode afm_compare_kern_pairs PSaux_Err_Out_Of_Memory secondHintEdge AFM_STREAM_STATUS_EOL stemWidthPer1000 bchar_index cf2_cmdHLINETO CF2_Locked cf2_cmdHINTMASK CF2_Err_Invalid_Stream_Handle outerTransform AFM_TOKEN_CHARACTERSET cf2_setError AFM_TOKEN_BLENDDESIGNMAP in_charstring_type CF2_ArrStackRec_ ps_builder_init PSaux_Err_Could_Not_Find_Context AFM_TOKEN_ENCODINGSCHEME yOffset3 CF2_Err_Invalid_Horiz_Metrics t1_builder_done glyphpath boost cf2_hintmap_isValid PSaux_Err_Too_Many_Caches hintmap cf2_stack_pop maskByte CF2_Err_Invalid_Post_Table_Format CF2_BufferRec_ CF2_GlyphPath op_callothersubr reverseWinding PSaux_Err_Invalid_Pixel_Size cf2_cmdHSBW hintOriginY AFM_TOKEN_ISFIXEDPITCH windingMomentum AFM_TOKEN_ENDKERNPAIRS decimal iSrc AFM_TOKEN_ENDKERNDATA cff_builder_done cf2_computeDarkening downMoveUp cf2_hintmap_init cf2_blues_init CF2_Err_Invalid_Glyph_Index reallocate_t1_table CF2_RenderingFlags PSaux_Err_Too_Few_Arguments op_dotsection CF2_Err_Invalid_Library_Handle psaux_driver_class upMinCounter CF2_Err_Bad_Argument AFM_TOKEN_WEIGHTVECTOR CF2_Err_Unknown_File_Format innerTransform maskPtr cf2_getBlueMetrics AFM_VALUE_TYPE_BOOL op_setcurrentpoint PSaux_Err_Raster_Negative_Height PS_Conv_Strtol cf2_hint_isBottom PS_Conv_ASCIIHexDecode cf2_stack_count AFM_TOKEN_ISBASEFONT doingSeac cf2_doBlend ps_parser_to_bytes cf2_builder_moveTo CF2_StackRec_ isCFF2 AFM_TOKEN_STARTFONTMETRICS cf2_getPpemY opIdx PSaux_Err_Invalid_Stream_Operation cf2_initGlobalRegionBuffer CF2_Err_Too_Many_Hints CF2_OutlineCallbacksRec_ cff_builder_close_contour iDst stemHint cf2_hint_isSynthetic ps_builder_check_points CF2_Err_Invalid_Frame_Read PSaux_Err_Invalid_CodeRange t1_cmap_custom_class_rec PSaux_Err_Nested_Frame_Access CF2_Err_Unimplemented_Feature blueValues cf2_hintmask_getMaskPtr cf2_glyphpath_lineTo prevElemP0 prevElemP3 cf2_escDROP code_to_sid cf2_cmdVVCURVETO CF2_ICF_Top t1_cmap_unicode_done CF2_NumberType ps_parser_to_token_array FT_UFast CF2_Err_Invalid_CodeRange CF2_Err_Raster_Uninitialized CF2_PathOp_ numElements embed PSaux_Err_Invalid_Size_Handle minDS indexStemHint cf2_cmdCLOSEPATH CF2_Err_Locations_Missing CF2_Font cf2_freeT1SeacComponent PSaux_Err_Too_Many_Drivers PSaux_Err_Too_Many_Hints opStack CF2_Err_Invalid_Outline cf2_cmdVSTEM cf2_getVStore CF2_ArrStack op_rmoveto PSaux_Err_Invalid_Library_Handle CF2_Err_Nested_Frame_Access CF2_Err_Missing_Size_Field CF2_Err_Table_Missing csBottomEdge ps_builder_add_point AFM_TOKEN_STARTKERNPAIRS0 cf2_escVSTEM3 CF2_Err_Divide_By_Zero initial_map_ready csFuzz CF2_Stack PSaux_Err_Cannot_Open_Stream cf2_glyphpath_hintPoint csUnitsPerPixel stemHintArray cf2_arrstack_getPointer cf2_glyphpath_moveTo t1builder T1_CMap_ClassesRec cf2_escHSTEM3 T1_CMapCustomRec_ cf2_arrstack_size CF2_Err_CMap_Table_Missing is_expert CF2_Err_Invalid_Character_Code CF2_OutlineCallbacks metrics_sets cf2_initLocalRegionBuffer op_pop cf2_stack_getReal t1_builder_start_point no_stem_darkening_driver cf2_cmdHSTEM cf2_cmdEXTENDEDNMBR AFM_Token_ PSaux_Err_Invalid_Character_Code numOtherBlues CF2_Err_Syntax_Error cf2_hintmask_read AFM_TOKEN_BLENDDESIGNPOSITIONS AFM_TOKEN_ENDCHARMETRICS PSaux_Err_Invalid_Table num_elements start_idx callbacks AFM_TOKEN_KPH AFM_TOKEN_KPX AFM_TOKEN_KPY afm_parse_track_kern PSaux_Err_Invalid_Version CF2_Err_Stack_Overflow lastVal CF2_Err_Invalid_CharMap_Handle ps_parser_skip_PS_token PS_Conv_ToFixed op_hstem3 CF2_Err_Missing_Encoding_Field prevElemOp AFM_TOKEN_ENDDIRECTION prevElemP2 cff_decoder_prepare CF2_Err_Name_Table_Missing t1_decoder cf2_getStdHW t1_cmap_custom_char_index ps_parser_to_coord_array cf2_getFamilyBlues PSaux_Err_Missing_Font_Field cf2_getFamilyOtherBlues CF2_Err_Could_Not_Find_Context PSaux_Err_Invalid_Cache_Handle cf2_cmdRLINECURVE fractionalTranslation counterHintMap CF2_HintMoveRec_ initialMap t1_decoder_init op_sbw CF2_OutlineRec_ prevP1 CF2_MAX_HINT_EDGES old_cur PSaux_Err_Max cf2_interpT2CharString cf2_cmdVLINETO CF2_OutlineRec N_AFM_TOKENS ft_char_table syntheticEmboldeningAmountX syntheticEmboldeningAmountY CF2_Err_Invalid_Slot_Handle PSaux_Err_Invalid_Stream_Skip acur AFM_TOKEN_UNDERLINEPOSITION old_base cf2_getUnitsPerEm factor1 t1_builder_init AFM_TOKEN_FULLNAME cff_builder_add_contour useIntersection op_hmoveto AFM_TOKEN_CHARWIDTH AFM_ValueRec PSaux_Err_Ok CF2_Err_Missing_Bbx_Field psaux_interface cf2_cmdVMOVETO cf2_cmdCALLSUBR op_vlineto cf2_hint_isLocked cf2_escRESERVED_38 AFM_TOKEN_TRACKKERN counterMask flexStore scaledStem cf2_getSubfont AFM_TOKEN_ISFIXEDV hintMap ps_builder_add_point1 newSize downMoveDown CF2_Err_Invalid_Cache_Handle AFM_VALUE_TYPE_NAME CF2_CallbackParamsRec CF2_Err_Hmtx_Table_Missing cf2_escPOP cf2_cmdRETURN PSaux_Err_Missing_Property CF2_PathOpMoveTo cf2_escRESERVED_13 readFromStack AFM_TOKEN_ENDFONTMETRICS PSaux_Err_Invalid_Driver_Handle cf2_cmdRMOVETO PS_Conv_ToInt T1_Operator_ csTopEdge gr_idx cf2_escSQRT CF2_Err_Missing_Bitmap op_callsubr PSaux_Err_Ignore newHintMap t1_cmap_custom_char_next cf2_outline_close CF2_Err_Missing_Property newPtr miterLimit cf2_getMaxstack cf2_escDOTSECTION AFM_TOKEN_KP cf2_escINDEX CF2_Err_Too_Many_Drivers prevElemP1 cf2_cmdHSTEMHM scaleC CF2_Err_Raster_Corrupted PSaux_Err_Array_Too_Large CF2_HintMapRec_ op_rlineto cf2_stack_init free_callback CF2_Err_Raster_Overflow cf2_escRESERVED_25 byteCount CF2_Err_Invalid_Glyph_Format PSaux_Err_Too_Many_Extensions max_bytes achar cf2_escFLEX AFM_TOKEN_ESCCHAR CF2_CallbackParamsRec_ afm_parser_init CF2_StemHintRec cf2_escSUB summand2 cf2_arrstack_setCount cf2_doFlex CF2_Err_Invalid_Frame_Operation t1_decoder_parse_metrics cff_compute_bias PSaux_Err_Invalid_Handle cf2_glyphpath_init afm_parser_skip_section CF2_Matrix CF2_HintMap cf2_buf_readByte cf2_stack_pushInt CF2_StemHint PSaux_Err_Corrupted_Font_Glyphs moveIsPending numFamilyOtherBlues CF2_Err_Cannot_Render_Glyph cf2_escRESERVED_31 CF2_PathOpCubeTo translation isHFlex PSaux_Err_CMap_Table_Missing CF2_Err_Nested_DEFS PSaux_Err_Horiz_Header_Missing PSaux_Err_Invalid_Stream_Handle cf2_getDefaultWidthX quadTo sid_to_string ps_parser_done PSaux_Err_Unlisted_Object delimiters CF2_BlueRec afm_parser_done t1_cmap_expert_class_rec cf2_glyphpath_finalize hintOrigin hasVariations CF2_HintRec_ AFM_TOKEN_BLENDAXISTYPES boldenX CF2_Err_DEF_In_Glyf_Bytecode nextP0 midpoint cf2_glyphpath_pushMove AFM_TOKEN_STDHW fieldrec CF2_Err_Array_Too_Large AFM_TOKEN_CHARACTERS dividend PSaux_Err_Invalid_Glyph_Format cf2_getWindingMomentum AFM_TOKEN_FONTBBOX pnum_bytes pnum_tokens zoneHeight PSaux_Err_Invalid_File_Format savedMove CF2_Err_Invalid_Composite ps_builder_close_contour CF2_Err_Horiz_Header_Missing cff_check_points max_values stemhint CF2_Err_Unlisted_Object cond1 ps_tocoordarray afm_stream_skip_spaces Store_Integer cf2_hintmap_insertHint CF2_Err_Out_Of_Memory cf2_checkTransform cf2_escHFLEX1 AFM_TOKEN_STDVW CF2_Err_Invalid_Stream_Seek AFM_TOKEN_UNKNOWN cf2_cmdHVCURVETO CF2_Err_Invalid_Size_Handle AFM_TOKEN_B needExtraSetup cf2_escOR CF2_ArrStackRec advWidth boldenAmount t1_args_count CF2_Err_Too_Few_Arguments stemDarkened CF2_OutlineCallbacksRec subrStack firstHintEdge integral cf2_arrstack_getBuffer bchar ps_parser_to_token maxScale hintMoves PSaux_Err_Raster_Uninitialized ps_decoder /home/computerfido/Desktop/freetypetest2/freetype/src/psaux/psaux.c AFM_TOKEN_AXISLABEL minuend AFM_TOKEN_ENDTRACKKERN AFM_TOKEN_UNDERLINETHICKNESS CF2_FontRec_ cf2_escRESERVED_32 cff_lookup_glyph_by_stdcharcode cf2_escSBW cf2_getStdVW cf2_cmdENDCHAR PSaux_Err_Invalid_Opcode lenNormalizedV PSaux_Err_Stack_Overflow afm_tokenize PSaux_Err_No_Unicode_Glyph_Name PSaux_Err_Missing_Startfont_Field cf2_stack_setReal suppressOvershoot op_vstem AFM_STREAM_STATUS_EOF CF2_Err_Raster_Negative_Height CF2_Err_No_Unicode_Glyph_Name CF2_HintMapRec AFM_TOKEN_DESCENDER AFM_ValueRec_ CF2_CallbackParams upMoveUp PSaux_Err_Post_Table_Missing ps_parser_init pathIsOpen PSaux_Err_Invalid_CharMap_Handle PSaux_Err_Code_Overflow T1_Operator AFM_VALUE_TYPE_INDEX CF2_Err_Invalid_Driver_Handle CF2_GlyphPathRec_ byte2 cf2_escHFLEX numFamilyBlues cf2_setGlyphWidth darken PSaux_Err_Divide_By_Zero lastIndex cf2_escAND indexInsert isT1 op_return op_vstem3 byte4 CF2_Err_Invalid_File_Format CF2_Err_Too_Many_Function_Defs AFM_Value CF2_Err_Execution_Too_Long CF2_Frac CF2_F16Dot16 CF2_Err_Cannot_Open_Stream AFM_TOKEN_VV byte3 AFM_TOKEN_W0 AFM_TOKEN_W1 AFM_TOKEN_ASCENDER CF2_Err_Invalid_Argument ps_parser_load_field t1_cmap_unicode_init PSaux_Err_Invalid_CharMap_Format cf2_glyphpath_pushPrevElem cf2_hintmap_adjustHints hasWidthArg PSaux_Err_Invalid_Frame_Read subr_no idx2 T1_CMapCustom AFM_TOKEN_WX AFM_TOKEN_WY byte1 CF2_HintMaskRec cf2_freeSeacComponent PSAux_ServiceRec CF2_Err_Missing_Fontboundingbox_Field cf2_cmdRCURVELINE t1_cmap_custom_done cf2_cmdRESERVED_2 t1_cmap_standard_class_rec firstHintMap t1_cmap_std_done numBlueValues CF2_BluesRec_ PSaux_Err_Missing_Encoding_Field PSaux_Err_Invalid_Outline CF2_GlyphPathRec cf2_getLanguageGroup no_stem_darkening_font op_none cf2_escNEG PSaux_Err_Too_Many_Function_Defs skip_comment afm_parser_next_key PSaux_Err_Invalid_Composite saveEdge skip_string emBoxTopEdge t1_builder_add_point AFM_STREAM_STATUS_EOC AFM_ValueType_ alternate op_vmoveto CF2_Synthetic cf2_hintmask_setAll AFM_TOKEN_FAMILYNAME AFM_TOKEN_STARTCHARMETRICS PSaux_Err_Invalid_Offset cff_builder_add_point1 CF2_Err_Invalid_Post_Table cf2_decoder_parse_charstrings offsetStart0 cf2_stack_roll PSaux_Err_Missing_Size_Field No_Width CF2_ICF_Bottom cf2_doStems dsFlatEdge achar_index op_seac divider CF2_Hint lastSubfont PSaux_Err_Bbx_Too_Big cf2_hintmask_isValid moveDown CF2_PathOpLineTo maxDS PSaux_Err_Invalid_Horiz_Metrics AFM_TOKEN_STARTDIRECTION minDiff PSaux_Err_Invalid_Face_Handle PSaux_Err_Invalid_Stream_Read cf2_hintmask_setNew ps_tofixedarray AFM_TOKEN_MAPPINGSCHEME cffbuilder cf2_cmdRRCURVETO cf2_escSEAC cf2_glyphpath_computeOffset cf2_hint_initZero cf2_escEQ t1_builder_add_point1 AFM_STREAM_STATUS_NORMAL max_coords cf2_escEXCH CF2_Err_Max yOffset1 AFM_TOKEN_PCC cf2_cmdESC AFM_TOKEN_STARTTRACKKERN halfWidth dsNew bottomZone CF2_Err_Invalid_Stream_Skip AFM_TOKEN_VERSION CF2_NumberFixed PSaux_Err_Invalid_Vert_Metrics cf2_font_setup afm_parser_read_vals cf2_arrstack_setNumElements hintMask op_hvcurveto t1_cmap_unicode_class_rec subrNum T1_CMapStdRec_ CF2_Err_Invalid_Table cf2_hintmask_isNew darkenParams lastIsX cf2_hint_isTop t1_builder_close_contour cf2_escABS lastError cf2_escROLL CF2_Err_Invalid_Pixel_Size ps_builder_start_point cf2_stack_free blueScale glyphPath boldenY new_root hintMove cf2_escIFELSE CF2_Err_Ok maxZoneHeight t1_builder_check_points currentTransform cf2_hintmap_map cf2_cmdRESERVED_0 cf2_escRESERVED_19 CF2_StemHintRec_ ps_builder PSaux_Err_Nested_DEFS arg_cnt num_limit AFM_TOKEN_STARTKERNPAIRS CF2_Err_Invalid_Stream_Operation CF2_Err_Invalid_Reference downMinCounter cf2_outline_reset CF2_Err_Invalid_Vert_Metrics cf2_getNormalizedVector afm_parser_parse large_int CF2_Err_Too_Many_Caches nominalWidthX shift_elements cf2_escCALLOTHERSUBR cf2_getSeacComponent AFM_TOKEN_W1Y CF2_Err_Invalid_Offset CF2_BlueRec_ CF2_Err_ENDF_In_Exec_Stream AFM_TOKEN_ISCIDFONT unitsPerEm PSaux_Err_Unimplemented_Feature op_max darkened fracDown op_unknown15 cf2_hint_init CF2_Err_Lower_Module_Version cf2_stack_popFixed hinted nextP1 cf2_getGlyphOutline CF2_PairTop CF2_GhostBottom offsetStart1 t1_cmap_std_char_next tempHintMask PSaux_Err_Invalid_Frame_Operation totalSize CF2_Err_Ignore CF2_Err_Invalid_PPem familyOtherBlues CF2_Buffer AFM_TOKEN_WEIGHT cf2_blues_capture op_closepath component cff_builder_init cf2_escADD PSaux_Err_Hmtx_Table_Missing cf2_escDIV AFM_TOKEN_W t1_decoder_done PSaux_Err_Locations_Missing cf2_arrstack_clear stemWidth blueShift csCoord t1_cmap_unicode_char_next PSnames_Err_Invalid_CodeRange pscmaps_services NextIter PSnames_Err_Unknown_File_Format PSnames_Err_Unimplemented_Feature pscmaps_interface PSnames_Err_Too_Many_Extensions compare_uni_maps PSnames_Err_Invalid_PPem ft_adobe_glyph_list PSnames_Err_Syntax_Error PSnames_Err_Invalid_Post_Table ps_get_macintosh_name PSnames_Err_Missing_Bbx_Field PSnames_Err_Too_Many_Function_Defs t1_standard_encoding PSnames_Err_Name_Table_Missing PSnames_Err_Nested_DEFS PSnames_Err_Invalid_Slot_Handle PSnames_Err_Invalid_Cache_Handle PSnames_Err_Glyph_Too_Big PSnames_Err_Ignore PSnames_Err_Corrupted_Font_Glyphs PSnames_Err_Invalid_Composite ft_extra_glyph_names ft_sid_names ft_standard_glyph_names PSnames_Err_Missing_Chars_Field PSnames_Err_No_Unicode_Glyph_Name PSnames_Err_Corrupted_Font_Header PSnames_Err_Code_Overflow PSnames_Err_Invalid_Post_Table_Format PSnames_Err_Too_Many_Hints PSnames_Err_Bbx_Too_Big PSnames_Err_Cannot_Open_Resource PSnames_Err_Missing_Module map1 map2 ft_extra_glyph_unicodes PSnames_Err_Invalid_Version PSnames_Err_Invalid_Argument PSnames_Err_Invalid_Vert_Metrics PSnames_Err_Invalid_Frame_Read PSnames_Err_Invalid_Reference PSnames_Err_Missing_Encoding_Field PSnames_Err_Out_Of_Memory free_glyph_name PSnames_Err_Too_Many_Instruction_Defs /home/computerfido/Desktop/freetypetest2/freetype/src/psnames/psnames.c PSnames_Err_Invalid_Stream_Seek PSnames_Err_Raster_Negative_Height PSnames_Err_Post_Table_Missing ft_mac_names PSnames_Err_Missing_Startchar_Field PSnames_Err_Max PSnames_Err_Invalid_Offset PSnames_Err_Missing_Startfont_Field PSnames_Err_Ok PSnames_Err_Stack_Overflow NotFound PSnames_Err_Bad_Argument PSnames_Err_Invalid_Stream_Operation PSnames_Err_CMap_Table_Missing PSnames_Err_Unlisted_Object PSnames_Err_Invalid_Handle PSnames_Err_Invalid_File_Format PSnames_Err_Invalid_Library_Handle PSnames_Err_Nested_Frame_Access PSnames_Err_Invalid_Pixel_Size PSnames_Err_Missing_Bitmap PSnames_Err_Invalid_Opcode FT_Service_PsCMapsRec PSnames_Err_Invalid_Size_Handle unicode1 PSnames_Err_Raster_Corrupted PSnames_Err_Missing_Font_Field PSnames_Err_DEF_In_Glyf_Bytecode PSnames_Err_Invalid_Glyph_Index PSnames_Err_Invalid_Table PSnames_Err_Lower_Module_Version PSnames_Err_Invalid_CharMap_Handle ft_extra_glyph_name_offsets psnames_get_service ps_unicodes_char_index PSnames_Err_Divide_By_Zero ps_unicode_value PSnames_Err_Array_Too_Large PSnames_Err_Invalid_Glyph_Format PSnames_Err_Could_Not_Find_Context unicode2 PSnames_Err_Invalid_Horiz_Metrics PSnames_Err_Invalid_Character_Code PSnames_Err_Too_Many_Drivers base_glyph PSnames_Err_Invalid_Frame_Operation PSnames_Err_Cannot_Open_Stream PSnames_Err_Table_Missing PSnames_Err_Invalid_CharMap_Format PSnames_Err_Invalid_Face_Handle PSnames_Err_Missing_Fontboundingbox_Field ps_check_extra_glyph_unicode ft_get_adobe_glyph_index PSnames_Err_Horiz_Header_Missing extra_glyphs PSnames_Err_Invalid_Stream_Skip PSnames_Err_Stack_Underflow PSnames_Err_Execution_Too_Long PSnames_Err_Missing_Property PSnames_Err_Invalid_Stream_Read PSnames_Err_Missing_Size_Field PSnames_Err_Hmtx_Table_Missing PSnames_Err_Locations_Missing PSnames_Err_Invalid_Stream_Handle ps_unicodes_char_next uni_char PSnames_Err_Raster_Overflow PSnames_Err_Too_Few_Arguments ps_unicodes_init ps_get_standard_strings PSnames_Err_Debug_OpCode extra_glyph_list_states PSnames_Err_Cannot_Render_Glyph t1_expert_encoding PSnames_Err_Too_Many_Caches PSnames_Err_Invalid_Outline PSnames_Err_ENDF_In_Exec_Stream PSnames_Err_Invalid_Driver_Handle PSnames_Err_Raster_Uninitialized ps_check_extra_glyph_name malloc /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftsystem.c ft_ansi_stream_close fseek ft_realloc fopen ft_alloc fread fclose ft_free ftell ft_ansi_stream_io ft_bitmap_assure_buffer target_pitch_sign xstr bit_last xStrength /home/computerfido/Desktop/freetypetest2/freetype/src/base/ftbitmap.c yStrength target_size FT_Bitmap_Copy FT_Bitmap_Embolden source_pitch_sign null_bitmap ft_gray_for_premultiplied_srgb_bgra FT_GlyphSlot_Own_Bitmap FT_Bitmap_New new_pitch ypixels xpixels old_target_pitch ystr /home/computerfido/Desktop/Lemon/LibC/build syscall arg0 arg4 ../sysdeps/lemon/generic/syscall.c GNU C17 8.2.0 -mtune=generic -march=x86-64 -g -fno-builtin -fPIC arg3 _ZNK3frg8optionalIiE9has_valueEv _millis sys_anon_allocate stack_buffer_logger<mlibc::InfoSink, 128> _ZN3frg8optionalIiEC2Ev sys_exit _ZN5mlibc14sys_libc_panicEv message _ZNSt17integral_constantIbLb0EE5valueE format_integer<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg14format_optionsC2ERKS0_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4EPS3_ _ZSt18is_constructible_vIiJON3frg8optionalIiEEEE _fmt_basics alt_conversion wchar_t _ZN3frg14format_options15with_conversionENS_17format_conversionE print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> assertion absv _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD4Ev null_opt_type _ZNKSt17integral_constantIbLb0EEcvbEv _sink _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC4ERKS4_ _ZN3frg8optionalIiEptEv operator() endlog operator std::integral_constant<bool, true>::value_type _ZN3frg8optionalIiE13storage_unionD4Ev _ZNSt17integral_constantIbLb1EE5valueE has_value sys_anon_free _ZNSt16is_constructibleIiJON3frg8optionalIiEEEE5valueE ~storage_union _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc _ZN3frg14format_optionsC4ERKS0_ append format<char const*, frg::stack_buffer_logger<mlibc::PanicSink>::item> format_conversion _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic long long unsigned int _ZN3frg8optionalIiEcvbEv ~item _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc _ZN5mlibc17sys_anon_allocateEmPPv _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemaSERKS4_ __cxa_atexit _ZN5mlibc8sys_exitEi _ZN5mlibc12sys_libc_logEPKc _ZN3frg8optionalIiE13storage_unionD2Ev format_object<frg::stack_buffer_logger<mlibc::PanicSink>::item> _ZN3frg8optionalIiEdeEv _Z19__frigg_assert_failPKcS0_jS0_ _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc9PanicSinkclEPKc _ZNKSt17integral_constantIbLb1EEclEv _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ operator std::integral_constant<bool, false>::value_type _emit _emitted _ZN5mlibc10sys_getpidEv with_conversion _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ clock operator<< <char const*> _ZN3frg8optionalIiED4Ev minimum_width sys_clock_get _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZNSt16is_constructibleIiJRKN3frg8optionalIiEEEE5valueE _ZN3frg14format_optionsD4Ev mlibc PanicSink time_t GNU C++17 8.2.0 -mtune=generic -march=x86-64 -g -std=c++17 -fno-builtin -fno-rtti -fno-exceptions -fPIC sys_getpid _ZN3frg8optionalIiEC4EOi _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEC4ES2_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv pid_t _ZN3frg14format_optionsD2Ev operator-> _ZNKSt17integral_constantIbLb1EEcvbEv operator* _pid _ZN3frg8optionalIiEC4ENS_13null_opt_typeE operator= _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ sys_libc_panic _ZN5mlibc11panicLoggerE format<unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> operator<< <unsigned int> endlog_t optional<int> _ZN3frg8optionalIiEC2ERKS1_ _stor _ZN5mlibc13sys_anon_freeEPvm _ZN5mlibc9PanicSinkC4Ev nanos _ZSt18is_constructible_vIiJRKN3frg8optionalIiEEEE small_digits _ZN3frg8optionalIiE13storage_unionC4Ev _ZN3frg8optionalIiED2Ev operator new operator<< sys_libc_log null_opt _ZN3frg8optionalIiEC4EOS1_ _ZNK3frg8optionalIiEcvbEv panicLogger _non_null plus_becomes_space _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE negative stack_buffer_logger ~format_options is_constructible<int, frg::optional<int>&&> _ZN3frg8optionalIiEC4ERKS1_ _ZN3frg8optionalIiE6_resetEv ~optional _ZN3frg14format_optionsC4Ev is_constructible<int, const frg::optional<int>&> radix operator bool max<int> _ZNKSt17integral_constantIbLb0EEclEv integral_constant<bool, false> stack_buffer_logger<mlibc::PanicSink, 128> left_justify _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev _to_string_impl _Z19__mlibc_do_finalizev _ZN3frg8optionalIiE13storage_unionC2Ev _ZN3frg8optionalIiEC4Ev function _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ fill_zeros _secs always_sign is_constructible_v print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, unsigned int> _ZnwmPv _ZN5mlibc13sys_clock_getEiPlS0_ _ZN5mlibc10infoLoggerE _ZN3frg8optionalIiEC4ERKi ../sysdeps/lemon/generic/lemon.cpp integral_constant<bool, true> __func__ _ZN3frg14format_optionsC2Ev _ZN3frg3maxIiEERKT_S3_S3_ __mlibc_do_finalize _ZNK3frg8optionalIiEdeEv _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic __frigg_assert_fail infoLogger _ZN3frg8optionalIiEaSES1_ InfoSink _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv _ZN5mlibc8InfoSinkC4Ev _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEC4ES2_ ../options/internal/generic/debug.cpp _ZN5mlibc8InfoSinkclEPKc format_integer<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> format<char const*, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4ERKS4_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic format<unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC4EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ ../options/internal/generic/ensure.cpp _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc __ensure_warn _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> format_object<frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD4Ev _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ __ensure_fail _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemaSERKS4_ print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, unsigned int> src_bytes ../options/internal/generic/essential.cpp dest_bytes ../options/internal/x86_64/setjmp.S GNU AS 2.32 mb_chr _ZN3frg11unique_lockI13AllocatorLockEC4EOS2_ size_to_bucket _ZN3frg7mt19937C2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC4Ev _ZN3frg11unique_lockI13AllocatorLockEC4ENS_11dont_lock_tERS1_ replacement _ZN3frg7mt199371nE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ mag01 _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ code_seq<char const> wseq mbstowcs lldiv _tree_mutex strtold _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ strtoll print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> lsbs get_root dont_lock_t __mlibc_rand_engine _is_locked _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg10bitop_implImE3clzEm _ZN5mlibc8code_seqIwEcvbEv operator<< <void*> _verify_integrity _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameaSERKS4_ _ZN3frg11unique_lockI13AllocatorLockED2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC4ERKS4_ tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE12huge_paddingE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14small_base_expE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ atof rotateRight _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ locale_t __cpoint _ZN5mlibc7strtofpIeEET_PKcPPc _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE12numUsedPagesEv endptr _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC4EPNS_9slab_poolIS1_S2_EE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11_find_frameEm _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ aggregate_node _usedPages atoi illegal_input address_ frame_hook _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC4ERS1_ wctomb _ZN3frg7mt199378matrix_aE insert_right left_ptr _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE23test_bucket_calculationEj _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ area_size _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ _ZN13AllocatorLock4lockEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ _ZN5mlibc7strtofpIfEET_PKcPPc type_ abort _ZN13AllocatorLockC4ERKS_ partial_hook slab_allocator tiny_sizes _ZN3frg11unique_lockI13AllocatorLockE9is_lockedEv num_buckets slabsize _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ 7lldiv_t pool_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameaSERKS4_ num_reserved insert_root rbtree successor huge_padding _ZN3frg9_redblack11hook_structC4ERKS1_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ bucket_mutex isRed _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ fix_insert _ZN3frg9_redblack11hook_structC4Ev llabs color_type mblen_state 5div_t _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ VirtualAllocator was_unavailable tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::_redblack::null_aggregator> deallocate predecessor mblen _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EaSERKSB_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE23_verify_frame_integrityEPNS3_5frameE _ZN3frg11unique_lockI13AllocatorLockE8protectsEPS1_ print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, long unsigned int> _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEaSERKS3_ check_invariant _frame_tree succ _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE9page_sizeE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14size_to_bucketEm replace_node _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EaSERKSB_ rand_r _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ Member frame_type AllocatorLock _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ strtoul cutlim atoll aggregate<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame> dot_end _ZN3frg11unique_lockI13AllocatorLockEaSES2_ strtofp<double> _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC4ES7_ grand frame_less format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _construct_large 6ldiv_t _Exit output_overflow _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ code_seq<wchar_t> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ get_right _ZN16VirtualAllocator3mapEm _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj frame_tree_type slab_frame length_ remove_half_leaf reallocate format<void*, frg::stack_buffer_logger<mlibc::InfoSink>::item> numUsedPages tree_crtp_struct<frg::_redblack::tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator>, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::frame::frame_hook, frg::_redblack::null_aggregator> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15max_bucket_sizeE _ZN3frg11unique_lockI13AllocatorLockE6unlockEv _ZN3frg11unique_lockI13AllocatorLockED4Ev _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg11unique_lockI13AllocatorLockEC4ERS1_ Mutex _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ _plcy _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm freelist child _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ _verify_frame_integrity bsearch _ZN3frg7mt19937C4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv slab_allocator<VirtualAllocator, AllocatorLock> _redblack _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE16_construct_largeEm mb_string input_underflow _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ wcstombs isBlack _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEv small_step_exp _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E15check_invariantEPS7_RiRSC_SE_ _ZN3frg11unique_lockI13AllocatorLockEC4ERKS2_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frame8containsEPv tree_crtp_struct _ZN3frg7mt199374lsbsE protects _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC4Emmi _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC2Ev _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10reallocateEPvm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ partial_tree _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14small_step_expE strtoull _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11num_bucketsE _ZN16VirtualAllocator5unmapEmm overhead _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE7reallocEPvm _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistaSERKS4_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ _ZN3frg3maxImEERKT_S3_S3_ enable_checking _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ _ZN13AllocatorLockaSERKS_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE17_verify_integrityEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ get_parent _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv _ZN3frg7mt199373msbE _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8slabsizeE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ max<long unsigned int> hook_struct head_slb _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8allocateEm strtofp<float> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5firstEv mb_limit mbtowc get_left rotateLeft null_aggregator _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15_construct_slabEi _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ quot parent_color _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4ERKSB_ u_bytes _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm wc_limit ULONG_MAX _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC4ERKS3_ _ZN3frg7mt199374seedEj slab_pool _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv _bkts new_pointer mktemp _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC4ERKSB_ bucket_guard unique_lock<AllocatorLock> matrix_a rbtree_hook at_quick_exit _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ small_base_exp aligned_alloc v_bytes index_ strtod strtof _GLOBAL__sub_I_stdlib_stubs.cpp right_ptr _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC4Ev tree_guard _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E15check_invariantEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC4ERKS4_ charcode_error Policy max_bucket_size aggregate_path _ZN3frg9_redblack11hook_structaSERKS1_ __progress strtofp<long double> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10tiny_sizesE unlock _ctr test_bucket_calculation srand partial_tree_type _ZN13AllocatorLockC4Ev tree_struct _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ _ZN3frg9_redblack11hook_structC2Ev ../options/ansi/generic/stdlib-stubs.cpp cutoff strtod_l ~unique_lock _find_frame bucket_to_size tree_struct<frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame, &frg::slab_pool<VirtualAllocator, AllocatorLock>::slab_frame::partial_hook, frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less, frg::_redblack::null_aggregator> aggregate<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame> _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _futex _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ contains insert_left page_size _ZN5mlibc7strtofpIdEET_PKcPPc _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC4ENS3_10frame_typeEmm __shift mt19937 _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE4freeEPv _ZN5mlibc8code_seqIKcEcvbEv _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ slab_pool<VirtualAllocator, AllocatorLock> wc_string dont_lock _construct_slab dirty _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10deallocateEPvm denom posix_memalign bitop_impl<long unsigned int> pred _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC4Ev _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN13AllocatorLock6unlockEv fix_remove _ZN3frg11unique_lockI13AllocatorLockEC4Ev _ZN3frg7mt199371mE _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN3frg7mt19937clEv srandom _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC4ERKS4_ _ZN5mlibc8code_seqIjEcvbEv iswlower iscntrl isalnum _ZN3frg17basic_string_viewIcE10find_firstEcm _ZNK3frg17basic_string_viewIcE4sizeEv isprint isdigit isspace ct_digit _ZN3frg17basic_string_viewIcEC2EPKc ct_space iswspace ispunct _ZN5mlibc13wide_charcode7promoteEwRj _ZNK3frg17basic_string_viewIcEneES1_ isupper ct_punct iswcntrl toupper generic_is_control iswdigit iswpunct isgraph iswprint ct_graph isalpha basic_string_view towupper ct_alpha _ZN5mlibc18generic_is_controlEj _ZNK3frg17basic_string_viewIcEixEm iswxdigit _ZN3frg17basic_string_viewIcEC4EPKc basic_string_view<char> _ZN3frg17basic_string_viewIcEC4EPKcm ct_alnum isblank sub_string ct_blank codepoint _ZNK3frg17basic_string_viewIcEeqES1_ ct_cntrl iswblank find_first ct_upper iswalpha find_last iswctype _ZN3frg17basic_string_viewIcEC4Ev iswupper tolower operator== ct_print operator!= ct_xdigit wint_t towlower isascii _ZN5mlibc20polymorphic_charcode7promoteEcRj promote _ZNK3frg17basic_string_viewIcE4dataEv iswgraph ct_count isxdigit ct_null _ZN3frg17basic_string_viewIcE9find_lastEc iswalnum islower code_seq<unsigned int> _ZN3frg17basic_string_viewIcE10sub_stringEmm wctype_t ct_lower ../options/ansi/generic/ctype-stubs.cpp unsetenv self _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ _ZN3frg10escape_fmtC4EPKvm update_vector _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED4Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEaSES6_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ES5_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv new_capacity push_back get_vector _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm move<char*&> remove_reference<char*&> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4EOS6_ ../options/ansi/generic/environment.cpp _ZSt4swapIPcEvRT_S2_ unassign_variable operator<< <frg::escape_fmt> remove_reference<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv escape_fmt _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ remove_reference_t _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv ~vector _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backEOS1_ _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ empty_environment overwrite _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ES5_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE9push_backERKS1_ _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEENSt16remove_referenceIT_E4typeEOS7_ _ensure_capacity format<frg::escape_fmt, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4ERKS6_ move<frg::slab_allocator<VirtualAllocator, AllocatorLock>&> vector<char*, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv putenv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv swap<char*> _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3endEv _ZN3frg10escape_fmtC2EPKvm new_array _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5beginEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5frontEv start_from _ZN3frg17basic_string_viewIcEC2EPKcm find_environ_index _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5emptyEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ ../options/ansi/generic/errno-stubs.cpp _ZN5mlibc13abstract_file5closeEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE4backEv default_list_hook _ZN5mlibc13abstract_file9_save_posEv _ZN5mlibc13abstract_file7io_readEPcmPm _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ _vptr.abstract_file format_integer<int, frg::stack_buffer_logger<mlibc::InfoSink>::item> intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*> _init_bufmode _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC4Ev _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ __vtbl_ptr_type _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> pipe_like whence erased remove_reference<int&> stdout_file forward<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > ssize_t rewind _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ ~fd_file fileno _write_back destruct<mlibc::abstract_file, frg::slab_allocator<VirtualAllocator, AllocatorLock> > _ZN5mlibc7fd_fileD2Ev _ZN3frg3minImEERKT_S3_S3_ _ZN5mlibc13abstract_file14determine_typeEPNS_11stream_typeE _ZN5mlibc13abstract_file6_resetEv composition<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > ~<lambda> _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8pop_backEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN5mlibc13abstract_file8io_writeEPKcmPm _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ _save_pos _init_type _ZN5mlibc13abstract_file10_init_typeEv _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ fileno_unlocked unknown _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN5mlibc13abstract_file13_init_bufmodeEv abstract _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5emptyEv OwnerPointer _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE _void_impl determine_bufmode intrusive_traits<mlibc::abstract_file, mlibc::abstract_file*, mlibc::abstract_file*> _ZN5mlibc13abstract_fileC4EPFvPS0_E __closure stream_type format<char, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN5mlibc13abstract_file7disposeEv fdopen _ZN3frg6formatIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN5mlibc13abstract_fileD4Ev file_like update_bufmode _ZN5mlibc7fd_fileC4EiPFvPNS_13abstract_fileEE _ZN5mlibc13abstract_file4seekEli _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ setvbuf io_read _GLOBAL__sub_I_file_io.cpp _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic new_offset line_buffer io_size operator<< <int> intrusive_list Locate _ZN5mlibc13abstract_fileaSERKS0_ _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE10push_frontES6_ unget _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ __for_range _ensure_allocation print_digits<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> has_plus _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _ZN5mlibc13abstract_file5purgeEv _ZN5mlibc13abstract_file5ungetEc _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _current _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6spliceENS9_8iteratorERS9_ _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE _ZN5mlibc13abstract_file18_ensure_allocationEv io_write format<int, frg::stack_buffer_logger<mlibc::InfoSink>::item> _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE _ZN5mlibc7fd_file2fdEv _ZN5mlibc13abstract_fileD0Ev _ZN5mlibc7fd_fileD4Ev print_int<frg::stack_buffer_logger<mlibc::InfoSink>::item, int> borrow_pointer _ZN5mlibc7fd_file5closeEv _ZN5mlibc13abstract_file7io_seekEliPl push_front BorrowPointer _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEi _ZN5mlibc13abstract_fileC4ERKS0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv forward<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > _ZN5mlibc7fd_fileC4ERKS0_ __for_begin _ZN5mlibc13abstract_file11_write_backEv off_t _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev previous __fpurge _ZN5mlibc13abstract_file4readEPcmPm current_offset ~abstract_file globallyDisableBuffering global_file_list _ZN5mlibc13abstract_file5flushEv _ZN5mlibc13abstract_fileC2EPFvPS0_E intrusive_list_hook _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ min<long unsigned int> stderr_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC4ES6_ io_seek _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIiEERS4_T_ actual_size __for_end _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE full_buffer _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv _ZN5mlibc7fd_fileD0Ev <lambda(mlibc::abstract_file*)> remove_reference<fopen(char const*, char const*)::<lambda(mlibc::abstract_file*)> > _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE6insertENS9_8iteratorES6_ operator void (*)(mlibc::abstract_file*) move<mlibc::abstract_file*&> args#1 _result_of_impl splice owner_pointer determine_type locate_tag remove_reference<fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > args#0 _ZN5mlibc13abstract_file5writeEPKcmPm decay _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5frontEv pop_front _ZN5mlibc7fd_file7io_seekEliPl operator<< <char> remove_reference<mlibc::abstract_file*&> operator++ borrow _ZN5mlibc7fd_fileC4EOS0_ buffer_mode _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ _do_dispose pop_back _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC4Ev remove_reference<frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>&> intrusive_list<mlibc::abstract_file, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > ungetc erase no_buffer flush_line get<frg::_list::locate_tag, frg::locate_member<mlibc::abstract_file, frg::_list::intrusive_list_hook<mlibc::abstract_file*, mlibc::abstract_file*>, &mlibc::abstract_file::_list_hook> > construct<mlibc::fd_file, frg::slab_allocator<VirtualAllocator, AllocatorLock>, int&, fdopen(int, char const*)::<lambda(mlibc::abstract_file*)> > seek_offset global_stdio_guard ../options/ansi/generic/file-io.cpp _ZN5mlibc7fd_file7io_readEPcmPm _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic in_list ~stdio_guard _ZN5mlibc13abstract_file4tellEPl stdin_file _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ _ZN5mlibc13abstract_fileD2Ev _ZN5mlibc13abstract_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc7fd_file8io_writeEPKcmPm iterator_to forward<int&> _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE fflush _FUN fflush_unlocked _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9pop_frontEv print_int<StreamPrinter, long int> _ZN3frg17basic_string_viewIwE9find_lastEw do_printf_ints<StreamPrinter> fgetc printf_format<PrintfAgent<StreamPrinter> > print_int<StreamPrinter, long unsigned int> fgets _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev vfprintf _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN11PrintfAgentI14LimitedPrinterEclEc _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_digits<BufferPrinter, long int> vswscanf fread_unlocked print_digits<ResizePrinter, long unsigned int> _ZN13ResizePrinter6expandEv BufferPrinter renameat fputws _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev vasprintf _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _vsp putchar __mlibc_intmax print_digits<BufferPrinter, long long unsigned int> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev is_constructible<int, int&&> print_int<ResizePrinter, long long unsigned int> fgetpos _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ clearerr _ZN13ResizePrinterC4Ev _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic SCANF_TYPE_INT print_int<ResizePrinter, long int> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ fputs_unlocked _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic ftrylockfile SCANF_TYPE_SIZE_T vfscanf _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN13StreamPrinter6appendEPKc print_digits<BufferPrinter, long unsigned int> do_scanf<sscanf(char const*, char const*, ...)::<unnamed class> > swap<int> _ZN3frg4swapERNS_8optionalIiEES2_ _ZNK3frg17basic_string_viewIwEneES1_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ print_digits<LimitedPrinter, long int> bytes_read feof_unlocked print_int<BufferPrinter, unsigned int> default_size print_int<ResizePrinter, long unsigned int> _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ vscanf _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN3frg17basic_string_viewIwEC2EPKw PrintfAgent _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ filename <lambda(auto:1)> fgetwc getwchar _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ print_int<LimitedPrinter, long int> fgetws vwprintf _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ do_printf_chars<LimitedPrinter> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE native_size _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ __builtin_va_list do_scanf<vfscanf(FILE*, char const*, __va_list_tag*)::<unnamed struct> > _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ do_printf_floats<LimitedPrinter> __gnuc_va_list handler _ZNK3frg17basic_string_viewIwE4sizeEv clearerr_unlocked _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZN11PrintfAgentI13StreamPrinterEC4EPS0_PN3frg9va_structE move<bool&> _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic print_int<BufferPrinter, long unsigned int> fwrite_unlocked _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE print_digits<StreamPrinter, long unsigned int> do_printf_chars<BufferPrinter> _ZN13BufferPrinterC2EPc _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic ungetwc fp_offset new_limit _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg8optionalIiEC4IRivEEOT_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ vsnprintf _ZN11PrintfAgentI13BufferPrinterEclEc new_path _ZSt4swapIiEvRT_S1_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ new_buffer vswprintf szmod _ZNK3frg17basic_string_viewIwEixEm print_int<LimitedPrinter, long unsigned int> fwide _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic _ZN14LimitedPrinter6appendEPKcm funlockfile _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _ZSt18is_constructible_vIiJRiEE putchar_unlocked _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic print_int<StreamPrinter, unsigned int> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE putwchar print_int<ResizePrinter, unsigned int> _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ SCANF_TYPE_PTRDIFF _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN3frg17basic_string_viewIwE10find_firstEwm print_digits<StreamPrinter, long int> rename _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ print_digits<ResizePrinter, long int> <lambda(auto:2)> do_printf_ints<BufferPrinter> print_digits<LimitedPrinter, long long unsigned int> _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ ferror vfwprintf _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic print_int<StreamPrinter, long long unsigned int> unused _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ _ZN13ResizePrinter6appendEc _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic _ZNSt16is_constructibleIiJOiEE5valueE _ZN3frg17basic_string_viewIwEC4Ev _ZN11PrintfAgentI13ResizePrinterEC4EPS0_PN3frg9va_structE _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE PrintfAgent<ResizePrinter> _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic printf_size_mod second printf_format<PrintfAgent<BufferPrinter> > StreamPrinter _ZN3frg8optionalIiEC2EOi PrintfAgent<StreamPrinter> _ZN13StreamPrinter6appendEPKcm _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN11PrintfAgentI13BufferPrinterEC4EPS0_PN3frg9va_structE SCANF_TYPE_SHORT _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN11PrintfAgentI13ResizePrinterEclEc gp_offset _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE vprintf _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN11PrintfAgentI13BufferPrinterEclEPKcm perror move<int&> consume fputc_unlocked _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev _ZN14LimitedPrinter6appendEc _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4ERKS8_ _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN11PrintfAgentI13StreamPrinterEclEc _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE agent optional<int&> _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN13ResizePrinter6appendEPKcm overflow_arg_area _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev operator()<long unsigned int> fsetpos _ZN14LimitedPrinter6appendEPKc _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZN13BufferPrinterC4EPc <lambda(auto:3)> SCANF_TYPE_LL setbuf feof _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE print_int<BufferPrinter, long int> intmax_t LimitedPrinter expand __opts _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic olddirfd _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg8optionalIiEC2IRivEEOT_ swap<bool> va_struct _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE fgets_unlocked num_consumed _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13ResizePrinterEclEPKcm _ZN3frg17basic_string_viewIwEC4EPKwm reg_save_area getdelim _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN14LimitedPrinterC2EPcm _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN13StreamPrinter6appendEc _ZN11PrintfAgentI14LimitedPrinterEC4EPS0_PN3frg9va_structE _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev getchar_unlocked print_int<LimitedPrinter, unsigned int> old_path print_digits<BufferPrinter, unsigned int> _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic match_count ~<constructor> _ZNSt16is_constructibleIiJRiEE5valueE print_int<BufferPrinter, long long unsigned int> _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic __formatter _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev longlong_size _ZN14LimitedPrinterC4EPcm remove_reference<bool&> vsscanf do_printf_ints<ResizePrinter> ../options/ansi/generic/stdio-stubs.cpp SCANF_TYPE_CHAR _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ fputs vwscanf _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev getline _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev _ZN13BufferPrinter6appendEPKc _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZSt4swapIbEvRT_S1_ do_printf_ints<LimitedPrinter> _ZNK3frg17basic_string_viewIwEeqES1_ _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4Ev _ZN3frg17basic_string_viewIwE10sub_stringEmm print_int<LimitedPrinter, long long unsigned int> _ZNK3frg17basic_string_viewIwE4dataEv freopen print_digits<StreamPrinter, long long unsigned int> _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ print_digits<ResizePrinter, long long unsigned int> tmpnam _ZN13ResizePrinter6appendEPKc SCANF_TYPE_INTMAX scanset newdirfd look_ahead tmpfile print_digits<StreamPrinter, unsigned int> auto:2 auto:3 _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN13BufferPrinter6appendEc ferror_unlocked print_digits<ResizePrinter, unsigned int> SCANF_TYPE_L _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4EOS8_ do_printf_floats<StreamPrinter> fputc auto:1 do_printf_chars<StreamPrinter> print_digits<LimitedPrinter, long unsigned int> _ZN13BufferPrinter6appendEPKcm _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE fpos_t _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4ERKS8_ PrintfAgent<LimitedPrinter> fgetc_unlocked _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4Ev basic_string_view<wchar_t> _ZN3frg17basic_string_viewIwEC4EPKw fputwc _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_D4Ev typed_dest store_int is_constructible<int, int&> PrintfAgent<BufferPrinter> _ZN13StreamPrinterC2EP17__mlibc_file_base vfwscanf _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ printf_format<PrintfAgent<ResizePrinter> > _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_C4ERKS8_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_D4Ev _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E_D4Ev vsprintf do_printf_floats<BufferPrinter> _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4Ev ResizePrinter _ZN13StreamPrinterC4EP17__mlibc_file_base _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E0_C4EOS8_ flockfile do_printf_floats<ResizePrinter> do_printf_chars<ResizePrinter> printf_format<PrintfAgent<LimitedPrinter> > _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZSt18is_constructible_vIiJOiEE operator()<unsigned int> _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENUlS2_E1_C4EOS8_ typedef __va_list_tag __va_list_tag fwrite print_digits<LimitedPrinter, unsigned int> getchar _ZN13ResizePrinterC2Ev wcsrchr strchrnul pattern wmemmove wmemcmp wcsncat bufsz wmemset wcstod wcscpy wcstof wcsncpy stpcpy wcstok wcstold wcstoull wcstol chrs wcstoll strerror ../options/ansi/generic/string-stubs.cpp delimiter strtok_r wcspbrk wcschr mempcpy wcsncmp wcsstr b_byte strtok wcscspn wcscat wcslen s_bytes strchr strncat strcspn wcstoul wcscmp strerror_r strcoll a_byte strxfrm wmemchr strspn wcscoll wcsspn saved wcsxfrm wmemcpy strpbrk sys_access sys_close written sys_read _ZN5mlibc8sys_openEPKciPi _ZN5mlibc10sys_accessEPKci ../sysdeps/lemon/generic/filesystem.cpp sys_write sys_open _ZN5mlibc8sys_seekEiliPl sys_errno _ZN5mlibc9sys_writeEiPKvmPl _ZN5mlibc9sys_closeEi sys_seek _ZN5mlibc8sys_readEiPvmPl _ZN3frg15aligned_storageILm456ELm8EEC2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC2ERS1_ remove_reference<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less&> _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC4IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _ZN3frg15aligned_storageILm1ELm1EEC2Ev heap Align _ZN3frg7eternalI16VirtualAllocatorE3getEv aligned_storage<8, 8> aligned_storage eternal<> _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC4IJRS2_EEEDpOT_ eternal<VirtualAllocator&> _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEE3getEv move<frg::slab_pool<VirtualAllocator, AllocatorLock>::frame_less&> remove_reference<frg::slab_pool<VirtualAllocator, AllocatorLock>*> _ZSt7forwardIPN3frg9slab_poolI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ eternal<frg::slab_allocator<VirtualAllocator, AllocatorLock> > MemoryAllocator getAllocator _ZSt4moveIRN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ _ZN3frg15aligned_storageILm8ELm8EEC4Ev forward<VirtualAllocator&> aligned_storage<456, 8> _ZN3frg7eternalI16VirtualAllocatorEC4IJEEEDpOT_ eternal<frg::slab_pool<VirtualAllocator, AllocatorLock>*> eternal<VirtualAllocator> virtualAllocator forward<frg::slab_pool<VirtualAllocator, AllocatorLock>*> _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2EPNS_9slab_poolIS1_S2_EE _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv _Z12getAllocatorv eternal<frg::slab_pool<VirtualAllocator, AllocatorLock> > _ZN3frg15aligned_storageILm8ELm8EEC2Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE aligned_storage<1, 1> _ZN3frg15aligned_storageILm456ELm8EEC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev _ZN13AllocatorLockC2Ev _ZN3frg15aligned_storageILm1ELm1EEC4Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC2Ev singleton ../options/internal/generic/allocator.cpp remove_reference<VirtualAllocator&> global_wide_charcode code_seq<unsigned int const> _ZN5mlibc16current_charcodeEv _ZN5mlibc8code_seqIKwEcvbEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate promote_wtranscode has_shift_states_ _ZN5mlibc20polymorphic_charcodeC2Ebb platform_wide_charcode _ZN5mlibc20polymorphic_charcodeD4Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED4Ev preserves_7bit_units _ZN5mlibc20polymorphic_charcodeC4ERKS0_ decode_wtranscode utf8_charcode code_seq<char> _ZN5mlibc13utf8_charcode16has_shift_statesE _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4Ev decode_wtranscode_length _ZN5mlibc20polymorphic_charcode17decode_wtranscodeERNS_8code_seqIKcEERNS1_IwEER15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode6decodeERNS_8code_seqIKcEERNS1_IjEER15__mlibc_mbstate _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4ERKS2_ auto has_shift_states _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE encode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate polymorphic_charcode_adapter<mlibc::utf8_charcode> _ZN5mlibc13utf8_charcode20preserves_7bit_unitsE code_seq<wchar_t const> _ZN5mlibc8code_seqIcEcvbEv _ZN5mlibc13utf8_charcode12decode_stateC4Ev global_charcode _ZN5mlibc20polymorphic_charcodeD2Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE ../options/internal/generic/charcode.cpp decode_nseq _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _vptr.polymorphic_charcode current_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN5mlibc20polymorphic_charcode24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc20polymorphic_charcode17encode_wtranscodeERNS_8code_seqIcEERNS1_IKwEER15__mlibc_mbstate ~polymorphic_charcode _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13utf8_charcode12decode_state6cpointEv encode_wtranscode _ZN5mlibc13utf8_charcode12decode_stateC2Ev _ZN5mlibc13utf8_charcode12decode_state8progressEv preserves_7bit_units_ ~polymorphic_charcode_adapter _ZN5mlibc8code_seqIKjEcvbEv _ZN5mlibc22platform_wide_charcodeEv _ZN5mlibc20polymorphic_charcodeC4Ebb _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC4EOS2_ _ZN5mlibc20polymorphic_charcodeD0Ev _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev encode_state _ZN5mlibc20polymorphic_charcode18promote_wtranscodeEcRw decode_state _ZN5mlibc7charset8is_blankEj is_graph _ZN5mlibc7charset8is_alphaEj is_alpha _ZN5mlibc7charset8is_spaceEj is_alnum is_blank _ZN5mlibc7charset8is_printEj is_upper _ZN5mlibc7charset8is_lowerEj _ZN5mlibc7charset8is_upperEj _ZN5mlibc15current_charsetEv _ZN5mlibc7charset8is_graphEj _ZN5mlibc7charset9is_xdigitEj ../options/internal/generic/charset.cpp is_lower _ZN5mlibc7charset8to_lowerEj _ZN5mlibc7charset8is_alnumEj to_lower _ZN5mlibc7charset8to_upperEj _ZN5mlibc7charset17is_ascii_supersetEv _ZN5mlibc7charset8is_digitEj global_charset is_ascii_superset is_punct _ZN5mlibc7charset8is_punctEj is_print is_xdigit current_charset to_upper Guard _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic __mlibc_int64 ../options/internal/gcc/guard-abi.cpp _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ complete _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ print_int<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> print_digits<frg::stack_buffer_logger<mlibc::PanicSink>::item, long unsigned int> _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ __cxa_guard_acquire __cxa_guard_release format<void*, frg::stack_buffer_logger<mlibc::PanicSink>::item> format_integer<long unsigned int, frg::stack_buffer_logger<mlibc::PanicSink>::item> __cxa_pure_virtual _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_       �      �       U�      �       �U��      �       U                  �      �       S                          �      �       U�      H       \H      K       �U�K      q       \q      t       �U�                                     P      J       ]J      W       PW      Z       ]                        �             P             SK      Z       SZ      n       P                        4       V                                 
 �-H     �      '       S'      ,       sx�,      4       S                        @       J        UJ       �       S�      �       �U��      �       S                  V       j        P                                  _       �        P�       �        T�       /       R/      �       V�      �       P�      �       P�      �       T�      �       R�      �       V                        �       (       T(      }       R�      �       T�      �       R                                    �       �        Q�       �        U�       �        Q�       �        0��       �        P�       �        U      
       P(      /       0�/      @       P@      D       TW      \       P                                      U       2        V2       3        �U�                                    
 �-H     �               S       $        sx�$       1        S                      ��      ��       U��      ׯ       �U�ׯ      �       U                            ��      ��       T��      ǯ       Vǯ      ʯ       �T�ʯ      ԯ       Vԯ      ׯ       �T�ׯ      �       T                            ��      ��       Q��      ɯ       \ɯ      ʯ       �Q�ʯ      ֯       \֯      ׯ       �Q�ׯ      �       Q                        ��      ��       U��      ��       S��      ��       Uʯ      ׯ       U                     ��      ��       0���      ʯ       Pʯ      �       0�                    ��      ��       S��      Ư       S                    �      �       P�      �       P                      @�      c�       Uc�      g�       u�g�      ��       U                    @�      g�       Tg�      ��       T                    @�      R�       QR�      {�       �Q�                         �      �       U�      +�       V+�      1�       U1�      2�       �U�                         �      �       T�      *�       S*�      1�       T1�      2�       �T�                         �      �       Q�      -�       \-�      1�       R1�      2�       �Q�                   �      1�       Q                        ��      ��       U��      Ѭ       �U�Ѭ      �       U�      ��       �U�                          ��      ��       T��      ̬       V̬      Ѭ       �T�Ѭ      �       T�      ��       V                          ��      ��       Q��      ˬ       Sˬ      Ѭ       �Q�Ѭ      �       Q�      ��       S                          ��      ��       R��      ά       \ά      Ѭ       �R�Ѭ      �       R�      ��       \                 ��      ��       �&�                            ��      ��       Q��      ˬ       Sˬ      Ѭ       �Q�Ѭ      �       Q�      ��       S                       ��      ��       U��      Ѭ       �U�Ѭ      �       U�      ��       �U�                       ��      ��       0���      ��       PѬ      �       0��      ��       P                                  ��      ��       U��      ��       Z��      ł       �U�ł      �       Z�      �       �U��      ,�       Z,�      @�       �U�@�      V�       ZV�      u�       �U�                                ��      ��       T��      ł       �T�ł      ��       T��      �       �T��      &�       T&�      @�       �T�@�      D�       TD�      u�       �T�                                  ��      ��       Q��      ��       U��      ł       �Q�ł      ��       U��      �       �Q��      )�       U)�      @�       �Q�@�      O�       UO�      u�       �Q�                            ��      ��       R��      ł       �R�ł      �       R�      �       �R��      ,�       R,�      u�       �R�                                    ��      ��       X��      �       X�      �       �X��      �       P�      ,�       X,�      4�       �X�4�      ?�       S?�      @�       P@�      V�       XV�      u�       w                                   ��      ��       Y��      ł       �Y�ł      �       Y�      �       w �      ,�       Y,�      >�       w >�      @�       �`@�      V�       YV�      u�       �h                             ��      ��       0���      Ă       SĂ      ł       y ł      1�       0�1�      ?�       S?�      @�       y @�      u�       0�                  W�      u�       P                   �      ,�       X,�      @�       �X�                   �      ,�       Z,�      @�       �U�                    ��      ��       U��      �       �U�                          ��      ��       T��      ��       V��      ΃       �T�΃      ��       V��      �       �T�                        ��      ��       Q��      ˃       ]˃      ΃       �Q�΃      �       ]                          ��      ��       R��      ��       S��      ΃       �R�΃      Ӄ       SӃ      �       �R�                            ��      ��       X��      ��       �X���      ��       P��      ̓       ^̓      ΃       P΃      �       ^                        ��      ��       Y��      Ƀ       \Ƀ      ΃       �Y�΃      �       \                        @q      Sq       USq      {q       �U�{q      �q       U�q      �q       �U�                            @q      Sq       TSq      yq       Syq      {q       �T�{q      �q       S�q      �q       T�q      �q       S                          @q      Sq       QSq      zq       Vzq      {q       �Q�{q      �q       Q�q      �q       V                 @q      �q       ��                              @q      Sq       TSq      yq       Syq      {q       �T�{q      �q       S�q      �q       T�q      �q       S                       @q      Sq       USq      {q       �U�{q      �q       U�q      �q       �U�                         @q      Wq       0�Wq      hq       P{q      �q       0��q      �q       P�q      �q       R                  q      ?q       P                      �p      �p       U�p      �p       �U��p      q       U                        �p      �p       T�p      �p       u �p      �p       �T��p      q       T                      �p      �p       Q�p      �p       �Q��p      q       Q                        p      Lp       ULp      �p       �U��p      �p       U�p      �p       �U�                          p      Up       TUp      �p       S�p      �p       �T��p      �p       T�p      �p       S                          p      Yp       QYp      �p       V�p      �p       �Q��p      �p       Q�p      �p       V                      `p      dp       Pdp      �p       \�p      �p       \                           ip      wp       Uwp      �p       w �p      �p       U�p      �p       U�p      �p       u ��p      �p       u �ɚ�r@J$" %��p      �p       w �ɚ�r@J$" %��p      �p       U                  ip      �p       1��p      �p       1��p      �p       	��                           o      @o       U@o      �o       �U��o      �o       U�o      �o       �U��o      �o       U                        Mo      Qo       PQo      ~o       S~o      �o       r ��o      �o       S                           Vo      do       Qdo      oo       u oo      oo       Q�o      �o       Q�o      �o       q ��o      �o       q �ɚ�r@J$" %��o      �o       u �ɚ�r@J$" %��o      �o       Q                  Vo      oo       1��o      �o       1��o      �o       	��                            �m      �m       U�m      �n       S�n      �n       �U��n      �n       S�n      �n       �U��n      �n       U                        �m      �m       T�m      n       Zn      �n       �T��n      �n       T                        n      n       Pn      �n       V�n      �n       V�n      �n       R                 Tn      �n       1v$�                           n      #n       Q#n      3n       u 3n      3n       T�n      �n       Q�n      �n       q ��n      �n       q �ɚ�r@J$" %��n      �n       u �ɚ�r@J$" %��n      �n       T                  n      3n       1��n      �n       1��n      �n       	��                         3n      An       QAn      Ln       �XLn      Ln       Q�n      �n       Q�n      �n       q ��n      �n       q �ɚ�r@J$" %��n      �n       �X�ɚ�r@J$" %��n      �n       Q                 3n      Ln       1��n      �n       1��n      �n       	��                      `m      �m       U�m      �m       u �m      �m       �U�                      `m      �m       T�m      �m       t �m      �m       �T�                      �l      �l       U�l      �l       T�l      Xm       �U�                      �l      �l       U�l      �l       T�l      �l       �U�                  �l      �l       W                      m      %m       P%m      *m       R*m      Sm       w                      m      m       1�m      m       	��m      'm       T'm      *m       t �*m      Sm       T                 m      ;m       Q                        m      %m       P%m      *m       R*m      /m       P/m      Sm       R                    Fm      Sm       PSm      Xm       q �                 Fm      Sm       P                      �l      �l       U�l      �l       T�l      �l       �U�                      �l      �l       U�l      �l       T�l      �l       �U�                  �l      �l       W                      �l      �l       U�l      �l       T�l      �l       �U�                      �l      �l       U�l      �l       T�l      �l       �U�                  �l      �l       W                            �i      j       Uj      |j       V|j      �j       �U��j      l       Vl      6l       U6l      �l       V                          �i      �i       T�i      j       s|��j      �j       s|��k      �k       Sl      l       Sl      6l       T                            �i      j       Qj      ~j       \~j      �j       �Q��j      l       \l      6l       Q6l      �l       \                              j      7j       0�7j      Yj       PYj      ^j       �L�j      �j       0��j      �k       0��k      �k       P�k      l       0�6l      �l       0�                          �i      j       0�j      �j       ]�j      �j       ]�j      �k       ]�k      �k       1��k      l       ]l      6l       0�6l      �l       ]                                           j      7j       Q�j      �j       Q�j      �j       q��j      k       Qk      k       q�k      0k       Q0k      8k       q�8k      =k       Q=k      Hk       q�Hk      Qk       QQk      `k       q�`k      xk       Qxk      �k       q��k      �k       Q�k      �k       q��k      �k       Q�k      l       Ql      l       X6l      [l       Qbl      �l       Q�l      �l       Q                                 �j      �j       P�j      �j       P)k      0k       P2k      =k       PLk      Qk       Psk      xk       P�k      �k       P�k      �k       P�k      l       P                         �j      �j       8��j      �j       R)k      0k       8�2k      =k       0�Lk      Qk       0�sk      xk       @��k      �k       @��k      �k       H�                        �j      �j       R�k      l       R6l      Pl       s~�
��| "�bl      nl       s~�
��| "��l      �l       s~�
��| "�                          j      7j       s}���l      l       s}���6l      Pl       s}���bl      nl       s}����l      �l       s}���                 <j      vj       V                 Cj      Yj       v8                  Gj      Yj       T                  Gj      Yj       v8                        Pi      �i       U�i      �i       S�i      �i       �U��i      �i       S                            Pi      ci       Tci      �i       V�i      �i       �T��i      �i       V�i      �i       �T��i      �i       V                       Pi      �i       0��i      �i       Q�i      �i       q��i      �i       0��i      �i       s t "��i      �i       Q                     Pi      �i       0��i      �i       P�i      �i       0�                        �f      $g       U$g      Gg       SGg      `g       �U�`g      lg       S                            �f      g       Tg      Hg       VHg      Ig       �T�Ig      _g       V_g      `g       �T�`g      lg       V                       �f      4g       0�4g      4g       Q4g      :g       q�Ig      `g       0�`g      hg       s t "�hg      lg       Q                     �f      :g       0�:g      Ig       PIg      lg       0�                        `f      �f       U�f      �f       S�f      �f       �U��f      �f       S                            `f      sf       Tsf      �f       V�f      �f       �T��f      �f       V�f      �f       �T��f      �f       V                       `f      �f       0��f      �f       Q�f      �f       q��f      �f       0��f      �f       s t "��f      �f       Q                     `f      �f       0��f      �f       P�f      �f       0�                        �e      f       Uf      /f       S/f      Hf       �U�Hf      \f       S                            �e      �e       T�e      0f       V0f      1f       �T�1f      Gf       VGf      Hf       �T�Hf      \f       V                       �e      f       0�f      f       Qf      "f       q�1f      Hf       0�Hf      Xf       s t "�Xf      \f       Q                     �e      "f       0�"f      1f       P1f      \f       0�                        b      Db       UDb      ob       Sob      �b       �U��b      �b       S                            b      #b       T#b      pb       Vpb      qb       �T�qb      �b       V�b      �b       �T��b      �b       V                       b      Tb       0�Tb      Tb       QTb      bb       q�qb      �b       0��b      �b       s t "��b      �b       Q                     b      bb       0�bb      qb       Pqb      �b       0�                            �a      �a       U�a      �a       S�a      �a       �U��a      �a       S�a      �a       �U��a      b       S                            �a      �a       T�a      �a       V�a      �a       �T��a      �a       V�a      �a       �T��a      b       V                  b      b       P                    ta      �a       Q�a      �a       q��a      �a       Q                   pa      �a       0��a      �a       P                    Ta      `a       Q`a      fa       q�fa      oa       Q                   Pa      ja       0�ja      oa       P                    $a      0a       Q0a      ;a       q�;a      Na       Q                    a      Ia       0�Ia      Na       P                    �`       a       Q a      a       q�a      a       Q                   �`      a       0�a      a       P                    �`      �`       Q�`      �`       q��`      �`       Q                   �`      �`       0��`      �`       P                 �`      �`       0�                              �^      _       U_      v_       Sv_      |_       �U�|_      �_       S�_      �_       �U��_      �_       U�_      `       S                                    �^      _       T_      w_       Vw_      |_       �T�|_      �_       T�_      �_       V�_      �_       �T��_      �_       T�_      �_       �T��_      �_       T�_      `       V                      �^      m_       0�m_      q_       P|_      �_       0��_      �_       P�_      �_       0��_      `       @�                       B_      S_       PS_      q_       ]�_      �_       P�_      �_       ]                 �^      _       u8                  _      )_       �   |_      �_       �   �_      �_       �                       _      _       T_      )_       V|_      �_       T�_      �_       V                  _      )_       0�|_      �_       0��_      �_       0��_      �_       @�                    _       _       0� _      )_       P|_      �_       0��_      �_       P�_      �_       0�                 G_      S_       T                    �^      �^       U�^      �^       �U�                      �^      �^       T�^      �^       S�^      �^       �T�                   �^      �^       u8�^      �^       P                  �^      �^       T                    �^      �^       u8�^      �^       P                       `      0`       U0`      R`       SR`      T`       �U�                     `      0`       T0`      T`       �T�                       `      0`       Q0`      S`       VS`      T`       �Q�                  1`      T`       P                        @^      o^       Uo^      w^       Sw^      �^       �U��^      �^       S                            @^      m^       Tm^      o^       Qo^      �^       �T��^      �^       T�^      �^       X�^      �^       �T�                            @^      j^       Qj^      o^       Ro^      �^       �Q��^      �^       Q�^      �^       R�^      �^       �Q�                               @^      s^       0�s^      w^       V�^      �^       0��^      �^       Y�^      �^       sp ��^      �^       ss��^      �^       Q�^      �^       V                          �]      �]       U�]      �]       V�]      ^       �U�^      ^       U^      -^       V                        �]      �]       T�]      �]       S�]      ^       �T�^      -^       S                        �]      �]       Q�]      ^       �Q�^      *^       P*^      -^       �Q�                          �]      �]       R�]      �]       ]�]      ^       �R�^      *^       R*^      -^       ]                   �]       ^       0� ^      ^       U�^      -^       0�                    �]      �]       \^      -^       \                        ��      �       U�      %�       �U�%�      H�       UH�      �       �U�                    ��      ݪ       Tݪ      �       �T�                      ��      �       Q�      �       S�      %�       �Q�%�      �       S                      ��      �       U�      �       �U�%�      H�       UH�      �       �U�                   ��      �       V%�      �       V                  ,�      �       \                  ;�      �       ]                   a�      |�       _ի      ۫       _�      �       _                   a�      |�       ]ի      ۫       ]�      �       ]                  a�      |�       0�ի      ۫       0��      �       0�                  ��      ��      	 v �
���                  ��      ��       Q                    ��      ��       U��      ��       ]                 ��      ��       v                 ��      ��       \                        �      p�       Up�      ��       �U���      ө       Uө      ��       �U�                    �      X�       TX�      ��       �T�                        �      T�       QT�      ��       V��      ��       �Q���      ��       V                 ��      ��       0�                       ;�      p�       Up�      ��       �U���      ө       Uө      ��       �U�                    [�      ��       S��      ��       S                  ��      ��       \                  Ʃ      ��       ]                   �      �       _:�      @�       _s�      s�       _                   �      �       ]:�      @�       ]s�      s�       ]                  �      �       0�:�      @�       0�s�      s�       0�                   �      $�       R                   �      $�       s                     �      $�       U$�      %�       ]                 H�      W�       s                 H�      X�       \                          �q      r       Ur      Er       SEr      �r       �U��r      �r       S�r      �r       �U�                            �q      r       Tr      br       Vbr      jr       Tjr      �r       �T��r      �r       V�r      �r       �T�                          �q      r       Qr      �r       \�r      �r       �Q��r      �r       \�r      �r       �Q�                           �q      2r       0�2r      Ir       PIr      �r       S�r      �r       P�r      �r       S�r      �r       P                      Mr      jr       Pjr      �r       ]�r      �r       P                  qr      �r       V�r      �r       V                   r      1r       } p "�                    `v      �v       U�v      �v       �U�                      `v      zv       Tzv      �v       ���v      �v       �T�                          `v      uv       Quv      �v       V�v      �v       �Q��v      �v       V�v      �v       �Q�                 `v      �v       0�                          �v      �v       P�v      �v       S�v      �v       P�v      �v       S�v      �v       P                        �v      �v       V�v      �v       �Q��v      �v       V�v      �v       �Q�                    �v      �v       �+�   �v      �v       �+�                       �v      �v       �T��v      �v       �T�                    �v      �v       U�v      �v       U                    �v      �v       �U��v      �v       �U�                  �v      �v        ��v      �v        �                �v      �v       0�                �v      �v       V                 �v      �v       \                 �v      �v       V                 �v      �v       V                 �v      �v       \                              �v      w       Uw      Kw       VKw      Rw       �U�Rw      bw       Vbw      iw       �U�iw      {w       V{w      �w       �U�                    �v      �v       T�v      �w       �T�                      �v      �v       Q�v      w       Tw      �w       �Q�                              �v      w       Rw      Ow       ]Ow      Rw       �R�Rw      fw       ]fw      iw       �R�iw      w       ]w      �w       �R�                              �v      w       Xw      Qw       ^Qw      Rw       �X�Rw      hw       ^hw      iw       �X�iw      �w       ^�w      �w       �X�                            w      -w       P-w      Aw       SAw      Rw       0�Rw      aw       Saw      fw       } fw      iw       �Riw      yw       P                      .w      @w       P@w      Rw       �LRw      iw       P                      w      Mw       \Rw      dw       \iw      }w       \                 6w      Aw       S                 6w      Aw       \                              �w      �w       U�w      �w       V�w      �w       �U��w      x       Vx      	x       �U�	x      x       Vx      "x       �U�                    �w      �w       T�w      "x       �T�                      �w      �w       Q�w      �w       T�w      "x       �Q�                              �w      �w       R�w      �w       ]�w      �w       �R��w      x       ]x      	x       �R�	x      x       ]x      "x       �R�                              �w      �w       X�w      �w       ^�w      �w       �X��w      x       ^x      	x       �X�	x      !x       ^!x      "x       �X�                            �w      �w       P�w      �w       S�w      �w       0��w      x       Sx      x       } x      	x       �R	x      x       P                      �w      �w       P�w      �w       �L�w      	x       P                      �w      �w       \�w      x       \	x      x       \                 �w      �w       S                 �w      �w       \                    �r      �r       U�r      s       �U�                    �r      �r       T�r      s       �T�                      �r      �r       Q�r      �r       T�r      s       �Q�                          �r      �r       R�r      �r       V�r      �r       �R��r      s       Vs      s       �R�                          �r      �r       X�r      �r       S�r      �r       �X��r      s       Ss      s       �X�                        �r      �r       P�r      �r       v �r      �r       �R�r      s       P                 �r      �r       u                     s      's       U's      Ts       �U�                    s      s       Ts      Ts       �T�                      s      s       Qs      +s       T+s      Ts       �Q�                          s      +s       R+s      Ds       VDs      Es       �R�Es      Ss       VSs      Ts       �R�                          s      +s       X+s      Cs       SCs      Es       �X�Es      Rs       SRs      Ts       �X�                        ,s      7s       P7s      Ds       v Ds      Es       �REs      Qs       P                 s      s       u                         �s      �s       U�s      Kt       _Kt      Lt       �U�Lt      �t       _                    �s      t       Tt      �t       �T�                        �s      t       Qt      Et       \Et      Lt       �Q�Lt      �t       \                        �s      t       Rt      It       ^It      Lt       �R�Lt      �t       ^                        �s      t       Xt      Gt       ]Gt      Lt       �X�Lt      �t       ]                     �s      3t       0�3t      ;t       PLt      ]t       P                 t      2t                              t      2t       P2t      ;t       SLt      it       S                        `s      hs       Uhs      �s       _�s      �s       �U��s      �s       _                    `s      �s       T�s      �s       �T�                        `s      �s       Q�s      �s       \�s      �s       �Q��s      �s       \                        `s      �s       R�s      �s       ^�s      �s       �R��s      �s       ^                        `s      �s       X�s      �s       ]�s      �s       �X��s      �s       ]                     `s      �s       0��s      �s       P�s      �s       P                 �s      �s                              �s      �s       P�s      �s       S�s      �s       S                              0x      Sx       USx      �x       V�x      �x       �U��x      �x       V�x      �x       �U��x      �x       V�x      �x       �U�                    0x      5x       T5x      �x       �T�                      0x      :x       Q:x      Wx       TWx      �x       �Q�                              0x      Wx       RWx      �x       ]�x      �x       �R��x      �x       ]�x      �x       �R��x      �x       ]�x      �x       �R�                              0x      Wx       XWx      �x       ^�x      �x       �X��x      �x       ^�x      �x       �X��x      �x       ^�x      �x       �X�                            Xx      mx       Pmx      �x       S�x      �x       0��x      �x       S�x      �x       } �x      �x       �R�x      �x       P                      nx      �x       P�x      �x       �L�x      �x       P                      Px      �x       \�x      �x       \�x      �x       \                 vx      �x       S                 vx      �x       \                    �h      �h       U�h      i       �U�                        �h      i       Ti      i       Ui      i       �T�i      i       T                      �h      i       Qi      i       �Q�i      i       Q                      �h      i       Ri      i       �R�i      i       R                      �h      i       Xi      i       �X�i      i       X                      �[      �[       U�[      |\       _|\      }\       �U�                      �[      �[       T�[      z\       ^z\      }\       �T�                    �[      �[       Q�[      }\       ��                    �[      �[       R�[      }\       �R�                      �[      �[       X�[      x\       ]x\      }\       �X�                      �[      �[       Y�[      v\       \v\      }\       �Y�                       �[      �[       0��[      1\       S1\      5\       s�;\      `\       S`\      d\       s�                 �[      \       0�R\      R\       0�                 �[      \       ^R\      R\       ^                 �[      \       0�R\      R\       0�                        p�      ��       U��      e�       �U�e�      r�       Ur�      �       �U�                        p�      ��       T��      [�       S[�      e�       �T�e�      �       S                              p�      ��       Q��      T�       _T�      e�       �Q�e�      r�       Qr�      ��       �Q���      ��       _��      �       �Q�                        p�      ��       R��      e�       ��e�      r�       Rr�      �       ��                                p�      ��       X��      T�       ^T�      e�       �X�e�      r�       Xr�      =�       ^=�      @�       �X�@�      O�       ^O�      �       �X�                        p�      ��       Y��      e�       �Y�e�      r�       Yr�      �       �Y�                        �      ��       0���      T�       V��      5�       V@�      O�       V                                 !�      =�       0�=�      Ȑ       \ؐ      �       \4�      @�       \�      ��       0���      ��       Q��      ��       q�đ      ё       \�      �       0�                        Ԏ      �      	 p 0$0&��      T�       \y�      8�       \@�      O�       \                      �      &�      	 p 0$0&�&�      <�       ���0$0&���      �       ���0$0&�                          ��      �       P�      <�       ]P�      T�       P��      �       ]@�      O�       ]                      '�      <�      	 p 0$0&���      ��      	 p 0$0&���      =�       _@�      O�       _                          ��      ��       P��      ��       u ��      e�       ��e�      r�       u r�      �       ��                        u�      ��       P��      Đ       _4�      @�       _đ      ё       _                         ��      T�       0�e�      �       0�4�      w�       0�w�      đ       Pđ      �       0�                             ��      T�       0�e�      �       0��      &�       P&�      +�       ]+�      4�       0�4�      @�       ]@�      O�       0�O�      �       ]                    ��      ��       Q��      ��       _e�      r�       Q                    ��      ��       T��      ��       Se�      r�       S                  ��      ��       0�e�      r�       0�                  Ǐ      �       _@�      O�       _                  Ǐ      �       S@�      O�       S                  Ǐ      �       0�@�      O�       0�                   =�      Y�       2��      �       2�                   =�      Y�       S�      �       S                    =�      ��       ^��      �       ^                        =�      ؐ       S��      �       S4�      @�       Sđ      ё       S                       =�      ؐ       0���      �       0�4�      @�       0�đ      ё       0�                   }�      ��       4�4�      @�       4�                   }�      ��       S4�      @�       S                      ��      ؐ       ^4�      @�       ^đ      ё       ^                      ��      ؐ       S4�      @�       Sđ      ё       S                     ��      ؐ       0�4�      @�       0�đ      ё       0�                 �      +�       ]                 �      +�       ��                        �b      �b       U�b      �e       �U��e      �e       U�e      �e       �U�                                �b      �b       T�b      De       SDe      Le       �T�Le      de       Sde      ne       �T�ne      �e       S�e      �e       �T��e      �e       S                              �b      �b       Q�b      d       \d      ne       �Q�ne      e       \e      �e       �Q��e      �e       Q�e      �e       �Q�                                  �b      �b       R�b      Ke       ^Ke      Le       �R�Le      me       ^me      ne       �R�ne      �e       ^�e      �e       �R��e      �e       R�e      �e       ^                                  �b      �b       X�b      Ie       ]Ie      Le       �X�Le      ke       ]ke      ne       �X�ne      �e       ]�e      �e       �X��e      �e       X�e      �e       ]                :e      =e       0�                        }c      .d       U.d      e       \Le      Ze       \ne      e       U�e      �e       \                    �c      d       Qne      e       Q                    �c      d       Pne      e       P                  �d      �d       T                    �d      �d       R�e      �e       R                    �d      �d       P�d      �d       p�                  e      e      	 p 0$0&�                    �b      �b       Q�b      �b       \�e      �e       Q                    �b      �b       T�b      �b       S�e      �e       S                
  �b      �b       0��e      �e       0�                 �b      �b       @�                   �b      �b       Q�b      �b       ���                   �b      �b       U�b      �b       S                  .d      Vd       \Le      Ze       \                  .d      Vd       SLe      Ze       S                  .d      Vd       0�Le      Ze       0�                 wd      ~d       @�                   wd      {d       Q{d      ~d       �@�                   wd      {d       U{d      ~d       S                   �d      �d       8��e      �e       8�                   �d      �d       S�e      �e       S                    �d      e       V�e      �e       V                   �d      =e       S�e      �e       S                  �d      =e       0��e      �e       0�                   e      :e       \�e      �e       \                   e      :e       S�e      �e       S                  e      :e       0��e      �e       0�                    �Z      �Z       U�Z      �[       X                  �Z      [       T                    �Z      �Z       U�Z      �[       X                 W[      �[       x� �                 W[      �[       Q                  T[      W[       R                 T[      W[       Q                  I[      L[       R                 I[      L[       Q                            0X      KX       UKX      �Y       \�Y      �Y       �U��Y      �Y       \�Y      �Y       �U��Y      �Z       \                  0X      SX       T                              0X      7X       Q7X      qX       ^qX      �X       �Q��X      �X       ^�X      �Y       �Q��Y      �Y       ^�Y      �Z       ^                    0X      <X       R<X      �Z       �R�                            FX      KX       UKX      �Y       \�Y      �Y       �U��Y      �Y       \�Y      �Y       �U��Y      �Z       \                     �X      �X       }d��X      �X       ^�X      yY       ^                  �X      yY       Q                   �X      TY       ~TY      yY       X                  �X      yY       P                   �X      TY       ~TY      yY       Z                   �X      TY       ~TY      yY       R                   �X      TY       ~TY      yY       Y                   �X      TY       ~TY      yY       T                 �X      TY       ~                  qX      �X       ^                   �Y      �Y       ^�Y      �Y       �Q�                   rZ      �Z       ^�Z      �Z       ^                 �Z      �Z       ^                  �Z      �Z       P                 dZ      rZ       ^                    CZ      CZ       PCZ      MZ       p  $0 $+( ��Z      �Z       P                 �Z      �Z       ^                            �S      #T       U#T      8T       S8T      QT       �U�QT      wT       SwT      �W       ���W      �W       U                        �S      T       TT      	T       R	T      �W       ���W      �W       T                            �S      T       QT      #T       P#T      QT       ��QT      YT       PYT      �W       ���W      �W       Q                    fT      �T       ^�T      �W       \                     fT      wT       0�wT      [W       ��~zW      �W       ��~                           fT      wT       0�wT      �T       _�T      �T       V�T      jW       ��jW      zW       _zW      �W       ��                        �T      �T       Y�T      aW       ^aW      zW       YzW      �W       ^                      (T      6T       P6T      8T       ��YT      �W       ��                  �T      �T       0��0��/U      :U      
 ������                           �T      �T       0��0���T      GU      
 ��~���~�GU      �U      
 ��~���~��U      �U       ��~���U      jW      
 ��~���~�zW      �W      
 ��~���~�                                     !V      !V       U��!V      (V       U�P�(V      bV       U����bV      gV       U����gV      �V       U���V      �V       P��W      W       �P��W      �W       U�����W      �W       U���W      �W       �P��W      �W       U���W      �W       P��                        wT      �T       0��T      /U       ]/U      :U       Z:U      {V       ]PW      �W       ]                       U      GU       ZxU      }U       ��~}U      PW       ZzW      �W       Z                   wT      �T       0��T      �W       ��~                    {V      W       ]�W      �W       ]                       bV      gV      L ��y ��y ?&#��"@& $ &��~� $ &{ ��~� $ &{ ?&"#��@& $ &�gV      W       ��~�W      �W       R�W      �W       ��~                                �U      �V       X�V      �V       ���V      W       XW      W       ��zW      �W       X�W      �W       ���W      �W       X�W      �W       ��                       �T      �T       Y�T      9W       S9W      =W       q�=W      �W       S                  �T      �W       V                     �T      �T       	���T      �U       ��~�U      �W       ��~                �U      �U       ��                �U      �U       P                 �U      �U       T�U      �U       t ��"#���                �U      �U       t ?&�                �U      �U       ��                �U      �U       U                   �U      �U       X�U      �U      
 r x "#���                  �U      �U       x ?&��U      �U       R                {V      �V       ��~                {V      �V       Y                {V      �V       ��~                {V      �V       ��                   �V      �V       P�V      �V      
 p r "#���                  �V      �V       p ?&��V      �V       R                 �V      �V       X                 �V      �V       ]                 �V      �V       X                 �V      �V       ]                �V      �V       ��~                �V      �V       ��                �V      �V       ��~                �V      �V       ��                   �V      �V       R�V      �V      
 q r "#���                  �V      �V       r ?&��V      �V       Q                     T      #T       U#T      (T       SQT      YT       S                   T      8T       0�QT      �W       0�                     X      X       UX      X       �U�                     X      X       TX      X       �T�                      @S      tS       UtS      zS       �U�zS      �S       U                      @S      tS       TtS      zS       �T�zS      �S       T                        @S      TS       QTS      tS       w tS      zS       �Q�zS      �S       Q                        �R      �R       U�R      S       VS      S       �U�S      7S       U                        �R      �R       T�R      �R       q�R      S       �T�S      7S       T                        �R      �R       Q�R      S       \S      S       �Q�S      7S       Q                         �R      �R       C��R      
S       P
S      S       C�S      S       P0S      7S       C�                     �R      �R       X�R      S       rS      S       X                        �R      S       SS      S       RS      S       S0S      5S       S                 �R      S       ��                    �R      S       ltuo�                 �R      S       V                    �R      S       RS      S       S                 �R      S       0�                      �R      �R       X�R      S       rS      S       X                      �Q      �Q       0��Q      fR       XmR      yR       X                      �Q      �Q       0��Q      ER       RmR      yR       R                  R      yR       Y                   R      R       QR      0R       qp�0R      9R       Q                    R      R       PR      0R       p�0R      =R       P                    R      R       Z��R      5R       Z�T�                    =R      RR       PRR      ]R       p�]R      iR       P                    @R      VR       QVR      ]R       q�]R      qR       Q                  KR      bR       R                      PQ      XQ       UXQ      ]Q       �U�]Q      fQ       U                      PQ      \Q       T\Q      ]Q       �T�]Q      fQ       T                        �P      �P       U�P      +Q       V+Q      ,Q       �U�,Q      FQ       U                        �P      �P       T�P      *Q       S*Q      ,Q       �T�,Q      FQ       T                  �P      �P       T                    �P      �P       U�P      �P       V                 �P      �P       T                 �P      �P       V                 �P      �P       T                 �P      �P       V                          �O       P       U P      AP       SAP      CP       �U�CP      YP       UYP      �P       S                              �O       P       T P      BP       VBP      CP       �T�CP      YP       TYP      rP       VrP      �P       T�P      �P       V                   )P      5P       v �1�5P      CP       Q                    0E      TE       UTE      �E       �U�                    9E      zE      	 t 0$0&�zE      �E      	 t0$0&�                  =E      �E      	 x 0$0&�                    `E      lE       RlE      �E       Q�E      �E       R                      `E      dE       RdE      �E       Q�E      �E       R                  `E      lE       PlE      pE       p�                      ��      ��       U��      ��       �U���      �       U                      ��      ��       T��      ��       �T���      �       T                      ��      ��       Q��      ��       �Q���      �       Q                      ��      ��       R��      ��       �R���      �       R                                    p@      �@       U�@      �A       ��~�A      B       �U�B      �D       ��~�D      �D       �U��D      �D       ��~�D      �D       U�D      �D       �U��D      �D       U�D      .E       ��~                                    p@      �@       T�@      �A       w �A      B       �T�B      �D       w �D      �D       �T��D      �D       w �D      �D       T�D      �D       �T��D      �D       T�D      .E       w                                     p@      �@       Q�@      �A       ��~�A      B       �Q�B      �D       ��~�D      �D       �Q��D      �D       ��~�D      �D       Q�D      �D       �Q��D      �D       Q�D      .E       ��~                                +A      0A       S��0A      <A       S�Y�<A      @A       [�Y�@A      CA       [�S�CA      KA       {  ��S�KA      fA       {  ��s  ��B      B       {  ��s  ��B      B      
 �s  ��                                 KA      �A       ^�A      �A       P�A      �A       ^B      ]C       ^]C      iC       PiC      SD       ^�D      �D       ^�D      E       ^E      .E       ^                          �@      �A       \B      �D       \�D      �D       \�D      �D       |��D      �D       \�D      .E       \                                           NA      oA       ZoA      �A       ��~�A      �A       _�A      �A       SB      ^B       Z^B      ]C       S]C      iC       _C      �C       S�C      @D       �@D      HD       _HD      jD       S�D      �D       Z�D      E       SE      E       �E      .E       s�                                  {A      �A       P�A      �A       P�B      �B       POC      ]C       PzC      C       P4D      CD       PHD      VD       PjD      wD       P)E      .E       P                               �@      �@       0��@      �A       ��~B      �D       ��~�D      �D       p��D      �D       P�D      �D       ��~�#��D      �D       ��~�D      .E       ��~                     �@      �@       0��@      NA       Z�D      �D       Z                               UA      fA      	 r 8$8&��A      �A       q 38$8&��A      �A       s �38$8&�B      B      	 r 8$8&�^B      tB       s �38$8&��B      �B      	 t 8$8&�C      GC      	 t 8$8&�C      �C       s �38$8&�                        �@      �A       VB      �D       V�D      �D       V�D      .E       V                                  �@      �A       _�A      �A       ]B      ^B       _^B      iC       ]iC      C       _C      jD       ]jD      �D       _�D      �D       _�D      �D       _�D      .E       ]                            �@      �@      	 p 0$0&��@      �A       ��~�0$0&�B      �D       ��~�0$0&��D      �D      	 s 0$0&��D      �D       ��~�0$0&��D      .E       ��~�0$0&�                   �?      O@       6�O@      W@       0�W@      f@       6�                  @      W@       Z                      �?      �?       U�?      �?       �U��?      �?       U                     �?      �?       0��?      �?       P�?      �?       0�                  �?      �?       P                  �?      �?       P                          >      m>       Um>      '?       \'?      8?       0�8?      A?       UA?      V?       \V?      \?       U                      j>      m>       Pm>      8?       ��A?      V?       ��                 j>      m>       0�                          m>      �>       0��>      �>       v��>      �>       V�>      �>       v�A?      V?       0�                    �>      �>       S�>      �>       S                  �>      �>       ~                 ?      '?       \                 ?      '?       ��                     �=      �=       0��=      �=       Y�=      
>       0�                     �=      �=       0��=      �=       X�=      
>       0�                     �=      �=       0��=      �=       P�=      
>       0�                        �t      �t       U�t      �t       S�t      �t       �U��t      �t       U                        �t      �t       T�t      �t       V�t      �t       �T��t      �t       T                       �t      �t       0��t      �t       P�t      �t       Q�t      �t       0�                    �=      �=       U�=      �=       �U�                    �=      �=       T�=      �=       �T�                    �=      �=       Q�=      �=       �Q�                    �=      �=       R�=      �=       �R�                    �=      �=       U�=      �=       �U�                    �=      �=       T�=      �=       �T�                    �=      �=       Q�=      �=       �Q�                    �=      �=       R�=      �=       �R�                    p=      }=       U}=      ~=       �U�                    p=      }=       T}=      ~=       �T�                    p=      }=       Q}=      ~=       �Q�                    p=      }=       R}=      ~=       �R�                        �;       <       U <      A=       �U�A=      N=       UN=      k=       �U�                            �;      7<       T7<      l<       Sl<      v<       �T�v<      A=       SA=      N=       TN=      k=       S                      �;      �;       P�;      <       P<      <       px�<      2<       P                              �;      �;       Q�;       <       Q <      I<       U�<      �<       U)=      A=       UN=      R=       UR=      a=       qx�                     +<      e<       Se<      v<       0�v<      A=       SN=      k=       S                      /<      q<       ]v<      A=       ]N=      k=       ]                     /<      s<       ^v<      A=       ^N=      k=       ^                     /<      o<       \v<      A=       \N=      k=       \                 [<      e<       S                 [<      e<       ]                 v<      �<       S                  �<      �<       S                  �<      �<       Q                  �<      �<      
  ;@     �                      �<      �<       s ��<      �<       U�<      �<       s �                    �<      )=       SN=      k=       S                    �<      )=       \N=      k=       \                   �<      �<       | N=      a=       |                       �<      �<       V�<      )=       0�N=      g=       Vg=      k=       0�                 �<      �<       S                 �<      �<       |��                  �<      �<       V                   �<      )=       SN=      k=       S                 �<      �<       V                 �<      �<       |��                   �<      )=       \g=      k=       \                  �<      =       0�g=      k=       0�                  �<      =       ltuo�g=      k=       ltuo�                  �<      =       \g=      k=       \                   �<      =       Pg=      k=       P                	   �<      =       0�g=      k=       0�                    �<      	=       Q=      =       Q                    �:      �:       U�:      �:       �U�                    �:      �:       T�:      �:       �T�                    �:      �:       P�:      �:       P                    `:      �:       U�:      �:       �U�                      `:      �:       T�:      �:       \�:      �:       �T�                 ~:      �:       S                  �:      �:       ]                              p      �       U�      ��       V��      ��       �U���      ր       Uր      �       V�      /�       U/�      J�       V                              p      �       T�      ��       w ��      ��       ����      ր       Tր      �       w �      /�       T/�      J�       w                       !�      ��       ]ր      �       ]"�      J�       ]                                   p      �       0��      �       _�      0�       _H�      L�       PL�      ��       S��      ր       0�ր      �       S�      �       0��      �       S�      /�       0�/�      J�       S                    �      �       0��      /�       0�                 t�      x�       S                 �      �       S                   ր      ��       SɁ      Ձ       S/�      J�       S                   ր      ��       VɁ      Ձ       V/�      J�       V                    ڀ      ��       \Ɂ      Ձ       \/�      J�       \                             ڀ      �       0��      �       P�      u�       _u�      ��       T��      ��       _Ɂ      Ձ       _/�      6�       T6�      J�       _                   ��      Ձ       S/�      J�       S                      ��      0�       Q0�      V�       ��Ɂ      Ձ       ��                 Z�      i�       _                   Z�      a�       v��a�      i�       U                   i�      ��       V/�      6�       V                  i�      ��       0�/�      6�       0�                  i�      ��       ltuo�/�      6�       ltuo�                  i�      ��       V/�      6�       V                   p�      ��       P/�      6�       P                   i�      ��       0�/�      6�       0�                    z�      ��       Q��      ��       Q                      ��      ��       T��      Ɂ       _Ɂ      Ձ       _6�      J�       _                    ��      Ɂ       \Ɂ      Ձ       \6�      J�       \                 �      �       S                 �      �       ]                           :      <:       U<:      E:       PE:      F:       �U�F:      U:       PU:      V:       U                         :      A:       TA:      E:       QE:      F:       �T�F:      V:       T                 1:      E:       r�#                               9      �9       U�9      �9       ]�9      �9       U�9      :       ]:      :       �U�:      :       ]:      :       �U�:      :       U                               9      �9       T�9      �9       V�9      �9       T�9      �9       V�9      :       �T�:      :       V:      :       �T�:      :       T                               9      �9       Q�9      �9       \�9      �9       Q�9       :       \ :      :       �Q�:      :       \:      :       �Q�:      :       Q                             9      �9       0��9      �9       7��9      �9       P�9      �9       0��9      �9       7��9      �9       7�:      :       0�                         �9      �9       X�9      �9       X�9      �9       r�9      �9       X�9      �9       X                           69      �9       0��9      �9       S�9      �9       R�9      �9       0��9      �9       S:      
:       S                 O9      �9       �P�                    O9      �9       P                 O9      �9       U                  _9      �9       S                 O9      �9       0�                    i9      y9       X}9      �9       X                  �9      �9       �P�                     �9      �9       Y                  �9      �9       ]                  �9      �9       R                 �9      �9       0�                      �9      �9       X�9      �9       r�9      �9       X                          ��      Į       UĮ      �       X�      X�       �U�X�      v�       Xv�      ��       U                                  ��      ��       T��      0�       V0�      5�       �T�5�      @�       V@�      E�       �T�E�      S�       VS�      X�       �T�X�      v�       Vv�      ��       T                          ��      �       Q�      �       YE�      X�       QX�      v�       Yv�      ��       Q                        ��      �       R�      /�       S5�      ?�       SE�      ��       R                    ߮      �       TX�      v�       T                             ��      �       0��      �       P�      &�       0�&�      *�       P5�      E�       0�E�      X�       6�X�      ��       0�                      ��      *�       ]5�      D�       ]o�      v�       ]                  Į      ߮       V                  Į      ߮       U                 Į      ߮       T                  �8      9       0�9      9       0�                  �8      9       T9      9       T                  �8      9       U9      9       U                    �8      9       Q9      9       Q                  �8      9       0�9      9       0�                      �8       9       P 9      	9       q	9      9       P9      9       P                        88      P8       PP8      Q8       u Q8      ]8       P]8      ^8       u                            5      <5       U<5      j5       Sj5      k5       �U�k5      y5       Sy5      ~5       U                 O5      [5       P                   55      ?5       Q?5      N5       s                   <5      N5       U                   <5      O5       0�O5      [5       P                            �4      �4       U�4      �4       S�4      �4       �U��4      5       S5      5       �U�5      5       U                 �4      �4       P                   �4      �4       P�4      �4       u                   �4      �4       Q                   �4      �4       0��4      �4       P                             4      \4       U\4      4       S4      �4       �U��4      �4       S�4      �4       �U��4      �4       U                             4      U4       TU4      �4       V�4      �4       �T��4      �4       V�4      �4       �T��4      �4       T                             4      a4       Qa4      �4       \�4      �4       �Q��4      �4       \�4      �4       �Q��4      �4       Q                             4      a4       Ra4      �4       ]�4      �4       �R��4      �4       ]�4      �4       �R��4      �4       R                   b4      y4       P�4      �4       P                    74      a4       Y�4      �4       Y                       74      b4       0�b4      y4       P�4      �4       P�4      �4       0�                                �3      �3       U�3      �3       S�3      �3       U�3      �3       �U��3      �3       U�3      4       S4      4       �U�4      4       U                                �3      �3       T�3      �3       V�3      �3       T�3      �3       �T��3      �3       T�3      4       V4      4       �T�4      4       T                                �3      �3       Q�3      �3       \�3      �3       Q�3      �3       �Q��3      �3       Q�3      	4       \	4      4       �Q�4      4       Q                                �3      �3       R�3      �3       ]�3      �3       R�3      �3       �R��3      �3       R�3      4       ]4      4       �R�4      4       R                                �3      �3       X�3      �3       ^�3      �3       X�3      �3       �X��3      �3       X�3      4       ^4      4       �X�4      4       X                   �3      �3       P�3      4       P                    �3      �3       Y4      4       Y                       �3      �3       0��3      �3       P�3      4       P4      4       0�                               3      M3       UM3      f3       Sf3      h3       Uh3      i3       �U�i3      w3       Sw3      y3       �U�y3      �3       U                               3      F3       TF3      g3       Vg3      h3       Th3      i3       �T�i3      x3       Vx3      y3       �T�y3      �3       T                   S3      \3       Pi3      v3       P                  23      R3       Q                     23      S3       0�S3      \3       Pi3      v3       P                                  �2      �2       U�2      �2       S�2      �2       U�2      �2       �U��2      �2       S�2      �2       �U��2      �2       S�2      3       U3      3       S                   �2      �2       P�2      �2       0��2      �2       P                         �2      �2       P�2      �2       P�2      �2       0��2      �2       P3      3       P                   �2      �2       U�2      �2       U                      �2      �2       0��2      �2       0��2      �2       P3      3       P                                �1      �1       U�1      �1       S�1      �1       U�1      �1       �U��1      2       S2      2       �U�2      &2       U&2      �2       S                                  �1      �1       T�1      �1       V�1      �1       T�1      �1       �T��1      �1       T�1      2       V2      2       �T�2      L2       TL2      �2       V                            �1      �1       Q�1      �1       �Q��1      �1       Q�1      2       �Q�2      Q2       QQ2      �2       w                             �1      �1       R�1      �1       �R��1      �1       R�1      2       �R�2      Q2       RQ2      �2       �\                    �1      �1       P�1      2       0�j2      o2       P                        �1      �1       P�1      2       0�&2      :2       PR2      w2       P                    �1      �1       U72      Q2       U                     �1      �1       0�72      R2       0�R2      w2       P                                �0      1       U1      1       S1      1       U1      1       �U�1      #1       U#1      J1       SJ1      L1       �U�L1      �1       S                                �0      1       T1      1       V1      1       T1      1       �T�1      C1       TC1      K1       VK1      L1       �T�L1      U1       TU1      �1       V                   1      1       PC1      C1       0�g1      i1       P                       �0      1       P#1      21       PC1      C1       0�W1      w1       P                   /1      C1       UL1      V1       U                    /1      C1       0�L1      W1       0�W1      w1       P                            �7      �7       U�7      8       S8      8       �U�8      8       S8      8       �U�8      #8       U                            �7      �7       T�7      8       V8      8       �T�8      8       V8      8       �T�8      #8       T                    �7      8       P8      8       P                 �7      8       P                   �7      8       s�8      8       T                            p7      �7       U�7      �7       S�7      �7       �U��7      �7       S�7      �7       �U��7      �7       U                            p7      �7       T�7      �7       V�7      �7       �T��7      �7       V�7      �7       �T��7      �7       T                    �7      �7       P�7      �7       P                 �7      �7       P                   �7      �7       s��7      �7       T                            07      @7       U@7      Y7       SY7      _7       �U�_7      c7       Sc7      d7       �U�d7      k7       U                    E7      ^7       P_7      b7       P                 J7      ^7       P                   J7      Y7       s�Y7      ^7       T                      �6      �6       U�6      !7       �U�!7      %7       U                          �6      �6       T�6      7       S7      7       �T�7      !7       S!7      %7       T                          �6      �6       Q�6      7       V7      7       �Q�7      !7       V!7      %7       Q                    �6      7       	��7      7       P7      %7       	��                    �6      7       P7      7       P                 7      7       P                          p6      �6       U�6      �6       S�6      �6       �U��6      �6       S�6      �6       �U�                          p6      �6       T�6      �6       V�6      �6       �T��6      �6       V�6      �6       �T�                          p6      �6       Q�6      �6       \�6      �6       �Q��6      �6       \�6      �6       �Q�                    �6      �6       P�6      �6       P                       �6      �6       s��6      �6       T�6      �6       s��6      �6       �U#�                 �6      �6       P                   0      $0       T                     0      [0       Q[0      �0       Q                    0      �0       0��0      �0       7�                        /      :/       U:/      `/       V`/      d/       Ud/      y/       �U�                        /      :/       T:/      `/       �T�`/      d/       Td/      y/       �T�                          /      :/       Q:/      `/       \`/      d/       Qd/      x/       \x/      y/       �Q�                   /      d/       0�d/      y/       Q                       /      :/       0�O/      `/       P`/      d/       0�d/      t/       P                  :/      `/       S                      �/      �/       U�/      �/       S�/      �/       �U�                      �/      �/       T�/      �/       V�/      �/       �T�                       �/      �/       0��/      �/       P�/      �/       0��/      �/       P                 �/      �/       0��/      �/       0�                 �/      �/       S�/      �/       S                   �/      �/       0��/      �/       P�/      �/       0��/      �/       P                 �/      �/       U                            ��      Ԋ       UԊ      O�       SO�      b�       �U�b�      |�       U|�      ��       S��      ��       �U�                        ��      ̊       T̊      b�       ��b�      |�       T|�      ��       ��                          ��      ъ       Qъ      Y�       VY�      b�       �Q�b�      |�       Q|�      ��       V                          ��      ؊       R؊      [�       \[�      b�       �R�b�      |�       R|�      ��       \                   ��      ]�       ]|�      ��       ]                   ��      a�       _|�      ��       _                            ��      ܊       0�܊      ��       P��      _�       ^b�      |�       0�|�      ��       ^��      ��       T��      ��       0���      ��       ^                   |�      ��       ^��      ��       T                 |�      ��       ~                 |�      ��       ~                  ��      ��       S                   ��      ��       ^��      ��       T                 ��      ��       S                              @�      ��       U��      ��       �U���      ��       U��      Z�       VZ�      _�       �U�_�      a�       Ua�      v�       V                      V�      ��       \��      \�       \a�      v�       \                   V�      ��       |���      ɉ       |�                           V�      y�       0�y�      ��       P��      ��       S��      ��       p���      ��       P��      ��       0�                    ߉      J�       Qa�      v�       Q                    ŉ      ^�       ]a�      v�       ]                 .�      T�       VT�      _�       0�                 .�      J�       v                 .�      J�       v                   9�      Y�       S                 K�      T�       V                 K�      T�       S                          }.      �.       0��.      �.       P�.      �.       q��.      �.       Q�.      �.       0�                              �5      �5       U�5      �5       \�5      �5       �U��5      �5       U�5      �5       \�5      �5       �U��5      6       U                                �5      �5       T�5      �5       V�5      �5       �T��5      �5       T�5      �5       V�5      �5       |��5      �5       �U#��5      6       T                        �5      �5       S�5      �5       S�5      �5       u� �5      �5       S                    �5      �5       P�5      �5       P                      �-      d.       Td.      e.       �T�e.      n.       T                        .      (.       P).      A.       Pe.      m.       Pm.      n.       u�                   .      A.       R                              P-      �-       U�-      �-       S�-      �-       U�-      �-       �U��-      �-       S�-      �-       �U��-      �-       U                              P-      w-       Tw-      �-       ]�-      �-       T�-      �-       �T��-      �-       ]�-      �-       �T��-      �-       T                              P-      �-       Q�-      �-       V�-      �-       Q�-      �-       �Q��-      �-       V�-      �-       �Q��-      �-       Q                              P-      �-       R�-      �-       \�-      �-       R�-      �-       �R��-      �-       \�-      �-       �R��-      �-       R                   �-      �-       P�-      �-       P                    a-      �-       X�-      �-       X                       a-      �-       0��-      �-       P�-      �-       P�-      �-       0�                              `+      �+       U�+      �,       S�,      �,       �U��,      �,       S�,      �,       �U��,      �,       U�,      M-       S                                `+      �+       T�+      �,       �T��,      �,       T�,      �,       �T��,      �,       T�,      �,       �T��,      �,       T�,      M-       �T�                        `+      �+       Q�+      �,       �Q��,      �,       Q�,      M-       �Q�                              `+      �+       R�+      �,       \�,      �,       �R��,      �,       \�,      �,       �R��,      �,       R�,      M-       \                              `+      �+       X�+      �,       V�,      �,       �X��,      �,       V�,      �,       �X��,      �,       X�,      M-       V                         `+      �+       0��+      �+       P�+      �,       T�,      �,       0��,      M-       T                      y+      �+       P�+      �+       u��,      �,       u�                       ,      Q,       RQ,      Y,       v -      /-       R/-      M-       v                        ,      ,       U,      �,       X�,      �,       v�,      M-       U                  #,      U,       I�-      M-       I�                    #,      ',       p 
���',      U,      	 y�
���-      M-      	 y�
���                      #,      Q,       RQ,      U,       v -      /-       R/-      M-       v                   #,      U,       1�-      -       1�-      M-       	��                    #,      ',       p 
���',      U,      	 y�
���-      M-      	 y�
���                  #,      U,       I�-      M-       I�                       0,      A,       p�-I�-� �A,      D,       p �-I�-� �D,      U,       z �-I�-� �-      5-       <p �-I�-� �5-      M-       <y�
��v �-I�-� �                 	   U,      U,       R-      5-       <p �-I�-� �5-      M-       <y�
��v �-I�-� �                  d,      �,       I��,      -       I�                    d,      h,       p 
���h,      �,      	 y�
����,      -      	 y�
���                      d,      ,       U,      �,       X�,      �,       v�,      -       U                  d,      �,       1��,      �,       1��,      -       	��                    d,      h,       p 
���h,      �,      	 y�
����,      -      	 y�
���                  d,      �,       I��,      -       I�                       q,      �,       p�-I�-� ��,      �,       p �-I�-� ��,      �,       u �-I�-� ��,      -       <p �-I�-� �-      -       <y�
��u �-I�-� �                    �,      �,       X�,      -       <p �-I�-� �-      -       <y�
��u �-I�-� �                  �+      �+       y                   �+      �+       v                  �+      �+       y                  �+      �+       v                       �+      �+       P�+      �+      
 p q "#����+      �+       R                       �+      �+       p ?&��+      �+       Q�+      �+       p ?&��+      �+       v � $ &y � $ &?&�                 �+      
,       y(                 �+      
,       v                 �+      ,       y(                 �+      ,       v                     �+      �+       P�+       ,      
 p q "#��� ,      ,       U                   �+      �+       p ?&��+      ,       Q                      �*      O+       UO+      U+       �U�U+      Y+       U                        �*      +       T+      )+       Q)+      .+       �Q�U+      Y+       Q                          �*      �*       Q�*      +       �Q�+      )+       Q)+      .+       �Q�U+      Y+       Q                      `*      �*       U�*      �*       �U��*      �*       U                      `*      p*       T�*      �*       T�*      �*       �T�                          `*      p*       Qp*      �*       �Q��*      �*       �Q��*      �*       �Q@+( ��*      �*       Q�*      �*       �Q@+( �                            `*      �*       R�*      �*       R�*      �*       X�*      �*       �X��*      �*       R�*      �*       X                          `*      �*       X�*      �*       X�*      �*       X�*      �*       �X��*      �*       X                          �)      �)       U�)      �)       S�)      �)       �U��)      �)       U�)      _*       S                            �)      �)       T�)      �)       �T��)      )*       T)*      <*       �T�<*      W*       TW*      _*       �T�                        �)      �)       0��)      �)       P�)      **       0�**      9*       P<*      _*       0�                     �)      �)       s�#�)      )*       s�#<*      W*       s�#                     *      "*       �h�"*      **       R<*      G*       �h�                   *      **       0�<*      G*       0�                     *      )*       T)*      **       �T�<*      G*       T                   *      **       S<*      G*       S                            @%      h%       Uh%      �%       S�%      �%       U�%      P'       SP'      Z'       UZ'      )       S                                    @%      �%       T�%      C&       RC&      �&       �T��&      �&       R�&      Z'       �T�Z'      �'       R�'      �(       �T��(      �(       R�(      �(       �T��(      )       R                        U%      �%       \�%      S'       \S'      Z'       TZ'      )       \                                        a%      �%       0��%      �%       0��%      �%       T�%      �%       T�&      �&       0�Z'      s'       0�s'      {'       T{'      �'       0��'      �'       T�'      �'       0��'      �'       T�(      �(       0��(      )       0�                                              a%      �%       0��%      �%       0��%      �%       Y�%      �&       Y�&      �&       0�Z'      s'       0�s'      {'       T{'      �'       0��'      �'       T�'      �'       0��'      �'       Y�'      (       Y
(      �(       Y�(      �(       0��(      �(       Y�(      )       0�                                         a%      �%       0��%      '&       0�'&      �&       [�&      �&       0�''      /'       [/'      ='       {`�Z'      �'       0��'      �'       [�'      �'       P�'      �(       [�(      �(       0��(      �(       [�(      )       0�                                         a%      �%       0��%      W&       0�W&      �&       Z�&      �&       0�+'      3'       Z3'      A'       z`�Z'      �'       0��'      (       Z(      
(       P
(      �(       Z�(      �(       0��(      �(       Z�(      )       0�                   `&      �&       T6(      p(       T                   `&      �&       [6(      p(       [                   `&      �&       1�6(      6(       1�6(      p(       	��                   `&      �&       [6(      6(       [6(      p(       { �                   `&      �&       T6(      p(       T                      s&      �&       t 1%{ @$"�-t �-� ��&      �&       PP(      p(       { @$t 1%"�-t �-� �                    s&      �&       t 1%{ @$"�-t �-� ��&      �&       PP(      p(       { @$t 1%"�-t �-� �                     �&      �&       Yp(      �(       Y�(      �(       Y                     �&      �&       Zp(      �(       Z�(      �(       Z                     �&      �&       1�p(      p(       1�p(      �(       	���(      �(       1�                     �&      �&       Zp(      p(       Zp(      �(       z ��(      �(       Z                     �&      �&       Yp(      �(       Y�(      �(       Y                      �(      �(       z @$y 1%"�-y �-� ��(      �(       y 1%z @$"�-y �-� ��(      �(       P                    �(      �(       z @$y 1%"�-y �-� ��(      �(       y 1%z @$"�-y �-� ��(      �(       P                  �&      ''       v                     �&      '       P'      ''      
 s��
���                 �&      '       U                 �&      ''      
 s��
���                      '      '       U'      '      
 q u "#���'      ''       [                   '      '       u ?&�'      ''       Q                 ''      +'       v(                 ''      +'      
 s��
���                		 ''      ''       X''      +'       Z                 ''      +'       P                   �'      �'       Y
(      6(       Y                   �'      �'       Z
(      6(       Z                   �'      �'       1�
(      
(       1�
(      6(       	��                   �'      �'       Z
(      
(       Z
(      6(       z �                   �'      �'       Y
(      6(       Y                    �'      �'       y 1%z @$"�-y �-� �(      6(       z @$y 1%"�-y �-� �                  �'      �'       y 1%z @$"�-y �-� �(      6(       z @$y 1%"�-y �-� �                    �#      �#       T�#      >%       �T�                            �#      m$       r�m$      n$       Tn$      %       r�%      %       T%      =%       r�=%      >%       T                           �#      "$       T"$      m$       �T5$u� "�n$      �$       �T5$u� "��$      �$       T�$      %       �T5$u� "�%      =%       �T5$u� "�                    $      "$      
 u��
���"$      0$       Tn$      �$       T                    $      0$       Qn$      �$       Q�$      �$       �T5$u� "#                  $      0$       1�n$      n$       1�n$      �$       	��                    $      0$       Qn$      n$       Qn$      �$       q ��$      �$       �T5$u� "#�                   "$      0$       Tn$      �$       T                          0$      7$       t 1%q @$"�-t �-� �7$      B$       t 1%�T5$u� "#@$"�-t �-� �B$      O$       P|$      �$       q @$t 1%"�-t �-� ��$      �$       �T5$u� "#@$t 1%"�-t �-� �                   0$      0$       t 1%q @$"�-t �-� �|$      �$       q @$t 1%"�-t �-� ��$      �$       �T5$u� "#@$t 1%"�-t �-� �                      F$      a$       T�$      �$       T�$      %       T%      2%       T2%      5%      
 u��
���                          F$      V$       YV$      a$       �T5$u� "#�$      �$       Y�$      �$       P�$      %       Y%      #%       Y#%      5%       �T5$u� "#                    F$      a$       1��$      �$       1��$      %       1�%      %       1�%      5%       	��                           F$      V$       YV$      a$       �T5$u� "#�$      �$       Y�$      �$       P�$      %       Y%      %       Y%      #%       y �#%      5%       �T5$u� "#�                      F$      a$       T�$      �$       T�$      %       0�%      2%       T2%      5%      
 u��
���                            O$      V$       t 1%y @$"�-t �-� �V$      a$       t 1%�T5$u� "#@$"�-t �-� �a$      m$       P%      #%       y @$t 1%"�-t �-� �#%      2%       �T5$u� "#@$t 1%"�-t �-� �2%      =%      - �T5$u� "#@$u��
��1%"�-u��
���-� �                      a$      a$       P%      #%       y @$t 1%"�-t �-� �#%      2%       �T5$u� "#@$t 1%"�-t �-� �2%      5%      - �T5$u� "#@$u��
��1%"�-u��
���-� �                       7       t                           (       u��0$0&�(      0       Q0      7       u��0$0&�                       7       t                       7       u��0$0&�                   0      7       Q7      7      
 p q "#���                  0      7       q ?&�7      7       P                [      b       t                [      b       u��0$0&�                [      b       t                [      b       u��0$0&�                  [      b       Qb      b      
 p q "#���                  [      b       q ?&�b      b       P                w      �       t                    w             u��0$0&�      �       P�      �       u��0$0&�                w      �       t                w      �       u��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       t                    �      �       u��0$0&��      �       P�      �       u��0$0&�                �      �       t                �      �       u��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                      `#      �#       T�#      �#       �T��#      �#       T                      d#      z#       Qz#      }#       u}#      �#       X                            0"      �"       U�"      �"       S�"      �"       �U��"      �"       U�"      #       S#      '#       U                   _"      �"       0��"      #       0�                          V"      �"       \�"      �"       \�"      �"       u #��"      #       \#      '#       \                     _"      �"       |�"      �"       |�"      �"      	 u #�#                          F"      �"       V�"      �"       V�"      �"       u �"      #       V#      '#       V                     �"      �"       R�"      �"       0��"      #       0�                   _"      �"       U�"      �"       U                     _"      �"       v���"      �"       v���"      �"       u #��                    f"      �"       R�"      �"       R                 �"      �"       R                 �"      �"       v��                          0~      �~       U�~      �~       S�~      �~       �U��~      E       SE      f       U                          0~      �~       T�~      �~       \�~      �~       �T��~      E       \E      f       T                    x~      �~       V�~      E       V                 q~      �~       P                   q~      �~       ^�~      E       ^                           0~      �~       0��~      �~       P�~      �~       ]�~      �~       P�~      E       ]E      f       0�                               0~      �~       0��~      �~       0��~      �~       0��~      �~       P�~      �~       _�~      �~       P�~      7       _7      E       TE      f       0�                           0~      �~       0��~      �~       0��~      �~       0��~             P             }� E      f       0�                �~      �~       ]                �~      �~       V                 �~      �~       _                 �~      �~       V                 2      E       T                 2      E       U                        �!      �!       U�!      "       S"      "       �U�"      &"       U                   �!       "       #� "      "       0�"      &"       #�                 �!      "       V                 �!      �!       v                   �!      �!       R�!      "       0�                 �!      �!       U                 �!      �!       v �                  �!      �!       R                 �!      �!       R                 �!      �!       v �                        �x      �x       U�x      4y       V4y      �y       �U��y      �y       U                        �x      y       Ty      Qy       SQy      �y       �T��y      �y       T                      y      
y       P
y      -y       7�-y      ^y       P^y      cy       �L                      �x      y       \�y      �y       \�y      �y       u�                   
y      y       |y       y       P                  By      xy       V                   By      ^y       �Xty      xy       0�                  Qy      xy       S                 Qy      ^y       �X                 ky      ty       S                      �y      �y       U�y      �y       �U��y      �y       U                        �y      �y       T�y      �y       �H�y      �y       �T��y      �y       T                                                                    ��      @�       U@�      ��       S��      -�       �U�-�      ?�       S?�      S�       ��|S�      ��       �U���      Ŝ       ��|Ŝ      Ϝ       �U�Ϝ      �       S�      ��       ��|��      ��       U��      ǝ       �U�ǝ      x�       ��|x�      ��       �U���      ��       ��|��             S      ՟       �U�՟      �       ��|�      ��       S��      p�       ��|p�      s�       �U�s�      ��       ��|��      )�       �U�)�      8�       ��|8�      ��       �U���      �       ��|                                                        ��      @�       T@�      S�       VS�      ��       �T���      Ŝ       VŜ      Ϝ       �T�Ϝ      ��       V��      ��       T��      ǝ       �T�ǝ      x�       Vx�      ��       �T���      k�       Vk�      s�       _s�      �       V�      )�       _)�      8�       V8�      Y�       _Y�      ��       �T���      ��       _��      ޢ       Vޢ      �       �T�                              ��      '�       Q'�      j�       ��|j�      ��       �Q���      ��       ��|��      ��       Q��      ǝ       �Q�ǝ      �       ��|                          ��      @�       R@�      ��       ��|��      ��       R��      ǝ       �R�ǝ      �       ��|                                                  ��      @�       X@�      S�       ^S�      ��       �X���      Ŝ       ^Ŝ      Ϝ       �X�Ϝ      ��       ^��      ��       X��      ǝ       �X�ǝ      x�       ^x�      ��       �X���      .�       ^.�      s�       �X�s�      �       ^�      )�       �X�)�      8�       ^8�      ��       �X���      �       ^                                                      ��      m�       0�m�      ��       [��      Ě       ��|Ě      -�       _-�      ?�       0�?�      S�       [��      ��       ��|��      ��       [Ϝ      ��       0���      |�       _|�      ��       [��      ��       _��      ��       0�ǝ      M�       _M�      n�       [n�      }�       ��|��             [�      ��       [��      �       _��      ��       _��      Ȣ       0�Ȣ      �       _                                                 ��      U�       0�U�      X�       PX�      ��       s ��      -�       ��|-�      ?�       0�?�      ��       ��|��      Ϝ       ��|Ϝ      �       s �      ��       ��|��      ��       ��|��      ��       0�ǝ      ��       ��|��             s       �       ��|�      ��       s ��      ��       ��|��      �       ��|                                 ��      ؚ       0�ؚ      �       P�      �       T-�      ��       0���      ��       0�ǝ      ��       0�	�      �       P�      ��       0���      �       0�                                <�      S�       ]��      Ŝ       ]Ϝ      ��       ]ǝ      x�       ]��      ]�       ]s�      �       ])�      8�       ]��      �       ]                            �      ��       Sǝ      J�       S��      ��       S��      ��       S��      Ȣ       ��|#�Ȣ      ͢       S                        �      ��       \ǝ      M�       \��      ��       \��      �       \                     y�      ��       0���      ��       X�      ��       0�                     y�      ��       0���      ��       Y�      ��       0�                     ��      �       0��      �       X��      ��       0�                   ��      �       0���      ��       0�                  ՝      �       0�5�      =�       0�                       ՝      �       X�      ��       ��|5�      =�       X=�      =�       ��|                 ՝      �       0�5�      =�       0�                  ͢      ��       ]                  ͢      ��       S��      ��       0�                  ޢ      ��       V                 ޢ      �       S                 �      ��       S                 �      ��       V                  ��      ��       0�                   ��      ɛ       P֛      -�       P                    ��      �       P��      ��       P                   ��      �       P�      �       T                 ��      �       x�# �                 S�      X�       ]                  S�      X�       ��|��      ��       0�                  `�      ��       V                 ~�      ��       V                                M�      g�       V՟      ۟       V��      k�       Vk�      s�       _s�      ��       V�      )�       _)�      8�       V8�      Y�       _Y�      ��       �T���      ��       _                      M�      g�       ��|՟      ۟       ��|��      ��       ��|�      ��       ��|��      ��       ��|                      M�      g�       ��|՟      ۟       ��|��      ��       ��|�      ��       ��|��      ��       ��|                 M�      n�       ��|                       M�      g�       ��|՟      ۟       ��|��      p�       ��|s�      ��       ��|)�      8�       ��|                        I�      g�       P՟      ۟       U���      �       U���      ��       P)�      8�       P��      ��       0�                 M�      I�       ��|                 M�      I�       ��|                 M�      n�       ��|                 M�      I�       ��|                   ��      ��       0���      ��       P                        0�      3�      	 q  $ &�3�      7�       Q7�      ;�       q��;�      C�      , ���H0H%�$!0)( 8/�� $ &�                       0�      7�       q  $ &#	�#��7�      ;�       q� $ &#	�#��;�      ?�      4 ���H0H%�$!0)( 8/�� $ &#	�#��?�      C�       Q                V�      ��       0�                 V�      n�       ��|                V�      ��       0�                 ��      ��       ��                     ��      ��       ��~���      ��       P��      ��       ��|                           #�      k�       Vk�      s�       _�      )�       _8�      Y�       _Y�      ��       �T���      ��       _                      #�      s�       ��|�      )�       ��|8�      ��       ��|��      ��       ��|                      #�      s�       ��|�      )�       ��|8�      ��       ��|��      ��       ��|                           #�      G�       PG�      p�       Sp�      s�       ^�      )�       ^8�      R�       ^��      ��       ^                         .�      c�       ^c�      s�       ��|�      )�       ��|8�      ��       ��|��      ��       ��|                                  .�      p�       2�p�      ��       P��      �       P�      �       P�      �       ��|;�      s�       PM�      Y�       PY�      ��       \��      ��       0���      ��       P                            H�      p�       0�p�      ;�       \;�      ?�       |�V�      s�       \�      )�       \M�      Y�       0���      ��       \                        p�      ;�       Sd�      s�       1��      )�       S��      ��       S                         .�      p�       0�p�      s�       V�      )�       V8�      E�       V��      ��       V                 �      )�       0�                    �      �       T�      �       ��|                    ��      �       Q�      �       ��|                   ��      �       T�      �       ��|                 �      $�       T                 �      $�       Q                         p�      V�       ^V�      s�       ^�      )�       ^8�      R�       ^��      ��       ^                 V�      d�       \                 i�      o�       T                 i�      p�       ^                x�      ��       ]                 x�      ��       ��|                 ��      ��       V                 ��      ��       ��|                 ��      ��       V                  ǟ      ՟       ]                  ǟ      ՟       S                     �      
�       U
�      �       �U�                     �      
�       T
�      �       �T�                     �      
�       Q
�      �       �Q�                     �      
�       R
�      �       �R�                                                    �      $�       U$�      ,�       V,�      A�       �U�A�      ה       Vה      m�       ��~m�      ��       �U���      ѕ       Vѕ      o�       ��~o�      �       �U��      j�       Vj�      u�       ��~u�      ��       �U���      ��       V��      ��       �U���      Ә       VӘ      [�       �U�[�      ��       V��      ��       �U�                                          �      $�       T$�      ,�       S,�      A�       �T�A�      m�       Sm�      ��       �T���      ��       S��      �       �T��      ��       S��      ��       �T���      ޘ       Sޘ      [�       �T�[�      ��       S��      ��       �T�                    �      $�       Q$�      ��       �Q�                                �      �       R�      ,�       \,�      A�       �R�A�      Ȓ       \Ȓ      ��       �R���      ��       \��      ˔       |�˔      ��       �R�                    �      �       X�      ��       ��~                                 �      $�       P$�      3�       w 3�      A�       ��~A�      [�       w [�      {�       ��~{�      ��       w ��      ��       ��~��      ��       w                                            (�      ,�       PA�      v�       Pw�      ��       P��      ��       P��      �       Z�      �       ��~T�      ^�       ����      Ŕ       Pm�      r�       Z��      ��       Z��      ɕ       ���      4�       1�4�      >�       Z>�      C�       ^��      Ә       0�                        Œ      ��       Q��      �       �R~ ���      ��       Q4�      C�       Q                           Œ      T�       ��~��      ��       ��~4�      >�       ��~C�      j�       ��~��      ��       ��~��      ��       ��~[�      ��       ��~                            Œ      ϒ       Qϒ      �       \��      ��       \4�      >�       \C�      `�       \��      ��       \��      ��       \                       Œ      ��       R��      �       ~ ��      ��       R4�      >�       R                       Œ      ��       T��      �       ����      ��       T4�      >�       T                           Œ      T�       S��      ��       S4�      >�       SC�      j�       S��      ��       S��      ��       S[�      ��       S                           Œ      T�       V��      ��       V4�      >�       VC�      j�       V��      ��       V��      ��       V[�      ��       V                             Œ      �       v �      T�       ��~��      ��       v 4�      >�       v C�      j�       ��~��      ��       ��~��      ��       ��~[�      ��       ��~                               Œ      �       0��       �       P �      T�       \��      ��       0�4�      >�       0�C�      `�       0���      ��       0���      ��       0�[�      ��       \                           �      ��       ]��      T�       }|���      ��       ]C�      M�       }|���      ��       ]��      ��       ][�      ��       }|�                            <�      q�       Pq�      T�       _C�      M�       _`�      j�       _��      ��       P��      ��       _[�      ��       _                	           Œ      ��       0���      ѕ       0�4�      j�       0���      ��       0���      Ә       0�[�      ��       0�                  �      "�       ]��      ��       ]                  �      "�       S��      ��       S                  �      "�       0���      ��       0�                   ��      Ǔ       ]C�      M�       ]                   ��      Ǔ       SC�      M�       S                  ��      Ǔ       0�C�      M�       0�                 ��      �       _                   ��       �       P �      �       \                   ��       �       U �      �       S                 [�      ��       \                 [�      ��       ��~                      Y�      ^�       T��      ɕ       ��>�      C�       } Ř      Ә       T                      Y�      t�       w ��      ɕ       w >�      C�       w Ř      Ә       w                             ��      m�       ��~ѕ      �       ��~j�      ��       ��~��      ��       ��~Ә      [�       ��~��      ��       ��~                      ��      m�       _ѕ      �       _j�      ��       _                                  ��      g�       ^ѕ      ݕ       ^�      R�       ^R�      �       ��~j�      u�       ^��      ��       ��~��      ��       ��~Ә      [�       ��~��      ��       ��~                                  ��      m�       Sѕ      ��       S��      �       �T�j�      ��       S��      ��       �T�Ә      ޘ       Sޘ      [�       �T���      ��       S��      ��       �T�                                  ��      ה       Vה      m�       ��~ѕ      o�       ��~o�      �       �U�j�      u�       ��~u�      ��       �U���      ��       �U�Ә      [�       �U���      ��       �U�                               ��      ה       v ה      m�       ��~ѕ      �       ��~j�      u�       ��~��      ��       ��~��      ��       ��~Ә      [�       ��~��      ��       ��~                                 ��      m�       0�ѕ      �       0��      B�       PB�      
�       _
�      �       0�j�      ��       0���      ��       _��      ��       _Ә      [�       _��      ��       _                                          ��      ה       0�ה      ?�       ]?�      O�       }�O�      m�       ]ѕ      �       ]�      ;�       }�;�      o�       0�o�      ��       \��      ԗ       |�ԗ      ��       \j�      u�       }���      ��       \Ә      �       |���      ��       \                             ;�      o�       1�o�      g�       ��~g�      ��       P��      �       ��~��      ��       ��~��      ��       ��~Ә      [�       ��~��      ��       ��~                  ٖ      �       P                                   ;�      o�       0�o�      g�       ^g�      ��       R��      �       ^��      ��       ^��      ��       ^Ә      ��       ^��      >�       R>�      S�       ^��      ��       ^��      ��       R                                  ��      ה       0�ה      m�       \ѕ      J�       \J�      �       ��j�      u�       \��      ��       ����      ��       ��Ә      [�       ����      ��       ��                                 ;�      o�       6�o�      b�       Vb�      k�       v�k�      s�       ]s�      y�       v�y�      �       v��      ��       v���      ��       Q��      ��       V��      ��       VӘ      �       V�      ��       P��      �       p��      M�       Q��      ��       V��      ��       P��      ��       p���      ��       Q                                 ;�      o�       2�o�      k�       ]k�      s�       t}�s�      �       ]��      ��       ]��      ��       ]Ә      ��       ]��      [�       S��      ��       ]��      ��       S                              ��      і       Pі      �       ��~�      ��       R��      ��      ( ��~20��~#������������������+( ���      ��       R��      ��       R��      ��      ( ��~20��~#������������������+( �                    
�      C�       Pѕ      �       P                  ה      ��       VW�      b�       V                  ה      ��       SW�      b�       S                 ה      ��       0�W�      b�       0�                      o�      ��       X��      ��       ��~ݗ      ��       X                   o�      ��       Sݗ      ��       S                  o�      ��       0�ݗ      ��       0�                   ��      ��       R��      ��      ( ��~20��~#������������������+( �                   ��      ��        q "���      ��       Q                 ��      ��       S                 ��      
�       _                 ��      
�       ��~                  m�      r�       ���      4�       ^                  m�      ��       w �      4�       w                                 P�      ��       U��      '�       ]'�      ,�       �U�,�      ^�       ]^�      c�       �U�c�      ��       ]��      ��       �U���      ��       U                                P�      s�       Ts�      #�       V#�      ,�       �T�,�      Z�       VZ�      c�       �T�c�      ~�       V~�      ��       �T���      ��       T                                P�      ��       Q��      )�       ^)�      ,�       �Q�,�      `�       ^`�      c�       �Q�c�      ��       ^��      ��       �Q���      ��       Q                                P�      ��       R��      !�       w !�      ,�       ��~,�      <�       w <�      c�       �R�c�      k�       w k�      ��       �R���      ��       R                      P�      ��       X��      ��       ��~��      ��       X                                P�      ��       Y��      %�       \%�      ,�       �Y�,�      \�       \\�      c�       �Y�c�      ��       \��      ��       �Y���      ��       Y                           ̣      �       0��      @�       P@�      D�       w k�      |�       w |�      ��       ��~��      ��       6�                     P�      ̣       0�̣      "�       S,�      Y�       Sc�      ��       0�                   P�      [�       u ��      ��       u                   P�      ̣      
 P@     �c�      k�      
 P@     �                  P�      ̣       �=  c�      k�       �=                      P�      ��       Q��      ̣       ^c�      k�       ^                    P�      s�       Ts�      ̣       Vc�      k�       V                    P�      ��       U��      ̣       ]c�      k�       ]                
      P�      ��       0���      ��       P��      ̣       Sc�      k�       S                ��      ģ       ^                ��      ģ       V                ��      ģ       S                 ,�      G�       S                 G�      Y�       S                    k�      ~�       V~�      ��       �T���      ��       0�                 ��      ��       u                       �             U             S             �U�                 �      �       u8                  �             T                      ��      �       U�      �       �U��      ��       U                        ��      ͨ       Tͨ      �       ���      �       �T��      ��       T                        ��      ը       Qը      �       �@�      �       �Q��      ��       Q                        ��      ��       R��      �       P�      �       �R��      ��       R                        ��      Ũ       XŨ      �       R�      �       �X��      ��       X                      �      ;�       U;�      A�       �U�A�      N�       U                        �      '�       T'�      ;�       �H;�      A�       �T�A�      N�       T                      �      ;�       Q;�      A�       �Q�A�      N�       Q                      �      ;�       R;�      A�       �R�A�      N�       R                             |      R|       UR|      �|       _�|      �}       �U��}      �}       _�}      ~       �U�~      .~       _                         |      L|       TL|      �}       \�}      �}       �T��}      .~       \                     |      O|       QO|      .~       �Q�                     |      `|       R`|      .~       ��                         |      `|       X`|      �}       ]�}      �}       �X��}      .~       ]                     |      `|       Y`|      .~       ��                    ?|      �}       S�}      .~       S                    ;|      �}       V�}      .~       V                                 |      h|       0�h|      �|       P�|      }       ^}      �}       0��}      �}       P�}      �}       ^�}      �}       U�}      ~       ^~      ~       P~      .~       ^                            |      �|       0��|      �|       P�|      ^}       _q}      �}       0��}      �}       0��}      ~       _~      .~       0�                  �}      �}       P                 �|      �|       0�                    J}      U}       S�}      �}       S�}      ~       S                        J}      U}       ^�}      �}       P�}      �}       ^�}      ~       U~      ~       ^                  c}      q}       _)~      .~       0�                  c}      q}       S)~      .~       S                 q}      }       ^                 q}      }       S                  t      �       T                        �      �       R�      �       P�      �       R�      �       R                          �      �       U�      �        V�       �        U�       �        �U��       �        V                          �      �       T�      �        S�       �        T�       �        �T��       �        S                      �      �       Q�      E        ]E       �        �Q�                  �      7        \                 �      �       ]                 �      �       V                 �      �      
 p@     �                     �      �       s���      �       U�      �       s��                        !        V                        !        S                      7       S        s
 0.��S       ]        } 
 0.���       �        } 
 0.��                    7       ]        \�       �        \�       �        0�                    J       ]        ^�       �        ^                 J       T        \                 �       �        \                 �       �        ^                 x       |        T                 x       }        V                     �       �        S�       �        T�       �        �T�                     �       �        V�       �        U�       �        �U�                              )       U)      d       Vd      g       Ug      h       �U�                              *       T*      c       Sc      g       Tg      h       �T�                            *       Q*      f       \f      h       �Q�                  B      O       T                  B      T       V                     \      c       Sc      g       Tg      h       �T�                     \      d       Vd      g       Ug      h       �U�                          �O      �O       U�O      �O       S�O      �O       U�O      �O       �U��O      �O       U                      �O      �O       T�O      �O       �T��O      �O       T                          �O      �O       Q�O      �O       V�O      �O       Q�O      �O       �Q��O      �O       Q                     �O      �O       T�O      �O       �T��O      �O       T                   �O      �O       T�O      �O       �T�                 �O      �O       S                     �O      �O       0��O      �O       P�O      �O       T                 �O      �O       U                                      �E      �E       U�E      �G       \�G      �H       �U��H      I       UI      
K       \
K      K       UK      ]K       \]K      �K       �U��K      �L       \�L      �L       �U��L      �L       \                                        �E      �E       T�E      JG       ^JG      �H       �T��H      I       TI      #I       �T�#I      sJ       ^sJ      
K       �T�
K      K       TK      L       �T�L      �L       ^�L      �L       �T��L      �L       ^                                  �E      �E       Q�E      sF       VsF      �F       �Q��F      �F       V�F      �F       v :!��F      �F       p �Q�Q
  $0.( :!��F      �H       V�H      I       QI      
K       V
K      K       QK      �L       V                                            !G      JH       PfH      jH       PjH      oH       ��oH      �H       P�H      �H       P�H      �H       ��I      #I       P�I      �I       PJ      ?J       P@J      
K       PK      vK       P�K      L       P�L      �L       P�L      �L       ��                         �F      G       Q#I      wI       QL      -L       Q-L      �L       ���L      �L       ��                           �E      �H       S�H      �H       U�H      �H       S�H      �H       }�~�I      
K       SK      �L       S                     �F      G       q#I      wI       qL      -L       q                       �F      JG       _#I      oJ       _L      �L       _�L      �L       _                                     �E      �E       U�E      �G       \�G      �H       �U��H      I       UI      
K       \
K      K       UK      ]K       \]K      �K       �U��K      �L       \�L      �L       �U��L      �L       \                      )L      -L       P-L      �L       ���L      �L       ��                    UL      \L       0��L      �L       0�                 J      J       P                   �I      J       [J      2J       ��                 �I      J       ��                        �G      �G       r��G      �G       |�#�K      =K       r�=K      ]K       |�#�                   �G      �G       @�K      =K       @�                   �G      �G       UK      =K       U                       �G      �G       Q�G      �G       s� K      .K       Q.K      =K       s�                    �G      �G       1��G      �G       1�K      K       1�K      =K       	��                  �G      �G       QK      K       Q                  �G      �G       U�G      �G       u �K      =K       U                  �G      �G       @�K      =K       @�                      �G      �G       t 6%��G      �G       Q5K      8K       Q8K      =K       q �                    �G      �G       Q5K      8K       Q8K      =K       q �                   �G      �G       @�=K      ]K       @�                   �G      �G       T=K      ]K       T                       �G      �G       Q�G      �G       s� =K      NK       QNK      ]K       s�                     �G      �G       1��G      �G       1�=K      =K       1�=K      IK       	��IK      ]K       	��                  �G      �G       Q=K      =K       Q                  �G      �G       T�G      �G       t �=K      IK       TIK      ]K       t �                  �G      �G       @�=K      ]K       @�                      �G      �G       r 6%��G      �G       QUK      XK       QXK      ]K       q �                    �G      �G       QUK      XK       QXK      ]K       q �                      �G      oH       \]K      �K       \�L      �L       \                    FH      WH       U]K      �K       0��L      �L       0�                     �G      oH       S]K      �K       S�L      �L       S                   �G      H       QH      FH       s]K      ]K       s                    
H      "H       Q"H      FH      	 s#�#]K      ]K      	 s#�#                    H      =H       U=H      FH       qFH      FH       U]K      ]K       0�                     H      FH       0�]K      �K       0��L      �L       0�                     H      FH       R]K      vK       R�L      �L       R                       H      "H       Q"H      FH      	 s#�#]K      vK      	 s#�#�L      �L      	 s#�#                   "H      FH       Q]K      ]K       Q                     H      FH       0�]K      �K       0��L      �L       0�                    ,H      =H       UAH      FH       q                 fH      oH       \                 fH      oH       U                  �K      �K       X                  �K      �K       Y                  �K      �K       s��                     �K      �K       0��K      �K       R�K      �K       R                  �K      �K       Q                 �L      �L       \                   �L      �L       U�L      �L       ]                          �H      �H       t ?��H      �H       T�H      �H       v @&?��H      �H       T�H      �H       T                 �E      �F       S                   cJ      
K       Y�K      L       Y                   cJ      
K       S�K      L       S                   cJ      
K       s0��K      L       s0�                     �J      �J       r  "#?	���J      �J       Q�J      �J       r  "#?	��                     �J      �J       ��~ "#?	���J      �J       Q�J      �J       ��~ "#?	��                    �       !       T!      *!       �T�*!      Q!       T                   �       �        Q!      P!       Q                    �       !       P!      Q!       P                                 h       Uh      �       S�      �       T�      �       �U��      �       U                              5       q�5      h       u#�h      i       s#��      �       q�                          %      R       VR      S      	 u#�#S      �       V�      �       U�      �       V                        %      5       0�5      D       RG      L       RS      \       R�      �       0�                         %      5       R5      D       rG      G       RG      L       rS      \       r�      �       R                     r      �       S�      �       T�      �       �U�                   r      �       V�      �       U                              pz      �z       U�z      �z       S�z      �z       �U��z      �{       S�{      �{       �U��{      �{       U�{      |       S                              pz      �z       T�z      �z       V�z      �z       �T��z      �{       V�{      �{       �T��{      �{       T�{      |       V                 �z      �z       P                 �z      �z       p                      �z      �z       ]�z      �{       ]�{      |       ]                              pz      �z       0��z      �z       P�z      �z       \�z      �{       \�{      �{       �T�{      �{       0��{      �{       \�{      �{       0��{      |       \                   �z      U{       \�{      �{       \�{      |       \                    �z      U{       _�{      �{       _�{      |       _                      
{      {       P{      U{       w �{      �{       w �{      |       w                    
{      U{       ^�{      �{       ^�{      |       ^                           
{      !{       0�!{      4{       P4{      <{       X�{      �{       X�{      �{       ���{      |       ��                  �{      �{       ���{      �{       ��                    �{      �{       U�{      �{       ^�{      �{       ^                    �{      �{       0��{      �{       P�{      �{       P                 �{      �{       \                 �{      �{       ]                        �      �       U�      ,       S,      0       �U�0      M       S                    �      -       V0      M       V                 �      �       v                    �      /       \0      M       \                              s�                               \                  3      <       U                        �y      &z       U&z      Tz       STz      Xz       �U�Xz      hz       S                        �y      z       Tz      Wz       \Wz      Xz       �T�Xz      hz       T                    z      Uz       VXz      hz       V                  z      (z       T                  z      )z       V                      �      �       U�      �       S�      �       �U�                      �      �       T�      �       V�      �       �U#�                        P      b       Ub      ~       S~      �       �U��      �       S                              P      �       T�      y       \y      �       �T��      �       T�      �       \�      �       T�      �       \                            P      �       Q�      �       �Q��      �       Q�      �       �Q��      �       Q�      �       �Q�                              b      �       U�      ~       s��~      �       �U#���      �       U�      �       s���      �       U�      �       s��                     b      ~       s��~      �       �U#���      �       s��                           �      y       U�      �       U�      �       5��      -       6�-      �       1��      �       U�      �       1�                     b      �       0��      �       V�      �       0�                   b      �       0��      �       0�                             y       Z�      �       Z�      �       Z                      $      y       Y�      �       Y�      �       Y                      (      y       P�      �       P�      �       P                      ,      y       Q�      �       Q�      �       Q                      F      y       R�      �       R�      �       R                   �      �       W�      �       W                     �      �       U�      �       U�      �       s��                         u      ;u       U;u      v       �U�v      Fv       UFv      Zv       �U�                             u      8u       T8u      �u       S�u      �u       �T��u      v       Sv      Fv       TFv      Zv       S                             u      3u       Q3u      �u       \�u      �u       �Q��u      v       \v      Fv       QFv      Zv       \                     .u      �u       ^�u      v       ^Fv      Zv       ^                                u      Hu       0�Hu      Su       PSu      �u       V�u      �u       V�u      �u       0��u      v       Vv      	v       Tv      Fv       0�Fv      Zv       V                 [u      �u       P                 [u      �u       s                 [u      �u       V                 �u      �u       V                 �u      �u       ^                     �u      �u       V v      v       Vv      	v       T                   �u      �u       ^ v      v       ^                    �              U              �U�                      �      �       T�              u�               �T�                   �              U              �U�                        `      y       Uy      �       S�      �       �U��      �       U                            `      �       T�      �       V�      �       �T��      �       V�      �       �T��      �       T                     `      �       0��      �       P�      �       0�                     `      y       Uy      �       S�      �       U                    0      :       U:      S       �U�                    0      :       T:      S       �T�                   0      :       U��:      S       �U���                    6      :       T:      S       �T�                  ;      E       P                                  U      !       �U�                                  T      !       �T�                                 U�      !       �U��                                 T      !       �T�                  	             P                    `�      f�       Uf�      g�       �U�                    `�      f�       Tf�      g�       �T�                    `�      f�       Qf�      g�       �Q�                    `�      f�       Rf�      g�       �R�                    P�      T�       UT�      U�       �U�                    P�      T�       TT�      U�       �T�                    P�      T�       QT�      U�       �Q�                    P�      T�       RT�      U�       �R�                     �      1�       UK�      U�       \}�      ��       \                                �      �       T�      K�       ]K�      \�       �T�\�      ��       ]��      ��       �T���      �       ]�      G�       �T�G�      N�       ]                        �      1�       Q1�      R�       SR�      \�       �Q�\�      N�       S                        �      1�       R1�      Y�       ^Y�      \�       �R�\�      N�       ^                          @�      K�       P\�      q�       Pr�      ��       P��      ��        ��      ��                                =�      @�       P@�      K�       _\�      ��       _��      ��       _                 ;�      G�       P                   ��      /�       ^G�      N�       ^                   ��      /�       SG�      N�       S                    ��      /�       _G�      N�       _                      ߍ      �       _�      !�       \G�      N�       _                  �      �       P                    ߍ      �       0�G�      N�       0�                   ��      �       \G�      N�       \                  �      ;�       _G�      N�       _                  �      ;�       ^G�      N�       ^                        �      �       U�      �       ]�      �       �U��      �       U                        �      �       T�      �       V�      �       �T��      �       T                    �      �       P�      �       u                  �      �       S                 �      �       0�                  �      �       T                  �      �       V                 �      �       }                  �      �       V                      ��      �       U�      5�       S5�      6�       �U�                      ��      ��       T��      '�       U'�      6�       �T�                     �      ��       T��      '�       U'�      ,�       �T�                 �      ,�       1�                   �      �       U�      ,�       S                       �      
�       U
�      U�       SU�      V�       �U�                       �      �       T�      G�       UG�      V�       �T�                     
�      �       T�      G�       UG�      L�       �T�                 �      L�       0�                   �      
�       U
�      L�       S                      �       �        T�              V             �T�                   �       �        0��       �        P                  �       
       \                    �              S             P                    �      �       U�             �U�                    �      �       T�             �T�                      C       j        Qj       n        Rn       �        u � $ &�                              F       S        PS       V        q ��V       c        Pc       j        q �5$q 	�$"q ��j       n        r �5$r 	�$"r ��n       t        u ��Ou � $ &	�$"�t       �        R                         1        T                                    0�       +        P+       1        0�                        ��      �       U�      ��       S��       �       �U� �      Q�       S                        ��      �       T�      ��       \��       �       �T� �      Q�       \                        �      �       P �      �       P�      &�       R&�      Q�       ��                       ކ      �       _ �      ��       _��      �       _�      "�       V                   ކ      ��       ] �      Q�       ]                 
�      Q�       s�                 
�      Q�       |�                   z�      ��       Sȇ      �       S'�      Q�       S                   z�      ��       s�ȇ      �       s�'�      Q�       s�                   z�      ��       s� �ȇ      �       s� �'�      Q�       s� �                 %      t       u�                 %      t       u� �                    1      T      	 p 0$0&�T      Z       u� �0$0&�                 1      s      	 r 0$0&�                 D      Z       0�                 �             u� �                 �              U                 �             u�                 �             u� �                               U                               u�                               u� �                          `�      ��       U��      ��       �U���      ��       U��      ވ       Vވ      ߈       �U�                    `�      �       T�      ߈       �T�                    u�      ��       Z��      ��       Z                          �      ��       T��      ��       T��      ݈       S݈      ވ       vވ      ߈       �U#                   �      ��       Q��      ��       Q                         }�      ��       u���      ��       �U#���      ��       u���      ވ       v�ވ      ߈       �U#�                         }�      ��       u� ���      ��       �U#`���      ��       u� ���      ވ       v� �ވ      ߈       �U#`�                   ƈ      ވ       Vވ      ߈       �U�                   ƈ      ވ       v�ވ      ߈       �U#�                   ƈ      ވ       v� �ވ      ߈       �U#`�                                ��      τ       Uτ      Ԅ       SԄ      ބ       �U�ބ      -�       S-�      7�       �U�7�      J�       SJ�      T�       �U�T�      ��       S                    ��      ��       T��      ��       �T�                            ��      ��       Q��      Ą       \Ą      ބ       �Q�ބ      x�       \x�      e�       �Q�e�      ��       \                        ��      ل       ]ބ      2�       ]7�      O�       ]T�      ��       ]                               ��      τ       u�τ      Ԅ       s�Ԅ      ބ       �U#�ބ      -�       s�-�      7�       �U#�7�      J�       s�J�      T�       �U#�T�      ��       s�                               ��      τ       u� �τ      Ԅ       s� �Ԅ      ބ       �U#`�ބ      -�       s� �-�      7�       �U#`�7�      J�       s� �J�      T�       �U#`�T�      ��       s� �                        ��      τ       0�ބ      a�       0�a�      ��       1�Ņ      �       1�T�      e�       1�e�      ��       0�                                  ��      Ą       TĄ      ׄ       \ބ      �       T�      x�       Vx�      ��       \��      ��       |}���      �       \T�      e�       \e�      ��       V                           ��      ��       _��      τ       Qބ      p�       _p�      ��       QT�      e�       Qe�      ��       _                 ΅      �       S                 ΅      �       s�                 ΅      �       s� �                      ��      �       U�      �       S�      ��       �U�                 ��      �       u                 a�      z�       S                a�      z�       s�                a�      z�       s� �                      p      �       U�      N       SN      P       �U�                  �      O       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                 (      I       S                   (      N       s�N      P       �U#�                   (      N       s� �N      P       �U#`�                            P      b       Ub      e       �U�e      �       U�      �       �U?&�U'�U?&��             U             �U?&�U'�U?&�                              P      o       To      r       �T�r             T      �      
 �Ty 'y ��      �       �T?&�T'�T?&��             T            
 �Ty 'y �                            P      �       Q�      �       �Q��      �       Q�      �       �Q?&�Q'�Q?&��             Q             �Q?&�Q'�Q?&�                            P      �       R�      �       �R��      �       R�      �      
 �Ru 'u ��             R            
 �Ru 'u �                        W      �       P�      �       �U�Q"��      �       Y�             P                      [      �       X�      �       �T�R"��             X                      �      �       T�      �       T             T                  �      �       R                  �      �       P                    0      :       T:      J       �T�                    0      4       R4      J       �R�                    =      G       RG      J      
 �Ru t �                     C      �       R�      �       Y�      �       R                      G      �       Q�             P�      �       Q                  �      Z       R                         8       x x t t " ��8      W       q @<$�                      P      Y       RY      �       Y�             Y                        R      s       Qs             P�      �       P�             P                        |       X                          �       T      -       T                                  �      �       Q�      �       X�      �       Q�      �       P�      �       P�      �       Q�             X             Q      -       P                     G      Y       1�Y      _       	��_      �       Z�      -       Z                   G      s       1�s      �       [�      -       [                      �      �       S�      �       \�      *       \                        �      �       U�      %       S%      -       �U�-      1       U                      �      �       T�      -       [-      1       T                      �      �       Q�      -       �Q�-      1       Q                                    | p "�      (       \(      -       �U                                    v p "�       &       V&      -       �U#                       �      �       q @$��      �       Q�      -       Z-      1       q @$�                        �      �       U�      )       S)      �       �U��      �       U                      �      �       T�      �       [�      �       T                      �      �       Q�      �       �Q��      �       Q                  �      �      	 w ��"�                  	             v ��"�                  <      J      	 ���@"�                      `      v       ~ p "�v      �       ^�      �       {                       �      �       q @$��      �       Q�      �       Z�      �       q @$�                                 r z �      h       R                         n      �       T�             T6      h       T�      �       T�      �       T*      X       T                                   n      {       X{      �       u�             X             u6      C       XC      }       u�      �       u�      �       X�             u*      4       X4      h       u                 �      �       X                 �      �       T                �      �       X                �      �       T                   �      �       R�      �      
 r { "#���                  �      �       r ?&��      �       [                �      �       Y                �      �       Q                �      �       Y                �      �       Q                  �      �       P�      �      
 p z "#���                  �      �       p ?&��      �       Z                          5       R�      �       R�      �       R      *       R                              &       Q&      5       u�      �       Q�      �       u�      �       u      *       u                          5       1��      �       1��      �       	���      �       	���      �       1�             1�      *       	��                                &       Q&      5       u�      �       Q�      �       q ��      �       Q�      �       u��      �       u�      *       u                             5       R�      �       R�      �       R�      �       r �             R             r �      *       Z                              5      ;       q { "�-r �-� �;      E       u@${ "�-r �-� ��      �       P�      �       u�      �       q { "�-r �-� ��      �       u@${ "�-r �-� �%      *       P                 5      5       q { "�-r �-� ��      �       P�      �       q { "�-r �-� �%      *       P                   E      g       R�      �       R      2       R�      �       R                           E      R       YR      g       u�      �       Y�      �       u      $       Y$      2       u�      �       Y�      �       u                   E      g       1��      �       1��      �       	���      �       1�             1�      2       	���      �       1��      �       	��                            E      R       YR      g       u�      �       Y�      �       y ��      �       u�             Y      $       y �$      2       u��      �       Y�      �       y ��      �       u�                    E      N       R      2       R�      �       r �                g      g       P�      �       Y                     n      �       R�             R6      U       R�      �       R*      H       R                               n      {       X{      �       u�             X             u6      C       XC      U       u�      �       X�      �       u*      4       X4      H       u                     n      �       1��             1�             	��6      U       1��      �       1��      �       	��*      *       1�*      H       	��H      H       1�                                 n      {       X{      �       u�             X             x �             u�6      C       XC      U       u�      �       X�      �       x ��      �       u�*      *       X*      4       x �4      H       u�                �      �       PH      H       P                       �      �       R[      y       R�      �       R�             RK      h       R                       �      �       T[      h       T�      �       T�      �       TK      X       T                       �      �       1�[      v       1��      �       1��      �       	���      �       1��             	��K      T       1�T      h       	��                       �      �       T[      h       T�      �       T�      �       t ��      �       T�      �       t �K      T       TT      X       t �                      P      .       U.      �       �U��      �       U                     �      �      $ s  "#��@& $ &{ ~ "#��@& $ &"��      �       s @& $ &{ ~ "#��@& $ &"��      �       s @& $ &{ @& $ &"�                     ?      R      $ s x "#��@& $ &r u "#��@& $ &"�R      Z       x @& $ &r u "#��@& $ &"�Z      g       x @& $ &r @& $ &"�                 b      k       t                  b      k       u                    b      k       t k      �       X                 b      k       u                    �      �       S�      �      
 s  "#���                  �      �       s ?&��      �       _                �      �       t                �      �       u                �      �       t                �      �       u                  �      �       [�      �      
 { ~ "#���                  �      �       { ?&��      �       ^                �      �       t                �      �       t                �      �       t                �      �       u                �      �       t                �      �       u                �      �       Y�      �      
 p y "#���                �      �       P                �      �       u                �      �       t                 �      �       u                �      �       X�      �       x w "#���                �      �       x ?&�                ?      ?       t                ?      ?       �U#                ?      ?       t                ?      ?       �U#                �      ?       t                  �      .       u.      ?       �U#                !�      ?       t                !  �      .       u.      ?       �U#                         ?       R?      ?      
 r u "#���                        ?       r ?&�?      ?       U                ?      J       t                ?      J       �U#                ?      J       t                ?      J       �U#                  ?      J       PJ      J      
 p v "#���                  ?      J       p ?&�J      J       V                      �      �       U�      �       u ��      �       �U�                      �      �       T�      �       Y�      �       t ��      �       �T�                      �      �       Q�      �       X�      �       q ��      �       �Q�                       �      �       1��      �       	���      �       R�      �       r ��      �       R�      �       r ��      �       R                 �      �       U                      �      �       T�      �       Y�      �       T                        �      �       Q�      �       X�      �       Q�      �       X                    �      �       P�      �       q �                   �      �       P�      �       q �                      �o      �o       U�o      p       u p      
p       �U�                    �o      p       Tp      
p       �T�                                    �N      �N       U�N      O       SO      O       �U�O      8O       S8O      AO       UAO      BO       �U�BO      NO       UNO      gO       SgO      vO       �U�vO      �O       U                                      �N      �N       T�N      O       ]O      O       �T�O      #O       T#O      =O       ]=O      AO       TAO      BO       �T�BO      NO       TNO      qO       ]qO      vO       �T�vO      �O       T                                        �N      �N       Q�N      O       VO      O       �Q�O      O       QO      9O       V9O      AO       RAO      BO       �Q�BO      NO       QNO      mO       VmO      uO       RuO      vO       �Q�vO      �O       Q                                        �N      �N       R�N      O       \O      O       �R�O      #O       R#O      ;O       \;O      AO       XAO      BO       �R�BO      NO       RNO      oO       \oO      uO       TuO      vO       �R�vO      �O       R                    �N      �N       PO      #O       P                    �N      O       PNO      uO       P                     NO      gO       SgO      uO       u�~�uO      vO       �U�                     NO      mO       VmO      uO       RuO      vO       �Q�                 NO      vO       1�                     NO      oO       \oO      uO       TuO      vO       �R�                             M       QM      P       q���}�P      �       Q�      �       q�����      �       Q                    n      �       R�      �       R                                        #      6       R6      C       PC      F       RF      P       r �P      _       P_      w       Sz      �       S�      �       S�      �       u �      �       R�      �       S�      �       R�      �       P�      �       S�      �       R                                &      6       P6      C       [C      P       PP      S       RS      �       [�      �       P�      �       p ��      �       R�      �       P                               6      C       PC      _       Pw      �       S�      �       S�      �       u �      �       S�      �       P�      �       S                    n      �       X�      �       X                        n      t       p 3$ 0H     "�t      z       p3$ 0H     "�z      �       p3$0H     "��      �       p 3$ 0H     "��      �       p3$ 0H     "��      �       p3$0H     "�                                 :      ^       Sa      �       S�      �       sx��      �       S�      �       t �      �       ���}��      �       S�      �       S�      �       t                     :      P       Ra      �       R                                                  [       +       Q:      :       [:      G       { z "�G      ^       [a      t       [t      {       { z �{      �       [�      �       P�      �       [�      �       p ��      �       P�      �       { ��      �       [                                  +       Q:      ^       Qa      �       Q�      �       P�      �       p ��      �       [�      �       P�      �       Q                        G      ^       [{      �       [�      �       P�      �       [                      :      ^       Xa      �       X�      �       X                        :      D       p 3$ 0H     "�D      J       p3$ 0H     "�J      V       p3$0H     "�a      x       p 3$ 0H     "�x      ~       p3$ 0H     "�~      �       p3$0H     "�                              :       Y:      @       u D      R       YR      X       u                               =       X=      @       t D      U       XU      X       t                       +      5       Oq �5      D       q~�D      O       Oq �O      [       R[      \       P                            `      �       U�      M       �U�M      V       UV      y       �U�y      �       U�      �       �U�                                    `      �       T�              S       .       �T�.      C       SC      M       �T�M      V       TV      n       Sn      y       �T�y      �       T�      �       S                                        `      �       Q�      &       \&      -       T-      .       �Q�.      F       \F      M       �Q�M      V       QV      q       \q      x       Tx      y       �Q�y      �       Q�      �       \                                        `      �       R�      (       ](      -       Q-      .       �R�.      H       ]H      M       �R�M      V       RV      s       ]s      x       Qx      y       �R�y      �       R�      �       ]                            `      �       X�      M       �X�M      V       XV      y       �X�y      �       X�      �       �X�                            `      �       Y�      M       �Y�M      V       YV      y       �Y�y      �       Y�      �       �Y�                  �      �       ��                        �      ,       _.      L       _V      w       _�      �       _                                    �      �       R�      (       ](      -       Q-      .       �R�.      H       ]H      M       �R�V      s       ]s      x       Qx      y       �R��      �       ]                                    �      �       Q�      &       \&      -       T-      .       �Q�.      F       \F      M       �Q�V      q       \q      x       Tx      y       �Q��      �       \                                �      �       T�              S       .       �T�.      C       SC      M       �T�V      n       Sn      y       �T��      �       S                        �      �       U�      M       �U�V      y       �U��      �       �U�                       �      *       ^.      J       ^V      u       ^�      �       ^                        �      $       V.      D       VV      o       V�      �       V                    �             P.      4       P                                P.      4       P                            -       p 0)�4      9       p 0)�V      x       p 0)�                      �      �       T�      /       �T�/      6       T                      �      �       Q�      /       �Q�/      6       Q                      �      �       R�      /       �R�/      6       R                  �      /       U                 �      �       0�                     �      �       @��             @�      /       @�                     �      �       U�             U      /       U                           �      �       P�      �       t �      �       tx�      �       P�             t       /       t                      �      �       1��      �       1��      �       1��             	��             1�      /       	��                        �      �       P�      �       t �      �       P�      �       p ��             t �      /       t                    �      �       U�      �       u ��             U             U      /       u �                    �      �       @��             @�      /       @�                           �      �       p 6%��      �       p 6%��      �       P             P             p �-      /       P                   �      �       P             P-      /       P                        @      �       U�      %       �U�%      1       U1      D       �U�                    @      �       T�      D       �T�                    @      \       Q\      D       Z                          �      �       0��      �       u��             U             u�1      D       U                      x      �       Y�      �       y 	���      D       Y                        �      �       X�      �       x`��      /       X1      D       X                       �      �       tP��             tp�             tP�1      D       tp�                        P      f       Uf      �       �U��      �       U�      �       �U�                   m      �       U�      �       R                   m      �       R�      �       R                     m      |       U|      �       Y�      �       R                     m      |       R|      �       X�      �       R                  _      �       P                  m      �       Z                      �      �       Q�      �       p �      �       pp                  �      �       Q                    �      7	       T7	      l	       �T�                         ?	      O	      $ x z "#��@& $ &r t "#��@& $ &"�O	      S	       p @& $ &r t "#��@& $ &"�S	      ^	      $ x z "#��@& $ &r t "#��@& $ &"�^	      b	       x z "#��@& $ &p @& $ &"�b	      l	      $ x z "#��@& $ &r t "#��@& $ &"�                 �      �       t                  �      �       u                  �      �       t                    �      �       u �      	       R                   �      
	       P
	      
	      
 p s "#���                  �      
	       p ?&�
	      
	       S                
	      	       t                
	      	       u                
	      	       t                
	      	       u                  
	      	       Y	      	      
 y { "#���                  
	      	       y ?&�	      	       [                	      )	       t                	      )	       t                  	      )	       X)	      )	      
 x z "#���                	  	      )	       x ?&�)	      )	       Z                  )	      7	       t7	      ?	       �T#                )	      ?	       u                  )	      7	       t7	      ?	       �T#                )	      ?	       u                  )	      ?	       R?	      ?	      
 r t "#���                  )	      ?	       r ?&�?	      ?	       T                    p	      �	       U�	      �	       �U�                      p	      �	       T�	      �	       \�	      �	       �T�                  }	      �	       S                  �	      �	       V                 �	      �	       \                 �	      �	       S                        �	      �	       U�	      M
       [M
             �U�      %       [                    
      
       y p �
             Z                    ,
      /
       y p �/
             Y                     3
             V             }p�             �U#                           s
      y
       T��y
      �
       T�^��
      �
       �^��
      �
       Q�R��
             T�^�             T��                    �
      �
       Q���
      �
       Q�R�                 3
      S
       0�                 y
      �
       Q                     3
      S
       0�S
      �
       Q�
             Q                     3
      S
       0�S
      �
       U�
             U                  �	      �	       W                    �	      �	       U�	      �	       [                    b
             S             q�                      0      8       T8      K       QK      l       �T�                      p      �       U�      	       \	             �U�                      p      �       T�             ^             �T�                   p      �       0��      �       S                  �      �       V                �      �       V                 �      �       v                 �      �       v                  �      �       _                 �      �       V                 �      �       _                 �      �       |�                  �      �       ^                        8       P                  C      m       P                  G      m       Q                      p      �       U�      �       _�      �       �U�                      p      �       T�      �       ]�      �       �T�                      p      �       Q�      �       V�      �       �Q�                      p      �       R�      �       ^�      �       �R�                     �      �       S�      �       T�      �       0��      �       S                  �      �       \                 �      �       s                   �      �       S�      �       T                 �      �       V                             3       U3      8       u �8      |       �U�                             @       T@      E       YE      E       t �E      |       �T�                             M       QM      R       XR      R       q �R      |       �Q�                              3       1�3      8       	��8      B       RB      E       r �E      O       RO      R       r �R      |       R                        `       U                      #      @       T@      E       YE      |       T                          &      M       QM      R       XR      e       Qe      h       Ph      |       X                    n      {       P{      |       q �                   n      {       P{      |       q �                    �      �       U�              �U�                    �      �       T�              �T�                  �      �       T�      �       �T�                �      �       U                   �      �       T�      �      
 p t "#���                  �      �       t ?&��      �       P                                    U             u �      P       �U�                                   1�             	��      "       X"      %       x �%      P       X                        6       U                          %       T%      P       R                    A      O       PO      P       q �                   A      O       PO      P       q �                        d       u�                        d       u� �                        P      `       U`      p       Sp      r       Tr      s       �U�                    \      q       Vq      r       U                     a      p       Sp      r       Tr      s       �U�                   a      q       Vq      r       U                      �      �       U�      �       �U��      �       U                                    ,       U,      =       S=      A       TA      B       �U�B      I       SI      M       �U�M      Q       U                                  ,       T,      >       V>      B       �T�B      J       VJ      M       �T�M      Q       T                      &      @       \@      A       UB      L       \                   &      ,       U,      -       S                     1      =       S=      A       TA      B       �U�                   1      @       \@      A       U                        `      �       U�      �       S�      �       �U��      �       U                         �       u#��      �       s#�                       �       T                         �       u#��      �       s#�                    �      �       S�      �       �U�                      0#      C#       UC#      D#       �U�D#      V#       U                      0#      C#       TC#      D#       �T�D#      V#       T                      0#      C#       QC#      D#       �Q�D#      V#       Q                      )      E)       UE)      G)       �U�G)      �)       U                        )      F)       TF)      G)       �T�G)      x)       Tx)      �)       �T�                        $)      F)       TF)      G)       �T�f)      x)       Tx)      �)       �T�                      $)      E)       UE)      G)       �U�f)      �)       U                     $)      E)       u�#E)      F)      	 �U#�#f)      x)       u�#                        �.      �.       U�.      �.       S�.      �.       �U��.      /       U                      �.      �.       T�.      �.       �T��.      /       T                     �.      �.       0��.      �.       P�.      /       0�                 �.      �.       P                   6      ,6       Ti6      l6       T                   !6      Y6       VZ6      h6       V                     !6      ,6       T,6      X6       SZ6      g6       S                    |8      �8       R�8      �8       R                      �8      �8       P�8      �8       r�8      �8       P�8      �8       P                         ;      (;       U(;      ;       V;      �;       �U��;      �;       U                         ;      (;       T(;      �;       \�;      �;       �T��;      �;       T                           ;      (;       Q(;      �;       �Q��;      �;       Q�;      �;       �Q��;      �;       Q                      ;      );       0�);      ;;       P�;      �;       0�                  7;      y;       �Q�                  7;      y;       \                  7;      y;       V                     F;      i;       0�i;      n;       Pn;      y;       0�                    ;;      B;       PB;      K;       v                  ?;      y;       S                  F;      y;       ]                                    �L      pM       UpM      �M       \�M      N       UN      N       �U�N      (N       \(N      /N       �U�/N      gN       UgN      �N       \�N      �N       u�~��N      �N       �U�                                      �L      mM       TmM      �M       S�M      �M       �T��M      N       SN      N       �T�N      N       SN      /N       �T�/N      GN       SGN      gN       TgN      ~N       S~N      �N       �T�                                        �L      "M       Q"M      �M       _�M      �M       �Q��M      N       _N      N       �Q�N      N       _N      /N       �Q�/N      GN       _GN      gN       QgN      �N       _�N      �N       Q�N      �N       �Q�                                        �L      M       RM      �M       ]�M      �M       �R��M      N       ]N      N       �R�N      N       ]N      /N       �R�/N      GN       ]GN      gN       RgN      �N       ]�N      �N       R�N      �N       �R�                                        �L      eM       XeM      �M       V�M      �M       �X��M      N       VN      N       �X�N      N       VN      /N       �X�/N      GN       VGN      VN       XVN      �N       V�N      �N       T�N      �N       �X�                         M      (M       P(M      pM       u pM      qM       | �M      N       u /N      GN       u                                 M      N       ^N      ,N       ^,N      /N       �T�Q"�/N      GN       ^gN      �N       ^�N      �N       �T "��N      �N       �Tq "��N      �N       �T�Q"�                                AM      eM       XeM      �M       V�M      �M       �X�N      N       V/N      GN       VgN      �N       V�N      �N       T�N      �N       �X�                            AM      �M       ]N      N       ]/N      GN       ]gN      �N       ]�N      �N       R�N      �N       �R�                              AM      �M       _�M      �M       �Q�N      N       _/N      GN       _gN      �N       _�N      �N       Q�N      �N       �Q�                              AM      mM       TmM      �M       S�M      �M       �T�N      N       S/N      GN       SgN      ~N       S~N      �N       �T�                              AM      pM       UpM      �M       \N      N       \/N      GN       UgN      �N       \�N      �N       u�~��N      �N       �U�                           rM      �M       P�M      �M       0��M      �M       0��M      �M       PN      N       PgN      �N       P                    SM      qM       P/N      GN       P                     �M      �M       0��M      �M       1��M      �M       0�                  �M      �M       _                       N      N       \gN      �N       \�N      �N       u�~��N      �N       �U�                       N      N       ]gN      �N       ]�N      �N       R�N      �N       �R�                       N      N       _gN      �N       _�N      �N       Q�N      �N       �Q�                       N      N       VgN      �N       V�N      �N       T�N      �N       �X�                      pQ      ~Q       U~Q      Q       �U�Q      �Q       U                    �Q      �Q       U�Q      �Q       �U�                     �Q      �Q       0��Q      �Q       R�Q      �Q       R                  �Q      �Q       P                      �S      �S       T�S      �S       �T��S      �S       T                      �S      �S       U�S      �S       �U��S      �S       U                      �S      �S       T�S      �S       �T��S      �S       T                      X       X       U X      !X       �U�!X      +X       U                      �\      �\       U�\      �\       �U��\      �\       U                          �\      
]       U
]      ]       S]      ]       �U�]      0]       S0]      2]       �U�                            �\      
]       T
]      ]       V]      ]       �U#]      &]       T&]      1]       V1]      2]       �T�                              @]      f]       Uf]      x]       Vx]      y]       �U�y]      �]       U�]      �]       V�]      �]       �U��]      �]       U                          @]      e]       Te]      y]       �T�y]      �]       T�]      �]       �T��]      �]       T                        Y]      w]       Sw]      x]       vx]      y]       �U#y]      �]       S                            Y]      f]       Uf]      x]       Vx]      y]       �U�y]      �]       U�]      �]       V�]      �]       �U�                 Y]      �]       0�                    0^      >^       U>^      ?^       �U�                      0^      :^       T:^      >^       Q>^      ?^       �T�                      0^      6^       Q6^      >^       R>^      ?^       �Q�                      ``      z`       Uz`      �`       S�`      �`       �U�                   k`      z`       u8z`      |`       P                  n`      |`       T                    n`      z`       u8z`      |`       P                            pg      �g       U�g      �g       S�g      �g       �U��g      �h       S�h      �h       �U��h      �h       S                          pg      �g       T�g      �g       V�g      �g       �T��g      �g       V�g      �h       �T�                            pg      �g       Q�g      �g       \�g      �g       �Q��g      �h       \�h      �h       �Q��h      �h       \                 pg      �h       �{n  �                 pg      �h       �an  �                    �g      �g       P�g      �g       P                   pg      �g       0��g      �g       0�                      h      h       Ph      h       ^�h      �h       ^                      h      h       0�h      h       ]�h      �h       ]                    Wh      lh       P�h      �h       P                  �h      �h       V                     pg      �g       0��g      h       0��h      �h       0�                   �g      �g       @��h      �h       @�                   �g      �g       S�h      �h       S                    �g      h       V�h      �h       V                      �g      �h       S�h      �h       �U��h      �h       S                   h      5h       8�hh      h       8�                   h      5h       Shh      h       S                   h      =h       Vph      h       V                   h      =h       Sph      h       S                  h      =h       0�ph      h       0�                     i      #i       U#i      Fi       �U�                         i      7i       T7i      ;i       U;i      <i       �T�<i      Fi       T                       i      2i       Q2i      <i       �Q�<i      Fi       Q                       i      ;i       R;i      <i       �R�<i      Fi       R                       i      ;i       X;i      <i       �X�<i      Fi       X                      �m      �m       T�m      �m       �T��m      �m       T                      �q      �q       U�q      �q       S�q      �q       �U�                      �q      �q       T�q      �q       V�q      �q       �T�                   �q      �q       0��q      �q       P                      P�      [�       U[�      k�       �U�k�      ��       U                      P�      [�       T[�      k�       �T�k�      ��       T                        P�      [�       Q[�      j�       Sj�      k�       �Q�k�      ��       Q                       P�      g�       0�g�      k�       Rk�      }�       0�}�      ��       R                       P�      \�       0�\�      k�       Pk�      }�       0�}�      ��       P                          ��      F�       UF�      ��       V��      ��       �U���      ��       U��      �       V                          ��      %�       T%�      ��       ^��      ��       �T���      ��       T��      �       ^                          ��      .�       Q.�      ��       \��      ��       �Q���      ��       Q��      �       \                          ��      9�       R9�      ��       S��      ��       �R���      ��       R��      �       S                     6�      9�       R9�      ��       S��      �       S                   2�      ��       \��      �       \                   2�      ��       ^��      �       ^                     2�      F�       UF�      ��       V��      �       V                                  ��      ��       U��      ��       ]��      N�       �U�N�      ʥ       ]ʥ      ��       ����      ڦ       �U�ڦ      �       ]�      '�       ��'�      :�       �U�:�      ��       ��                          ��      ڤ       Tڤ      �       U�      :�       _:�      ;�       �T�;�      ��       _                        ��      Ѥ       QѤ      1�       S1�      ;�       �Q
���Q�Q0+( �;�      ��       S                    ��      �       R�      ��       ��                 ��      ��       �c�  �                 ��      ��       �V�  �                      ʤ      ͤ       Pͤ      �       } �      ��       ��                	                    ޤ      ��       0�N�      ե       0�ե      �       ^h�      |�       P|�      ��       ^��      ��       ~���      ��       ^ڦ      �       0��      �       ^�      �       ~��      '�       ^:�      ~�       ^�      ��       ^                
                        ޤ      ��       0�N�      ե       0�ե      �       P}�      ��       P��      ��       pj���      ��       Pڦ      �       0��      �       P�      �       ph��      '�       P:�      L�       PL�      ��       [��      ��       ��C�      V�       [�      ��       P                        ޤ      �       P�      .�       w .�      ;�       ��;�      ��       w                           ޤ      ��       0�N�      ե       0���      ��       1�ڦ      �       0��      '�       0��      ��       1���      ��       0�                               ʤ      ��       0�;�      G�       0�N�      ��       0�ڦ      ѧ       0�ѧ      ԧ       Pԧ      C�       VC�      V�       0�V�      �       V�      ��       0�                          ޤ      �       �W�  ;�      G�       �W�  N�      ��       �W�  ڦ      '�       �W�  :�      H�       �W�  �      ��       �W�                            ޤ      �       �=�  ;�      G�       �=�  N�      ��       �=�  ڦ      '�       �=�  :�      H�       �=�  �      ��       �=�                            ޤ      �       �0�  ;�      G�       �0�  N�      ��       �0�  ڦ      '�       �0�  :�      H�       �0�  �      ��       �0�                            ޤ      �       S;�      G�       SN�      ��       Sڦ      '�       S:�      H�       S�      ��       S                            ޤ      �       U�      �       _;�      G�       _N�      ��       _ڦ      '�       _:�      H�       _�      ��       _                              d�      l�       Pl�      ե       \ե      ��       ��ڦ      �       \�      '�       ��:�      H�       ���      ��       ��                            ��      ե       	��ե      ��       ]�      '�       ]:�      E�       ]�      ��       ]��      ��       ]                                �      �       PN�      \�       Pե      �       \�      "�       P"�      ��       \�      '�       \:�      H�       \�      ��       \                          ��      ե       0�ե      ��       V�      '�       V:�      H�       V�      ��       V                   h�      ��       6�ڦ      �       6�                   h�      ��       _ڦ      �       _                      p�      ��       V��      ե       ڦ      �       V                    p�      ��       _ڦ      ��       _                   p�      ��       0�ڦ      ��       0�                    �      L�       4��      �       4�                    �      L�       _�      �       _                    &�      h�       ^�      �       ^                        ե      �       _&�      ��       _�      '�       _:�      ��       _                       ե      �       0�&�      ��       0��      '�       0�:�      ��       0�                   Ѥ      ڤ       Tڤ      ޤ       U                *�      *�       0�                  ��      *�       w ��      Ʀ       w                   ��      *�       _��      Ʀ       _                  ��      *�       0���      Ʀ       0�                   ~�      ��       ^C�      V�       ^                   ~�      ��       _C�      V�       _                  ~�      ��       0�C�      V�       0�                 �      ��       V                 �      ��       _                 V�      �       V                 V�      �       ��                      `�      g�       Ug�      h�       �U�h�      q�       U                      `�      g�       Tg�      h�       �T�h�      q�       T                    ��      ��       P��      ��       P                    =�      U�       Pg�      v�       P                     =�      J�       tJ�      f�       Qg�      v�       Q                  R�      f�       T                  R�      f�       U                      �      ��       U��      ��       �U���      �       U                      �      ��       T��      ��       �T���      �       T                      �      ��       Q��      ��       �Q���      �       Q                      �      ��       R��      ��       �R���      �       R                                    U       #        �U�                                 U                                0�                        �=      >       U>      <>       S<>      B>       �U�B>      �>       S                          �=      >       T>      >       Q>      ?>       \?>      B>       �T�B>      �>       \                  7>      7>       0��>      �>       P                   >      7>       VB>      �>       V                      �>      �>       V�>      �>       v~��>      �>       V                  �>      �>       ]                            �      �       T�      )       Y)      2       T2      �       Y�      �       T�      �       Y                           �             0�      (       P)      P       0�P      �       P�      �       0��      �       P                               �             0�             P      )       X)      P       0�P      p       Pp      �       X�      �       0��      �       X�      �       P�      �       X                        �      �       T�             t�5      5       T5      X       t�X      p       t��      �       t��      �       t��      �       [                        �              Z5      M       r 1$x "�M      `       Z`      �      
 r 1$u�	"��      �       Z                    06      :6       U:6      ?6       �U�                 �      �       U                        �      H       UH      �       S�      �       �U��      �       S                            �      �       T�      �       �T��      �       T�      q       �T�q      �       T�      �       �T�                    �      �       V�      �       V                     �      H       u� �H      �       s� ��      �       s� �                  5      H       u� H      L       s�                 5      L       v��0$0&�                   E      L       PL      L      
 p u "#���                  E      L       p ?&�L      L       U                d      w       s�                 d      w       v��0$0&�                   p      w       Pw      w      
 p u "#���                  p      w       p ?&�w      w       U                �      �       s�                    �      �       v��0$0&��      �      	 p 0$0&�                   �      �       P�      �      
 p r "#���                  �      �       p ?&��      �       R                �      �       s�                 �      �       v��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                      p       x        Ux       �        S�       �        �U�                     p       x        Ux       �        S�       �        �U�                 �      �       U                      �      �       U�      h        Sh       j        �U�                     �      �       U�      h        Sh       j        �U�                 �      �       u                   �      i        V                          @'      c'       Uc'      g'       Qg'      �(       V�(      �(       �U��(      )       V                    @'      `'       T`'      )       �T�                    V'      �(       \�(      )       \                    ]'      �(       S�(      )       S                    h'      )       P)      )       P                 �'      �'       Q                 �'      �'       R                 �'      �'       2�                 �'      �'       S                 �'      �'       3�                 �'      �'       S                 �(      �(       V                 �(      �(       S                     �(      �(       0��(      �(       1��(      �(       2�                 �(      )       0�                 �(      )       2�                 �(      )       S                 �(      )       s��                        @6      ~6       U~6      N7       SN7      T7       �U�T7      Y7       U                       @6      ~6       U~6      N7       SN7      T7       �U�T7      Y7       U                  d6      S7       ]                  k6      O7       V                  r6      �6       \                 �6      �6       S                 �6      �6       s�                 �6      �6       S                 �6      �6       \                 �6      �6       |8                         �      1�       U1�      l�       ^l�      ١       s�?�      G�       ^��      ��       s�                                   �      )�       T)�      �       S�      ��       �T���      ��       S��      ��       �T���      ��       S��      ��       �T���      ��       S��      ��       �T�                     �      5�       Q5�      ��       ��~                                   �      5�       R5�      �       \�      ��       �R���      ��       \��      ?�       �R�?�      G�       \G�      ��       �R���      ��       \��      ��       �R�                                   �      5�       X5�      �       ]�      ��       �X���      �       ]�      ?�       �X�?�      G�       ]G�      ��       �X���      ��       ]��      ��       �X�                                                             N�      i�       Pi�      l�       Vl�      w�       Pw�      ܡ       Vܡ      �       P��      �       P�      ?�       VG�      ��       V��      ��       ��~l�      ݣ       ��~E�      h�       Ph�      ��       V��      ��       0���      ��       0�դ      %�       V%�      M�       ��~v�      ~�       P~�      ��       P��      ��       V��      ��       P��      ��       ��~��      ��       V��      Ш       PШ      ��       V��      
�       P\�      q�       P��      ��       V                  �      �       t�#                              6�      K�       PK�      �       _��      ?�       _?�      G�       PG�      ��       _��      ��       _��      ��       _                                  �      )�       T)�      �       S�      ��       �T���      ��       S��      ��       �T���      ��       S��      ��       �T���      ��       S��      ��       �T�                        ܤ      �       T�      %�       ��~�@%���      ��       T��      ֨       ��~�@%�                           ��      ?�       SG�      ��       S��      ��       �T���      ��       �T���      ��       S��      ��       �T�                         G�      ��       S��      ݣ       �T�%�      M�       �T���      ��       �T���      ��       S                           ��      ڢ       0�l�      ��       0���      ݣ       V%�      ��       V�      M�       0���      ��       V                             v�      ��       0���      ��       ��~l�      ݣ       ��~%�      -�       ��~2�      M�       ��~��      ��       ��~��      ��       0�                           v�      ��       0���      ��       ��~l�      ݣ       ��~%�      H�       ��~��      ��       ��~��      ��       0�                             v�      ��       0���      ��       ��~l�      u�       ��~��      ݣ       ��~%�      M�       ��~��      ��       ��~��      ��       0�                             v�      ��       0���      �       ��~�      ��       Pl�      ݣ       ��~%�      M�       ��~��      ��       ��~��      ��       0�                 ��      ��       0�                  ��      ��       X                   %�      �       ��~��      ��       ��~                     %�      ��       S��      ��       ��~��      ��       S                              ^�      ��       ]��      ��       S��      ��       s���      ��       S��      ѥ       ��~ѥ      ܥ       P��      ��       ]                     ^�      r�       Pr�      �       ��~��      ��       ��~                    s�      ��       P��      ��       P                       ^�      ��       0���      ܥ       Vܥ      �       ]��      ��       0�                        ��      ܥ       3�ܥ      �       V�      ��       v���      �       V                       �      �       SM�      v�       S��      ��       S
�      =�       S                        ��      �       \M�      v�       \��      ��       \
�      =�       \                        �      &�       0�&�      G�       TG�      T�       QT�      Y�       T                         ��      ��       p 
�����      �       Z�      Y�       ��~��      ��       p 
���
�      "�       Z                        ��      ��      , ��H$��@$!��8$!��!�������      ��      	 ~ �������      r�       ^��      ��      � �H0H%�$!0)( 8/��
���H0H%�$!0)( 8/���H0H%�$!0)( 8/����������+( �����
�      =�       ^                          u�      u�       _u�      u�       �u�      ��       ���      &�       �&�      3�       x r "�G�      Q�        r "#�Q�      Y�       x r "���      ��       �
�      =�       �                      u�      �      	  ��~"��      Y�        w "���      ��      	  ��~"�
�      "�      	  ��~"�                 Q�      ��       S֨      ��       S                    i�      ��       P��      ��       0�֨      �       P��      ��       P                	 ��      ��       S=�      \�       S                    ��      ��       P��      ��       0�=�      Y�       P\�      \�       P                 Ѥ      Ѥ       0�                      ۩      �       0��      T�       ^=�      ��       ^                        ۩      �       0��      �       ]#�      T�       ]=�      ��       ]                          ۩      �       0��      �       \�      #�       |�#�      4�       \:�      T�       1�=�      ��       1�                  R�      s�       P                 �      %�       S                      ��      ��       Sq�      ��       S��      ©       ST�      =�       S                           ܧ      �       P�      !�       V!�      ;�       P��      ��       Pq�      ��       P��      �       V                          A�      ]�       2�]�      s�       R��      ©       1�T�      g�       2�g�      z�       1�z�      ��       R                      ��      ��       T��      ��       ]�      =�       ]                   ��      ��       V�      =�       V                    ��      ��       \�      =�       \                    ��      �       P�      +�       P                       ��      ��       ������      ˪       RΪ      ��       R �      =�       R                   ��      ��       0���      ܪ       T                  ��      ܪ       Q                      �             U      t       St      {       �U�                  �      z       V                                                                    ��      �       U�      �       _�      �       U�      ��       _��      ��       �U���      ��       _��      �       U�      �       _�      ��       U��      M�       _M�      V�       UV�      n�       _n�      ��       U��      �       _�      !�       U!�      1�       _1�      C�       UC�       �       _ �      L�       UL�      l�       _l�      ��       U��      k�       _k�      ��       U��      w�       _w�      ��       U��      ��       _                             ��      �       0��      �       ]��      H�       ]H�      �       0��      �       ]�      ��       0���      ��       ]                  ��      �       T                      �      �       0��      �       Q�      $�       q�                                                                                   ��      ��       V��      ��       V��      ��      
 83$0"�V�      ��       Vڳ      .�       V*�      �       V�      �       q 3$x "��      �      	 83$x "�]�      ��       V��      �       V��      #�       V��      ��       V��      �       V�      ;�       q 3$x "�;�      K�      	 83$x "���      (�       V��      e�       Ve�      ��      	 83$x "���      �       V�      @�      
 83$0"�\�      ��       R��      X�       Vk�      ��       V��      e�       Vw�      ��       V �      F�       Vc�      |�      	 83$x "���      ?�       V��      ��       V��      ��       R��      ��      
 83$0"���      ��       Vn�      ��       V��      ��      	 83$x "�                                                                                                                                                                                                                   ��      ��       ���      ��       �V�      j�       �t�      ��       �ڳ      �       ���      �       ��      �       �*�      >�       �O�      c�       �x�      ��       ���      �       ���      �       ��      3�       �D�      ķ       �ʷ      �       ��      �       �+�      A�       �i�      ��       ���      ¸       �Ӹ      ڸ       ��      �       �]�      ��       ���      2�       ���      -�       �z�      ��       ���      �       ���      �       �v�      }�       ���      ׽       �ƾ      �       ���      ��       ��      �       �C�      w�       ���      ��       ���      ��       �J�      ��       ���      ��       ���      �       ��      d�       �u�      ��       ���      ��       ���      ��       ��      %�       �3�      C�       �T�      Y�       �j�      z�       ���      {�       ���      ��       ���      ��       ���      ��       ���      �       �,�      4�       �E�      ��       ���      ��       ���      �       �L�      [�       �q�      ��       ���      2�       ���      ��       ���      ��       ���      D�       �^�      ��       ���      K�       ���      ��       ���      ��       ��      #�       ���      ��       ���      W�       �d�      ��       ���      ��       ��      @�       �\�      \�       �\�      ��       	����      ��       ��      �       ���      ��       ���      ��       ��      �       �(�      =�       �B�      e�       ���      ��       � �      $�       ���      �       ��      0�       �:�      C�       �M�      ��       ���      8�       �E�      W�       ���      ��       ���      ��       �)�      F�       �c�      |�       ���      ��       ��      ?�       ���      #�       �a�      q�       ���      ��       ���      ��       	��n�      |�       ���      ��       �                 �      (�       V                       �      ��       _X�      a�       _��       �       _��      ��       _                       /�      ��       VX�      a�       V��       �       V��      ��       V                       /�      9�       1�9�      ^�       Sh�      ��       SX�      a�       S                      9�      Q�       Ty�      ��       TX�      a�       T                      ��      ��       P��      ��       ��
��p "���      ��       PX�      a�       P                          /�      9�       P9�      ��       \X�      a�       \��       �       \��      ��       \                                 9�      Q�       r 3$p "y�      ��       r 3$p "��      ��       r 3$0"��      ��       q 3$0"��      ��       ux���      ��       U��      ��       Q��      ��       q 6��
������$���      ��        p pp0*( 6��
������$�X�      a�       r 3$0"                   կ      �       V|�      ��       V                   կ      �       _|�      ��       _                      ٯ      �       P|�      ��       P��      ��       v                        ��      d�       V��      0�       V��      ��       Vn�      ��       V                       ��      d�       _��      0�       _��      ��       _n�      ��       _                       ��      W�       v��      #�       v��      ��       vn�      |�       v                          ��      %�       P%�      W�       v ��      #�       v ��      ��       v n�      |�       v                                       ��      ��       0���      ��       Q[�      _�       P_�      d�       Q0�      B�       0�'�      +�       P+�      0�       Q��      ��       P��      ��       Q}�      ��       P��      ��       Q                      ��      ��       P��      #�       v �
��4$� "�n�      |�       P                      ��      ��       Q��      #�       v�
��4$�"�n�      |�       v�
��4$�"�                ��      ��       Y                      ��      ��       t z ���      ��       P��      ��       t z ���      ��       v �
��4$� "�z �                   ��      ��       P��      ��      
 p t "#���                  ��      ��       p ?&���      ��       T                  ��      �       Q�      �      
 q r "#���                  ��      �       q ?&��      �       R                }�      ��       �                 }�      ��       P                   ��      ��       P��      ��      
 p q "#���                  ��      ��       p ?&���      ��       Q                  ��      ��       P                  ��      ��       R                 ��      ��       _                 ��      ��       V                     e�      ��       R��      ��       R��      ��      
 83$0"�                   e�      ��       _��      ��       _                        g�      ��       P��      ��       q ��      ��       P��      ��       q                      g�      ��       q��      ��       U��      ��       q                          v�      ��       0���      ��       p���      ��       P��      ��       p���      ��       0�                     t�      ~�       V �      ��       V0�      a�       V                     t�      ~�       _ �      ��       _0�      a�       _                    F�      ��       Z\�      a�       Z                       F�      U�       0�U�      v�       Yv�      z�       y���      ��       Y                 ڳ      �       V                 ڳ      �       _                 ��      �       V                 �      .�       V                   �      *�       _��      n�       _                	 �      �       v                 
 �      �       v                 �      �       v                    )�      ��       X��      �       v                   )�      ��       Q��      �       v                     E�      *�       V��      n�       V                          }�      ��       ��~p "���      ��       ��~u "���      ��       P��      �       ��~u "���      ��       ��~u "�                  �      �       r ��~�                      �      �       | �s "#��      �       | ��~���      �       | ��~�                       �      �       U�      *�       ��~��      n�       ��~                  �      �       ��~                 ��      ܴ       ��}                      ��      �       y | ��      �       ��~| ���      ��       ��~| �                  !�      n�       \                 *�      >�       _                 W�      x�       _                  W�      x�       V                 ��      ��       _                  ��      ��       V                 ��      Ҷ       _                 ��      Ҷ       V                ��      ��       �                ��      ��       v                    ��      ��       Q��      ��      
 q r "#���                  ��      ��       q ?&���      ��       R                 ֶ      �       _                 ֶ      �       V                 �      ��       _                  �      ��       V                 ��      �       V                    ��      �       P�      �       v                 �      +�       _                 +�      D�       V                 D�      ��       _                  O�      ��       P                  T�      ��       R                 D�      ��       �                 ��      ʷ       V                 ��      ʷ       _                  ��      ��       T��      ķ       P                   ��      ��      	 p 0$0&���      ķ       U                   ��      ��      	 t 0$0&���      ķ       T                     ��      ��       ����      ķ       Qķ      ʷ       ��                   ��      ��      	 t 0$0&���      ķ       T                   ��      ��      	 p 0$0&���      ķ       U                 ʷ      �       V                 ʷ      �       _                  ҷ      ҷ       Tҷ      �       P                   ҷ      �      	 p 0$0&��      �       U                   ҷ      �      	 t 0$0&��      �       T                     ҷ      �       ���      �       Q�      �       ��                   ҷ      �      	 t 0$0&��      �       T                   ҷ      �      	 p 0$0&��      �       U                 �      +�       V                 �      +�       _                 +�      i�       V                 +�      i�       _                 i�      ��       V                 i�      ��       _                    m�      ��       P��      ��       v                  ��      Ӹ       V                 ��      Ӹ       _                  ��      Ӹ       Q                   �      �       q 3$x "��      �      	 83$x "�                  �      ]�       _                 �      ]�       V                    #�      ,�       P,�      3�       S                  3�      C�       R                     ]�      ��       _��      ��       _E�      W�       _                          ��      ��       Q��      ��       �� $ &5$�"���      ��       r $ &5$�"���      ��       Q��      ��       �� $ &5$�"�                    ��      ��       q��      ��       Q                  ��      ��       T                  ��      ��       _                     ��      ��       V��      ��       V��      ��       V                       ��      n�       _n�      ��       U��      ��       _��      ��       _                     �      ^�       Q��      ��       Q��      ��       Q                      ޹      ��       Y��      ��       Y��      ��       Y                      �      /�       R��      ��       R��      ��       R                       ��      z�       V��      ��       V��      ��       Vq�      ��       V                       ��      z�       _��      ��       _��      ��       _q�      ��       _                        ��      �       R�      <�       v ��      ��       R��      ��       R                      +�      T�       QT�      h�       r $ &5$�"�q�      ��       r $ &5$�"�                            ��      Ⱥ      	 r (p "�Ⱥ      h�       P��      ��       P��      ��      	 r (p "���      ��       r (�"�q�      ~�       P~�      ��       r $ &5$�"#                    Һ      ��       T��      ��       T                    Q�      h�       ph�      m�       Qq�      y�       p                  Q�      m�       Tq�      y�       T                  Q�      m�       _q�      y�       _                 ~�      ��       V                  ~�      ��       _                 ~�      ��       Q                   ��      ��       	����      ��       R                 ��      һ       _                 һ      ��       _                    �      =�       VI�      ��       V                    ��      ��       P��      ��       p �                   ��      v�       V��      )�       V                   ��      v�       _��      )�       _                     ��      ��       0���      v�       S��      )�       S                  !�      >�       P                   ��      ƾ       V4�      X�       V                   ��      ƾ       _4�      X�       _                    �      ƾ       [4�      X�       [                    �      ƾ       Y4�      X�       Y                      ��      �       P9�      ��       P4�      N�       P                    ��      ƾ       Z4�      X�       Z                   Ӿ      ��       V��      �       V                    Ӿ      ��       _��      �       _                   Ӿ      S�       S��      �       S                    <�      b�       P��      �       P                    S�      ��       Z�      �       Z                       S�      b�       Pb�      ��       Y��      ��       y���      ��       Y                 ��      ¿       _                 ��      ¿       V                 ¿      ݿ       _                 ݿ      ��       _                 ��      �       _                 ��      �       V                  �      ��       V�      W�       V                   �      ��       _�      W�       _                   ��      .�       VW�      ��       V                    ��      .�       _W�      ��       _                   2�      ��       V��      ��       V                    2�      ��       _��      ��       _                   ��      ��       V��      &�       V                    ��      ��       _��      &�       _                       ��      �       V��      ��       V)�      F�       V��      ��       V                       ��      �       _��      ��       _)�      F�       _��      ��       _                        ��      }�       T}�      ��       v��      ��       T)�      F�       T                      ��      ��       P��      ��       r $ &5$�"���      ��       r $ &5$�"�                            �      �      	 t (q "��      ��       Q��      ��       r $ &5$�"#��      ��       Q)�      A�      	 t (q "�A�      F�       t (�"���      ��       Q                    (�      M�       U��      ��       U                     ��      ��       q��      ��       Q��      ��       q                   ��      ��       T��      ��       T                   ��      ��       _��      ��       _                      �      �       Y�      �       y p ��      C�       Y                   C�      ��       Va�      q�       V                   C�      ��       _a�      q�       _                      Z�      g�       x ��g�      ��       Ua�      q�       U                        g�      w�       1���      ��       P��      ��       p�a�      q�       1�                       ��      #�       VB�      e�       V��      !�       VW�      ��       V                       ��      ��       _B�      e�       _��      !�       _W�      ��       _                
     ��      ��       vB�      e�       v��      !�       v                            ��      ��       P��      ��       \B�      e�       P��      �       P�      !�       \W�      ��       \                      ��      ��       P��      ^�       SW�      ��       S                    #�      0�       P0�      ��       V                	         ��      ��       ���      ��       ��}B�      e�       ���      !�       �W�      ��       ��}                 ��      J�       _                    ��      ��       P�      C�       P                 J�      ��       V                 J�      ��       _                      a�      r�       x ��r�      ��       U��      ��       x ��                 y�      ��       0�                   ��      ��       _��      ��       _                 ��      ��       V                 ��      ��       V                 ��      �       V                 �      0�       _                 �      0�       V                 0�      A�       _                 0�      A�       V                 A�      R�       _                 A�      R�       V                 R�      u�       V                 u�      ��       V                 ��      ��       _                 ��      ��       _                 ��      ��       _                   ��      ��       V:�      M�       V                   ��      ��       _:�      M�       _                 ��      �       V                 ��      �       _                 �      3�       V                 �      3�       _                 3�      T�       V                 T�      j�       V                 j�      ~�       V                  n�      ~�       Q                  v�      ~�       P                 v�      z�       v                  ��      ��       _                 ��      ��       _                 ��      =�       V                 ��      =�       _                  ��      =�       T                 ��      �       v                           ��      ��      	 q  $ &���      ��       R��      ��      	 q  $ &���      �      
 q   $ &��      =�       1t�$ $ &�                 =�      [�       _                 [�      k�       V                 [�      k�       _                 k�      ��       V                 k�      ��       _                 ��      ��       V                 ��      ��       V                 ��      ��       V                   ��      �       _��      �       _                   ��      �       V��      �       V                 �      ,�       V                 ,�      E�       V                 I�      `�       _                 I�      `�       V                 `�      q�       _                 `�      q�       V                 q�      �       V                 ��      ��       V                 ��      ��       V                 ��      ��       V                 ��      ��       V                   ��      L�       Vk�      ��       V                     ��       �       _ �      L�       Uk�      ��       U                      �      L�       Yk�      k�       Yk�      o�       y�o�      ��       Y                          �      C�       0�C�      L�       Pk�      r�       0�r�      w�       Pw�      ��       0�                 L�      q�       V                 L�      q�       _                 q�      ��       V                 q�      ��       _                 ��      ��       V                   ��      ��       V��      ��       V                     ��      l�       _l�      ��       U��      ��       _                    ��      ��       Y��      ��       Y                    ��      \�       R��      ��       R                   ��      ��       V!�      E�       V                   ��      ��       _!�      E�       _                      ��      ��       P��      ��       v !�      8�       v                       ��      ��       P<�      @�       P@�      E�       Q                 ��      ��       V                 ��      ��       _                  ��      ��       T                   ��      ^�       VM�      |�       V                   ��      ^�       _M�      |�       _                  ;�      ^�       Q                  %�      ^�       R                    '�      D�       QD�      ^�       U                     ^�      ��       _��      ��       _��      ��       _                      ��      ��       P��      ��       P��      ��       q 3$x "                     ��      �       V�      ;�       q 3$x "�;�      K�      	 83$x "�                 ��      ��       _                  ��      ��       \                     ��      �       v�      ;�      	 q 3$x "#;�      K�      
 83$x "#                      j�      p�       Sp�      v�       Rv�      ��       s �                 ��      ��       V                 ��      ��       _                  ��      ��       Q                ��      ��       �                ��      ��       v                   ��      ��       P��      ��      
 p t "#���                  ��      ��       p ?&���      ��       T                 ��      �       V                 ��      �       _                   ��      �       V��      ��       V                   ��      �       _��      ��       _                       �      �       Q�      �       r� $ &3$ "#���      ��       Q��      ��       r� $ &3$ "#�                       �      �       P�      �       v ��      ��       P��      ��       v                    �      �       _��      ��       _                       �      �       q p "��      �       P�      �       r� $ &3$ "#�v "���      ��       p q ���      ��       P                       �      e�       Ve�      ��      	 83$x "�c�      |�      	 83$x "���      ��      	 83$x "�                     �      ��       _F�      ��       _��      ��       _                                        v�      ��       P��      ��       U��      ��       P��      ��       UF�      K�       PK�      ]�       Uc�      j�       Pj�      |�       U��      ��       U��      ��       P��      ��       U��      ��       P                                    �      ��       Q��      ��       P��      ��       Q��      ��       PF�      K�       QK�      ]�       Tc�      j�       Qj�      |�       T��      ��       P��      ��       Q��      ��       P��      ��       Q                      ��      ��       Q��      ��       Q��      ��       Q��      ��       Q                       �      e�       ve�      ��      
 83$x "#c�      |�      
 83$x "#��      ��      
 83$x "#                           �      Q�       QQ�      e�       v e�      ��       83$x "c�      |�       83$x "��      ��       83$x "                       �      ��       ���      ��       Sc�      |�       ���      ��       �                        X�      |�       T|�      ��       �| "�c�      |�       �| "���      ��       �| "�                        k�      y�       Qy�      ��       �v "�c�      |�       �v "���      ��       �v "�                            ��      ��       ����      ��       ��K�      c�       ��j�      ��       ����      ��       ����      ��       ����      ��       ����      ��       ��                      ��      ��       Pj�      |�       T��      ��       P��      ��       Q                      ��      ��       Uj�      |�       U��      ��       U��      ��       P                      ��      ��       \F�      c�       \��      ��       \                      ��      ��       VF�      c�       V��      ��       V                      ��      ��       ��K�      c�       ����      ��       ����      ��       ��                      ��      ��       PK�      ]�       T��      ��       P��      ��       Q                      ��      ��       UK�      ]�       U��      ��       U��      ��       P                 d�      ��       V                 d�      ��       _                  ��      ��       P                  h�      ��       S                 ��      �       V                 ��      �       _                  ��      ��       T                   	�      �       V��      ��       V                    	�      �       _��      ��       _                   	�      �       R��      ��       R                  ��      ��       S                 ��      ��       V                 ��      ��       _                   ��      ��       0���      ��       P                  ��      ��       t�                 ��      ��       _                 ��      ��       V                   ��      �       V��      ��       V                   ��      �       _��      ��       _                  ��      �       Q                  ��      �       R                    ��      ��       Q��      �       U                   �      ��       V��      ��       V                   �      ��       _��      ��       _                    �      ��       R��      ��       R                 ��      4�       V                 ��      4�       _                  �      4�       R                    �      &�       P&�      *�       p�                 �      ?�       V                 �      ��       _                   �      1�       s�~�1�      ��       s�                 5�      ?�       0�                   ?�      J�       _J�      ��       _                    ��      =�       Q=�      D�       �� $ &5$�"#                    ��      �       R�      D�       ������53$�"�                    �      0�       P0�      D�       �� $ &5$�"�                   -�      =�       q=�      E�       Q                 -�      E�       T                 -�      E�       _                     ߮      �       u��      �       ��      ��       u�                                                             ߮      �       U�      ��       _��      ��       �U���      H�       _�      �       _�      ��       U��      M�       _M�      V�       UV�      n�       _n�      ��       U��      �       _�      !�       U!�      1�       _1�      C�       UC�       �       _ �      L�       UL�      l�       _l�      ��       U��      k�       _k�      ��       U��      w�       _w�      ��       U��      ��       _                    �L      oM       PyM      �M       P                        �L      M       QM      oM       u������53$u�"�yM      �M       Q�M      �M       u������53$u�"�                  GM      bM       Q                     _M      oM       poM      pM       Q�M      �M       p                   _M      pM       T�M      �M       T                     _M      gM       XgM      pM       U�M      �M       U                            �      �       U�      |       S|      �       �U��             S             �U�      s       S                        �      �       T�      �       V�      j       �T�j      s       V                      �      �       ]�             ]      s       ]                           �      �       1��      :       \D      w       \�      �       \      j       \j      s       1�                          �      1       QU      w       Q�      �       Q�      �       Q      j       Q                                     T      )       s��
��t "�)      1       P�      �       P�      �       T                          �      �       P�      w       ^�             ^      j       ^j      s       P                                     �             u 3$p "      1       u 3$s0"U      w       u 3$p "�      �       t 3$s0"�      �       rx��      �       R�      �       T�      �      / u 3$s0"?7u 3$s0"?8u 3$s0"?80*( ��      �       R�      �       u 3$s0"      j       R                              @{      �{       U�{      >|       ^>|      }|       U}|      �|       �U��|      �|       U�|      I~       ^I~      ^~       U                      }{      �{       @��{      >|       ]�|      �|       8��|      I~       ]                   �{      &|       Z�|      �|       Z                    �{      >|       V�|      I~       V                 �|      I~       S                       �|      �|       S�|      �|       _�|      }       R}      I~       _                            �{      |       Z|      &|       S&|      >|       Z�|      �|       S�|      �|       P�|      I~       \                       �{      �{       0��{      &|       Y*|      >|       Y�|      �|       Y                      �|      }       \A}      L}       \L}      Q}       _                        �|      �|       _�|      }       RA}      H}       _H}      Q}       t�                      �|      }       Q}      }       |�A}      Q}       Q                    �|      }       TA}      Q}       T                        �|      �|       ����|      }       U}      }       ���A}      Q}       ���                  ]}      �}       S                  ]}      �}       _                  ]}      �}       V                    ]}      �}       T�}      �}       
���                      ]}      �}       ����}      �}       U�}      �}       ���                  �}      �}       S                  �}      �}       _                    �}      �}       Q�}      �}       s�                  �}      �}       Z                      �}      �}       ����}      �}       U�}      �}       ���                   �}      �}       ����}      I~       ���                    �}      �}       S�}      I~       S                    �}      �}       V�}      I~       V                      �}      �}       Z�}       ~       Z ~      0~       z  �                          �}       ~       Z ~      ~       z  �,~      5~       P5~      =~       p�=~      I~       P                      �}      �}      
 r u q "��}      �}       R�}      I~       R                            @      �       U�      =       S=      G       �U�G      �       S�      �       �U��      P       S                          �             ���      �       ��"      �       ��0      5       PK      P       P                                   P�      �       ��"      �       ��                      �             \�      �       \      P       \                      �             V�      �       V      P       V                        {      �       1�l      �       0�      "       1��      P       0�                                    t u "#��@& $ &���            ( t u "#��@& $ &��q r "#��@& $ &��            M s��
��4$s�"�y  $ &s�� $ &u "#��@& $ &��q r "#��@& $ &��            u s��
��4$s�"�y  $ &s�� $ &s��
��4$s�"�y  $ &s�� $ &?&"#��@& $ &��q r "#��@& $ &��      *      � s��
��4$s�"�y  $ &s�� $ &s��
��4$s�"�y  $ &s�� $ &?&"#��@& $ &��s��
��4$s�"#�x  $ &s�� $ &r "#��@& $ &��                  �      �       U�             s�                    �      �       t y ��      �       T�             s��
��4$s�"�y �                   �             T            
 t u "#���                  �             t ?&�             U                               Q            
 q r "#���                               q ?&�             R                      �      �       _�      �       p 3$�U#0""      �       _                          r      �       P�      �       ^d      i       Px      �       R�      �       ^                      �      �       Px      �       P�      �       ��                       4      8       p t "#��@& $ &���8      @      ( p t "#��@& $ &��q u "#��@& $ &��@      H      + p ?&p "#��@& $ &��q u "#��@& $ &��H      O      I p ?&p "#��@& $ &��s�r "#�z  $ &s�� $ &u "#��@& $ &��O      [      j p ?&p "#��@& $ &��s�r "#�z  $ &s�� $ &s�r "#�z  $ &s�� $ &?&"#��@& $ &��                      4       [                                t p �      -       T                   &      4       P4      4      
 p t "#���                  &      4       p ?&�4      4       T                  4      8       Q8      8      
 q u "#���                  4      8       q ?&�8      8       U                        �      �       U�             S             �U�      �       S                    �      �       T�      �       �T�                      �             ]             �U#�      �       ]                         �      �       t#��      3       t�      :      	 �T##�:      J       t�J      g       R                                  >      A       PA      �       _�      �       _:      g       0�g      x       _x      {       P{      �       _�      �       P�      �       _                    �      �       P�      �       P                          3      8       P8      �       R�      �       ��g      �       R�      �       R                            
       P
      �       ^g      �       ^                 �      �       u�                 �      �       u�                   g      �       t 3�#<3$s "#�      �       t 3�#<3$s "#                         g      x       _x      {       P{      �       _�      �       P�      �       _                   g      �       S�      �       S                        p      O       UO      �       S�      �       �U��      7       U                      p      C       TC      �       ���      7       T                            p      �       Q�      �       V�      �       �Q��      �       Q�      .       V.      7       �Q�                      p      O       RO      �       �R��      7       R                      p      O       XO      �       �X��      7       X                                                    �      �       Q��8�      �       Q�_��6�      �       Q�_�^�[��2�      �       Q�_�^�[�S�Y��(�      �       Q�_�^�[�u� �Y��(�      �       Q�_�^�[�u� �Y�Z�� �      �       Q�_�^�[����Y�Z�� �      -       r �_�^�[����Y�Z�� -      4       �_�^�[����Y�Z�� 4      O       �_�^�[����Y��(O      �       �_�^������0�      �       Q��8�      �       Q�_��6�      �       Q�_�^�[�����0�      �       Q�_�^�[����Y��(�      4       Q�_�^�[����Y�Z�� 4      6       Q�_��[����Y�Z�� 6      7       Q��[����Y�Z��                     �      1       P1      O       x              P                    e      i       Pi      �       ]                     
      
       T
      8
       �T�                     
      
       Q
      8
       �Q�                 
      )
       u��0$0&�                 
      )
       u��0$0&�                   
      "
       Q"
      )
       �Q�                 
      )
       T                     
      "
       R"
      )
       Q)
      )
      	 p q "#�@�                  "
      )
       q ?&�)
      )
       P                    �	      �	       T�	      �	       �T�                    �	      �	       Q�	      �	       �Q�                �	      �	       u��0$0&�                �	      �	       u��0$0&�                  �	      �	       Q�	      �	       �Q�                �	      �	       T                     �	      �	       R�	      �	       Q�	      �	      	 p q "#�@�                  �	      �	       q ?&��	      �	       P                                    `      �       T�      �       R�      	       �T�	      	       R	      (	       �T�(	      W	       RW	      q	       �T�q	      {	       R{	      �	       �T��	      �	       R                                  `      �       Q�      	       �Q�	      $	       Q$	      (	       �Q�(	      b	       Qb	      q	       �Q�q	      �	       Q�	      �	       �Q��	      �	       Q                           '       Q'      0       �Q�                                 Q             �Q�                    �      �       Q�             �Q�                    p      �       Q�      �       �Q�                            �      �       U�      �       V�      �       �U��      �       U�      1       V1      :       �U�                          �      �       T�      �       \�      �       �T��      3       \3      :       �T�                            �      �       Q�      �       S�      �       �Q��      �       Q�      
       S
      :       �Q�                            �      �       R�      �       ]�      �       �R��      �       R�      5       ]5      :       �R�                   �      �       T�             T                          @      �       U�      �       V�             �U�      '       U'      k       V                        @      _       T_      �       \�             �T�      k       \                          @      �       Q�      �       S�             �Q�      $       Q$      k       S                          @      �       R�             �R�      8       R8      O       ��O      k       �R�                        _      �       T�      �       T      8       TO      k       T                      �0      �0       U�0      �0       V�0      �0       �U�                      �0      �0       T�0      �0       S�0      �0       �T�                      �0      �0       Q�0      �0       \�0      �0       �Q�                      �0      �0       U�0      �0       S�0       1       �U�                      �0      �0       T�0      �0       \�0       1       �T�                      �0      �0       Q�0      �0       V�0       1       �Q�                       1      1       U1      #1       S#1      91       �U�                       1      1       T1      $1       V$1      91       �T�                  1      (1       P                     1      #1       v 3$s�"�#1      $1       v 3$�U#�"�$1      *1       �T3$�U#�"�                   (1      *1       P*1      *1      
 p q "#���                  (1      *1       p ?&�*1      *1       Q                      @1      H1       UH1      Q1       SQ1      f1       �U�                  I1      W1       P                     I1      Q1      
 s��
���Q1      Y1       q 
���Y1      Y1       �U#��
���                   W1      Y1       PY1      Y1      
 p q "#���                  W1      Y1       p ?&�Y1      Y1       Q                       0      z0       Uz0      �0       S�0      �0       �U�                    �0      �0      	 p  $ &��0      �0      	 x  $ &�                    �0      �0      	 p  $ &��0      �0       T                                 T      .       �T�                              !       T!      )      	 p t "#�@�)      -       P-      .       t ?&t "#�@�                           !       t ?&�!      )       P)      .       t ?&�                    ��      ��       U��      ��       �U�                    ��      ��       V��      ��       V                         ��      ��       0���      -�       P-�      ��       S��      ��       P��      ��       S                 �      ~�       V��      ��       V                   �      -�       P-�      ~�       S��      ��       S                          �#      :&       U:&      s&       Ss&      u&       �U�u&      2'       S2'      4'       �U�                          �#      H&       TH&      t&       Vt&      u&       �T�u&      3'       V3'      4'       �T�                      �#      ?&       Q?&      \&       s\&      4'       �Q�                     %      %       0�%      4%       1�4%      K%       2�K%      2&       3�                         �#      H&       t��H&      t&       v��t&      u&       �T#��u&      3'       v��3'      4'       �T#��                    ]&      ~&       P�&      4'       P                    �#      �#       U�#      �#       �U�                      �#      �#       T�#      �#       S�#      �#       �T�                    �#      �#       Q�#      �#       �Q�                      �#      �#       R�#      �#       \�#      �#       �R�                      �#      �#       X�#      �#       V�#      �#       �X�                     �#      �#       R�#      �#       \�#      �#       �R�                        P      n       Un      �       S�      �       T�      �       �U�                    ]      �       V�      �       U                        p!      �!       U�!      b#       ^b#      g#       �U�g#      y#       U                 p!      r!       u�                        !      [#       S[#      f#       Tg#      q#       Sq#      y#       u�	                  �!      "       0�                  �!      �!       V                    �       �        U�       n!       �U�                      �       �        T�       h!       Sh!      n!       �T�                  �       m!       ]                            �       �        0��       �        \�       �        |��       	!       \"!      +!       0�+!      9!       V9!      B!       v�B!      S!       V                          pU      �U       U�U      TV       ��~TV      fV       �U�fV      wV       UwV      �a       ��~                            pU      �U       T�U      'V       S'V      fV       �T�fV      wV       TwV      QW       SQW      �a       �T�                          pU      �U       Q�U      TV       ��}TV      fV       �Q�fV      wV       QwV      �a       ��}                          pU      �U       R�U      TV       ��~TV      fV       �R�fV      wV       RwV      �a       ��~                            �U      'V       ]fV      �X       ]�\      �\       ]	]      &]       ]ha      xa       ]�a      �a       ]                                  �U      'V       _fV      �X       _�X      �\       ��~�\      �\       _	]      &]       _&]      ha       ��~ha      xa       _xa      �a       ��~�a      �a       _                           �U      'V       ^fV      �X       ^�\      �\       ^	]      &]       ^ha      xa       ^�a      �a       ^                         �U      V       0�V      'V       P'V      4V       ��}4V      wV       0�wV      �V       P�V      �a       ��}                       �U      'V       0�'V      AV       ��}AV      �V       0��V      �V       P�V      �a       ��}                       �U      'V       0�'V      MV       w MV      �V       0��V      �V       P�V      �a       w                             UW      $X       s v �$X      0X       S�\      �\       s v �	]      &]       s v �ha      xa       s v ��a      �a       S                      �W      0X      
 ��~�
���ha      xa      
 ��~�
����a      �a      
 ��~�
���                                           �W      �Y       \�\      �\       ��~�]      �]       \�]      �]       P�]      �]       _�]      �]       \�]      �]       P�]      $^       __      i_       \i_      o_       Po_      �_       _ha      �a       \�a      �a       | q ��a      �a       \                            uY      yY       QyY      �\       ��~&]      �]       ��~$^      K_       ��~�_      ha       ��~�a      �a       S                          hX      �X       0��X      �\       ��~�\      �\       P&]      ha       ��~xa      �a       ��~                                                             0X      VX       0�Z      =Z       0�=Z      IZ       q v �VZ      yZ       0�yZ      �Z       R�[      �[       0��[      ,\       Q�]      �]       0��]      �]       V�]      �]       r��]      �]       0��]      ^       V^      $^       r��^      _       QK_      o_       0�o_      �_       V�_      �_       r��_      �_       QM`      _`       Q_`      �`       0��`      �`       Q�`      �`       q��`      ha       Q                           �U      fW       0�fW      �W       P�W      �\       ��~�\      �\       0��\      	]       ��~	]      &]       P&]      �a       ��~                            �U      �W       0��W      �W       P�W      �\       ��~�\      �\       0��\      �\       P	]      &]       0�&]      �a       ��~                          �U      �W       0��W      �W       P�W      �\       ��~�\      �\       0�	]      &]       0�&]      �a       ��~                                    �U      'V       0�fV      0X       0�0X      �\       ��~�\      �\       0�]      &]       0�&]      ha       ��~ha      xa       0�xa      �a       ��~�a      �a       0��a      �a       P�a      �a       ��~                                       �U      'V       0�fV      �X       0��X      C\       ��~C\      L\       0�L\      �\       ��~�\      �\       0�	]      &]       0�&]      <_       ��~<_      K_       PK_      ha       ��~ha      xa       0�xa      �a       ��~�a      �a       0�                      �Y      �Y       ��~�Y      �Z       S<_      K_       P_`      �`       S                                �Y      �Y       P�Y      yZ       \yZ      ^\       ��~^\      �\       0�&]      �]       ��~$^      _       ��~�_      _`       ��~_`      �`       \�`      ha       ��~                                �Y      �Y       P�Y      0Z       R0Z      k\       ��~k\      �\       0�&]      �]       ��~$^      _       ��~�_      _`       ��~_`      �`       R�`      ha       ��~                          �X      �X       p 
����X      UY      
 ��~�
����]      $^      
 ��~�
���K_      �_      
 ��~�
���xa      �a      
 ��~�
���                          �X      �X       p 
����X       Y       s 
���K_      f_       p 
���f_      �_      
 ��~�
���xa      �a       s 
���                        LY      PY       PPY      �Y       X_      *_       X*_      K_       ��~                          �`      �`       S�`      �`      / q 1$y "�0$0&p q 1$y "�0$0&p ?&"#��@&��`      %a       S%a      6a      / q 1$y "�0$0&p q 1$y "�0$0&p ?&"#��@&�6a      ha       S                          �`      �`       R�`      �`      / q 1$z "�0$0&p q 1$z "�0$0&p ?&"#��@&��`      Ba       RBa      Ra      / q 1$z "�0$0&p q 1$z "�0$0&p ?&"#��@&�Ra      ha       R                 �`      �`       q 1$y "�0$0&�                      �`      �`       R�`      �`      
 r s "#����`      �`       S                       �`      �`       r ?&��`      �`       S�`      �`       r ?&��`      �`       q 1$y "�0$0&p ?&�                 �`      �`       q 1$z "�0$0&�                      �`      �`       R�`      �`      
 r | "#����`      �`       R                     �`      �`       r ?&��`      �`       \�`      �`       q 1$z "�0$0&p ?&�                    �Z      �Z       U�Z      �Z       Q                  �Z      �Z       t 1$z "�0$0&��Z      �Z       r ����1$z "�0$0&�                   �Z      �Z       U�Z      �Z      
 u | "#���                  �Z      �Z       u ?&��Z      �Z       \                  �Z      �Z       T�Z      �Z      
 t u "#���                  �Z      �Z       t ?&��Z      �Z       U                          �[      �[       T�[      ,\       T�^      _       T�_      �_       TM`      _`       T                               �[      �[       R�[      �[       _�[      #\       R#\      ,\       _�^      _       R_      _       _�_      �_       RM`      _`       R                       �Z      ,\       ��}&]      �]       ��}$^      _       ��}�_      _`       ��}                               �Z      ,\       V&]      S]       VS]      X]       w X]      �]       S$^      -^       S-^      G^       w G^      _       V�_      _`       V                       �Z      ,\       ��}&]      �]       ��}$^      _       ��}�_      _`       ��}                       �Z      ,\       ��}&]      �]       ��}$^      _       ��}�_      _`       ��}                         #[      i[       ^&]      �]       ^$^      �^       ^�_      �_       ^�_      E`       ��~                              #[      �[       S&]      M]       SM]      X]       RX]      �]       \$^      G^       \G^      �^       S�_      M`       S                     )]      �]       ]$^      �^       ]�_      M`       ]                             )]      X]       ]X]      h]       Qk]      �]       Q�]      �]       u�$^      {^       Q{^      �^       _�_      M`       _                                      [      G[       ^G[      T[       QT[      _[       ]_[      b[       q�b[      i[       Qi[      �[       ^&]      )]       ^)]      -]       ]-]      X]       ZX]      k]       Vk]      o]       v�x]      �]       V                          [      i[       [m[      �[       [&]      X]       [X]      �]       ��$^      o^       ��                    X]      k]       ��}�]      �]       ��}                    X]      k]       ��}�]      �]       ��}                    X]      k]       V�]      �]       V                      X]      h]       Q�]      �]       Q�]      �]       u�                      X]      h]       Th]      k]       v��]      �]       T                    X]      h]       U�]      �]       U                  J^      �^       ��}                  J^      �^       ��}                  J^      �^       ]                    J^      {^       Q{^      �^       _                  J^      �^       S                    J^      {^       U{^      �^       �                  �^      �^       ��}                  �^      �^       ��}                  �^      �^       ]                  �^      �^       _                    �^      �^       T�^      �^       }�                  �^      �^       ^                 �_      E`       ��}                 �_      E`       ��}                 �_      E`       _                 �_      E`       S                   �_      �_       ^�_      E`       ��~                     �_      �_       ^�_      
`       ��~`      4`       �                                    `7      �7       U�7      �7       V�7      
8       �U�
8      �9       V�9      �;       ���;      �;       �U��;      R<       ��R<      j<       Vj<      H=       ��H=      �=       V                                  `7      �7       T�7      �7       Q�7      �7       \�7      
8       �T�
8      %9       \%9      )9       U)9      ]<       \]<      a<       Ua<      �=       \                              y7      �7       S
8      �9       S�9      �;       ���;      R<       ��R<      j<       Sj<      H=       ��H=      �=       S                      ;8      ?8       |� p �?8      v9      
 ��~��~�R<      j<      
 ��~��~�                        39      �9      
 ��~�
���R<      ]<      
 ��~�
���H=      V=      
 ��~�
����=      �=      
 ��~�
���                                                D9      v9       Rv9      �9       P�9      �:       ��~m;      �;       ��~�;      R<       ��~R<      ]<       Rj<      w<       ��~�<      �<       ��~1=      H=       ��~H=      Q=       PQ=      �=       ��~�=      �=       q p ��=      �=       Q�=      �=       ��~�=      �=       P�=      �=       ��~                              N:      S:       QS:      m;       ��~�;      �;       ��~j<      �<       ��~�<      1=       ��~w=      �=       Y�=      �=       ��~                          9      �9       0��9      w;       ��~{;      �;       P�;      R<       ��~j<      H=       ��~�=      �=       0�                                          �:      �:       0��:      �:       q��:      ;       Q;      %;       q��;      �;       0��;      <       S<      '<       0�'<      R<       V�<      �<       0��<      �<       V�<      �<       0��<      '=       T'=      1=       P                          y7      �7       0��7      �8       0��8      �8       P�8      �8       ^�8      �8       P�8      �=       ^                          y7      �7       0��7      �8       0��8      �8       P�8      �8       w �8      9       P9      �=       w                 	      y7      �7       0��7      9       0�9      )9       P)9      �=       _                
   y7      8       ]
8      �=       ]                                   �7      �7       0�
8      �9       0��;      �;       Z�;      �;       ��~�;      �;       ZR<      j<       0�H=      �=       0��=      �=       P�=      �=       Z�=      �=       0�                                     �7      �7       0�
8      �9       0��9      4;       ��~4;      =;       0�=;      �;       ��~�;      �;       ��~�;      R<       ��~R<      j<       0�j<      �<       ��~�<      �<       P�<      H=       ��~H=      �=       0�                        v:      �:       ���:      X;       S�;      �;       S�<      �<       P�<      1=       S                          �:      �:       P�:      J;       VJ;      m;       0��;      �;       P�;      �;       V�<      1=       V                          �9      �9       p 
����9      /:      
 ��~�
����;      R<      
 ��~�
����<      �<      
 ��~�
���1=      H=      
 ��~�
���                              �9      �9       p 
����9      :       s 
����;      �;       s 
����;      R<      
 ��~�
����<      �<       p 
����<      �<       s 
���1=      ;=       s 
���                        *:      <:       P<:      �:       Rj<      {<       R{<      �<       ��~                 �<      !=       p 1$u "�0$0&�                �<      =       p 1$v "�0$0&�                   
=      =       Q=      =      
 q y "#���                  
=      =       q ?&�=      =       Y                 �:      ;       q 1$s "�
���                  ;      ;       r 1$t "�0$0&�                ;      ;       q 1$v "�0$0&�                   ;      ;       P;      ;      
 p { "#���                  ;      ;       p ?&�;      ;       [                            ��      ��       U��      ��       S��      ��       �U���      '�       S'�      /�       �U�/�      w�       S                                ��      ��       T��      ��       V��      ��       �T���      �       V�      /�       �T�/�      Z�       VZ�      b�       Tb�      w�       V                             ��      ��       6���      ��       P�      �       P�      ;�       PT�      Z�       PZ�      g�       6�g�      w�       P                   ��      �       s�	��      �       s�	                     ��      ��       q��      �       ]/�      Z�       ]                   ��      �       s�@%���      �       s�@%�                    ȗ      �       \/�      Z�       \                 ȗ      �       s�                    ԗ      �       ^/�      Z�       ^                            ��      ��       U��      �       ]�      �       �U��      B�       ]B�      N�       UN�      ��       ]                          ��      ��       T��      �       S�      �       s��      �       �T��      ��       S                            ��      ��       Q��      �       \�      �       �Q��      B�       \B�      N�       QN�      ��       \                       ��      ��       0�B�      O�       0�O�      e�       Py�      ��       P                    ��      �       V�      B�       VZ�      ��       V                            ��      Ϙ       0�Ϙ      Ә       p�Ә      ۘ       Pۘ      �       p��      ��       R�      /�       0�                     ��      ��       S��      �       R�      B�       R                            �      E�       UE�      ��       ]��      ��       �U���      ��       ]��      �       U�      s�       ]                      �      E�       TE�      ��       S��      s�       S                                  �      E�       QE�      �       _�      ��       �Q���      �       _�      ��       �Q���      �       Q�      S�       _S�      X�       �Q�X�      s�       _                   E�      ^�       }�	�      6�       }�	                        I�      u�       V��      ��       V�      K�       VX�      s�       V                           ^�      t�       0�t�      {�       q�{�      ��       Q��      ��       q�Õ      ֕       T��      ��       TX�      i�       0�                   <�      ��       \��      s�       \                                  t�      {�      
 q 3$p "#�{�      ��       q 3$p "���      ��      
 q 3$p "#�Õ      ֕       P֕      �       p q "��      ��       p q "#���      ��       p q "���      Ֆ       PՖ      ٖ       px�ٖ      �       P                                 ^�      t�       _t�      {�      
 q 3$ "#�{�      ��       q 3$ "���      ��      
 q 3$ "#�Õ      ֕       X֕      �       x q "��      ��       x q "#���      ��       x q "�X�      i�       _                         <�      �       0��      #�       P#�      ��       _��      �       0��      ��       _��      s�       0�                                   <�      t�       0�t�      ��       U��      ��       1���      ��       UÕ      �       U�      �       1��      �       U�      u�       1���      ̖       U̖      і       1�і      �       U�      ��       1���      i�       0�i�      s�       U                   ��      ��       q @%���      ֕       }�@%�                   ��      ��       q @%����4$v"@���      ֕       }�@%����4$v"@�                  ��      �       Q                            ��      ��       U��      ,�       ],�      -�       �U�-�      R�       ]R�      ^�       U^�      ��       ]                          ��      ��       T��      ��       S��      ��       s���      -�       �T�-�      ��       S                            ��      ��       Q��      *�       \*�      -�       �Q�-�      R�       \R�      ^�       Q^�      ��       \                       ��      ��       0�R�      _�       0�_�      u�       P��      ��       P                    ��      "�       V-�      R�       Vj�      ��       V                            Й      ߙ       0�ߙ      �       p��      �       P�      ��       p���      �       R-�      ?�       0�                     ��      ƙ       Sƙ      "�       R-�      R�       R                                    `�      ��       U��      ŏ       \ŏ      ̏       �U�̏      ��       \��      ��       �U���      ��       \��      �       U�      ��       \��      ��       ^��      	�       \                                        `�      ��       T��      L�       S��             S��      3�       SQ�      ,�       S,�      \�       V\�      ��       S��      �       S�      "�       V"�      ��       S��      ��       \��      	�       S                                      `�      ��       Q��      �       ^�      ��       �Q���      ��       ^��      ��       �Q���      �       Q�       �       ^ �      ő       �Q�ő      m�       ^m�      ͓       �Q�͓      ��       ^��      	�       ��~                        `�      ��       R��      ��       �R���      �       R�      	�       �R�                    ��      �       |�	��      ��       |�	ő      �       |�	                         ��      U�       _��      ��       _Q�      ��       _��      œ       _͓      	�       _                               ��      Ԍ       0�.�      U�       0�U�      p�       Pp�      r�       p�r�      z�       P�      �       Q �      3�       P��      œ       0�                                      ��      !�       0�!�      `�       ��~��      ��       0���      ��       ��~��       �       0� �      3�       ��~Q�      ��       0���      ő       ��~ő      ��       0���      ��       ��~��      ͓       ��~͓      	�       0�                                ��      ��       P��      ��       w ��      ̏       ��~̏      ��       w ��      ��       ��~��      ��       w ��      �       P�      	�       w                           ��      ��       ��~̏      ��       ��~3�      Q�       ��~��      ��       ��~œ      ͓       ��~                            ��      �       Y�      �       1���      �       Y�      ��       1���      ��       Yœ      ͓       Y                        ʍ      ܍       r x "�܍      ��       r x "#���      �       r x "�А      �       P                        ��      ʍ       Pʍ      ܍       p x "�܍      ��       p x "#���      �       p x "�                     ��      ��       x @%���      ��       X��      �       |�@%�                       `�      ��       \̏      �       \��      ��       \��      ��       \                        `�      ��       ^̏      �       ^��      ��       ^��      ��       ^                        `�      ��       R��      ��       }��      ��       R��      ��       }                      `�      ��       S��      ��       s���      ��       S                         `�      m�       Pm�      ��       ��~̏      �       ��~��      ��       ��~��      ��       P                    T�      X�       pX�      ^�       P �      �       ��~#                      \�      ��       R�      �       R��      ��       R                	                       `�      o�       0�o�      s�       p�s�      {�       P{�      ��       p���      ��       R      �       0�\�      `�       0�`�      ��       P��      ��       p���      ��       P�      �       0���      ��       P��      ��       0�                          �      �       1��      6�       R6�      9�       T9�      >�       Ȑ      ڏ       R                        `�      `�       S`�      ׎       V׎      \�       ��~̏       �       ��~ �      �       V��      ��       V                           �       ]�      \�       _̏       �       _                 f�      k�       r�u �                 f�      k�       Q                   u�      |�       Q|�      |�      
 q t "#���                  u�      |�       q ?&�|�      |�       T                   ��      ��       u r����      ��       T                 ��      ��       Q                       ő      q�       \͓      ��       \��      ��       ^��      	�       \                      ͑      �       P�      q�       ��~͓      	�       ��~                 ͑      �       ��~                 ͑      �       |�	                      ,�      X�       S�      "�       S��      ��       V                      ��      ��       0���      ޔ       Sޔ      �       s��      �       S                  	�      �       ��~                       ʒ      
 ��~��~"�                                         �      r�       Ur�      Á       ]Á      �       �U��      -�       U-�      �       ]�      4�       �U�4�      ̆       ]̆      ��       �U���      n�       ]n�      Q�       ��~Q�      ҋ       ]ҋ      _�       �U�                         �      r�       Tr�      �       ��}�      (�       T(�      _�       ��}                          N�      Á       V�      �       V4�      ݆       V��      ҋ       V�      ��       V                        S�      r�       Pr�      �       ��}�      -�       P-�      _�       ��}                             ^�      r�       0�r�      Á       ^�      ��       0���      ��       P��      �       ^4�      ��       ^Q�      w�       ^                             ڄ      ��       0�$�      =�       0���      ��       0�!�      n�       0�n�      �       _�      �       ��      Q�       _Q�      w�       0�ǋ      ҋ       0�                  t�      ��       0���      ��       0�                               ^�      Á       0��      ��       P��      �       R�      �       0�4�      �       0��      ��       P��      ք       Uք      _�       ��~                    >�      ��       Uڄ      �       T                          !�      1�       P1�      n�       Rn�      *�       \9�      Q�       \ǋ      ҋ       P                              |�      �       Q�      �       p �      �       q{��      ��       Q�      4�       Q$�      a�       [Q�      ]�       []�      w�        ��}"��~"��~"��~"�                            o�      ��       P�      4�       P��      ��       ^��      ��       Sq�      ��       Q��      ��       qP���      ��       Q                              t�      ��       P��      ��       px���      ��       P��      Ǌ       ]Ǌ      Њ       }x�Њ      /�       ]9�      Q�       ]                                b�      t�       Pt�      ��       ��~�
��4$u"��      n�       Un�      ��       ^��      �       ~p��      Q�       ^��      ��       P��      ҋ       U                           ^�      r�       0�r�      Á       ��~�      ك       0�ك      �       s 
�� $| 
��2$# $)�4�      ��       ��~��      ��       ��~                          ��      ��       R��      Á       ��~4�      �       ��~��      ҋ       ��~�      ��       ��~                          o�      Á       \�      �       \4�      ��       \��      ��       ��~Q�      w�       \                          "�      '�       p �'�      ��       r ��      4�       r �Ʉ      ��       _��      i�       \i�      m�       |~�m�      {�       \Q�      w�       _                   ��       �        ��      _�        �                      ��      ��       P��       �       ��~�      _�       ��~                      ��      ��       P��       �       ��~�      _�       ��~                      ��      ��       P��       �       ��}�      _�       ��}                          ��      Á       PÁ       �       ��~�      4�       ��~4�      A�       PA�      _�       ��~                       ��      Á       | 5�����4�      ��       | 5�������      ��       ��~�5�����Q�      w�       | 5�����                     ^�      Á        0)��      �        0)�4�      ��        0)�                    ��      ��       P��      ҋ       ^                    ݆      ��       Vҋ      �       V                        �      #�       p ��$�      .�       p ��I�      U�       p ��ҋ      �       p ��                     ݆      .�       	��.�      ��       ^ҋ      �       	��                  >�      W�       0�|�      ��       0�                   ��      ��       ]��      _�       ]                    ��      ��       V��      _�       V                  ��      ��       ^                   ��      ��       _��      _�       _                     ��      ��       r���      �       s���      �       s�                      ��      ��       ^��      &�       ^&�      _�       Q                        ��      ��       P��      ��       ��~��      -�       ��~-�      _�       R                  ��      ��       ��~                    �      �       P�      �       ��~                  ��      ��       ��~                  Ɉ      ܈       ��~                  :�      B�       P                            p      �       U�      L       _L      M       �U�M      x       _x      y       �U�y             U                      p      �       T�      y       �T�y             T                            p      �       Q�      H       ]H      M       �Q�M      t       ]t      y       �Q�y             Q                            p      �       R�      F       \F      M       �R�M      r       \r      y       �R�y             R                      p      �       X�      y       ��y             X                           p      �       0��      4       ^4      9       ~�9      J       ^M      v       ^y             0�                           p      �       @<$��      �       P�      8       P9      n       Pn      y       0�y             @<$�                    P      X       UX      i       �U�                    P      ]       T]      i       �T�                   P      X       uX      a       �U#                                                                          `      �       U�      �       u�{��      4       U4      E       u�z�E      O       UO      `       u�{�`      �       U�      �       u�z��      �       U�      	       u�{�	      A       UA      R       u�z�R      �       U�      �       u�z��      �       U�      �       p�|��             u�|�             U             p�{�      (       u�{�(      7       U7      <       p�y�<      H       u�z�H      �       U�      �       u�z��      �       U�      �       p�{��      �       u�{��             U                                             �      �       P�      �       P�      �       P�      �       P             P1      2       PQ      R       Pq      r       P�      �       P�      �       P�      �       P�      �       P�      �       P�      �       P             P                    p�      y�       Uy�      z�       �U�                    p�      y�       Ty�      z�       �T�                    p�      y�       Qy�      z�       �Q�                    ��      ��       U��      ��       �U�                    ��      ��       T��      ��       �T�                    ��      ��       Q��      ��       �Q�                          P�      ��       U��       �       S �      &�       �U�&�      1�       U1�      k�       S                                  P�      ��       T��      ��       V��      ʞ       Tʞ      �       V�      &�       �T�&�      1�       T1�      G�       VG�      U�       TU�      k�       V                                  P�      ��       Q��      ��       ]��      Ξ       QΞ      �       ]�      &�       �Q�&�      1�       Q1�      G�       ]G�      Y�       QY�      k�       ]                                P�      ��       R��      ��       �R���      Ξ       RΞ      &�       �R�&�      1�       R1�      G�       �R�G�      Y�       RY�      k�       �R�                           P�      �       0�&�      =�       0�=�      ?�       P?�      E�       0�E�      G�       PG�      k�       0�                   ��      ��       V�      �       V                   ��      ��       0��      �       Q                  �      �       P                    ��      ��       T�      �       T                 �      �       V                     ��      ��       t��      ��       Q��      ��       t                          ��      $�       U$�      @�       ^@�      C�       �U�C�      Z�       UZ�      L�       ^                        ��      #�       T#�      C�       �T�C�      Y�       TY�      L�       �T�                    ��      1�       SC�      �       S                            �      1�       ]C�      �       ]�      �       U�      �       ]{�      �       U�      ��       ]                   �      :�       VC�      L�       V                    �      {�       ]��      L�       ]                 Ü      ˜       T                    ��      ��       P��      ˛       _                          {�      �       P�      E�       w {�      Ü       w ˜      �       w �      ��       w                       ˛      ��       P��      E�       _{�      ��       _                          �      �       P�      E�       S{�      �       P�      Ü       S˜      ߜ       S                 ��      L�       ]                  ��      Ü       } �˜      <�       } �                       ��      ��       t s "���      ��       T��      Ü       w s "�˜      ߜ       w s "�                  ��      Ü       ^˜      <�       ^                  ��      Ü       _˜      <�       _                        ��      ��       P��      Ü       ��˜      �       ���      ��       ��                 �      �       8�                      ߜ      �       S�      v�       Sv�      ~�       R                   .�      v�       s 
��4&3#�v�      ~�       r 
��4&3#�                   .�      v�       s ?
��#�v�      ~�       r ?
��#�                   .�      v�       1s ?
��#$1�v�      ~�       1r ?
��#$1�                    ��      ��       X)�      <�       X                      ��      ��       Y��      �       ���      1�       Y                      ��      ��       Q��      �       ���      �       Q                    ��      �       P�      ,�       t 2$u "                 �      1�       Q                        ��       P                    A      5A       U5A      F       �U�                        A      =A       T=A      `A       \`A      gA       �T�gA      F       \                        A      =A       Q=A      bA       ]bA      gA       �Q�gA      F       ]                    +A      ]A       SgA      F       S                    9A      ^A       VgA      F       V                    }A      �A       P�A      �A       P                      �A      �A       P�A      �B       ���B      �B       ��                                  B      B       0�B      *B       Q*B      GB       ��GB      MB       Q�B      �C       ���C      D       PD      ,D       ��,D      �E       w �E      F       w                                           OC      \C       0�\C      �C       w �C      �C       R�D      E       QE      6E       ��6E      IE       QlE      }E       R}E      �E       Q�E      �E       ���E      �E       Q�E      �E       R�E      �E       Q�E      	F       ��	F      F       Q                  �E      �E       x�                  �D      �D       ��                     9A      IA       ^gA      �B       ^�B      �B       ^                  KD      F       ^                       9A      IA       0�IA      TA       _TA      �A       0��A      B       PB      F       _                  OC      \C       ^                  iC      rC       ��                  �C      �C       ��                  �C      �C       P                  �E      �E       P                  �E      	F       P                    �>      0?       U0?      
A       �U�                      
?      >?       SH?      �?       S�?      
A       S                      "?      C?       ]H?      �?       ]�?      
A       ]                     "?      A?       \H?      �?       \�?      
A       \                    �?      �?       P�?      �@       _                      s?      w?       Pw?      �?       V�?      �?       V                              �?      �?       P�?      �?       ���?      �?       P�?      �?       Q�?      �?       ���?      �?       ^�?      
A       ��                      �?      �?       0��?      �@       w �@      �@       w �#��@      
A       w                           9@      B@       0�B@      R@       V�@      �@       P�@      �@       _�@      �@       v�                          �.      /       U/      }/       ^}/      �/       �U��/      0       ^0      0       �U�                    �.      �.       T�.      0       �T�                          �.      �.       Q�.      }/       V}/      �/       �Q��/      0       V0      0       �Q�                          �.      /       0�/      /       P/      }/       ]�/      0       ]0      0       T0      0       0�                      (/      F/       p ���/      �/       p ���/      �/       p ��                    //      }/       \�/      0       \                                /      /       0�/      _/       S_/      t/       Rt/      }/       S�/      �/       S�/      �/       R�/      �/       S�/      �/       P                                    ;/      F/       0�F/      W/       _W/      _/       �_/      }/       _�/      �/       0��/      �/       _�/      �/       ��/      �/       _�/      �/       0��/      �/       _                    �.      /       P/      0       ��                        �,      -       U-      .       \.      .       �U�.      �.       \                            �,      -       T-      t-       Vt-      .       �T�.      .       V.      �.       �T��.      �.       V                            �,      -       Q-      v-       Sv-      .       �Q�.      .       S.      �.       �Q��.      �.       S                         �,      c-       0�c-      g-       Pg-      �-       w .      �.       w �.      �.       0�                          -      2-       p ��2-      �-       ^.      �.       ^�.      �.       p ���.      �.       ^                          �-      �-       p ���-      �-        ���-      �-       P�-      �-       ��3.      3.        ��3.      G.       ��                                   r-      {-       0�{-      �-       S�-      �-       s��-      �-       s��-      �-       S�-      �-       s��-      �-       S.      (.       ](.      3.       S3.      N.       s�N.      l.       s�l.      .       S.      �.       s��.      �.       S                        �-      �-       0��-      �-       	��(.      3.       0�S.      l.       0�l.      �.       	��                     r-      {-       0�{-      �-       V.      �.       V                      -      {-       ].      .       ]�.      �.       ]                        p�      ��       U��      ��       ^��      ��       �U���      T�       ^                        p�      ��       T��      ��       V��      ��       �T���      T�       V                        p�      ��       Q��      ��       ]��      ��       �Q���      T�       ]                                          p�      ��       R��      ��       _��      ��       �R���      ��       _��      ��       �R���      ��       _��      #�       �R�#�      A�       _A�      ��       �R���      ��       _��      )�       �R�)�      A�       _A�      T�       �R�                                    ��      ��       0���      ��       P��      ��       S��      ,�       P,�      /�       S/�      I�       PI�      ��       S��      ��       S��      T�       S��      )�       SA�      T�       S                 �      Y�       v                    4�      H�       ��|�H�      Y�       XY�      Z�       ��|�                    4�      M�       ��{�M�      Y�       RY�      Z�       ��{�                4�      Z�       ]                 4�      Y�       v                       ��      ��       ^��      ��       ^��      ��       ^)�      A�       ^                     ��      ��       R��      ��       _��      ��       _)�      A�       _                     ��      ��       Q��      ��       ]��      ��       ])�      A�       ]                   ��      ��       V��      ��       V)�      A�       V                 ��      ��       U                	   ��      ��       u���      ��       P                
 ��      ��       u�                      ��      �       P�      ��       S��      ��       P)�      A�       S                 ��      �       \                3�      F�       ~� #�                3�      F�       ��}                   ?�      F�       QF�      F�      
 q r "#���                  ?�      F�       q ?&�F�      F�       R                e�      s�       ~� #�                e�      s�       ��~                   q�      s�       Ps�      s�      
 p q "#���                  q�      s�       p ?&�s�      s�       Q                          ��      O�       ]��      ��       ]��      #�       ]A�      b�       ]|�      ��       ]��      )�       ]                          ��      O�       \��      ��       \��      #�       \A�      b�       \|�      ��       \��      )�       \                            ��      ��       _��      ��       _��      #�       _A�      b�       _|�      ��       _��      )�       _                       �      G�       PG�      W�       ��{��      ��       P                             �      �       @<$��      O�       ��{��      ��       ��{��      #�       ��{A�      b�       ��{|�      ��       ��{��      )�       ��{                      �      G�       XG�      W�       ��{��      ��       X                      �      G�       RG�      W�       ��{��      ��       R                   �      �       �	p "��      �       P                   ��      ��       ]��      ��       ]��      �       }�                   ��      ��       z 
�����      �       z 
���                   ��      ��       _��      �       _                     ��      ��       0���      ��       P��      ��       0�                    ��      ��       0���      �       0��      �       �	p "�                  ��      ��       �	��      �       �	                   ��      ��       �	#���      )�       �	#�                         ��      ��       Y��      ��       Y$�      O�       Y��      ��       Y��      ��       ��{                             m�      ��       R��      ��       ��|��      ��       R��      +�       x� +�      O�       R]�      b�       R��      ��       R                    R�      ��       PA�      b�       P                    ��      ��       Q��      ��       �#h                    ��      ��       P��      ��       P                ��      �       ��{                 ��      ��       Y                   ��      �       Y�      �      
 p y "#���                  ��      �       y ?&��      �       P                $�      $�       ��{                $�      $�       _$�      $�       R                $�      $�       P                 O�      o�       \                        ��      ��       U��      0�       S0�      :�       �U�:�      a�       S                                  ��       �       T �      1�       V1�      :�       �T�:�      E�       TE�      q�       Vq�      ��       T��      ��       V��      ��       T��      a�       V                                      ��       �       Q �      :�       �Q�:�      E�       QE�      q�       �Q�q�      ��       Q��      ��       Z��      ��       �Q���      ��       Z��      ��       Q��      g�       ��g�      a�       �Q�                              ��      ��       R��       �       [:�      Q�       [Q�      q�       ��q�      ��       �R���      ��       [��      a�       �R�                                              ��       �       X �      :�       �X�:�      E�       XE�      q�       �X�q�      ��       X��      ��       ����      ��       �X���      ��       X��      ��       ����      ��       �X���      ��       ����      �       �X��      �       ���      ,�       �X�,�      a�       ��                   ��      3�       \:�      a�       \                   ��      7�       ^:�      a�       ^                    ��      �       P��      ��       P                                ��       �       { 	�� �      :�       �R	��:�      E�       { 	��E�      q�       �R	��q�      ��       { 	����      ��       �R	����      ��       { 	����      a�       �R	��                              ��      ��       P��       �       |�:�      E�       |�q�      ��       |���      ��       ��~��      ��       |���      a�       ��~                    ��      ��       _m�      ,�       _                                   ��      ��       1���      ��       { @&? $@M$.���      ��       ����      ��       1���      ��       0���      ��       ����      ��       1���      �       ���      �       1��      ,�       ��,�      a�       1�                    ��      ��       0�m�      ��       { @&? $@M$.��      �       { @&? $@M$.�                       ��      ��       0�y�      ��       ����      ��       ���      �       0�                           ��      0�       0�<�      ��       1���      ��       0���      ��       1���      ��       1���      �       0��      ,�       1�,�      a�       0�                     <�      Y�       0�Y�      ��       T��      ��       Q                Y�      w�       v�                Y�      w�       q 1$x "�0$0&�                   p�      w�       Pw�      w�      
 p r "#���                  p�      w�       p ?&�w�      w�       R                      ��      ��       { 	����      ��       { 	����      m�       �R	��,�      a�       �R	��                 ��      ��       T                          ��      ��       0���      ��       P��      }�       0�0�      ?�       P?�      V�       0�V�      m�       P,�      a�       0�                       ��      ��       { 	����      }�       �R	��?�      V�       �R	��,�      a�       �R	��                	     ��      �       _?�      V�       _��      a�       _                      ��      ��       P��      �       ����      a�       ��                     ��      �       ��?�      m�       ����      a�       ��                     *�      ��       v��?�      m�       v��,�      a�       v��                  ��      �       0���      \�       0�                  ��      �       ����      \�       ��                    ��      ��       U��      �       ����      \�       ��                     ��      ��       p��      ��       P��      �       �#                   �      }�       �R	��,�      ��       �R	��                     �      �       Q�      }�       V,�      ��       V                    �      }�       _,�      ��       _                    �      �       R�       �       ��,�      a�       ��                     �      1�       P�       �       0�h�      ��       P                     ��       �       r�� �      }�       ��#��,�      g�       r��g�      ��       ��#��                     ��       �       r�� �      }�       ��#��,�      g�       r��g�      ��       ��#��                 ��      ��       P                 ��      ��       Q                 ��      ��       1�                 ��      ��       R                 ��      ��       2�                 ��      ��       R                 ��      �       3�                 ��      �       R                  �      }�       V                  �      }�       R                     o�      o�       0�o�      v�       1�v�      }�       2�}�      }�       3�                 9�      \�       0�                 9�      \�       1�                 9�      \�       U                   9�      g�       u��g�      ��       ��#��                         ��      ��       0���      ��       R��      ��       Q��      �       0�C�      b�       0�                    ��      ��       P��      /�       v                 ��      ��       v�                ��      ��       q 1$x "�0$0&�                   ��      ��       P��      ��      
 p y "#���                  ��      ��       p ?&���      ��       Y                  Y�      q�       ]                                               b      b       Ub      �b       ]�b      �b       �U��b      �b       U�b      �e       ]�e      �e       �U��e      !r       ]!r      �t       S�t      �t       ]�t      u       Su      ru       ]ru      �u       S�u      �v       ]�v      w       Sw      �w       ]                                               b      Qb       TQb      �b       S�b      �b       �T��b      ^c       S^c      �d       �T��d      �e       S�e      �e       �T��e      �i       S�i      �l       �T��l      8p       S8p      u       �T�u      Uu       SUu      aw       �T�aw      pw       Spw      �w       �T�                                                             b      �b       Q�b      �b       V�b      �b       �Q��b      �b       Q�b      *d       V*d      �d       �Q��d      �e       V�e      �e       �Q��e      �i       V�i      �j       �Q��j      |l       ��}�1�|l      �l       �Q��l      !r       V!r      �t       ��}�1��t      �t       �Q��t      u       ��}�1�u      ru       Vru      w       ��}�1�w      @w       V@w      aw       ��}�1�aw      pw       Vpw      �w       ��}�1�                         b      ]b       R]b      �b       �R��b      �b       R�b      �w       �R�                                    rb      {b       R{b      �b       ��|�b      �b       ��|�b      �e       ��|�e      �j       ��|�l      !r       ��|�t      �t       ��|u      ru       ��|w      @w       ��|aw      pw       ��|                                 rb      {b       u#X#{b      �b       ��|�b      �e       ��|�e      �j       ��|�l      !r       ��|�t      �t       ��|u      ru       ��|w      @w       ��|aw      pw       ��|                       �b      �b       P�d      `e       0�`e      �e       P`g      �g       P                                           -b      �b       ^�b      �e       ^�e      �j       ^�j      |l       ��}�l      r       ^r      �t       ��}�t      �t       ^�t      u       ��}u      ru       ^ru      w       ��}w      @w       ^@w      aw       ��}aw      pw       ^pw      �w       ��}                                          2b      :b       P:b      b       ub      �b       }�b      �b       ��|�b      �b       u�b      �b       }�b      �e       ��|�e      �j       ��|�l      !r       ��|�t      �t       ��|u      ru       ��|w      @w       ��|aw      pw       ��|                                     2b      �b       0��b      �b       0��b      Fc       ��}Fc      �e       0��e      �e       1��e      `g       ��}`g      �g       0��g      �g       1��g      �i       ��}�i      �l       0��l      m       ��}m      u       0�u      Uu       ��}Uu      �w       0�                                                 2b      �b       0��b      �b       0��b      �d       _�d      �d       0��d      `e       1�`e      �e       _�e      �j       _�j      |l       ��}�l      r       _r      �t       ��}�t      �t       _�t      u       ��}u      ru       _ru      w       ��}w      @w       _@w      aw       ��}aw      pw       _pw      �w       ��}                                }i      �i       P�i      �i       ~��i      �i       ��}�l      �l       ~��l      !r       ��}u      ru       ��}w      @w       ��}aw      pw       ��}                          �j      |l       ��}�0$0&��l      �l      	 r 0$0&��l      �t       ��}�0$0&��t      u       ��}�0$0&�Uu      �w       ��}�0$0&�                          �j      |l       ��}�0$0&��l      �l      	 p 0$0&��l      �t       ��}�0$0&��t      u       ��}�0$0&�Uu      �w       ��}�0$0&�                          �j      |l       ��}m      m       Pm      �t       ��}�t      u       ��}Uu      �w       ��}                  .u      Ou       P                    �l      �l       Q�l      �l       P                             "n      -n       0�-n      Nn       QNn      Rn       q�Rn      ]n       q1$p "�#��n      �n       U�n      (o       Q(o      *o       t 1$p "bo      �o       0�aw      pw       0�                      ?m      um       Rum      �p       ��}aw      pw       ��}                            "n      9n       T9n      Nn       tP�Nn      an       Tbo      �o       Qaw      iw       Qiw      pw       T                       "m      �m       0��m      �m       P�m      �p       \aw      pw       \                       "m      �m       0��m      �m       P�m      jn       ��}iw      pw       ��}                     "m      �m       0��m      Fo       Piw      pw       P                   �q      !r       0�w      @w       0�                        s      s       [s      �s       ��|�t      �t       ��|ru      �u       ��|                               �q      !r       0�}r      �r       R�r      �r       0��r      s       ~�  "�'s      �s       R�t      �t       R�t      �t       ��|�u      v       Rw      @w       0�@w      Lw       R                                     �j      �j       V�q      !r       ��}�0$0&�!r      �r       V�r      �s       ��}�0$0&��s      �t       V�t      u       Vru      �u       ��}�0$0&��u      �v       V�v      w       Vw      @w       ��}�0$0&�@w      aw       V                    �q      !r       \w      @w       \                    �q      �q       Sw      @w       S                              �j      |l       ��}�q      �q       R�q      �q       }0�q      �t       ��}�t      u       ��}ru      aw       ��}pw      �w       ��}                            �j      |l       ��}�q      �q       R�q      �t       ��}�t      u       ��}ru      aw       ��}pw      �w       ��}                                        �j      |l       ���}���}��(!r      �r       ���}���}��(�r      �r      
 ]���}��0�r      �r       ]���}���}��(�r      �s       ]���}���}�\�� �s      �s       ]���}���}��(�s      �t       ���}���}��(�t      �t       ]���}���}��(�t      u       ���}���}��(ru      �u       ]���}���}�\�� �u      w       ���}���}��(@w      aw       ���}���}��(pw      �w       ���}���}��(                 �r      �r       ��|                 �r      s       ��|                     �s      �s       [�t      �t       [�t      �t       ��|                         !r      rr       ��}�0$0&��s      �t       ��}�0$0&��t      �t       ��}�0$0&��u      �u       ��}�0$0&��v      w       ��}�0$0&�                     �s      �s       R�t      �t       R�t      �t       ��|                         !r      rr       S�s      �t       S�t      �t       S�u      �u       S�v      w       S                        !r      [r       \�s      �s       \�t      �t       \�u      �u       \                   �s      �s       p 	���t      �t       p 	��                                 br      rr       \�s      �s      	 q  $ &��s      t       \=t      zt       \zt      ~t       |`�~t      �t       \�t      �t       \�v      �v       \w      w       \                                 fr      rr       ]�s      t      	 }  $ &�t      :t       ]St      �t       ]�t      �t       }`��t      �t       ]�t      �t       ]�v      �v      	 }  $ &�w      w       ]                       !r      'r       |�0$0&�'r      Gr       PGr      [r       |�0$0&��u      �u       P                       !r      Jr       QJr      Nr       PNr      fr       r���}�"��u      �u       Q                    !r      *r       ].r      _r       ]�u      �u       ]                  Ur      fr       P                  Xr      fr       Q                  t      �t       t                 t      �t       t                t      &t       t                 t      t       \                   t      &t       \&t      &t      
 p | "#���                  t      &t       | ?&�&t      &t       P                =t      Dt       t                  =t      Dt       ]Dt      Dt      
 p } "#���                  =t      Dt       } ?&�Dt      Dt       P                 ]t      �t       s                  ]t      �t       s #�                  �v      �v       ��|                  �v      �v       P                �v      �v       ��|                 �v      �v       \                   �v      �v       \�v      �v      
 q | "#���                  �v      �v       | ?&��v      �v       Q                       �j      |l       ��}�0$0&��u      �v       ��}�0$0&�@w      aw       ��}�0$0&�pw      �w       ��}�0$0&�                       �j      |l       ��}�0$0&��u      �v       ��}�0$0&�@w      aw       ��}�0$0&�pw      �w       ��}�0$0&�                         �j      |l       ]�u      �u       S�u      �v       ]@w      aw       ]pw      �w       ]                    �u      �v       s�@w      aw       s�                     Cl      El       0�El      Sl       QVl      {l       Q                      �j      �k       S�v      �v       Spw      �w       S                    �j      |l       Vpw      �w       V                     k      [k       } #�pw      �w       q��w      �w       } #�                  �k      Cl       ��}�0$0&�                  �k      Cl       ��}�0$0&�                    �k      &l       q�&l      Cl       }#�                  �k      Cl       }��                   }i      �i       V�i      �i       P                                           }i      �i       X�i      �i       ��}�i      �i       }���j      |l       }���l      �l       X�l      !r       }��!r      �t       s���t      u       s��u      !u       ��}!u      ru       }��ru      �u       s���u      �v       }���v      w       s��w      �w       }��                
       }i      �i       Q�i      �i       Q�l      �l       Q�l      �l       ��}                �p      �p       ��|                �p      �p       }�                    �p      �p       Q�p      �p      
 q r "#���                  �p      �p       q ?&��p      �p       R                #q      5q       ��|                #q      5q       }�                   .q      5q       Q5q      5q      
 q r "#���                  .q      5q       q ?&�5q      5q       R                �p      �p       ��|                �p      �p       }�                   �p      �p       Q�p      �p      
 q r "#���                  �p      �p       q ?&��p      �p       R                �p      q       ��|                �p      q       }�                   q      q       Qq      q      
 q r "#���                  q      q       q ?&�q      q       R                Kq      `q       ��|                Kq      `q       }�                   Yq      `q       R`q      `q      
 q r "#���                  Yq      `q       r ?&�`q      `q       Q                vq      �q       ��|                vq      �q       }�                   �q      �q       R�q      �q      
 q r "#���                  �q      �q       r ?&��q      �q       Q                       Fc      �d       ]�i      j       ]-j      �j       ]�t      �t       ]                        Jc      �d       \�i      j       \-j      �j       \�t      �t       \                           Jc      �c       0��c      d       Pd      �d       0��i      j       0�-j      �j       0��t      �t       0�                       Jc      �d       |� ��i      j       |� �-j      �j       |� ��t      �t       |� �                  Vc      �c       R                       3d      \d       |� \d      gd       Pgd      �d       pp��d      �d       P                            7d      Bd       t r "�Bd      �d       R�d      �d       t s "#@��i      j       t s "#@��j      �j       t s "#@��t      �t       t s "#@�                     7d      Jd       0�Jd      Vd       YVd      \d       p                     7d      Nd       0�Nd      Yd       XYd      \d       p                 7d      Nd       0�Nd      �d       1�                  \d      gd       p gd      rd       pp                   kd      rd       Qrd      rd      
 q z "#���                  kd      rd       q ?&�rd      rd       Z                   �d      �d       Q�d      �d      
 q z "#���                  �d      �d       q ?&��d      �d       Z                 -j      �j       0�                 -j      �j       |� �                 -j      �j       }��                ^f      mf       ��|                ^f      mf       }�                    kf      mf       Pmf      mf      
 p q "#���                  kf      mf       p ?&�mf      mf       Q                f      �f       ��|                f      �f       }�                   �f      �f       P�f      �f      
 p q "#���                  �f      �f       p ?&��f      �f       Q                �f      �f       ��|                �f      �f       }�                   �f      �f       P�f      �f      
 p q "#���                  �f      �f       p ?&��f      �f       Q                �f      �f       ��|                �f      �f       }�                   �f      �f       P�f      �f      
 p r "#���                  �f      �f       p ?&��f      �f       R                �f      g       ��|                �f      g       }�                   �f      g       Pg      g      
 p r "#���                  �f      g       p ?&�g      g       P                g      (g       ��|                g      (g       }�                   !g      (g       Q(g      (g      
 p q "#���                  !g      (g       q ?&�(g      (g       P                    �      �       0��             0�      "       q�                  �      �       0��             0�      "       q�                      �      �       0��      %       0�%      F       x q �U      W       x q �                     �      �       u #��             Q      \       u #�                             )      ])       U])      �*       S�*      �*       �U��*      1,       S1,      9,       �U�9,      y,       S                     )      8)       T8)      y,       �T�                  )      ")       u                       ?)      �*       V�*      2,       V9,      y,       V                           ?)      ])       u��])      �*       s���*      �*       �U#���*      1,       s��1,      9,       �U#��9,      y,       s��                     J)      �*       \�*      4,       \9,      y,       \                  �+      ,       P                   �*      �*       s�*      �*       P                  �*      ,       �^��                 �*      �*       \                 �*      �*       P                 �*      �*       3�                 �*      �*       U                 #+      �+       U                 #+      ?+       0�                 #+      ?+       3�                 #+      ?+       U                 #+      �+       u��                         F      KF       UKF      �G       \�G      �G       �U��G      TI       \                          KF      �F       T G      G       PG      �G       T�G      4I       T4I      OI       ��OI      TI       T                                      ;F      KF       ]KF      wF       XwF      |F       x�|F      �F       }��F      �F       X�F      (G       ](G      ;G       }�;G      �G       X�G      �G       X�G      �G       x��G      �G       ]�G      H       XH      H       x�H      "H       }�"H      PH       XPH      \H       x�\H      qH       XqH      �H       x��H      �H       x��H      �H       x��H      �H       ]�H      �H       X�H      �H       x��H      I       XI      TI       ]                    BF      �G       V�G      TI       V                    FF      �G       S�G      TI       S                      KF      �F       P G      �G       P�G      4I       P                           FF      KF       0�KF      �F       ^�F      �F       ��F      �F       _�F      �G       ^�G      I       ^I      TI       _                               �F      �F       @<$��F      �F       R�G      �G       @<$��G      �G       RdH      �H       @<$��H      �H       R�H      I       @<$�I      4I       R                             �F      �F       0��F      �F       Z�G      �G       0�dH      �H       0��H      �H       Z�H      I       0�I      4I       Z                                 �F      �F       @<$��F      �F       R�F      �F       U�G      �G       @<$��G      �G       UdH      �H       @<$��H      �H       U�H      I       @<$�I      ,I       U,I      4I       p(                             �F      �F       0��F      �F       Y�G      �G       0�dH      �H       0��H      �H       Y�H      I       0�I      4I       Y                           KF      VF       R_G      gG       2�gG      �G       R�G      �G       	�0y 0$0)( 	�#�@H      KH       RKH      PH       	�0y 0$0)( 	�#�                 0I      4I       U                                  p1      �1       U�1      �4       V�4      �4       U�4      �4       V�4      �4       �U��4      �4       U�4      �4       V�4      �4       U�4      .6       V                             *3      H3       P�3      �4       0��4      �4       P5      (5       P(5      y5       0�y5      �5       F��5      .6       0�                                                      �1      �1       R�1      2       r�"2      j2       S�2      )3       Z)3      v3       ���3      �3       Y�3      �3       T�3      4       U4      	4       T'4      A4       RA4      N4       XN4      |4       R|4      �4       X�4      �4       R�4      �4       R�4      �4       r��4      �4       R�4      �4       w (5      .5       T.5      =5       U=5      y5       Yy5      �5       Z�5      �5       R�5      �5       X�5      �5       R�5      6       X6      6       R6      .6       Y                    �1      �4       ]�4      .6       ]                    �1      �4       \�4      .6       \                    �1      �4       ^�4      .6       ^                     �3      �4       |� �(5      y5       |� ��5      .6       |� �                    �2      �4       S(5      .6       S                       j2      x2       0�x2      |2       �|2      �2       _�4      
5       0�                                       �3      �3       X�3      	4       P4      44       |� 44      \4       T\4      _4       t�_4      �4       T(5      y5       P�5      �5       T�5      �5       T�5      �5       t��5      6       T6      &6       X&6      .6       P                      �3      44       [(5      y5       [6      .6       [                             �3      �3       Q�3      �3       x �3      �3       p�3      �3       t �3      4       Q(5      y5       Q&6      .6       Q                    C5      b5       u &6      .6       u                      4      �4       Q�5      �5       Q�5      6       Q                      4      �4       Z�5      �5       Z�5      �5       q y "��5      �5         $ &4$q "�                          4      44       0�44      K4       Uh4      �4       U�5      �5       0��5      �5       U�5      �5       U                           �1      2       |� 2      2       X2      �2       Q�4      �4       X�4      �4       X�4      5       Q                          �1      �1       ~ 0$0&1$|� "��1      �1      
 p 1$|� "��1      �2       U�4      �4       X�4      �4       X�4      5       U                       �1      >2       P>2      a2       Ta2      j2       T�4      �4       P                           44      D4       0�D4      H4       RH4      N4       r �h4      |4       0�|4      �4       r ��8$r��!0$0&��4      �4       { 8$r��!0$0&��4      �4       { 8$x��!0$0&��4      �4       x~��8$x��!0$0&�                    44      T4       Pk4      �4       P                           �5      �5       0��5      �5       R�5      �5       r ��5      �5       0��5      �5       r ��8$r��!0$0&��5      �5       z 8$r��!0$0&��5      �5       z 8$x��!0$0&��5      �5       x~��8$x��!0$0&�                    �5      �5       P�5      6       P                    �       �        Q�              q�      "       q�"      9       q�9      P       q�P      p       Rp      q       u�                 �       q       u�                    �,      �,       U�,      �,       �U�                   �,      �,       u0�,      �,       U                          �,      �,       U�,      �,       V�,      �,       �U��,      �,       V�,      �,       �U�                    �,      �,       T�,      �,       �T�                    �,      �,       Q�,      �,       �Q�                          �,      �,       R�,      �,       \�,      �,       �R��,      �,       \�,      �,       �R�                    �,      �,       P�,      �,       P                    �,      �,       S�,      �,       S                        @       �        U�       �        S�       �        �U��       �        U                      @       �        T�       �        �T��       �        T                   @       `        u �       �        u                    @       �        0��       �        w �       �        0�                   @       �        0��       �        �`�       �        0�                  �       �        P                      J      9J       U9J      �J       S�J      �J       �U�                      J      J       TJ      �J       ]�J      �J       �T�                  1J      �J       V                  �J      �J       P                 1J      �J       \                    ZJ      aJ       PaJ      �J       ^                  ZJ      nJ       XnJ      oJ       �L�                    ZJ      fJ       �H�fJ      nJ       RnJ      oJ       �H�                ZJ      oJ       ]                ZJ      oJ       V                              `�      ��       U��      ��       T��      ��       �U���      �       U�      
�       T
�      �       �U��      V�       U                                      `�      g�       Tg�      ��       P��      ��       �T���      
�       P
�      �       �T��      5�       P5�      6�       �T�6�      E�       PE�      F�       �T�F�      U�       PU�      V�       �T�                          `�      ��       Q��      ��       �Q���      
�       Q
�      �       �Q��      V�       Q                              `�      ��       R��      ��       R��      ��       r 9!���      ��       x 9!���      ��       X��      ��       R��      
�       R�      V�       R                             `�      ��       U��      ��       T��      ��       �U���      �       U�      
�       T
�      �       �U��      V�       U                                      c�      g�       Tg�      ��       P��      ��       �T���      
�       P
�      �       �T��      5�       P5�      6�       �T�6�      E�       PE�      F�       �T�F�      U�       PU�      V�       �T�                                    g�      ��       T��      ��       u��      ��       t��      ��       T��      �       u�      
�       t�      �       u�      $�       T$�      ,�       u,�      V�       T                          �      �       U�      &       S&      '       �U�'      B       SB      C       �U�                        �             T      '       �T�'      4       T4      C       �T�                    �             U'      4       U                       �      &       S&      '       �U�'      B       SB      C       �U�                     �             0�      '       P'      C       0�                              u�                                    s�             Q      &       s�&      '       �U#�                              $        U$       .        �U�.       3        U                              $        T$       .        �T�.       3        T                              $        Q$       .        �Q�.       3        Q                                $        R$       -        S-       .        �R�.       3        R                             $        U$       .        �U�.       3        U                             $        P.       2        P2       3        u�                    `I      mI       UmI      �I       X                  `I      oI       T                    cI      mI       UmI      �I       X                   cI      mI       u� mI      �I       x�                  �I      �I       Q                      0      E       TE      K       PK      X       T                        0      @       Q@      E       �Q�E      P       QP      X       �Q�                  W      X       P                          �I      �I       U�I      �I       �U��I      �I       U�I      �I       �U��I      J       U                              �I      �I       T�I      �I       Q�I      �I       �T��I      �I       T�I      �I       �T��I      
J       T
J      J       �T�                      �I      �I       Q�I      �I       �Q��I      J       Q                          �I      �I       R�I      �I       �R��I      �I       R�I      �I       �R��I      J       R                      �I      �I       X�I      �I       �X��I      J       X                    �I      
J       T
J      J       �T�                  �I      J       X                  �I      J       R                  �I      J       Q                  �I      J       U                            �J      /K       U/K      aK       \aK      hK       �U�hK      �K       U�K      �K       \�K      �K       U                          �J      /K       T/K      hK       �T�hK      �K       S�K      �K       �T��K      �K       S                          �J      /K       Q/K      hK       �Q�hK      �K       Q�K      �K       �Q��K      �K       Q                    �J      �J       R�J      �K       �R�                          �J      /K       X/K      hK       �X�hK      �K       X�K      �K       �X��K      �K       X                    K      RK       0�RK      WK       1�                           �J      /K       U/K      aK       \aK      hK       �U�hK      �K       U�K      �K       \�K      �K       U                    hK      �K       �R��K      �K       �R�                      hK      �K       X�K      �K       �X��K      �K       X                      hK      �K       Q�K      �K       �Q��K      �K       Q                      hK      �K       S�K      �K       �T��K      �K       S                      hK      �K       U�K      �K       \�K      �K       U                    �K      �K       0��K      �K       1�                �K      �K       ^                �K      �K       ]                    �K      �K       S�K      �K       Q�K      �K       s�                �K      �K       \                       L      L       UL      <L       �U�<L      fL       U                       L      L       TL      <L       �T�<L      fL       T                       L      *L       Q*L      <L       �Q�<L      fL       Q                  <L      fL       U                  <L      fL       R                  <L      fL       X                  <L      fL       Q                  <L      fL       T                 pL      �L       t $ &#04$u "#�                        �M      �M       Q�M      �M       �Q��M      �M       Q�M      �M       �Q�                           �M      �M      	 p t "	���M      �M       q t "# 	���M      �M       �Qt "# 	���M      �M       P�M      �M       �Qt "# 	���M      �M       P                  �M      �M       U                    �M      �M       Q�M      �M       �Q�                  �M      �M       T                         �M      �M      
 p t 	���M      �M       q t # 	���M      �M       �Qt # 	���M      �M       P�M      �M       �Qt # 	��                        �M      �M       Q�M      �M       �Q��M      N       QN      N       �Q�                      �M      �M       p ��M      �M       P�M      �M       �Qt "	�# �                  �M      N       U                    �M      N       QN      N       �Q�                  �M      N       T                    N      N       PN      N       r q �                           N      .N       Q.N      7N       �Q�7N      HN       QHN      KN       PKN      ZN       �Q�                         %N      .N      	 t q "	��.N      2N      
 t �Q"	��2N      6N       P6N      7N      
 t �Q"	��YN      ZN       P                  7N      ZN       U                      7N      HN       QHN      KN       PKN      ZN       �Q�                  7N      ZN       T                         7N      HN      
 q t 	��HN      KN      
 p t 	��KN      RN       �Qt 	��RN      YN       PYN      ZN       �Qt 	��                        `N      qN       QqN      zN       �Q�zN      �N       Q�N      �N       �Q�                           iN      lN      	 p t "	��lN      qN       q t "#?	��qN      uN       �Qt "#?	��uN      yN       PyN      zN       �Qt "#?	���N      �N       P                  zN      �N       U                    zN      �N       Q�N      �N       �Q�                  zN      �N       T                         zN      �N      
 p t 	���N      �N       q t #?	���N      �N       �Qt #?	���N      �N       P�N      �N       �Qt #?	��                        �N      �N       Q�N      �N       �Q��N      �N       Q�N      �N       �Q�                           �N      �N      	 p t "	���N      �N       q t "#	���N      �N       �Qt "#	���N      �N       P�N      �N       �Qt "#	���N      �N       P                  �N      �N       U                    �N      �N       Q�N      �N       �Q�                  �N      �N       T                         �N      �N      
 p t 	���N      �N       q t #	���N      �N       �Qt #	���N      �N       P�N      �N       �Qt #	��                    �N      O       QO      2O       �Q�                    O      O       PO      O       p x "�O      O       r t "q x "�                  O      2O       �Q�                  O      2O       T                  O      2O       U                    $O      1O       P1O      2O       r q u��                        @O      fO       QfO      uO       �Q�uO      }O       Q}O      �O       �Q�                      mO      mO       PmO      pO       p x "�pO      tO       PtO      uO       u�t "x �Q"r r x "�                    uO      }O       Q}O      �O       �Q�                  uO      �O       T                  uO      �O       U                    �O      �O       P�O      �O       u�t u��Q"r r u��                   P      #P       T                   P      #P       U                      0P      �P       T�P      �P       �T��P      �P       T                    wP      �P       Q�P      �P       Q                    wP      �P       X�P      �P       X                    wP      �P       R�P      �P       R                    wP      �P       T�P      �P       T                    wP      �P       U�P      �P       U                        �P      QQ       UQQ      \R       S\R      fR       �U�fR      �S       S                     �P      �P       0��P      JQ       TfR      �R       T�R      �R       T                              gQ      �Q       _R      /R       P�R      �R       _AS      FS       PFS      SS       _{S      �S       P�S      �S       _                        �Q      �Q       P�Q      7R       ^�R      �R       ^bS      oS       ^                 �P      �P       u�                    TQ      [Q       T[Q      cQ       u�v "�                 TQ      cQ       P                     �R      �R       p 3�#<3$s "#�R      �R       s��3�#<3$s "#FS      oS       s��3�#<3$s "#                   �R      �R       _FS      SS       _                   �R      �R       SFS      oS       S                      �R      �R        q "��R      �R       ^FS      SS        q �SS      oS       _                      �R      �R       Q�R      =S       s�v "�oS      zS       s�v "�                     �R      S       PS      =S       s��
��4$s� "�oS      zS       P                       S      S       p t "#��@& $ &���S      #S      ( p t "#��@& $ &��q u "#��@& $ &��#S      +S      ; s�v "�z  $ &x p "#��@& $ &��q u "#��@& $ &��+S      2S      Y s�v "�z  $ &x p "#��@& $ &��s�v "#�y  $ &s�� $ &u "#��@& $ &��2S      =S      z s�v "�z  $ &x p "#��@& $ &��s�v "#�y  $ &s�� $ &s�v "#�y  $ &s�� $ &?&"#��@& $ &��                �R      S       X                    �R      �R       t z ��R      	S       T	S      S       s�v "�z �                   	S      S       TS      S      
 p t "#���                  	S      S       t ?&�S      S       P                  S      S       QS      S      
 q u "#���                  S      S       q ?&�S      S       U                {S      �S       s�                 {S      �S       P                   �S      �S       P�S      �S      
 p q "#���                  �S      �S       p ?&��S      �S       Q                        �S      �S       U�S      �S       P�S      �S       [�S      oU       �U�                    �S      �S       T�S      oU       ��                                �S      �S       Q�S      �S       ]�S      T       X6T      >T       Z>T      zT       ���T      U       XFU      jU       XjU      oU       Z                              �S      �S       R�S      T       Z6T      >T       X>T      zT       ���T      U       ZFU      gU       ZgU      oU       P                      �S      �S       X�S      �T       ^�T      oU       ^                          �S      �S       Y�S      >T       Y>T      zT       ���T      U       YFU      oU       Y                    hT      T       TT      �T       ��U      U       ��                 �S      �S       0�                          �T      �T       P�T      �T       PU      "U       P"U      AU       q AU      FU       P                         6T      kT       \kT      �T       S�T      aU       SaU      jU       x  $ &4$~ "jU      oU       z  $ &4$~ "                           6T      cT       ScT      nT       QnT      �T       \�T      ^U       \^U      gU       z  $ &4$~ "gU      oU       p  $ &4$~ "                         6T      >T       Q>T      zT       w �T      U       x  $ &4$y "FU      jU       x  $ &4$y "jU      oU       z  $ &4$y "                     �T      U       z  $ &4$y "FU      gU       z  $ &4$y "gU      oU       p  $ &4$y "                         6T      ZT       _ZT      zT       ]�T      U       x  $ &4$y "x  $ &4$~ "�FU      jU       x  $ &4$y "x  $ &4$~ "�jU      oU       z  $ &4$y "z  $ &4$~ "�                         6T      WT       ]WT      zT       R�T      U       z  $ &4$y "z  $ &4$~ "�FU      gU       z  $ &4$y "z  $ &4$~ "�gU      oU       p  $ &4$y "p  $ &4$~ "�                    hT      zT       PU      U       0�                   U      "U       p s �"U      )U       P                   )U      0U       P0U      0U      
 p { "#���                  )U      0U       p ?&�0U      0U       [                          �w      �w       T�w      �x       ]�x      �x       �T��x      hy       ]hy      yy       T                      �w      �w       Q�w      �w       P�w      yy       �Q�                      �w      �w       R�w      hy       �R�hy      yy       R                    �w      �w       Xhy      yy       X                    �w      �w       q 1$z "�hy      yy       q 1$z "�                           �w      �w       0��w      {x       _{x      �x       ��x      �x       _�x      hy       _hy      yy       0�                         �w      �w       0��w      Zx       \Zx      ix       |��x      Ly       \Ly      Zy       0�Zy      hy       \                         �w      �w       0��w      �w       R�x      �x       RLy      Zy       Rhy      yy       0�                   �x      �x       p s "#��@& $ &��x      �x       s ?&s "#��@& $ &�                     rx      wx       ��~ "1$z "�0$0&@$�wx      {x        ������"1$z "�0$0&@$�{x      �x       ������"1$z "�0$0&@$�                           �w      �w       @<$��w      Zx       S�x      y       S&y      4y       SLy      Zy       @<$�Zy      hy       S                      �w      �w       ~ 2$p "�w      �w       ~ 2$x"Ly      Zy       ~ 2$x"                    �w      �x       V�x      hy       V                  �x      �x       P                    rx      wx       ��~ "1$z "�0$0&@$�wx      {x        ������"1$z "�0$0&@$�{x      �x       ������"1$z "�0$0&@$�                 rx      �x       S                   �x      �x       S�x      �x      
 p s "#���                  �x      �x       s ?&��x      �x       P                        �y      �y       U�y      az       ^az      dz       �U�dz      <{       ^                          �y      �y       T�y      z       Sz      dz       �T�dz      |z       S|z      <{       �T�                        �y      �y       Q�y      ]z       \]z      dz       �Q�dz      <{       \                    �y      �y       R�y      �y       �R�                    �y      �y       X�y      �y       �X�                    �y      Zz       Sdz      <{       S                        �y      �y       Y�y      �y       P�y      z       Ydz      wz       Y                        �y      z       Zz      Uz       ��dz      |z       Z�z      <{       ��                    �y      _z       ]dz      <{       ]                        �y      z       Qz      Uz       _dz      �z       Q�z      <{       _                     �y      z       _z      z       Vdz      �z       _                            �y      �y       X�y      z       [z      Yz       w Yz      dz       ��dz      �z       [�z      <{       w                     �y      z       Rdz      �z       R                        �y      z       Xz      Uz       w  �dz      �z       X�z      <{       w  �                        �y      z       0�z      Uz       Z�z      {       Z#{      <{       P                          �y      z       0�z      Uz       [�z      �z       [�z      �z       1��z      {       [{      <{       1�                        z      2z       P<z      Uz       P�z      �z       P�z      {       P                �z      �z       Z                �z      �z       ~v "y �                   �z      �z       P�z      �z      
 p { "#���                  �z      �z       p ?&��z      �z       [                  wz      �z       Y                              `~      q~       Uq~      �~       S�~      �~       �U��~             S      #       �U�#      <       S<      B       �U�                                `~      �~       T�~      �~       \�~      �~       �T��~      �~       T�~      "       \"      #       �T�#      A       \A      B       �T�                             `~      q~       Uq~      �~       S�~      �~       �U��~             S      #       �U�#      <       S<      B       �U�                             `~      �~       0��~      �~       P�~      �~       V�~      �~       0��~      �~       V#      4       P4      ;       V                 w~      �~       U                 w~      �~       u�                    �~      "       \"      #       �T�                    �~             S      #       �U�                      �~      �~       P�~              V       #       P                  �~      �~       Q                        P      v       Tv      z       �T�z      �       T�      �       ��                          P      �       Q�      �       ]�      ��       �Q���      ̀       ]̀      �       �Q�                        P      m       Rm      ��       ^��      ��       �R���      �       ^                   P      �       U�      �       ��                    e      ��       V��      �       V                                       z      �       0��      �       _�      �       ��      �       _�      �       ��      "�       ��@�      ��       ]��      ̀       _̀      �       ]�      �       }��      �       ]�      �       S�      �       0�                          @�      u�       1�u�      ��       T��      ��       X��      ��       T̀      ڀ       T                       z      �       S�      �       sP��      �       S��      ̀       S                        @�      ��       \̀      �       \�      �       |p��      �       \�      �       ��#8                          �      �       U�      �       P�      �        3$} "�      �       U��      ��       U                      ��      ��       U��      ՚       S՚      ך       �U�                      ��      ��       T��      ֚       V֚      ך       �T�                    ��      ��       Q��      ך       �Q�                  ��      ך       P                  ��      К       �Q�                  ��      К       V                  ��      К       S                            ��      ן       Uן      ��       ^��      ��       u�~���      ��       �U���      ��       U��      ��       ^                   ��      ��       u�	��      ��       u�	                          ��       S��      ��       S                    ɟ      ��       V��      ��       V                      ן      �       _��      �       P�      �       _                  �      �       P                        �      ��       ^��      ��       u�~���      ��       �U���      ��       ^                       �      ��       ^��      ��       u�~���      ��       �U���      ��       ^                            ��      ��       U��      ��       \��      ��       �U���      �       \�      �       U�      �       �U�                            ��      ��       T��      ��       V��      ��       �T���      �       V�      �       T�      �       �T�                        ��      ��       P��      ��       S��      Ы       PЫ      �       S                      ��      �       V�      �       T�      �       �T�                      ��      �       \�      �       U�      �       �U�                  «      Ы       U                  ѫ      ٫       P                  ݫ      �       P                                 �      �       U�      1�       V1�      2�       �U�2�      X�       VX�      Y�       �U�Y�      k�       Vk�      l�       �U�l�      ~�       V                   �      �       T                           �      A�       QA�      l�       �Q�l�      u�       Qu�      {�       U{�      ~�       �Q�                     �      �       R�      ~�       �R�                               �      �       U�      1�       V1�      2�       �U�2�      X�       VX�      Y�       �U�Y�      k�       Vk�      l�       �U�l�      ~�       V                  ;�      ~�       �T�                    ;�      A�       Pl�      {�       P                            ;�      ?�       U?�      A�       QA�      l�       �Q�l�      u�       Qu�      {�       U{�      ~�       �Q�                          ;�      X�       VX�      Y�       �U�Y�      k�       Vk�      l�       �U�l�      ~�       V                          A�      V�       PY�      i�       Pi�      k�       v� k�      l�       �U#x|�      ~�       P                 ?�      A�       Q                     l�      u�       Qu�      {�       U{�      ~�       �Q�                      ��      ��       U��      ��       u ��      Ҭ       �U�                    ��      ��       T��      Ҭ       �T�                            �      :�       U:�      E�       �U�E�      e�       Ue�      |�       �U�|�      ��       U��      ��       �U�                            �      #�       T#�      E�       �T�E�      ^�       T^�      |�       �T�|�      }�       T}�      ��       �T�                            �       �       Q �      E�       �Q�E�      ^�       Q^�      |�       �Q�|�      }�       Q}�      ��       �Q�                        �      p�       Rp�      t�       Qt�      |�       �R�|�      ��       R                              �      :�       Y:�      =�       P=�      E�       U^�      e�       Yl�      t�       U}�      ��       Y��      ��       U                          &�      4�       Q4�      E�       Y^�      e�       Ql�      t�       T}�      ��       Q��      ��       Y                   4�      E�       Q��      ��       Q                                �      �       X�       �       q 
��4$u�"� �      :�       �Q
��4$u�"�:�      E�       �Q
��4$�U#�"�^�      e�       �Q
��4$u�"�e�      t�       �Q
��4$�U#�"�}�      ��       �Q
��4$u�"���      ��       �Q
��4$�U#�"�                                �      �       P�      #�       t 
��4$u�"�#�      :�       �T
��4$u�"�:�      E�       �T
��4$�U#�"�^�      e�       �T
��4$u�"�e�      t�       �T
��4$�U#�"�}�      ��       �T
��4$u�"���      ��       �T
��4$�U#�"�                           �      :�       u�:�      E�       �U#�E�      e�       u�e�      t�       �U#�|�      ��       u���      ��       �U#�                        :�      E�       Rl�      p�       Rp�      t�       Qt�      |�       �R���      ��       R                        :�      E�       Rl�      p�       Rp�      t�       Qt�      |�       �R���      ��       R                      :�      E�       Yl�      t�       T��      ��       Q��      ��       Y                        :�      =�       P=�      E�       Ul�      t�       U��      ��       Y��      ��       U                    E�      ^�       T|�      }�       T                    E�      ^�       Q|�      }�       Q                    E�      ^�       R|�      }�       R                    E�      ^�       U|�      }�       U                         %      (%       U(%      K%       VK%      P%       �U�P%      n%       V                         %      $%       T$%      J%       SJ%      P%       �T�P%      n%       S                         %      (%       Q(%      M%       \M%      P%       �Q�P%      n%       \                      ,%      0%       P0%      O%       ]P%      n%       ]                    `%      d%       Pd%      n%       Q                 �      (       U                    �Y      �Y       U�Y      p^       �U�                                �Y      �Y       T�Y      �\       S�\      �\       �T��\      k]       Sk]      v]       �T�v]      �]       S�]      �]       �T��]      p^       S                          �Y      �Y       Q�Y      -Z       V-Z      ]]       �Q�]]      o]       Vo]      p^       �Q�                    �Y      �Y       R�Y      p^       �R�                    �Y      �Y       X�Y      p^       �X�                               �Y      �Y       T�Y      �\       S�\      �\       �T��\      k]       Sk]      v]       �T�v]      �]       S�]      �]       �T��]      p^       S                                          Z      :Z       P:Z      \       ]\      \       P\      e\       0�e\      m\       Pm\      �\       0��\      �\       V�\      ]]       ]v]      �]       ]�]      �]       0��]      �]       6��]      �]       P�]      1^       ]1^      p^       0�                           �Y      �Y       P�Y      >\       \�\      q]       \v]      �]       \�]      �]       \�]      1^       \                             �Y      �Y       P�Y      �\       ^�\      ]]       ^]]      n]       Pn]      v]       �T#�v]      �]       ^�]      p^       ^                               �Y      �Y       t���Y      �\       s���\      �\       �T#���\      k]       s��k]      v]       �T#��v]      �]       s���]      �]       �T#���]      p^       s��                               �Y      �Y       t���Y      �\       s���\      �\       �T#���\      k]       s��k]      v]       �T#��v]      �]       s���]      �]       �T#���]      p^       s��                   �Y      �Y       t��Y      �Y       U                            �Y      �Y       P�Y      >\       \�\      q]       \v]      �]       \�]      �]       \�]      1^       \                       3Z      �\       S�\      ]]       Sv]      �]       S�]      p^       S                          �Z      	[       Q2]      @]       Q@]      D]       q�D]      P]       QP]      X]       q�X]      ]]       Q�]      ^       Q                     �Z      	[       R2]      ]]       R�]      ^       R                   �Z      �Z       1��]      ^       0�                     1\      �\       S�]      �]       S1^      p^       S                      >\      �\       \�]      �]       \1^      p^       \                       }\      �\       0��\      �\       U�]      �]       0��]      �]       U1^      O^       0�O^      T^       UT^      k^       0�k^      p^       U                        0      X       UX      w       Sw      y       �U�y      �       U                       0      X       UX      w       Sw      y       �U�y      �       U                  P      x       V                     P      X       u��X      w       s��w      y       �U#��                   �      w       s��w      y       �U#��                      @      i       Ui      �       S�      �       �U�                      J      ]       P]      i       ui      m       s                  Q      �       V                  n      x       P                  y      �       P                      �E      �E       U�E      F       SF      #F       �U�                      �E      �E       T�E      "F       \"F      #F       �T�                     �E      �E       U�E      F       SF      #F       �U�                    �E      �E       P�E       F       V                      0F      ;F       U;F      wF       SwF      xF       �U�                     0F      ;F       U;F      wF       SwF      xF       �U�                   0F      bF       0�bF      rF       P                    CF      EF       PEF      aF       R                  MF      aF       P                                        pL      �L       U�L      �M       ^�M      N       �U�N      O       ^O      )O       �U�)O      _U       ^_U      ]V       ��y]V      2W       ^2W      BW       ��yBW      �W       ^�W      �W       ��y�W      �W       �U��W      �Y       ^                     �L      uN       SuN      N       ��y�N      �Y       S                                       pL      �L       u���L      �M       ~���M      N       �U#��N      O       ~��O      )O       �U#��)O      _U       ~��_U      ]V       ��y#��]V      2W       ~��2W      BW       ��y#��BW      �W       ~���W      �W       ��y#���W      �W       �U#���W      �Y       ~��                                       pL      �L       u���L      �M       ~���M      N       �U#��N      O       ~��O      )O       �U#��)O      _U       ~��_U      ]V       ��y#��]V      2W       ~��2W      BW       ��y#��BW      �W       ~���W      �W       ��y#���W      �W       �U#���W      �Y       ~��                                  �L      �M       VN      O       V)O      �R       V]V      zV       V�V      �V       V�V      2W       ��yBW      �W       VNX      Y       ��yY      �Y       V                  �S      �S       0�                 X      *X       ~�                                &U      �U       0��U      �U       ��y�U      �U       \�U      �U       p��U      ]V       ��y�1�2W      BW       ��y�1��W      �W       ��yY      Y       0�                        �U      �U       0��U      �U       |��U      V       \2W      =W       |�                        &U      ]V       0�2W      BW       0��W      �W       0�Y      Y       0�                          &U      �U       0��U      XV       ��y2W      BW       ��y�W      �W       ��yY      Y       0�                      �U      �U       V�U      6V       V2W      BW       V                        �U      �U       ]�U      ]V       ]2W      BW       ]�W      �W       ]                                       �L      �L       U�L      �M       ^�M      N       �U�N      O       ^O      )O       �U�)O      _U       ^_U      ]V       ��y]V      2W       ^2W      BW       ��yBW      �W       ^�W      �W       ��y�W      �W       �U��W      �Y       ^                   �L      �L       ��y��L      �L       S                                 �L      �M       VN      O       V)O      �R       V]V      zV       V�V      �V       V�V      2W       ��yBW      �W       VNX      Y       ��yY      �Y       V                         �L      M       RM      �M       _N      O       _)O      PO       _kO      �O       _BW      �W       _                       �L      �M       \N      O       \)O      PO       \kO      �O       \BW      �W       \                       �L      �M       SN      O       S)O      PO       SkO      �O       SBW      �W       S                   �M      iN       SO      )O       S                   �M      iN       SO      )O       S                  �M      )N       V                   =N      iN       SO      )O       S                   =N      iN       VO      )O       V                           P      �R       V]V      zV       V�V      �V       V�V      2W       ��yNX      Y       ��yY      �Y       V                     P      QS       S]V      %W       SNX      Y       SY      �Y       S                       %P      NP       \NP      TP       ��{�V      %W       \NX      Y       \                         5P      �R       _]V      zV       _�V      %W       _NX      �X       _Y      �Y       _                               NP      TP       RTP      �P       \�P      �P       |v��P      �P       P�P      Q       PQ      2Q       s @Q      �R       ]mV      zV       \Y      �Y       ]                          RP      �P       P�P      ;Q       \@Q      �R       \]V      qV       \qV      zV       PY      �Y       \                      [Q      }Q       P}Q      �Q       ��y#Y      (Y       P                  �Q      �Q       P                     �V      �V       P�V      %W       ��yNX      Y       ��y                                     U        �$       ��                                        -        T-       "!       _"!      #!       �T�#!      $       _$      %$       U%$      ($       _($      .$       U.$      �$       _                            -        Q-       �$       �Q�                            -        R-       �$       �R�                                       -        T-       "!       _"!      #!       �T�#!      $       _$      %$       U%$      ($       _($      .$       U.$      �$       _                     +       !       S!      #!       �Q�R"�#!      �$       S                               K        0�K       !       V#!      �!       V�!      �!       ^�!      �$       V                                   K        0�K       �        \�       !       \#!      �!       \�!      j"       \�#      �#       \                                 K       �        ^�       !       ^#!      �!       ^�!      �!       ~s��!      j"       ^j"      �#       \�#      �#       ^�#      �#       \�#      �$       \                      �"      �"       Q�"      �#       ���#      �$       ��                            �"      �#       ^�#      $       ^$      %$       T%$      ($       ^($      .$       T.$      �$       ^                    �"      �"       X�"      9#       ��                              #      <#       P<#      �#      
 ��1#��#      �#      
 ��1#��#      $      
 ��1#�$      %$      
 u��1#�($      .$      
 u��1#�1$      �$      
 ��1#�                            F#      �#       ^�#      �#       ^�#      $       ^$      %$       T%$      ($       ^($      .$       T.$      �$       ^                            F#      �#       _�#      �#       _�#      $       _$      %$       U%$      ($       _($      .$       U.$      �$       _                    F#      �#       ���#      �#       ���#      �$       ��                     �#      �#       P&$      ($       P/$      1$       P                                      $      $       ���$      %$       Q($      .$       QA$      H$       ���H$      J$       Q[$      g$       ���g$      k$       Q�$      �$       Q�$      �$       Q�$      �$       ����$      �$       Q�$      �$       ����$      �$       Q�$      �$       ����$      �$       Q                                  $      $       0�$      %$       R($      .$       RA$      J$       0�[$      i$       0�i$      k$       R�$      �$       0��$      �$       0��$      �$       0��$      �$       0��$      �$       R�$      �$       0��$      �$       R                                R#      a#       Qa#      �#       P�#      �#       P�#      $       P1$      6$       PJ$      p$       P�$      �$       P�$      �$       P                            �&      �&       U�&      �*       \�*      �*       �U��*      1+       \1+      8+       �U�8+      7-       \                            �&      �&       T�&      �*       ^�*      �*       �T��*      5+       ^5+      8+       �T�8+      7-       ^                           �&      �&       T�&      �*       ^�*      �*       �T��*      5+       ^5+      8+       �T�8+      7-       ^                                   �&      �&       t���&      '       ~��'       '       P '      �*       ���*      �*       ~���*      �*       �T#���*      +       ��+      5+       ~��5+      8+       �T#��8+      7-       ��                                   �&      �&       t���&       '       ~�� '      ,'       P,'      �*       ���*      �*       ~���*      �*       �T#���*      +       ��+      5+       ~��5+      8+       �T#��8+      7-       ��                                     �&      �&       t���&      ,'       ~��,'      9'       P9'      �*       ���*      �*       ~���*      �*       �T#���*      +       ��+      5+       ~��5+      8+       �T#��8+      [+       P[+      7-       ��                      �&      �&       P�&      �&       t �&      7-       ��~                   +      %+       3�*-      7-       P                    �&      �&       P�&      7-       ��~                                   �&      9'       ]Z'      �'       _�'      #(       �#(      =(       Q=(      �(       �^)      "*       _�*      �*       ��*      +       _8+      I+       ]�+      �+       _�+      �+       ~                      �&      �)       S�*      %+       S8+      ,       S                      I'      �*       ]�*      +       ]�+      7-       ]                        �&      �&       P�&      �*       V�*      +       V8+      7-       V                           �&      I'       0�I'      �(       ���(      �*       ���*      +       ��8+      �+       0��+      7-       ��                         �&      I'       0�I'      �*       ���*      +       ��8+      �+       0��+      7-       ��                     �'      (         x "�(      #(      
   ��~�"�#(      7(      	 ��~�q �                     �(      �(       0��(      �(       P�(      U)       _U)      ^)       0�                 �)      �*      
 �1H     �                                @-      b-       Ub-      �/       V�/      �/       �U��/      0       V0      (0       �U�(0      70       V70      @0       �U�@0      z0       V                                  @-      i-       Ti-      �/       _�/      �/       �T��/      �/       U�/      '0       _'0      (0       �T�(0      ?0       _?0      @0       �T�@0      z0       _                                 @-      i-       Ti-      �/       _�/      �/       �T��/      �/       U�/      '0       _'0      (0       �T�(0      ?0       _?0      @0       �T�@0      z0       _                                 @-      i-       t��i-      �/       ���/      �/       �T#���/      �/       u���/      '0       ��'0      (0       �T#��(0      ?0       ��?0      @0       �T#��@0      z0       ��                        _-      �/       ^�/      %0       ^(0      =0       ^@0      z0       ^                              �-      �-       P�-      �-       ���-      �-       Q�-      �/       ��(0      -0       ��@0      H0       QH0      Q0      	 r 3&�                      .      ).       0�).      �/       \(0      -0       \                    g-      i-       Pi-      z0       ��                         ).      �.       S/      /       P/      �/       S�/      �/       S(0      -0       S                       ).      I.       0�I.      M.       PM.      �.       ]�.      �.       0�(0      -0       0�                                              �      �       U�      �       V�             �U�      �       V�      �       �U��      >       V>      G       �U�G      C       VC      �       ���      �       V�             �U�      /       V/             ��      *       �U�*      k       ��                                    �      �       T�             _             �T�      �       _�      �       �����      F       _F      G       �T�G             _             �T�      k       _                                   �      �       T�             _             �T�      �       _�      �       �����      F       _F      G       �T�G             _             �T�      k       _                                                       �      �       ^      �       ^0      D       ^D      F        F      G       �T�      ;       ^Q      �       V�      �       ]�      �       V      /       ^/      7       V7      <       ]<      c       Vc      �       ]�             V      *       ^*      8       V8      <       ]<      >       ^>      N       VN      k       ]                              �      �       S      �       S�      =       SG      �       S�      "       w �      �       S      /       S                           �      �       ]      �       ]�      B       ]G      �       ]�             ]      /       ]                                     �       v���      �       �U#���      C       v��C      �       ��#��      /       v��/             ��#��      *       �U#��*      k       ��#��                   3      7       P      /       
 �                              3      7       P7      �       \�      �       ���      Q       \Q      �       ��"      /       
 �/             ��*      k       ��                                   �      �       0��             S             T             s�      "       S"      Q       0�Q      �       w /      �       w �             w *      k       w                              �       ���      �       ���      �       ��      k       ��                                $       R$      �       w �      �       ���      �       w       /       R                         7       0�             0�      /       1�                 �      "      
 �1H     �                        ~      �       \/      K       w X      c       RN      k       \                     �      �       p } ��      �       P�      �       V                            �0      �0       U�0      1       S1      1       �U�1      ,1       S,1      .1       �U�.1      �1       S                          �0      �0       T�0      �0       V�0      1       �T�1      -1       V-1      �1       �T�                          �0      �0       T�0      �0       V�0      1       �T�1      -1       V-1      �1       �T�                            �0      �0       u���0      1       s��1      1       �U#��1      ,1       s��,1      .1       �U#��.1      �1       s��                           �0      �0       u���0      1       s��1      1       �U#��1      ,1       s��,1      .1       �U#��.1      �1       s��                           �0      �0       U�0      1       S1      1       �U�1      ,1       S,1      .1       �U�.1      �1       S                    �0      �0       q �.1      <1       q �                    �0      �0       P1      .1       P                                         U       t       St      ~       �U�~      �       S�      �       �U�                                         T       y       ]y      ~       �T�~      �       ]�      �       �T�                                         Q       {       ^{      ~       �Q�~      �       ^�      �       �Q�                                   R       �       �R�                    $      ,       P,      9       s                         U       V                    @      B       PB      o       _                      �      �       U�      �       S�      �       �U�                      �      �       T�      �       P�      �       �T�                            0      V       UV      �       V�      �       �U��      �       V�      3       �U�3      F       V                        0      [       T[      �       S�      �       �T��      F       S                         0      �       0��      �       P�      �       0��      �       P�      F       0�                        E      [       T[      �       S�      �       �T��      F       S                    S      �       _�      F       _                   �      �       \�              |h�                      �      �       0��             V             v�D      F       0�                    �      3       ^?      F       ^                        �      �       P�      �       s�      3       ��|D      F       P                             &       U&      �       S�             �U�                                 8       T8      @       U@      �       _�      �       �T��             _                         3      8       T8      @       U@      �       _�      �       �T��             _                    �      �       V�      �       s�                     �      �       0��      �       ��z�      �       P                      n      r       Pr      {        {      �       ��z                    w      {       P{      �       ��z                    =      @       P@             ��z                 �      �       ��z                   H      Y       0�d             ^                     Y      d       }h�d      s       ]s      �       }h�                      P      y       Uy      �       S�      �       ��{                          P      �       T�      �       U�      �       _�      �       �T��      �       _                    �      �       0�      9       ��{9      M       ��{                          U      �       T�      �       U�      �       _�      �       �T��      �       _                         U      :       0�:      M       PM      �       0��      �       P�      �       0�                   B      I       s�I      M       S                        �      �       P�      �        �      �       ��{�      �       ��{                        �      �       P�      �       �      �       ��{�      �       ��{                           �      �       0��             ��{      M       0��      �       P�      �       ��{�      �       ��{                   �      �       ��{�      �       ��{                   M      b       0�b      �       ]                   b      u       Vu      �       vh�                      p%      �%       U�%      �%       S�%      �&       �U�                          p%      �%       T�%      �%       U�%      �&       ]�&      �&       �T��&      �&       ]                     �%      �%       0��%      >&       VT&      n&       V                 n&      u&       3�                    �%      n&       \�&      �&       \                    �%      n&       ^�&      �&       ^                       �%      E&       _E&      T&       h�T&      n&       _�&      �&       h�                   &      &       T2&      I&       R                      �%      T&       Sj&      n&       S�&      �&       S                        `      �       U�      �       ]�      �       �U��      }       ]                 `      b       u�                    u      �       S�      }       S                    �      ~       ^�      }       ^                    �      �       V�      }       V                         �      �       1�       D       PD      H       p�r      �       0��      N       1�N      x       0�x      }       1�                   �      �       vx��      �       v`�                      P?      v?       Uv?      �?       �U��?      @       U                          P?      ?       T?      �?       \�?      �?       |��?      �?       �T��?      @       T                        P?      y?       Qy?      �?       ]�?      �?       �Q��?      @       Q                        c?      �?       V�?      �?       v�~��?      @       V@      @       u�                       �?      �?       0��?      �?       S�?      �?       s��?      �?       ^                   �?      �?       \�?      �?       ^                      �D      	E       U	E      @E       ]@E      CE       �U�                      �D      �D       T�D      <E       V<E      CE       �T4�T����4,( �                      �D      	E       Q	E      )E       ^)E      CE       �Q�                     �D      	E       0�	E      !E       S!E      %E       s�                    �E      �E       U�E      �E       �U�                    �E      �E       T�E      �E       �T�                              0C      xC       UxC      .D       ��~.D      @D       �U�@D      �D       ��~�D      �D       U�D      �D       ��~�D      �D       U                        0C      XC       TXC      .D       \@D      �D       \�D      �D       T                              0C      xC       QxC      .D       ].D      @D       �Q�@D      �D       ]�D      �D       Q�D      �D       ]�D      �D       Q                    D      .D       P�D      �D       P                    HC      =D       ^@D      �D       ^                         gC      xC       0�xC      �C       S�C      �C       s�@D      �D       S�D      �D       0�                          �C      �C       0��C      �C       P�C      �C       X�C      �C       P@D      CD       PnD      �D       P                      �C      �C       U@D      HD       UiD      �D       U                      �C      D       PFD      HD       P�D      �D       P                     xC      �C       V�C      .D       vh�@D      �D       V                    �C      �C       Y@D      �D       Y                        �C      �C       [@D      CD       [CD      HD       vHD      �D       [                          �C      �C       	���C      �C       X�C      �C       	���C      �C       X@D      CD       XHD      nD       	��nD      �D       X                    �C      �C       	��@D      CD       	��HD      nD       	��nD      �D       P                          �C      �C       y �C      �C       R�C      �C       y @D      CD       RnD      tD       RtD      xD       y q "8                      �>      �>       U�>      9?       �U�9?      L?       U                          �>      �>       T�>      	?       [	?      ?       {�?      9?       �T�9?      L?       T                        �>      �>       Q�>      7?       S7?      9?       �Q�9?      L?       Q                      �>      8?       V9?      K?       VK?      L?       u�                       �>      �>       0��>      �>       P�>      �>       p� ?      ?       Q                     �>      �>       [�>      ?       Q?      8?       v��Tv��T����,( �                     @      I@       UI@      B       �U�                             @      E@       TE@      [@       V[@      b@       �T�b@      gA       VgA      nA       �T�nA      B       V                    9@      R@       Zb@      �@       Z                           9@      R@       0�b@      �@       0��@      �@       P�@      iA       \iA      nA       �TnA      B       \                    �@      �@       0��A      �A       0��A      �A       ]                        @@      Z@       Sb@      ZA       SnA      �A       S�A      �A       s�~�                          �1      �1       U�1       2       �U� 2      (2       U(2      m2       �U�m2      w2       U                        �1      A2       TA2      H2       UH2      m2       �T�m2      w2       T                    �1      �1       1�m2      w2       1�                      `      �       U�      �       �U��      �       U                  g      �       R                   |      �       0��      �       Q                   �      �       p t "#��      �       p t "@�                   �      �      	 r p "#���      �      	 r p "#��                                  �      �       U�      �       V�      �       �U��      �	       V�	      5
       v�z�5
      �
       �U��
      �
       U�
      �
       V�
      .       �U�                            �      �       T�      �       \�      �       �T��      
       \�
      �
       T�
      .       \                              �      �       Q�      �       ]�      �       �Q��      c
       ]c
      w
       s�
      �
       Q�
      �
       ]�
      �
       s                         �      �       S�      |
       S�
      �
       S�
      �
       P�
      .       S                      �      �       _�      �
       _�
      .       _                 �      �       3�                 �	      �	       2�                  �
             1�                        p      �       U�      !       S!      +       �U�+      %       S                                      p             T      �       ]�      ?       �T�?      l       Tl             ]      +       �T�+      B       ]B      P       TP      �       �T��             ]      %       �T�                                  p      �       Q�             ^      ?       �Q�?      H       QH      l       ^l      +       �Q�+      B       ^B      P       QP      %       �Q�                             p      �       R�      w       _?      D       RD      �       _+      B       _B      P       R�      %       _                       p      �       U�      !       S!      +       �U�+      %       S                                  \      j       Pj      �       \�              P       ?       \l      �       \�             0�+      5       P5      B       \P      %       \                    �      "       V+      %       V                                           
 p 3 $0)�      &      
  3 $0)�&      .       R.      ?       s�?      ?       ��gl             ��g+      B      
  3 $0)�P      %       ��g                                     p  1�      w         1�l      �         1�+      B         1��      %         1�                   �      "       v��+      %       v��                     �      �       v�?      l       v�B      P       v�                             �      �       P�      �       v�#�      �       ��g?      l       v�#l      �       ��g+      B       ��gB      P       v�#                       8      =       ��g�^�=      ?       �^�l             �^�P      %       �^�                     �      d       0�d      @       1�@             0�+      B       1�B      %       0�                         �      �       0��      ?       1�?      l       0�l             1�+      P       0�P      %       1�                       �       ]                   ^      ?       s0�P      %       s0�                  \      w      	 q 0$0&�                   �      �       ��hP      �       ��h                         �      �       ��h#P      w       ��h#w      �       P�      �       pp��      �       P                   �      �       s�P      w       s�                   �      �       s�P      w       s�                �      �       s�                    �      �       T�      �      
 p t "#���                  �      �       t ?&��      �       P                �      �       s�                    �      �       R�      �      
 p r "#���                  �      �       r ?&��      �       P                  w      �       p �      �       pp                   �      �       Q�      �      
 q x "#���                  �      �       q ?&��      �       X                   �      �       Q�      �      
 q x "#���                  �      �       q ?&��      �       X                             ��g                             s�                                 P            
 p q "#���                               p ?&�             Q                1      <       ��g                1      <       s�                    :      <       P<      <      
 p q "#���                  :      <       p ?&�<      <       Q                                 s       Us      t       Tt      7       ]7      G       �U�G      t       U                               V       TV      �       V�      G       �T�G      t       T                               Z       QZ      �       \�      G       �Q�G      t       Q                           6       R6      t       �R�                                 e       Xe      �       S�      G       �X�G      \       S\      t       X                                s       Us      t       Tt      7       ]7      G       �U�G      t       U                                s       u��s      t       t��t      7       }��7      G       �U#��G      t       u��                        "       u�                         �             0�             1�      2       0�2      7       1�G      \       0�                      u      �       P�             P      )       P                               J       UJ      K       TK             V             �U�                             *       T*             \             �T�                      S      a       Pa             ]             P                   �      �       0��              S                              J       u��J      K       t��K             v��             �U#��                                ^                      �      �       U�      �       S�      �       �U�                    �      �       T�      �       �T�                   �      �       P�      �       �L                 �      �       s                        �             U      @       S@      J       �U�J      �       S                          �             T      E       ]E      J       �T�J      f       ]f      �       T                            �             Q      I       _I      J       �Q�J      f       _f      w       Qw      �       _                      �             R      f       ��kf      �       R                    �      A       VJ      �       V                   �      A       v��J      �       v��                             �             0�      #       Pm      u       P�      �       P      J       Pa      f       Pf      �       0�                    �      G       ^J      �       ^                        �      �       P�      ?       w ?      J       ��kJ      �       w                     �      C       \J      �       \                    �<      =       U=      �=       �U�                    �<      
=       T
=      �=       �T�                    �<      =       Q=      �=       �Q�                   �<      =       U=      �=       �U�                       �<      =       P=      =       u�=      g=       �U#�j=      �=       �U#�                       �<      =       P=      =       u�=      g=       �U#�j=      �=       �U#�                   �<      g=       Rj=      �=       R                      �<      =       Q=      g=       �Q�j=      �=       �Q�                      �<      
=       T
=      g=       �T�j=      �=       �T�                   =      g=       Xj=      �=       X                      =      ,=       PG=      g=       Pj=      x=       P                      =      =       x p "�=      /=       TY=      g=       T                      =      g=       Qj=      t=       Qt=      �=       �T����@$�Q����!�                      =      /=       UT=      g=       Uj=      �=       U                    �2      �2       U�2      �2       �U�                    �2      �2       T�2      �2       �T�                                      `3      �3       U�3      �3       �U��3      k4       Uk4      �4       �U��4      b6       Ub6      �6       \�6      �6       �U��6      &7       U&7      37       \37      a7       �U�a7      �<       U                    `3      �3       T�3      �<       �T�                                      `3      �3       Q�3      o4       Qo4      �4       �Q��4      k6       Qk6      w6       �Q�w6      |6       p �6      *7       Q*7      a7       �Q�a7      �7       Q�7      �7       P�7      �<       Q                                        `3      �3       R�3      �3       �R��3      o4       Ro4      �4       �H�4      k6       Rk6      |6       �H|6      �6       �R��6      *7       R*7      @7       �H@7      V7       RV7      a7       �Ha7      �<       R                                  `3      �3       X�3      �3       �X��3      o4       Xo4      �4       �X��4      k6       Xk6      �6       �X��6      *7       X*7      a7       �X�a7      �<       X                                                                                                                       `3      �3       0��3      �3       0��3      �3       2��3      �3       0��3      �3       2��3      �3       0��3      '4       2�'4      '4       0�'4      U4       1�U4      p4       0�p4      y4       p�y4      �4       V�4      �4       0��4      5       8�5      5       0�5      75       8�75      I5       0�I5      s5       2�s5      s5       0�s5      �5       1��5      �5       0��5      �5       4��5      �5       0��5      �5       1��5      �5       0��5      6       2�6      6       0�6      G6       2�G6      �6       0��6      �6       V�6      �6       P�6      �6       0��6      �6       4��6      +7       0�+7      77       p�77      a7       Va7      a7       0�a7      �7       4��7      �7       0��7      �7       V�7      �7       0��7      8       4�8      8       0�8      E8       4�E8      `8       0�`8      �8       1��8      �8       0��8      �8       8��8      �8       0��8      �8       1��8      �8       0��8      9       8�9      )9       0�)9      [9       8�[9      [9       0�[9      �9       1��9      �9       0��9      �9       1��9      �9       0��9      �9       2��9      �9       0��9      :       1�:      :       0�:      =:       4�=:      =:       0�=:      _:       8�_:      o:       0�o:      �:       2��:      �:       0��:      �:       1��:      �:       0��:      ;       2�;      ;       0�;      A;       2�A;      A;       0�A;      m;       1�m;      m;       0�m;      �;       4��;      �;       0��;      �;       2��;      �;       0��;      �;       1��;      <       0�<      )<       2�)<      C<       1�C<      R<       2�R<      b<       4�b<      �<       8�                              v3      �3       S�3      �3       �X0�X0*( ��3      �6       S�6      �6       �X0�X0*( ��6      :<       S:<      C<       x 0x 0*( �C<      �<       S                                     v3      �3       U�3      �3       �U��3      k4       Uk4      �4       �U��4      b6       Ub6      �6       \�6      �6       �U��6      &7       U&7      37       \37      a7       �U�a7      �<       U                                     v3      �3       u���3      �3       �U#���3      k4       u��k4      �4       �U#���4      b6       u��b6      �6       |���6      �6       �U#���6      &7       u��&7      37       |��37      a7       �U#��a7      �<       u��                               )9      V9       0�V9      [9       Pb<      i<       0�i<      n<       Pn<      u<       0�u<      z<       Pz<      �<       0��<      �<       P                               �8      �8       0��8      �8       P�<      �<       0��<      �<       P�<      �<       0��<      �<       P�<      �<       0��<      �<       P                   �3      �3       0�G6      w6       0�w6      |6       1�                  l6      |6       P                      �      �       U�      �       �U��               U                            �      �       T�      �       V�      �       �T��      �       V�      �       �T��               T                           �      �       0��      �       s��      �       S�      �       P�      �       s��               0�                 �      �       s 3$| "                    �<      �<       U�<      �<       �U�                    �<      �<       T�<      �<       �T�                      �<      �<       Q�<      �<       P�<      �<       �Q�                      �<      �<       R�<      �<       Q�<      �<       �R�                      �2      �2       U�2      C3       �U�C3      \3       U                          �2      �2       T�2      3       ^3      "3       �T�"3      C3       ^C3      \3       T                          �2      �2       Q�2      3       ]3      "3       �Q�"3      C3       ]C3      \3       Q                          �2      �2       R�2      !3       _!3      "3       �R�"3      C3       _C3      \3       R                      �2      3       \"3      U3       \U3      \3       u�                      �2      �2       0��2      3       S"3      C3       S                      �2      �2       V�2      3       V"3      C3       V                        pG      �G       U�G      �G       S�G      �G       �U��G      �K       S                        pG      �G       T�G      �G       _�G      �G       �T��G      �K       _                       =H      }H       ]�H      �H       ]�I      �J       ]pK      |K       ]                    �G      �G       \�G      �K       \                           �G      �G       0��G      �G       P�G      �G       V�G      �G       P�G      }I       V}I      �I       0��I      �K       V                       �G      �G       U�G      �G       S�G      �G       �U��G      �K       S                       �G      �G       u���G      �G       s���G      �G       �U#���G      �K       s��                       eH      }H       � �I      J       QJ      ]J       � pK      |K       �                  �I      �K       V                   �I      cK       _pK      �K       _�K      �K       _                   �I      cK       SpK      �K       S�K      �K       S                          �I      �I       P�I      ]J       8]J      cK       ��~pK      |K       8|K      �K       ��~�K      �K       ��~                	     �I      J       QJ      ]J       � pK      |K       �                 
         �I      JJ       RJJ      ]J       � �J      cK       ]pK      |K       R�K      �K       ]                           �I      �I       q� ��I      �I       P�I      �I       p� J      'J       P'J      *J       ~~�*J      �J       ^�J       K       ~|� K      cK       ^�K      �K       ^                         sJ      vJ       PvJ      �J       Q�J       K       ��~ K      9K       Q�K      �K       Q�K      �K       ��~                       �I      �I       q� ��8$q� ��!
����I      �I       p 8$q� ��!
����I      J       q� ��8$q� ��!
���J      *J       � #d��8$� #c��!
���                          �J      �J       P�J      �J       s��J      cK       ��~�K      �K       s��K      �K       ��~                       �J      �J       0��J      �J       T�J      �J       p �J      �J       T�K      �K       T                 �J      �J       0�                         )        U                         )        T                         )        R                           %        Q%       )        t �����@$t�����!�                              $       U$      [       V[      _       U_      `       �U�                                      T       Z       SZ      _       T_      `       �T�                    �=      G>       Ql>      �>       Q                    �=      G>       Tl>      �>       T                    �=      G>       Ul>      �>       U                           B      EB       TEB      HB       �T�HB      yB       TyB      (C       Z(C      .C       T                    B      yB       U(C      .C       U                         HB      yB       0��B      �B       V�B      
C       v�
C      C       y�C      C       v�                          �B      �B       0��B      �B       u��B      �B       R�B      �B       U�B      �B       u�                        B      yB       0��B      �B       �G�B      �B       1��B      C       �G(C      .C       0�                          �B      �B       @<$��B      �B       T�B      �B       T�B      �B       P�B      �B       T                    �B      �B       u 3$q "�B      �B       P                 �B      �B       P                 �B      �B       T                    �B      �B       P�B      �B       p����B      �B       P                 �B      �B       0�                      PE      ^E       U^E      E       SE      �E       �U�                      PE      bE       TbE      �E       V�E      �E       �T�                    PE      kE       QkE      �E       �Q�                  cE      �E       P                    gE      kE       QkE      ~E       �Q�                  gE      ~E       V                  gE      ~E       S                 �E      �E       U                    �E      �E       S�E      �E       S                    �E      �E       P�E      �E       P                        �F      �F       U�F      �F       S�F      �F       �U��F      �F       U                       �F      �F       U�F      �F       S�F      �F       �U��F      �F       U                      �F      �F       U�F      �F       S�F      �F       �U�                  �F      �F       P                        �F      �F       U�F      EG       ^EG      WG       �U�WG      eG       ^                        �F      �F       T�F      EG       ��EG      WG       �T�WG      eG       ��                    �F      �F       Q�F      eG       �Q�                   �F      �F       Q�F      eG       �Q�                        �F      �F       0��F      G       s�G      EG       SWG      eG       s�                     �F      G       VG      EG       VWG      eG       V                          �K      �K       U�K      �K       S�K      �K       �U��K      bL       SbL      fL       �U�                          �K      �K       T�K      �K       \�K      �K       �T��K      eL       \eL      fL       �T�                          �K      �K       Q�K      �K       V�K      �K       �Q��K      cL       VcL      fL       �Q�                         �K      	L       P
L       L       P!L      /L       P0L      BL       P]L      fL       P                 4L      ]L       V                 4L      ]L       \                 4L      ]L       S                      4L      TL       0�TL      XL       PXL      ]L       �L]L      ]L       P                 �      (       U                         1      I1       UI1      �3       V�3      �3       �U��3      �3       U                        1      I1       UI1      �3       V�3      �3       �U��3      �3       U                  B1      �3       ^                 B1      I1       P                  Q1      �3       S                 Z1      ~3       S                  e1      ~3       \                    �1      �1       ]�1      �1       }�                  �1      �1       T                  �1      �1       \                 �1      2       s��                 
2      2       P                  
2      `2       s�
�                 
2      `2       ]                 
2      �3       s�
�                 
2      12       ]                     e2      l2       s��l2      s2       Ts2      t2       s��                 e2      t2       \                 t2      �2       s                 t2      �2       s�&�                 �3      �3       V                  �3      �3       P                                                                            pI      �I       U�I      �J       S�J      K       �U�K      �O       S�O      P       \P      [R       S[R      �T       �U��T      =U       S=U      �X       �U��X      8Y       S8Y      MY       �U�MY      �Z       S�Z       \       �U� \      \       S\      �^       �U��^      Ij       SIj      wj       ]wj      �j       S�j      �j       \�j      �k       S�k      �k       ]�k      �m       S�m      �m       ]�m      =o       S=o      ho       \ho      vo       Svo      �o       \�o      �o       S�o      �o       \�o      �o       S                                                                  pI      �I       T�I      �J       ]�J      K       �T�K      �N       ]�N      ZQ       �T�ZQ      �Q       ]�Q      �T       �T��T      =U       ]=U      �X       �T��X      8Y       ]8Y      MY       �T�MY      �Z       ]�Z       \       �T� \      \       ]\      �^       �T��^      h_       ]h_      �_       �T��_      T`       ]T`      �j       �T��j      �k       ]�k      l       ��}l      �m       �T��m      �m       ]�m      �m       ��}�m      �o       �T�                                                                  pI      �I       Q�I      �J       ^�J      K       �Q�K      �N       ^�N      ZQ       �Q�ZQ      �Q       ^�Q      �T       �Q��T      =U       ^=U      �X       �Q��X      8Y       ^8Y      MY       �Q�MY      �Z       ^�Z       \       �Q� \      \       ^\      �^       �Q��^      h_       ^h_      �_       �Q��_      T`       ^T`      �j       �Q��j      �k       ^�k      �l       ��}�l      �m       �Q��m      �m       ^�m      �m       ��}�m      �o       �Q�                              pI      �I       R�I      �J       w �J      K       �R�K      DK       w DK      ZQ       �R�ZQ      �Q       w �Q      �o       �R�                                  pI      �I       X�I      �J       ��}�J      K       �X�K      `K       ��}`K      ZQ       �X�ZQ      �Q       ��}�Q      �T       �X��T      U       ��}U      �o       �X�                                                                 pI      �I       T�I      �J       ]�J      K       �T�K      �N       ]�N      ZQ       �T�ZQ      �Q       ]�Q      �T       �T��T      =U       ]=U      �X       �T��X      8Y       ]8Y      MY       �T�MY      �Z       ]�Z       \       �T� \      \       ]\      �^       �T��^      h_       ]h_      �_       �T��_      T`       ]T`      �j       �T��j      �k       ]�k      l       ��}l      �m       �T��m      �m       ]�m      �m       ��}�m      �o       �T�                   �J      �J       ;��X      �X       P                          �I      �I       P�I      �J       \K      @K       \ZQ      �Q       \�T      U       \                         �I      �I       P�I      �J       ��}K      �K       ��}ZQ      �Q       ��}�T      U       ��}                          �I      �I       P�I      �J       ��}K      �K       ��}ZQ      �Q       ��}�T      U       ��}                  �I      J       P                          J      $J       P$J      �J       ��}K      �K       ��}ZQ      �Q       ��}�T      U       ��}                	           pI      �J       1��J      �J       w K      DK       1�DK      �K       w ZQ      ZQ       1�ZQ      �Q       0��T      U       w                 
                                                                 pI      �J       0��J      �J       1�K      DK       0�DK      �N       \�N       Q       ��~ZQ      �Q       0��Q      �Q       \�T      U       0�U      =U       \�X      8Y       \MY      �Z       \ \      \       \�^      h_       \h_      �_       ��~�_      T`       \T`      qa       ��~-c      7c       ��~�f      Ig       ��~fg      �h       ��~[i      mi       ��~�i      �j       ��~�j      �j       ��~�j      �j       ��~�j      �k       \�k      �k       ��~�k      �k       ^�k      l       ��~l      �l       \�l      �m       ��}�m      �m       \�m      �m       ^�m      �m       ��~�m      En       ��}En      �o       ��~                         pI      yJ       0�yJ      �J       1�K      DK       0�DK      �K       ��~ZQ      �Q       1��T      U       1�                          �I      �J       VK      �L       VZQ      �Q       V�T      U       VMY      tY       V                 �I      �I       U                          �I      �I       P�I      �J       ��}K      �K       ��}ZQ      �Q       ��}�T      U       ��}                  J      J       }�                           J      $J       P$J      �J       ��}K      �K       ��}ZQ      �Q       ��}�T      U       ��}                           DK      pK       0�pK      �K       P�K      �K       R�K      �K       [�K      YL       ��}MY      `Y       ��}                   (R      cR       {��cR      �R       ��}#��                    `K      dK       PdK      �K       ��}                           �V      �V       
��V      W       PW      $W       0�$W      dW       s ��dW      �W       S�W      �W       S�W      �W       }                      S      S       PS      S       {�S      -S       s                  3R      cR       }�                   3R      cR       }�cR      �R       S                   3R      ER       ~ @%�ER      �R       ^                          �R      �T       V=U      �X       V8Y      MY       V�Z       \       V\      �^       V                           �R      �R       {���R      �T       v0�=U      �X       v0�8Y      MY       v0��Z       \       v0�\      �^       v0�                           �R      �R       {���R      �T       v(�=U      �X       v(�8Y      MY       v(��Z       \       v(�\      �^       v(�                    �R      S       S=[       \       S                      -S      �S       \�S      �T       \=U      HU       \                     -S      �S       }���S      �T       }��=U      HU       }��                     �S      �S       |� �1T      �T       |� �=U      HU       |� �                     �S      �S       |� �1T      �T       |� �=U      HU       |� �                     �S      �S       |� �1T      �T       |� �=U      HU       |� �                      �S      �S       ^QT      �T       ^=U      HU       ^                  bS      �S       ^                       YU      �V       0�F\      �]       0��]      ^       0�^      !^       P!^      �^       \                  _\      �\       P                 �\      �\       P                  �\      �\       U�\      �\       ��}                 �\      �\       P                  uV      �V       P                           uV      �V       P�\      �\       P�\      �\       p��\      �\       P�\      �\       p��\      �\       P�]      �]       P�]      ^       P                        yV      �V       T�\      �\       T�]      �]       T�]      ^       T                 ^      ^       T                  ^      ^       U^      ^       ��}                 ^      ^       P                   ^      !^       P!^      �^       \                 ^      �^       S                  (^      �^       ^                  8^      �^       P                                  >^      n^       1�n^      x^       2q �^      �^       2q ��^      �^       r��^      �^       R�^      �^       p��^      �^       P�^      �^       P�^      �^       R                  �]      �]       P                 �]      �]       P                �]      �]       ��}                 �]      �]       P                  )W      BW       P                �V      �V      
 �BH     �                  �V      �V       U�V      �V       ��}                 �V      �V       P                         �\      �\       P�\      �\       U�\      ]       X]      P]       RP]      z]       X                         �\      ]       0�]      %]       q x #�)]      6]       q x �6]      E]       q x #�E]      P]       7�P]      X]       r x #�                  �\      z]       U                         �\      ]       1�]      %]       Z)]      6]       Z6]      @]       0�@]      c]       Zc]      o]       1�                        �W      �W       Q�W      X       }� X      X       RX      4X       }�                        �W      �W       0��W      4X       QcX      �X       S[      [       0��]      �]       S                  �W      �W       {��[      [       {��                   �X      �X      
 �gH     �A\      F\      
 �gH     ��]      �]      
 �gH     �                                                                         �K      �N       \�N       Q       ��~�Q      �Q       \U      =U       \�X      Y       \MY      �Z       \�^      B_       \]_      h_       \h_      �_       ��~�_      T`       \T`      qa       ��~-c      7c       ��~�f      Ig       ��~fg      �h       ��~[i      mi       ��~�i      �j       ��~�j      �j       ��~�j      �j       ��~�j      �k       \�k      �k       ��~�k      �k       ^�k      l       ��~l      �l       \�l      �m       ��}�m      �m       \�m      �m       ^�m      �m       ��~�m      En       ��}En      �o       ��~                 �K      �K       w                                                  �K      �N       ]�N      7Q       �T��Q      �Q       ]U      =U       ]�X      Y       ]MY      �Z       ]�^      B_       ]]_      h_       ]h_      �_       �T��_      T`       ]T`      �j       �T��j      �k       ]�k      l       ��}l      �m       �T��m      �m       ]�m      �m       ��}�m      �o       �T�                         �K      �K       P�K      �K       R�K      �K       [�K      YL       ��}MY      `Y       ��}                                                 �K      �N       ^�N      7Q       �Q��Q      �Q       ^U      =U       ^�X      Y       ^MY      �Z       ^�^      B_       ^]_      h_       ^h_      �_       �Q��_      T`       ^T`      �j       �Q��j      �k       ^�k      �l       ��}�l      �m       �Q��m      �m       ^�m      �m       ��}�m      �o       �Q�                                                             �K      �O       S�O      P       \P      7Q       S�Q      �Q       SU      =U       S�X      Y       SMY      �Z       S�^      B_       S]_      Ij       SIj      wj       ]wj      �j       S�j      �j       \�j      �k       S�k      �k       ]�k      �m       S�m      �m       ]�m      =o       S=o      ho       \ho      vo       Svo      �o       \�o      �o       S�o      �o       \�o      �o       S                   �K      �L       VMY      tY       V                 �K      �K       ��}                                              �K      L       PL       Q       ��}�Q      �Q       ��}U      =U       ��}�X      Y       ��}MY      �Z       ��}�^      B_       ��}]_      qa       ��}-c      7c       ��}�f      Ig       ��}fg      �h       ��}[i      mi       ��}�i      �j       ��}�j      �j       ��}�j      �o       ��}                   �K      YL       ��}#��MY      `Y       ��}#��                                           �M      �M       R�M       Q       ��~�X      Y       ��~�^      �^       0� _      9_       R9_      B_       ��}]_      qa       ��~-c      7c       ��~�f      Ig       ��~fg      �h       ��~[i      mi       ��~�i      �j       ��~�j      �j       ��~�j      �o       ��~                          ZN      UO       0�UO      sO       P�O      �O       v�3$s "�_      T`       0��j      �m       0��m      �o       0�                            sO      {O       R{O      O       r��O      �O       R�O      �O       V�O      �O       Q�O      1P       V                    aN      �N       P�_      �_       P                         aN      �N       ��}�_      �_       ��}�_      T`       ��}�j      �m       ��}�m      �o       ��}                                             aN      �N       S�_      �_       S�_      T`       S�j      �k       S�k      �k       ]�k      �m       S�m      �m       ]�m      �m       S�m      =o       S=o      ho       \ho      vo       Svo      �o       \�o      �o       S�o      �o       \�o      �o       S                      aN      �N       {�'��_      �_       {�'��_      �_       ��}#�'�                             ~N      �N       R�N      �N       ��}�_      �_       ��}�_      �_       R�_      T`       ��}�j      �m       ��}�m      �o       ��}                                      ~N      �N       0��N      �N       ��}�N      �N       T�N      �N       ��}�N      �N       0��_      �_       0��_      T`       0��j      tk       0�tk      �k       P�k      �m       ��}�m      �m       0��m      �m       ��}�m      �o       ��}                                    �k      �l       V�l      �m       ��~�m      �m       V�m      n       ��~n      In       PIn      tn       ��~tn      ho       ��}ho      vo       Pvo      �o       ��}�o      �o       ��}                           
m      ^m       \�m      �m       \=o      ho       Svo      |o       S|o      �o       T�o      �o       S                      "`      T`       ��}�j      �l       ��}�m      �m       ��}                  '`      >`       p 
���                      k      *k       P*k      �l       ��~�m      �m       ��~                    �l      �m       ]�m      
n       ]                 m      �m       V                  m      -m       ��~                  >m      Nm       ��~                  cm      �m       P                  �n      �n      
 v 4$��}"�                  1P      5P       T                      1P      5P       U5P      �P       S�m      �m       S                    1P      �P       V�m      �m       V                    1P      �P       ��}#�&��m      �m       ��}#�&�                    ZP      �P       P�m      �m       P                    �P      �P       p 
����P      �P       P                  mY      �Y       P                                �`      �`       p ����
��.w �0.��`      qa       ��}�
��.w �0.�-c      7c       ��}�
��.w �0.��f      Ig       ��}�
��.w �0.�fg      �h       ��}�
��.w �0.�[i      mi       ��}�
��.w �0.��i      �j       ��}�
��.w �0.��j      �j       ��}�
��.w �0.�                              �`      qa       ��}�
��.w �0.�-c      7c       ��}�
��.w �0.��f      Ig       ��}�
��.w �0.�fg      �h       ��}�
��.w �0.�[i      mi       ��}�
��.w �0.��i      �j       ��}�
��.w �0.��j      �j       ��}�
��.w �0.�                        �`      .a       P�f      g       Pfg      �g       P�i      �i       P                              �`      qa       ��}-c      7c       ��}�f      Ig       ��}fg      �h       ��}[i      mi       ��}�i      �j       ��}�j      �j       ��}                          �`      �a       S-c      Yc       S�f      Gi       S[i      Ij       SIj      wj       ]wj      �j       S                      �`      �a       \-c      Yc       \�f      Gi       \[i      �j       \                              �`      qa       ��}-c      7c       ��}�f      Ig       ��}fg      �h       ��}[i      mi       ��}�i      �j       ��}�j      �j       ��}                                          �`       a       R a      .a       U.a      qa       ��}-c      7c       ��}�f      �f       R�f      Ig       ��}fg      kg       Rkg      �h       ��}[i      mi       ��}�i      �i       ��}�i      �i       R�i      �j       ��}�j      �j       ��}                          Lh      ah       Pah      �h       ^�h      �h       ~ r "��h      �h       P�h      �h       ^                          -h      �h       ]�h      �h       }��h      �h       ]�i      j       ]cj      gj       v�                        mh      �h       P�h      �h       T�h      �h       P�h      �h       P                   �h      �h       0��h      �h       R                          b      cb       Qcb      �b       {��c      �c       Q�c      �c       {��c      �c       Q                         b      vb       ��}Yc      dc       ��}�c      �c       ��}�c      �d       ��};f      �f       ��}                        b      -c       SYc      kc       Swc      �c       S�c      �f       S                        b      -c       \Yc      kc       \wc      �c       \�c      �f       \                          b      �b       {���b      -c       ��}#���c      �c       {���c      �d       ��}#��;f      If       ��}#��                                  wc      c       ��}Hd      �d       p ���d      Ne       v ��[e      �e       v ���e      �e       P�e      ;f       ��};f      Tf       p ��Tf      �f       v ���f      �f       ��}                                    �b      �b       p��b      �b       Pc      -c       p�wc      c       R�d      �d       0��d      Ee       ��}[e      {e       ��}�e      ;f       ��}mf      vf       1�vf      �f       Q�f      �f       ��}                    �e      ;f       P�f      �f       P                           �d      �d       Q�d      e       ��}e      Ne       Q�e      	f       v ��vf      �f       t p "����f      �f       t r "1���                          �b      �b       R�b      �b       Q�b      �b       p 1${ "#��
���c      c       Rc       c       p 1${ "#��
���                   �b      �b       0��b      �b       q 
���c      c       0�                    �b      �b       R�b      �b       Q�b      �b       p 1${ "#��
���                  �b      �b       0��b      �b       q 
���                  �d      e       P                       wd      �d       1��d      @e       ��}@e      Ne       U[e      {e       ��}                  e      Ne       R                     f      f       0�f      ;f       R�f      �f       R                        mf      vf       Tvf      vf       t p "�vf      �f       t p "#��f      �f       t r "��f      �f       t p "�                      0      `       U`      {       S{      �       �U�                      :      T       PT      `       u`      d       s                   :      T       p�T      d       Q                  H      �       V                  e      o       P                  p      {       P                          �      �       U�      �       V�      �       �U��      �       V�      �       �U�                          �      �       T�      ,       S,      �       �T��      �       S�      �       �T�                         �      �       U�      �       V�      �       �U��      �       V�      �       �U�                    �      �       P�      �       ]                 �      �       U                 �      �       u�                 �             v                   	      �       ^                        �       _                        �       \                  %      2       P                   2      J       P�      �       ~ s "#�                      2      J       RJ      j       ���      �       R                       [      b       Pb      j       w j      ~       Y�      �       Y                    j      ~       Q�      �       Q                                    U      �       V�      �       �U�                                  T      �       �T�                                   U      �       V�      �       �U�                    &      6       P6      �       ]                 2      ^       v                   J      �       ^                  Q      �       _                  X      �       \                  f      s       P                   s      �       P�      �       ~ s "#�                      s      �       R�      �       ���      �       R                       �      �       P�      �       w �      �       Y�      �       Y                    �      �       Q�      �       Q                        �      �       U�      O       VO      X       �U�X             V                       �      �       U�      O       VO      X       �U�X             V                                       P      C       \X      �       \�      �       P             \                        0       P                      ,      C       ]X      �       ]             ]                           ,      >       0�>      C       PX      p       Pp      �       _�      �       ��}             ��}                 ,      0       U                  �      �       P                 �      �       } s "#�                    �      �       U�             Q                    �      �       u���             q��                                              �      �       0��      �       P�      �       p��      �       0��      �       P�      �       p�              0�             P      !       p�0      6       0�6      M       PM      Q       p��      �       0��      �       P�      �       p��      �       0��      �       P�      �       p�                            �      �       U�      �       U       ,       U0      �       U�      �       U�             U                                    U      v       �U�v      �       U                               u #�                                   U      v       �U�v      �       U                               u                                u #�                              m       Vm      u       Tv      �       V�      �       p                     /      :       P:      o       \                    A      H       PH      M       s�                        pE      F       UF      �G       ^�G      �G       �U��G      lI       ^                                        pE      �E       T�E      =G       V=G      DG       �T�DG      lG       VlG      �G       �T��G      RH       VRH      �H       �T��H      I       VI      +I       �T�+I      :I       V:I      bI       �T�bI      lI       V                          pE      �E       Q�E      VF       ��~VF      DG       �Q�DG      lG       ��~lG      lI       �Q�                        pE      �E       R�E      �G       \�G      �G       �R��G      lI       \                          pE      �E       X�E      VF       ��~VF      DG       �X�DG      lG       ��~lG      lI       �X�                      pE      	F       Y	F      &F       ��&F      lI       �Y�                    pE      VF       � DG      lG       �                     pE      VF       �DG      lG       �                                                     BF      BF       RBF      	G       0�	G      G       PG      DG       _aG      �G       _�G      �G       P�G      �G       0��G      �G       P�G      �G       _�G      �G       P�G      �G       0��G      �G       P�G      H       _H      +H       P+H      �H       _�H      �H       P�H      �H       _�H      �H       P�H      �H       _�H      bI       _bI      lI       P                       �E      F       UF      �G       ^�G      �G       �U��G      lI       ^                       �E      F       u��F      �G       ~���G      �G       �U#���G      lI       ~��                        �E      �E       P�E      &F       �#�&F      VF       ��~DG      lG       ��~                   �E      �G       s  $0)��G      lI       s  $0)�                        �E      BF       _BF      DG       	�0s  $0)( 
�#`�DG      XG       _XG      �G       	�0s  $0)( 
�#`��G      lI       	�0s  $0)( 
�#`�                  :I      bI       V                  �E      BF       0�DG      aG       0�                    �E      BF       _DG      XG       _XG      aG       	�0s  $0)( 
�#`�                    �E      F       QF      &F       p                     �E      F       UF      BF       ^DG      aG       ^                      �E      	F       Y	F      &F       ��&F      BF       �Y�DG      aG       �Y�                  �E      BF       ��~�DG      aG       ��~�                  �E      BF       ]DG      aG       ]                   G      'G       V�H      I       V                   G      'G       ]�H      I       ]                 �H      I       v                  lG      �G       ��~�                 lG      xG       ��~                          9      n9       Un9      �9       t��9      �:       ]�:      �:       �U��:      �;       ]                            9      :       T:      E:       z�E:      �:       \�:      �:       �T��:      �:       T�:      �;       \                              9      �9       Q�9      :       t�:      E:       z�E:      �:       �Q��:      �:       Q�:      �:       t��:      �;       �Q�                              9      q9       Rq9      �9       Y�9      :       t�:      E:       z�E:      �:       �R��:      �:       t��:      �;       �R�                                     9      v:       0�v:      �:       P�:      �:       V�:      �:       P�:      �:       V�:      �:       P�:      !;       0�!;      9;       P9;      ?;       V?;      C;       PC;      �;       V                           9      :       T:      E:       z�E:      �:       \�:      �:       �T��:      �:       T�:      �;       \                           9      :       t��:      E:       z�#��E:      �:       |���:      �:       �T#���:      �:       t���:      �;       |��                      *9      K9       SS9      �:       S�:      �;       S                    �9      �9       a��:      �:       R                    :      :       t�:      E:       zn                    :      :       t�:      E:       zl                  :      `:       V�:      ;       V                    :      :       Q:      E:       ��                      :      :       t��:      E:       z�#��E:      `:       |���:      ;       |��                    :      2:       U2:      E:       ��                  :      `:       ����:      ;       ���                 :      `:       ^�:      ;       ^                �:      �:       \                 �:      �:       ���                 �:      �:       ��                    p      y       Uy      z       �U�                    p      y       Ty      z       �T�                    p      y       Qy      z       �Q�                    p      y       Ry      z       �R�                    p      y       Xy      z       �X�                 p      y       u�                    p      �       U�      �       �U�                    p      �       T�      �       �T�                    p      �       Q�      �       �Q�                    p      �       R�      �       �R�                            �      �       U�      �       �U��      =       U=      �       ]�      �       X�      �       �U�                        �      �       T�      �       �T��      B       TB      �       ��                        �      �       Q�      �       �Q��             Q      �       ��                        �      �       R�      �       �R��      J       RJ      �       ��                 �      �       3�                    �      �       P�      �       ��                        M      Q       RQ      �       S�              ��~�#�4      0       ��~�#�                   �      �       ~�'��      �       ~�'�                           U       PU      �       ��~                       h      �       0��      �       V�      �       v��      �       V�      �       v�4      0       V                 J      U       0�                   �      �       P4      U       P                  �      �       p ����3$z�'"�4      U       p ����3$z�'"�                        c      s       Us      �        s "��              s "�"      0        s "�                        "       P                 �      �       t                    �      �       Q�      �      
 p q "#���                  �      �       q ?&��      �       P                      p      �       U�             S      %       �U�                      p      �       T�      $       ]$      %       �T�                            �      �       0��      �       V�      �       v��      �       V�      �       0��      �       \�      �       |��      
       \                          �      �       U�      +       V+      4       �U�4      O       UO      d       V                          �      �       T�      +       \+      4       �T�4      L       TL      d       \                            �      �       Q�      �       Z�      4       �Q�4      G       QG      U       ZU      d       �Q�                    �      �       0�4      d       0�                        "       Q                     �      �       0��      "       S4      d       0�                         �      F       0�F      G       PG      T       0�T      U       PU      [       0�[      i       P                       �      �       Q�      �       q��      �       q��             R             r�      <       RU      i       R                    �      <       ZU      i       Z                      �             P             r       <       PU      i       P                        �             X      /       Y/      2       QU      [       X[      i       Y                                 +       Y+      2       Q2      <       YU      [       Y[      ^       Q                                �       �        U�       �        S�       �        �U��       !       S!      !       �U�!      !       S!       !       �U� !      4!       S                    �       �        T�       4!       �T�                                 �       �        u8��       �        U�       �        s8��       �        �U#8��       !       s8�!      !       �U#8�!      !       s8�!       !       �U#8� !      4!       s8�                 �       �        V                               �       �        0��       �        P�       �        V�       �        P�       !       0�!      !       V!       !       P !      4!       V                       �       �        s8��       �        �U#8�!      !       s8�!       !       �U#8�                       �       �        s8��       �        �U#8�!      !       s8�!       !       �U#8�                       �       �        �P�!      !       �P�!      !       T!       !       �P�                 !      !       s8                            �      �       U�      H       SH      W       �U�W      �       S�      �       �U��      t        S                          �      �       T�      �       V�      �       v  �W      c       V�      (        V                              �      �       Q�      H       ^H      W       �Q�W      �       ^�      �       �Q��      �       Q�      t        ^                          �             R      �       �R��      �       R�      �       ���      t        �R�                  [       `        P                      �      H       _W      �       _�      t        _                        �      H       \W      �       \�      �       P�      t        \                                 �      �       0��      �       P�             P      )       PW      t       0��      �       0��              P       (        P`       t        P                 �      �       s��v �����                        �      �       U�      �       S�      �       �U��      �       S                            �      �       T�      �       ^�      �       �T��      ^       ^^      �       T�      �       ^                                �      �       Q�      ^       �Q�^      �       Q�      �       Z�      �       ���      �       �Q��             ��      �       �Q�                            �      �       R�      �       w �      �       ���      ^       w ^      �       R�      �       w                        �      �       \�      x       \^      �       \�      �       \                                 �      �       0��             0�             P      ^       ��^      �       0��      �       ���             0�      	       ��	      �       0�                               �      �       0��      D       0�D      H       PH      e       _^      �       0��             0�      	       _	      �       0�                   �      �       } ����s("��             } ����s("�                            ]      z       1�z             ]      &       }�&      ?       ]�      �       ]�      �       1�      	       1�                         Z      Z       s01�Z      z       0�z      �       T�      ?       T�      �       T�      �       s01��      �       0�      	       0�                          N      z       0�z      �       R�      �       ���      ?       R�      �       R�      �       0�      	       0�                      Z      z       Y�      �       Y      	       Y                         z      �       V       	       V	      .       T�      �       V�      �       T                     e      �       S�      �       S�      �       S	      �       S                     m      �       _�      �       _�      �       _	      �       _                     m      �       \�      �       \�      �       \	      �       \                        �      �       P�      �       ���      �       ���      �       ��	      �       ��                            �      �      	 p �r ��      �       ����v ��      �       }����������      !       ����v �!      �       }����������      �       }���������	      �       }���������                                   C      �       P	             P      #       p~�#      D       PD      L       p r "�L      P       p r "#�P      Z       p r "�Z      n       Pn      ~       p}�~      �       P                          G      �       T�      �       � v "�	      D       TD      Z       p v "�Z      �       T                                        C      t       Qt      |       qx�|      �       Q	             Q      /       qx�/      D       QD      L       r 3$q "�L      P      
 r 3$q "#�P      Z      
 r3$q "#�Z      r       Qr      �       qx��      �       Q                               C       UC      l       Sl      n       �U�n      q       U                 -      G       P                  :      m       V                                @!      �!       U�!      �!       S�!      �!       �U��!      �!       S�!      �!       �U��!      �"       S�"      �"       �U��"      �"       S                                  @!      �!       T�!      �!       V�!      �!       �T��!      �!       V�!      �!       �T��!      "       U"      �"       V�"      �"       �T��"      �"       V                    @!      �!       Q�!      �"       �Q�                    @!      �!       R�!      �"       �R�                        b!      �!       ]�!      �!       ]�!      �"       ]�"      �"       ]                           �!      �!       P�!      �!       \�!      �!       \"      "       p 
���"      �"       \�"      �"       \                    ("      C"       PC"      c"       s                         R"      ["       T["      c"       s�#����p �"      �"       P�"      �"       T�"      �"       T                    p      �       U�      �       �U�                            �5      �5       U�5      �6       \�6      �6       �U��6      �8       \�8      �8       �U��8      9       \                    �5      �5       T�5      9       �T�                      �5      �5       Q�5      �5       P�5      9       ��                                                       �5      �5       T�5      6       ^$6      �6       ^�6      ,7       ^,7      ?7       ~�?7      �7       ^�7      �7       Q�7      �7       ^�7      �7       ~��7      �7       q #��7      V8       ^V8      Z8       ~�Z8      _8       q #�_8      _8       ^_8      h8       ~�h8      v8       Pv8      �8       ~��8      �8       p��8      �8       ~��8      �8       p~��8      �8       p��8      �8       ^�8      �8       ~��8      9      	 |(8#�                      �5      �6       0��6      f7       0�f7      o7       Po7      9       0�                 �5      �5       u                                         �5      6       P(6      c6       P�7      �7       P�7      �7       PV8      h8       Pv8      �8       p 4%���8      �8       p ?���8      �8      
 ~�?���8      �8       |(8#�?���8      �8       q 4%���8      �8       q ?���8      �8      
 p�?���8      �8      
 ~�?���8      �8       |(8#�?��                           Z6      c6       Pc6      h6       |4�p !�h6      �6       P�6      �6       Po7      }7       P�7      �7       P�7      �7       P                               W6      �6      
 |(| 8��6      7      
 |(| 8�?7      O7      
 |(| 8�_7      e7      
 |(| 8�o7      �7      
 |(| 8��7      �7      
 |(| 8��7      �7      
 |(| 8��7      �7       T                             c6      ~6      
  ZH     �~6      �6       S�6      7       S?7      Y7       S_7      o7       So7      }7      
  ZH     ��7      V8       S                           7      "7       PP7      _7       P�7      �7       P�7      �7       0��7      V8       _�8      �8       P                        �6      o7       Vu7      �7       V�7      V8       V�8      �8       V                   �7      �7       s�����p "��7      �7       q ����p "�                   �7      �7       | �7      V8       ]                 �6      7       |                  �6      7       3�                 �6      7       \                 ?7      O7       |                  ?7      P7       \                        �;      �;       U�;      �;       up��;      <       �U�<      <       U                      �;      <       S<      <       S<      <       u8                     �;      �;       u �;      �;       u #��;      �;       p�<      <       u                    �;      <       0�<      <       3�                              �=      �=       U�=      �?       _�?      �?       �U��?      @       _@      @       �U�@      �@       _�@      �@       U                      �=      �=       P�@      �@       P�@      �@       u8                     �=      �?       ^�?      @       ^@      �@       ^                        �=      P>       SP>      �?       ~���?      @       ~��@      �@       ~��                  >      ->       P                   �=      >       P�?      �?       ���?      @       P                   &>      �>       V@      �@       V                    &>      �?       _�?      �?       _@      �@       _                    &>      �?       ^�?      �?       ^@      �@       ^                                  �>      �>       P�>      �>       Q�>      �>       ���>      ?       Q?      ?       Y?      ?       ��?      0?       Y�?      �?       Y@      @       ��                 �>      �>       S                       �>      �>       0��>      �?       0��?      �?       1�@      @       0�                   �>      �>       1�@      @       1�                        q>      �>       [�>      �>       v 2$v "�@      R@       [R@      �@       ��                	     &>      �?       ~���?      @       ~��@      �@       ~��                    D>      �>       U@      R@       U                    L>      �>       ]@      �@       ]                    \>      �>       S@      �@       S                        �>      �>       V�>      �>       v|�?      �?       V@      @       V                        �>      �>       X�>      ?       ��?      �?       X@      @       X                    '@      R@       ZR@      �@       ��                    I@      R@       PR@      �@       ��                  �@      �@       P                   �@      �@        �@      �@       Q                        �;      �;       U�;      �;       up��;      �;       �U��;      �;       U                      �;      �;       S�;      �;       S�;      �;       u8                     �;      �;       u �;      �;       u #��;      �;       p��;      �;       u                  �;      �;       q��                 �;      �;       0�                       <      F<       UF<      }<       sp�}<      �<       �U�                  <      "<       u8                  -<      C<       VC<      Z<       v�Z<      }<       v�                 -<      {<       ��{<      }<       0�                      �<      �<       U�<      �<       S�<      =       �U�                 �<      �<       u8                �<      �<       ��                    �<      �<       P�<      =       R                      =      ?=       U?=      m=       sp�m=      �=       �U�                 =      =       u8                        =      )=       V)=      ,=       u ,=      <=       V<=      n=       v�q=      =       v�                   =      j=       ��j=      q=       0�q=      �=       ��                        D=      \=       P]=      l=       Pl=      p=       |�q=      ~=       P                      `4      �4       U�4       5       S 5      5       �U�                 `4      b4       u8                 `4      b4       u8#��                  m4      4       V4      �4       v��4      �4       v��4       5       v�                 m4      �4       ���4       5       0�                 4      �4       V�4      �4       v��4      �4       v��4       5       v�                   4      �4       U�4      �4       S                 �4      �4       v��4      �4       v��4       5       v�                 �4      �4       S                 �4      �4       v��4       5       v�                 �4      �4       S                 �4       5       v�                 �4      �4       S                            �@      >A       U>A      �B       ]�B      �B       �U��B      �C       ]�C      �C       �U��C      ED       ]                 �@      �@       u8                 �@      �@       u8#@�                 �@      �@       u8#p�                 �@      �@       u8#h�                                A      >A       _>A      �A        ~ "#��A      �A        ~ "��A      2B        ~ "#�2B      �B        ~ "��B      �C        ~ "��C      �C        ~ "#��C      �C        ~ "��C      ED        ~ "#�                   A      A       ��A      �B       0��B      ED       0�                       9A      >A      
 ��������>A      �B       V�B      �C       V�C      ED       V                         9A      >A      
 �       �>A      ?B       S?B      �B       s ��B      �C       S�C      ED       S                 9A      >A       0�                                �B      �B       P�B      �B       � r "�C      BC       PBC      KC       � r "��C      �C       P�C      �C       � r "��C      �C       P�C      �C       � r "�                      �B      �B       T'C      MC       T�C      �C       T                                �B      �B       Q�B      �B       t 1&�-C      DC       QDC      MC       t 1&��C      �C       Q�C      �C       t 1&��C      �C       Q�C      �C       t 1&�                         >A      �A       ]�A      �B       ]�B      �C       ]�C      �C       �U��C      ED       ]                       >A      �A        ~ "��A      2B        ~ "��C      �C        ~ "��C      ED        ~ "�                          >A      �A       P�A      �A       U�A      B       PB      /B       U�C      ED       P                                  >A      LA       5�LA      XA       6�XA      dA       7�dA      pA       8�pA      �A       9��C      �C       5��C      D       6�D      -D       7�-D      ED       8�                    p      �       U�      o       �U�                                        p      �       T�      	       �T�	      G       TG      t       �T�t      �       T�      �       �T��      �       T�             �T�             T      J       �T�J      m       Tm      o       �T�                            p      �       Q�      	       �Q�	      }	       Q}	      
       �Q�
      1       Q1      o       �Q�                        p      �       R�      	       V	      	       �R�	      o       V                           p      �       U	      _       Ut      �       U�      �       U      =       UJ      o       U                            �      �       P	      z	       P
      
       PB
      �
       P�
      �
       P             P                                �      �       4��      �       R�      �       R	      ?
       RB
      �
       R�
      g       Rt      �       R�      �       R      A       RJ      o       R                                             �      �       0��      �       X�      	       p �	      	
       0�	
      
       X
      o       0�o      t       Pt      �       0��      �       P�      �       0��      �       P�             X      E       0�E      J       PJ      o       0�                                                     �      �       0��      �       X	      ,	       X1	      <	       XF	      �	       X�	      �	       X�	      �	       P
      
       Q
      	
       X
      s
       X}
      7       X<      g       Xt      �       X�      �       X�      �       X      
       X
             P&      &       QJ      `       X`      e       Pe      o       X                                        �      �       0�	      z	       0��	      �	       ]�	      �	       Z�	      
       ^
      
       Z
      �
       0��
      �
       Z�
      �
       Z�
             z �             Z             0�      1       Zt      �       ]      o       ]                       p      �       0��      	       S	      	       S	      o       S                             p      �       0�	      z	       0�
      �
       0��
      �
       ^�
             ^             0�      1       ^                             �      �       0��      �       Y	      g       Yt      �       Y�      �       Y      A       YJ      o       Y                    �      �       0�1	      B	       {�B	      K	       [                                           �      �       0�	      \	       0�\	      �	       \�	      
       [
      
       0�
      1       \<      g       [t      t       \t      �       | } ��      �       \�      �       | ��      �       [�      �       [      &       \&      &       9�J      S       | } �`      o       \                  �	      �	       P                  �	      �	       Q                        �#      �#       U�#      $       S$      $       �U�$      }.       S                                          �#      �#       T�#      �#       \�#      $       �T�$      ^$       T^$      �)       \�)      �)       T�)      !+       \!+      �,       �T��,      �,       \�,      Q-       �T�Q-      m-       \m-      �-       �T��-      }.       \                              �#      �#       Q$      $       Q$      �)       ]�)      �)       Q�)      �+       ]�,      �,       ]Q-      m-       ]�-      }.       ]                                        �#      �#       R�#      �#       V$      D$       RD$      )       V)      �)       �R3!�R�R
  $0.( ��)      �)       R�)      s-       Vs-      �-       �R3!�R�R
  $0.( ��-      .       V.      Q.       �R3!�R�R
  $0.( �Q.      `.       V`.      }.       �R3!�R�R
  $0.( �                                                     �%      �%       P�%      �%       Y�%      �%       P�%      &       P&      L&       ��hL&      L&       0��&      '       P`(      p(       Pp(      G)       YG)      x)       ��h�)      �)       P�)      �)       Y�)      �)       P�-      .       ��h.      .       0�.      8.       ��h8.      Q.       YQ.      `.       P`.      }.       ��h                          �#      �#       ^$      �+       ^�,      �,       ^Q-      m-       ^�-      }.       ^                            .%      Z%       RZ%      �%       ��i&      m'       ��i�)      �)       ��i�)      �)       0��)      .       ��iQ.      `.       ��i                       .%      m'       v  1��)      s-       v  1�s-      .       ��i�1�Q.      `.       v  1�                                   �#      �#       0�$      �$       0��$      �%       ��h&      m'       ��hm'      %(       0�%(      *(       1�*(      �)       0��)      �)       ��h�)      �)       1��)      .       ��h.      Q.       0�Q.      `.       ��h`.      }.       0�                        �#      �#       _$      '       _m'      �)       _�-      }.       _                       �#      �#       ~�$      �$       ~�*(      P(       ~��)      �)       ~�                       �#      �#       ~�#P$      �$       ~�#P*(      P(       ~�#P�)      �)       ~�#P                               �$      m'      
 ��h���h��'      �'       T���'      �'       T�P��'      �'       ��h�P��'      *(      
 ��h���h��)      �-      
 ��h���h��-      .      
 ��h���h�Q.      `.      
 ��h���h�                     q$      �$       | *(      H(       QH(      X(       |                      q$      �$       | #�*(      H(       q�H(      P(       | #�                     q$      �$       | #�*(      H(       q�H(      X(       | #�                      x)      �)       1�.      8.       0�`.      }.       0�                    �'      �'       R�'      (       ��h                    �'      �'       X�'      *(       ��i                  '      �'       P�'      �'       q�                 �-      .       �
�                  .'      m'       P                 �)      �-       s0�                      �*      �*       1��,      �,       0��-      �-       0�                  �,      �,      	 q 0$0&�                   �+      5,       s���,      Q-       s��                         �+      �+       s��,      �,       s��,      -       P-      G-       pp�G-      Q-       P                   �+      �+       s��,      �,       s�                   �+      �+       s��,      �,       s�                �+      ,       s�                    �+      ,       R,      ,      
 p r "#���                  �+      ,       r ?&�,      ,       P                ,      #,       s�                    ,      #,       T#,      #,      
 p t "#���                  ,      #,       t ?&�#,      #,       P                  �,      -       p -      -       pp                   -      -       Q-      -      
 q x "#���                  -      -       q ?&�-      -       X                   --      4-       Q4-      4-      
 q x "#���                  --      4-       q ?&�4-      4-       X                D+      X+       ��i                D+      X+       s�                    V+      X+       PX+      X+      
 p q "#���                  V+      X+       p ?&�X+      X+       Q                o+      y+       ��i                o+      y+       s�                    w+      y+       Py+      y+      
 p q "#���                  w+      y+       p ?&�y+      y+       Q                   �#      �#       �
��)      �)       �
�                    �#      �#       ]�)      �)       ]�)      �)       Q                    �#      �#       0��)      �)       0��)      �)       ]                    `      i       Ui      j       �U�                 `      i       u�                    P      X       UX      Y       �U�                    P      X       TX      Y       �T�                    P      X       QX      Y       �Q�                 P      X       u�                    @      I       UI      J       �U�                    @      I       TI      J       �T�                 @      I       u�                    0      9       U9      :       �U�                    0      9       T9      :       �T�                    0      9       Q9      :       �Q�                 0      9       u�                           )       U)      *       �U�                           )       T)      *       �T�                           )       Q)      *       �Q�                        )       u�                                 U             �U�                                 T             �T�                              u�                           	       U	      
       �U�                           	       T	      
       �T�                           	       Q	      
       �Q�                        	       u�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                 �      �       u�                      �      �       R�      �       u��      �       R                       �      �       t ����1$r�
"�
����      �       t ����1$r "�
����      �       t 1$r "�
����      �       t 1$u�#�
"�
���                   �      �       r���      �       u�#��                  w      �       P                       �       p��                    �      �       U�      _       �U�                          �      �       T�             ]      #       �T�#      2       T2      _       ]                          �      �       Q�             \      #       �Q�#      9       Q9      _       \                          �      �       R�             V      #       �R�#      9       R9      _       V                     �             0�#      /       6�/      _       0�                    �             S#      _       S                   �             s��#      _       s��                              �      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U��      �       U                              �      �       T�      �       V�      �       T�      �       �T��      �       V�      �       �T��      �       T                             �      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U��      �       U                   �      �       u �      �       u                    �      �      	 u #�#�      �      	 u #�#                  �      �       P                  �      �       P                                          U      +       �U�+      C       UC      l       Sl      n       Un      o       �U�                          *       V+      m       V                                  u�+      C       u�C      G       s�                 :      G       p                  H      V       P                  W      _       P                        �      �       U�      �       �U��      �       U�      �       �U�                          �      �       T�      �       V�      �       �T��      �       T�      �       V                    �      �       \�      �       \                 �      �       |��                     �      �       0��      �       P�      �       S                   �      �       u��      �       U                               P                           5       P5      L       }y�                    6      �       P�      �       P                    ;      �       ]�      �       ]                        `      �       U�      �       �U��      �       U�      �       �U�                        `      �       T�      �       S�      �       �T��      �       S                    q      �       \�      �       \                 �      �       |��                     �      �       0��      �       P�      �       V                   �      �       u��      �       U                                p      �       U�      �       V�             �U�      K       VK      a       �U�a      t       Vt      y       Uy      z       �U�                            p      �       T�      [       S[      a       �T�a      s       Ss      y       Ty      z       �T�                    �      `       ]a      x       ]                   �      `       }�
�a      x       }�
�                   �      �       P�             V                    �      �       T             P                        �      �       U�      �       p 1$q "�      �       | ����1$q "             U                    �      �       0��             \                         $       u$      -       U                  .      <       P                  =      F       P                 �      �       v�                    �      �       P�             V                 �      �       ]                  �      �       U                                �.      T/       UT/      �/       \�/      �/       �U��/      �/       U�/      0       \0      0       �U�0      P0       UP0      �0       \                              �.      
/       T
/      T/       ST/      �/       �T��/      �/       S�/      0       �T�0      P0       SP0      �0       �T�                            �.      T/       QT/      �/       �Q��/      �/       Q�/      0       �Q�0      P0       QP0      �0       �Q�                              �.      T/       RT/      �/       �R��/      �/       R�/      �/       R�/      0       ]0      P0       RP0      �0       �R�                              �.      T/       XT/      �/       �X��/      �/       X�/      �/       V�/      0       �X�0      P0       XP0      �0       �X�                             ?/      �/       0��/      �/       1��/      �/       0��/      �/       1��/      0       0�70      {0       0�{0      �0       1�                         �.      �/       0��/      �/       P�/      �/       0��/      0       P0      �0       0�                          �.      J/       _J/      T/       u��/      0       _0      F0       _F0      P0       u�                       /      T/       UT/      �/       \0      P0       UP0      �0       \                              �.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U                              �.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T                              �.      �.       Q�.      �.       �Q��.      �.       Q�.      �.       �Q��.      �.       Q�.      �.       �Q��.      �.       Q                              �.      �.       R�.      �.       �R��.      �.       R�.      �.       �R��.      �.       R�.      �.       �R3!��.      �.       R                             �.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U                             �.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T                             D       UD      N       �U�N      S       U                             D       TD      N       �T�N      S       T                             D       QD      N       �Q�N      S       Q                               D       RD      M       SM      N       �R�N      S       R                            D       UD      N       �U�N      S       U                      '      D       PN      R       PR      S       u�                                  U             �U�                                  T             �T�                               u                                u #�                              
 u #�#�&                    �       �        U�       �        �U�                    �       �        T�       �        �T�                 �       �        u                  �       �        u #�                 �       �       
 u #�#�&                      @      R       UR      g       Sg      h       �U�                 @      A       u                  @      A       u #�                        �       �        U�       �        T�       �        �U��       �        T                    �       �        T�       �        �T�                    �       �        Y�       �        Y                    �       �        U�       �        U                       �       �        P�       �        y��       �        P�       �        y�                       �       �        p�
��       �        y�#�
��       �        p�
��       �        y�#�
�                      �       �        R�       �        y�#�&�       �        R                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  �      �       U                 �      �       u�
�                     �      �       t ����1$u�
"�
����      �       t 1$u�
"�
����      �       �T����1$u�
"�
���                     P       t        0�t       x        Px       �        0��       �        P                  R       i        Q                     b       i        q�i       x        Qx       |        q��       �        Q                    0       D        TD       E        �T�                 0       D        0�                                 u                                  u #�                                 u #�#��                      �      �       U�      �       �U��      �       U                    �      �       P�      �       P                 �      �       U�      9       u�                                  �      �       Q�      �       u ����      �       Q�      �       u ����      �       Q�             u ���      +       Q+      2       q��2      9       u ���                             �      �       0��      �       P�      �       0��             0�             P      8       0�8      9       P                 �      �       T                 �      �       U                 �      �       P                      @      b       Ub      d       �U�d      �       U                            @      c       Tc      d       �T�d      n       Tn      �       �T��      �       T�      �       �T�                    d      n       Tn      �       �T�                  d      �       U                 n      �       U                  n      �       T                 �      �       U                 �      �       u�                    �      �       S�      �       S                    �      �       P�      �       P                             /       Q/      p       Vp      q       �Q�                      9      n       Pn      p       v p      q       �Q                        8       U                            H       0�H      Y       Q`      q       Q                    ?      H       0�H      ]       R                        �"       #       U #      #       �U�#      '#       U'#      :#       �U�                        �"      #       T#      #       �T�#      2#       T2#      :#       �T�                            �"      #       Q#      #       S#      #       �Q�#      2#       Q2#      8#       S8#      :#       �Q�                            �"      #       R#      #       V#      #       �R�#      2#       R2#      9#       V9#      :#       �R�                  #      #       P                    #      2#       R2#      3#       V                    #      2#       Q2#      3#       S                    #      2#       T2#      3#       �T�                    #      '#       U'#      3#       �U�                     #      '#       u�'#      .#       U.#      2#       u�u�                        @#      [#       U[#      q#       �U�q#      �#       U�#      �#       �U�                        @#      b#       Tb#      q#       �T�q#      �#       T�#      �#       �T�                        @#      k#       Qk#      q#       �Q�q#      �#       Q�#      �#       �Q�                    q#      �#       Q�#      �#       �Q�                    q#      �#       T�#      �#       �T�                    q#      �#       U�#      �#       �U�                  #      �#       P                 #      �#       p�
�                   #      �#       T�#      �#       �T�                 �#      �#       p�
                      �0      �0       U�0      1       V1      1       �U�                      �0      �0       T�0      1       S1      1       �T�                          �3      �3       Q�3      54       X54      D4       QD4      E4       �Q�E4      ]4       X                          �3      �3       P�3      4       R4      4       P4      54       RE4      ]4       R                          PD      ZD       UZD      sD       \sD      tD       �U�tD      �D       \�D      �D       �U�                            PD      cD       TcD      qD       VqD      tD       �T�tD      �D       V�D      �D       T�D      �D       �T�                        gD      lD       PlD      pD       SpD      �D       P�D      �D       S                      }D      �D       V�D      �D       T�D      �D       �T�                    }D      �D       \�D      �D       �U�                  �D      �D       U                  �D      �D       P                                �D      �D       U�D      	E       V	E      E       �U�E      FE       VFE      KE       �U�KE      iE       ViE      nE       UnE      oE       �U�                            �D      �D       T�D      �D       S�D      E       �T�E      E       TE      BE       SBE      oE       �T�                                  �D      �D       Q�D      E       ]E      E       �Q�E      $E       Q$E      JE       ]JE      KE       �Q�KE      mE       ]mE      nE       QnE      oE       �Q�                                  �D      �D       R�D      E       \E      E       �R�E      $E       R$E      HE       \HE      KE       �R�KE      kE       \kE      nE       RnE      oE       �R�                      �D      �D       UE       E       U E      $E       v�                  �D       E       P                   �D      �D       s ����1$u�
"�D      �D       �T����1$u�
"                          E      $E       R$E      9E       \KE      kE       \kE      nE       RnE      oE       �R�                          E      $E       Q$E      9E       ]KE      mE       ]mE      nE       QnE      oE       �Q�                      E      9E       SKE      hE       ShE      nE       T                        E      9E       VKE      iE       ViE      nE       UnE      oE       �U�                 E      $E       v�#                  %E      3E       P                    4E      9E       PKE      SE       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 `      �       u��                    �              P             u�                 `       �        U                        P      �       U�      -       S-      3       �U�3      9       U                       P      �       U�      -       S-      3       �U�3      9       U                  t      2       ]                     b      �       u���      -       s��-      3       �U#��                     b      �       u���      -       s��-      3       �U#��                      y      �       0��      �       \�      �       |�                  �      �       V                      �      �       U�      #       S#      $       �U�                    �      �       T�      $       �T�                               P                      0      ;       U;      �       S�      �       �U�                     0      ;       U;      �       S�      �       �U�                   0      s       0�s      �       P                    C      E       PE      r       X                    M      p       Qp      r       s                    M      p       q
Pq�"�p      r       r 
Ps #�"�                   M      p       q
Pq�"�p      r       r 
Ps #�"�                      �      �       U�      �       S�      �       �U�                      �      �       P�      �       u�      �       s                  �      �       V                  �      �       P                  �      �       P                              /        U/       D        �U�D       K        U                                        T       1        Q1       D        �T�D       K        T                  ,       C        S                        �      �       U�              \       #       �U�#      �       \                    �      �       T�      �       �T�                       �      �       u���              |��       #       �U#��#      �       |��                    �             V#      �       V                    �      "       ]#      �       ]                      �      �       P�             S#      �       S                 ]      |       0�                   |      �       q|��      �       q�}�                      @      �       U�             V             �U�      �       V                      @      �       T�      �       P�      �       �T�                  w             s  $ &
P| "�      �       s  $ &
P| "�                     @      �       U�             V             �U�      �       V                   �             ]      �       ]                  w             s  $ &
P| "#��      �       s  $ &
P| "#��                  w             s  $ &
P| "#��      �       s  $ &
P| "#��                    �      �       P�      �       Q                        �      �       U�      ^       S^      s       �U�s      E       S                              �      )       T)      #
       ]#
      s       �T�s      �       T�      �       ]�      *       �T�*      E       ]                                �             Q      �       ^�      s       �Q�s             Q      �       ^�      �       �Q��      �       ^�      E       �Q�                                  �             R      P       VP      ^       ��g� �s      {       R{      �       V�      �       ��g� ��             V      *       ��g� �*      E       V                       �      �       U�      ^       S^      s       �U�s      E       S                                    �      �       P�      �       _�      �       P�      ^       _�      �       _�      �       0��      �       P�      %       _%      *       0�*      E       _                    �      �	       \s      �       \                             p      �      
 v 3 $0)��      	       P	      "	       s�"	      ^       ��g�      �       ��g�      �      
 v 3 $0)��      E       ��g                             p      	       v  1�	      	       P	      "	       s�"	      ^       ��g�      �       ��g�      �       v  1��      E       ��g                   �      :       |�s      �       |�                       	      	       ��g�^�	      ^       �^��      �       �^��      E       �^�                       �      �       0��      #	       1�#	      ^       0�s      �       0��      �       1��      E       0�                  �      �       V                   A	      ^       s0��      E       s0�                  x
      �
      	 q 0$0&�                   S
             ��h�             ��h                         S
      �
       ��h#�
      �
       P�
      �
       pp��
      �
       P�             ��h#                   S
      �
       s��             s�                   S
      �
       s��             s�                  �
      �
       p �
      �
       pp                   �
      �
       Q�
      �
      
 q y "#���                  �
      �
       q ?&��
      �
       Y                   �
      �
       Q�
      �
      
 q y "#���                  �
      �
       q ?&��
      �
       Y                �
      �
       s�                    �
      �
       U�
      �
      
 p u "#���                  �
      �
       u ?&��
      �
       P                �
             s�                                 T            
 p t "#���                               t ?&�             P                �	      �	       ��g                �	      �	       s�                    �	      �	       P�	      �	      
 p q "#���                  �	      �	       p ?&��	      �	       Q                
      
       ��g                
      
       s�                    

      
       P
      
      
 p q "#���                  

      
       p ?&�
      
       Q                                   ]       U]      �       V�      �       �U��      �       V�      �       U�      �       V                               f       Tf      �       ��k�             T      �       ��k                                �       _�      �       _�             _             U�      �       _                               �       ���      �       ���             ��             u���      �       ��                            �      �       P�      �       P`      v       Qv      �       x� �      �       P�      �       P�      �       P�      �       Q                    �      &       S�      �       S�      �       S                      *      f       X�      "       X"      ?       ��k                                   2      �       0��      �       ]�      �       0��      �       ]�      �       0��      �       P�      �       ]�      ^       0�^      b       Pb      �       ]�      �       0�                        6      =       P=      �       w �      �       ��k�      �       w                                   6      �       0��      �       ��k�      �       0��      �       ��k�      �       0��      �       P�      �       ��k�      ;       0��      �       0��      �       0�                          B      I       PI      f       �f      �       ��k�      "       �"      �       ��k                           B      �       0��      �       \�      �       0��      �       \�      z       0�z      �       1��      �       0�                    M      �       ^�      �       ^                   �      �       T�      �       T                  �      �       ���  �      �       ���                       �      �       0��      �       S�      �       0�                   �      �       P�      �       P                    
      n       S�      �       S                   �             R      @       ��k                  �      6       \�      �       0�                   `      �       T�      �       T                  `      �       ���  �      �       ���                       `      v       0�v      �       S�      �       0�                    `      �       Q�      �       q��      �       Q�      �       Q                     �      �       Q�      �       ��      �       Q                   �      �       ���  �      �       ���                      �      �       0��      �       R�      �       0�                    �      �       P�      �       p��      �       P�      �       P                �      �       �                �      �       ���                    �      �       0��      �       \                  �      �       P�      �       p��      �       P                      <      �       S�      �       S�      &       S                    �             P      &      
 s 4$�"�                     w      �       P�      �       ��k�      �       P                 �      �       U                    �      �       S�      �       S                    �      �       P�      �       P                        �      �       U�      �       S�      �       �U��      �       U                       �      �       U�      �       S�      �       �U��      �       U                      �      �       U�      �       S�      �       �U�                  �      �       P                                    �             U             S      4       �U�4      �       S�      �       �U��      �       S�      e       �U�e      �       S�             �U�             S      �$       �U�                                                          �             T             ]      4       �T�4      �       ]�      �       �T��      �       ]�      F       ��{F      X       �T�X      �       ��{�      �       �T��      &       ��{&      e       �T�e      t       Tt      �       ]�      �       ��{�             �T�             ]      6       �T�6      E       ��{E      �       �T��      �       ��{�      �$       �T�                        �             Q      e       ��{e      |       Q|      �$       ��{                        �             R      e       �R�e      |       R|      �$       �R�                        �             X      e       �X�e      |       X|      �$       �X�                                                         �             T             ]      4       �T�4      �       ]�      �       �T��      �       ]�      F       ��{F      X       �T�X      �       ��{�      �       �T��      &       ��{&      e       �T�e      t       Tt      �       ]�      �       ��{�             �T�             ]      6       �T�6      E       ��{E      �       �T��      �       ��{�      �$       �T�                                     P4      ?       P?             X9      K       6�                         �             t�e      t       t�t      |       }�}      �       P             P                                  t��      �       }��      �       P                          4      �       S�      �       �U��      �       S�      e       �U��             �U�      �$       �U�                      4      e       �R��             �R�      �$       �R�                      4      e       �X��             �X�      �$       �X�                      4      e       ��{�             ��{      �$       ��{                                              4      �       ]�      �       �T��      �       ]�      F       ��{F      X       �T�X      �       ��{�      �       �T��      &       ��{&      e       �T��      �       ��{�             �T�      6       �T�6      E       ��{E      �       �T��      �       ��{�      �$       �T�                                  �       X�      �       X9      e       X�      F       XF      K       ��{�             X                           4             ��{�      �       ��{�      9       ��{�      �       ��{K      �       ��{      �$       ��{                                           4      �       ]�             �T��      �       ]�      F       ��{F      X       �T�X      �       ��{�      &       ��{&      9       �T��      �       ��{K      �       �T�      6       �T�6      E       ��{E      �       �T��      �       ��{�      �$       �T�                               v             U      e       ^�      �       ^�      �       U�             ^              ^               U       �$       ^                                   v             R      �       ��{�      �       ��{�      9       ��{�      �       ��{K      �       ��{      �        ��{)#      ]#       ��{g#      y#       ��{8$      <$       ��{                       �       0�                                             v      �       }���      �       �T#���      �       }���      F       ��{#��F      X       �T#��X      �       ��{#���      �       �T#���      &       ��{#��&      e       �T#���      �       ��{#���             �T#��      6       �T#��6      E       ��{#��E      �       �T#���      �       ��{#���      �$       �T#��                            �       U       ,        U,       x       	 }��                         �       z { " $ &�       x        z { " $ &�                                             v      �       ]�      �       �T��      �       ]�      F       ��{F      X       �T�X      �       ��{�      �       �T��      &       ��{&      e       �T��      �       ��{�             �T�      6       �T�6      E       ��{E      �       �T��      �       ��{�      �$       �T�                	v      v       U                   v      ~       Q~             }�                           v             R      �       ��{�             ��{X      �       ��{�      &       ��{�      �       ��{6      E       ��{�      �       ��{                           v      �       V�      �       U�             VX      �       V�      &       V�      �       V6      E       V�      �       V                           v             U      �       ^�             ^X      �       ^�      &       ^�      �       ^6      E       ^�      �       ^                                  �      �       P�      �       2��      �       0�B      W       P�      �       P�      ;       P             0��      �       P�      �       P             3�@      E       3��      �       0�                            �      �       P�      �       ��{�             ��{X      �       ��{�      &       ��{�      �       ��{6      E       ��{�      �       ��{                                        �       ]�      �       P�             w X      �       ]�      �       P�      �       ]�      �       }�~��      �       ]�      &       w �      �       w 6      ;       ]�      �       w                           �             S      ;       ��};            	 w ��{��      &      	 w ��{��      �      	 w ��{��      �      	 w ��{�                        i      �       _�      �       Q�      �       _�      �       ~                                \      �       Yd      �       \�      �       ��{�             |	�X      �       Y�      &       |	��      �       }�6      E       Y�      �       |	�                          5      ;       X;      �       ��{�      �       X�      �       S�      	       X�      &       X                      N      �       S�      �       _�             S�      &       S�      �       S                        �             
	�      :       S:      �       _X      �       _�      �       
 �                         �             0�      �       w X      �       w �      �       w �      �       9�6      E       w                             �             ��}�      \       \\      p       P�      �       P�      �       P�      �       ��}��      �       \6      @       P                    *      3        p �3      :       _                 �      �       P                 �              ^                 �              ^                 �              ^                 �      �       ��|                  &      F       ��}                  &      F       \                                  &      �       ^K      �       ^�      �       U�             ^�              ^               U               ^)#      T#       ^g#      y#       ^                  &      F       ]                                   &      X       ^K      �       ^�      �       U�             ^      �       ^      6       ^E      �       ^�              ^               U       �$       ^                                       B      {       \�      �       \�      �       \�      �       VK      ]       \]      �       V�      �       v��      �       P�      �       v��             V�              v�               v�)#      T#       v�g#      y#       v�                               B      F       SF      �       w #�K             w #��      �       w #��              w #�               w #�)#      T#       w #�g#      y#       w #�                    t      �       PT      i       P                            �      �       Q�      �       ��{�              ��{               ��{)#      T#       ��{g#      y#       ��{                                    �      b       Sb      �       _�      �       T�      �       _�      �       S�              _               T               _)#      T#       _g#      y#       _                    �      ]       ]�      �       ]                      !      9       1�9      I       PP      U       P                             ]      �       _�      �       T�      �       _�              _               T               _)#      T#       _g#      g#       _                             ]      �       ^�      �       U�      �       ^�              ^               U               ^)#      T#       ^g#      g#       ^                       ]      �       ]�              ]               ])#      T#       ]g#      g#       ]                      �      �       P               P7#      <#       Pg#      g#       ��                             ]      �       ^�      �       U�      �       ^�              ^               U               ^)#      T#       ^g#      g#       ^                        �      �       P               PC#      H#       PO#      T#       P                       ]      �       }���              }��               }��)#      T#       }��g#      g#       }��                  �              P                             �      �       ]�      X       w       �       w       6       w E      b       w                w T#      ]#       w                   �      �       T                  �      �       \                    �      �       P�      �       V                         �      X       S      �       S      6       SE      b       S               ST#      X#       S                      �      �       Ph      w       Pb      b       0�T#      X#       P                                      �      �       ��}��      �       P�             Q             q�      X       Q      7       Qp      �       ��}��      �       R�      �       Q      (       QE      U       QU      Y       q�Y      b       Q               Q                     �      �       ��}��      �       P�      �      
 � p "
P�                                  �      �       V�             U      X       V      '       V'      ,       U,      �       V      6       VE      ^       V               VT#      X#       V                          �      X       \      �       \      6       \E      b       \               \T#      X#       \                      �      �       RT      X       R      #       R                                 �      �       1��      
       ]
             R      X       ]      �       ]      ,       ]E      b       ]               ]T#      X#       ]                                �      �       0��             T      X       0�      ,       T,      �       0�      6       0�E      ^       0�               0�T#      X#       0�                     ?      T       PT      �       _T#      X#       _                     ?      B       q p �B      c       Qc      g       s �                        /      r       Rr      �       }��      �       r�}��      �       r�z��      �       }�                       H       )#       ]]#      g#       ]y#      /$       ]8$      �$       ]                     H       )#       }��]#      g#       }��y#      �$       }��                          o       x        Ux       )#       w ]#      g#       w y#      /$       w 8$      �$       w                        o       )#       _]#      g#       _y#      /$       _8$      �$       _                                    �       #       ��{#      $#       ��{�#�]#      g#       ��{y#      �#       ��{�#      �#       0��#      �#       \<$      p$       ��{p$      y$       0�y$      ~$       P~$      �$       ��{                        �       #       ��{]#      g#       ��{y#      $       ��{<$      �$       ��{                             o       �        0��       )#       ��{]#      g#       ��{y#      $       ��{8$      <$       0�<$      �$       ��{�$      �$       R                                   o       �        0��       -!       \-!      =!       P=!      )#       \]#      g#       \y#      �#       \�#      ($       S($      /$       0�8$      <$       0�<$      p$       \p$      y$       Sy$      �$       \�$      �$       S                          t       x        Px       )#       ��{]#      g#       ��{y#      /$       ��{8$      �$       ��{                          �       `"       S]#      g#       Sy#      �#       S�$      �$       S�$      �$       }�{ "�                                 �       !!       s!!      #       ��{]#      g#       ��{y#      $       ��{<$      y$       ��{~$      �$       ��{�$      �$       s�$      �$      	 }�{ "#�$      �$       ��{                            �!      �!       0��!      �!       T�!      �!       1��"      �"       p��"      �"       p�]#      g#       TI$      d$       S                            �       )#       V]#      g#       Vy#      �#       V�#      $       ��{�1�<$      y$       V~$      �$       V                 ."      A"       ��{                     �!      �!       P�!      �!       X]#      g#       P                      �       !!       P!!      =!       ��{�$      �$       P                    �!      �!       s�]#      g#       s�                   �!      �!       ��  ]#      g#       ��                       �!      �!       0��!      �!       Q]#      g#       0�                    �!      �!       P�!      �!       p��!      �!       P]#      g#       P                 �"      �"       p3$| "p 3$| "�                   I$      d$       s3$| "s 3$| "�d$      f$       s 3$| "s3$| "�                         #      �       }���      �       }��9      e       }���      9       }���             }��                         #      �       }���      �       }��9      e       }���      9       }���             }��                          �      �       T9      H       TH      L       t�L      X       TX      `       t�`      e       T�             T                     �      �       Q9      e       Q�             Q                        �             U             �U�      �       U�      �       �U�                            �      �       T�             T      (       0�d      w       0��      �       T�      �       �T1�                              �             Q             Q      &       Q&      (       �Q�d      q       Qq      s       �Q�s      }       Q�      �       0�                              �      �       R�             \             �R�      (       R(      d       \d      n       Rn      �       \                       �             U             �U�      �       U�      �       �U�                           �             0�      �       0��      �       P�      �       P�      �       �L�      �       P                       �             u��             �U#��      �       u���      �       �U#��                        /      =       p t "=      @       V@      d       u�t "�      �       u�t "                       /      =       p q "=      d       u�q "�      �       u�q "�      �      
 �U#�q "                    B      d       V�      �       V                   B      d       S�      �       S                     B      d       u��      �       u��      �       �U#�                      �             Q      �       s����      �       s���                    �      �       X�      �       X                                   R      �      2 @K$Os��(  / 0@K$(	 1$#/��O'�%��      �      2 @K$Os��(  / 0@K$(	 1$#/��O'�%�                          �       T�      �       T                                      q r �             Q             s��r �      �      : s��@K$Os��(  / 0@K$(	 1$#/��O'�%��      �      : s��@K$Os��(  / 0@K$(	 1$#/��O'�%�                             8       U8      �       }� �      �       U�      �       }�                          �       Y�      �       Y                         �       [�      �       [                                             ,       Q,      F       ZF      V       QV      `       Zl      �       Q�      �       Z�      �       }� �      �       Z�      �       Q�      �       Z�      �       }� �      �       Z                            0      F       QX      `       R�      �       R�      �       Q�      �       Q�      �       Q                  �      �       R                                        @      �       U�      �       V�      �       �U��      ;       U;      �"       V�"      �"       �U��"      �$       V�$      %       �U�%      *%       V*%      �%       �U��%      �%       V�%      W&       �U�                              @      �       T�      �       _�      �       �T��      @       T@      �$       _�$      %       �T�%      �%       _�%      W&       �T�                                      @      Z       QZ      �       S�      �       �Q�Q $0.��      �       S�      �       �Q�Q $0.��      �       S�      �       �Q�Q $0.��      L"       SL"      �"       �Q�Q $0.��"      �$       S�$      W&       �Q�Q $0.�                                        @      �       R�             ^      �       �R��      �       R�      �       ^�      �       �R��      v"       ^v"      �"       �R��"      �$       ^�$      %       �R�%      �%       ^�%      W&       �R�                                       @      �       U�      �       V�      �       �U��      ;       U;      �"       V�"      �"       �U��"      �$       V�$      %       �U�%      *%       V*%      �%       �U��%      �%       V�%      W&       �U�                             @      �       T�      �       _�      �       �T��      @       T@      �$       _�$      %       �T�%      �%       _�%      W&       �T�                                     P      �       \�      �       \�$      %       0�                        T      �       ]�      ?       ]?      t       ��      -       ��                    �      �       S�      �       S                                       T      �       u���      �       v���      �       �U#���      ;       u��;      �"       v���"      �"       �U#���"      �$       v���$      %       �U#��%      *%       v��*%      �%       �U#���%      �%       v���%      W&       �U#��                      �      �       Q�      �       ���      �       ��                         �       v0��      �       v0�                      �      �       P�      �       P�      �       P                 �      �       Q                 �      �       T                          �       ~  $0)��      �       ~  $0)�                 �      �       0�                 �      �                         �      �       (                      �      �       P�      ?       pp�?      U       P                  �      �       p �      
       pp                         
       Q
      
      
 q y "#���                        
       q ?&�
      
       Y                   %      ,       Q,      ,      
 q y "#���                  %      ,       q ?&�,      ,       Y                D      Y       X                   N      Y       UY      Y      
 p u "#���                  N      Y       u ?&�Y      Y       P                  k      r       Tr      r      
 p t "#���                  k      r       t ?&�r      r       P                    �      �       X�             ��~                  �             \                    �      �       Q�             ��                    �      �       T�             w                       �              v��              U             v��                               �      �       r @B$ $0.��      �       ~ @B$ $0.��      v"       ~ @B$ $0.�v"      �"       �R@B$ $0.��"      �$       ~ @B$ $0.��$      �$       �R@B$ $0.�%      �%       ~ @B$ $0.��%      W&       �R@B$ $0.�                           �      �       S�      L"       SL"      �"       �Q�Q $0.��"      �$       S�$      �$       �Q�Q $0.�%      W&       �Q�Q $0.�                         �      @       T@      �       _�      �$       _�$      �$       �T�%      �%       _�%      W&       �T�                                   �      ;       U;      �       V�      �"       V�"      �"       �U��"      �$       V�$      �$       �U�%      *%       V*%      �%       �U��%      �%       V�%      W&       �U�                                        |      �       P�      �       P�      
       0��              P       !        P!       �        \�       �!       0��!      '"       P'"      �"       \�"      	#       0�	#      �$       \�$      �$       \�$      �$       0�%      W&       \                     �      ?       ]?      t       ��      -       ��                 �      {       }�                     �      ?       }��?      t       ��#��      -       ��#��                    {      �       \�$      �$       \                        �      
       ��T      �!       ���"      �$       ���$      �$       ��                 �      {       s ����4$}�"�                      �      8       \8      t       ��      -       ��                 �             0�                         /      Q       4�Q      g       Qg      w       |�1r  $0)#�w      {       Q{      �       ��~                     �      �       ��:        {       ��:  �$      �$       ��:                       �      �       ��:        {       ��:  �$      �$       ��:                       �      �       Y      {       Y�$      �$       Y                     �      8       |�8      t       ��#�      -       ��#�                   �      �       T      -       T                     �      �       [      {       [�$      �$       [                      �      �       U-      {       U�$      �$       U                          �      �       T�      �       Q�      �       T-      {       T�$      �$       T                       �      �       4��      �       X      {       X�$      �$       X                     �             u 1�      �       ��~�1�      -       ��~�1�                            �      �       \�      �       R�      �       \-      j       \j      v       |��$      �$       \�$      �$       |��$      �$       \                            ?       [?      t       Q      -       Q                          �       U      -       U                      ?      O       Pe      t       P      -       P                             ?       	��?      ?       R?      O       PO      t       R      -       P                          �      �       Q�      �       Q-      3       Q3      {       u t "1%��$      �$       u t "1%�                      �      �       P�      �       P-      8       P                       �      
       [�      �        0��       �!       [�"      	#       [	#      �$       0�                       �      
       ���      �        0��       �!       ���"      	#       ��	#      �$       0�                                 �      
       ��~�      �       P�      �       P�      �       P�      �        ��~�       �!       ��~�"      E$       ��~J$      y$       ��~~$      �$       ��~                         �      
       Q�      �        0��       '!       Q'!      �!       v��"      	#       Q	#      �$       0�                         �      
       P�      �        0��       a!       Pa!      �!       v��"      	#       P	#      �$       0�                              �      
       z ���      �        0��       �!       z ���!      �"      	 ��~����"      	#       z ��	#      �$       0��$      �$      	 ��~���%      W&      	 ��~���                                             �      
       Y!       h        Ph       �        t� �       �        w #@�       �!       Y�!      �"       ���"      	#       Y	#      �#       w #@�#      �#       P�#      �#       t� �#      �#       P�#      �#       w #@�#      $       P$      &$       t� &$      �$       w #@�$      �$       ��%      W&       ��                   %       �        �A=  	#      �$       �A=                     %       �        �=  	#      �$       �=                     %       �        �4=  	#      �$       �4=                     %       �        �'=  	#      �$       �'=                     %       �        �=  	#      �$       �=                     %       �        � =  	#      �$       � =                          %       �        ��~	#      E$       ��~J$      y$       ��~~$      �$       ��~                               %       �        R�       �        w #H	#      7$       R7$      J$       w #HJ$      `$       R`$      ~$       w #H~$      �$       R�$      �$       w #H                   %       �        �N=  	#      �$       �N=                    %       �        0�	#      �$       0�                                 6       �        Z�       �        z 2%��       �        T�       �        z 2%��       �        z 4%��       �        T�       �        z 4%��       �        w #@�4%�	#      �#       z 2%��#      &$       Z&$      �$       z 4%�                           h       n        Pn       u        [u       �        t� ##      "#       P"#      %#       Q%#      -#       t                                      %       2        P2       9        Q9       d        p�d       �        Y	#      #       Y#      -#       T-#      :#       Y:#      U#       y�U#      X#       u~�X#      e#       Ue#      r#       Yr#      v#       y�v#      �#       T�#      �#       p��#      �#       p��#      �#       Y�#      �#       p��#      �#       p��#      �#       Y�#      �#       p��#      $       p�$      $       t� #�$      3$       Y3$      J$       TJ$      W$       YW$      ~$       T~$      �$       Y�$      �$       T                                6       }        0�}       �        [	#      �#       [�#      �#       0��#      �#       [�#      �#       0��#      �#       [�#      $       0�$      �$       [                                  6       �        0��       �        P�       �        ��	#      �#       ���#      �#       0��#      �#       P�#      �#       0��#      �#       P�#      !$       0�!$      &$       P&$      �$       ��                              6       �        0��       �        ��~	#      E$       0�E$      J$       UJ$      y$       0�y$      ~$       U~$      �$       0��$      �$       U                                  6       �        0��       �        Q	#      (#       0�(#      -#       Q-#      X#       0�X#      e#       Qe#      v#       0�v#      �#       Q�#      &$       0�&$      �$       Q                                6       �        0��       �        P	#      (#       0�(#      -#       P-#      `#       0�`#      e#       Pe#      {#       0�{#      �#       P�#      &$       0�&$      �$       P                            "      �"       v���"      �"       �U#���$      �$       �U#��%      *%       v��*%      �%       �U#���%      �%       v���%      W&       �U#��                     "      p"       }��2�%      #%       }��2��%      �%       }��2�                    "      �"      	 ��~����$      �$      	 ��~���%      W&      	 ��~���                            "      �"       Y�"      �"       ���$      �$       ��%      *%       Y*%      �%       ���%      �%       Y�%      W&       ��                    "      �"       0��$      �$       0�%      W&       0�                                               '"      -"       P��-"      B"       P�R��B"      H"      
 P�v���H"      H"      
 P�v���H"      �"       P�R���"      �"       ]�R���"      �"       P�R���"      �"       ]�R���$      �$       ]�R��%      *%       P�R��*%      0%       [�R��0%      >%       P�R��>%      �%       [�R���%      �%       P�R���%      �%       ]�R���%      �%       P�R���%      W&       ]�R��                 "      P"       }��2�                 "      P"       v��                 "      P"       ��>                     �"      �"       Y�$      �$       Y                   �"      �"       S�$      �$       S                   �"      �"       X�$      �$       X                   �"      �"       U�$      �$       U                       �"      �"       V�"      �"       v ���"      �"       V�$      �$       V                       �"      �"       [�"      �"       T�"      �"       [�"      �"       {��"      �"       [�$      �$       [                    �"      �"       P�"      �"       P�$      �$       P                       �"      �"       z 1%��"      �"       ���"      �"       Z�"      �"       z 1%��"      �"       Z�"      �"       ���$      �$       Z                     �"      �"       ^�"      �"       0��"      �"       ^�"      �"       0��$      �$       ^                   %      N%       YN%      V%       y�V%      �%       Y                 %      �%       ��>                      %      %       Q%      �%       U                  (%      �%       S                       %      *%       T*%      ,%       Z,%      >%       T>%      b%       Zb%      f%       z�f%      �%       Z                  %      0%       P0%      �%       P                         %      *%       ��*%      ,%       x 1%�,%      >%       ��>%      b%       Xb%      k%       x 1%�k%      o%       Xo%      }%       ��}%      �%       X                   %      *%       0�*%      �%       ]                       %      *%       0�*%      0%       Q0%      >%       0�>%      o%       Qo%      }%       0�}%      �%       Q                      �%      �%       Y�%      &       Y&      &       y�&      B&       Y                         �%      �%       [&      &       1�&      &       [-&      -&       0�-&      @&       [B&      W&       [                     �%      &       X-&      :&       XB&      W&       X                        �%      �%       �^��%      &&       �^�-&      2&       �^�2&      B&       �^�                  �%      W&       U                      �%      �%       V�%      �%       v ���%      W&       V                      �%      �%       S�%      �%       T�%      �%       S�%      �%       s��%      W&       S                   �%      �%       P�%      W&       P                        �%      �%       z 1%��%      �%       ���%      �%       Z�%      �%       z 1%��%      �%       Z�%      &       ��&      W&       Z                      �%      �%       _�%      �%       0��%      �%       _�%      &       0�&      W&       _                       &      #&       x ��#&      )&       { ��)&      -&       ~ ��-&      -&       y���                      �      �       U�             S             �U�                     �      �       U�             S             �U�                   �      �       u���      �       s��                  �      �       V                            %       U%      P       PP      X       �U�                           %       U%      P       PP      X       �U�                  %      P       U                 %      P       U                   %      P       p��P      Q       �U#��                                        (      -(       U-(      2(       V2(      A(       �U�A(      �-       V�-      �.       ���.      �1       �U��1      �1       ���1      2       �U�2      2       ��2      �4       �U��4      +5       V+5      R5       �U�                                        (      %(       T%(      2(       S2(      A(       �T�A(      �-       S�-      �4       �T��4      �4       S�4      5       ��~5      
5       �T�
5      5       ��~5      5       �T�5      +5       ��~+5      R5       �T�                              (      -(       Q-(      2(       \2(      A(       �Q�A(      �)       \�)      �+       �Q��+      
,       \
,      R5       �Q�                    (      -(       R-(      R5       �R�                    (      -(       X-(      R5       �X�                                        #(      %(       T%(      2(       S2(      A(       �T�A(      �-       S�-      �4       �T��4      �4       S�4      5       ��~5      
5       �T�
5      5       ��~5      5       �T�5      +5       ��~+5      R5       �T�                 ,      
,       8�                  )       )       Q,      
,       0�                 �(      )       �D  �+      ,       �D                     �(      �(       s��(      )       ]�+      ,       ]                 �(      )       V�+      ,       V                      �(      �(       q 
����(      	)       R	)      )       q 
����+      ,       q 
���                   �(      )       0�)      )       q 
����+      ,       0�                   �.      �1       s���1      2       s��                   �.      
/       0�
/      "/       P                 @1      K1       0�                 1      �1       V                     61      T1       QT1      r1       q`�r1      �1       Q                      @1      X1       UX1      r1       uX�r1      �1       U                 1      "1       s�#8                     �0      �0       0��0      �0       Q2      2       0�                        �0      �0       Q�0      �0       s�2      	2       Q	2      2       s�                    �0      1       P2      2       P                    #(      -(       U-(      2(       VA(      w(       V                    #(      %(       t��%(      2(       s��A(      w(       s��                       .(      2(       PA(      [(       P\(      f(       Pw(      w(       0�                w(      �(       s��                w(      �(       1�                    K)      �+       }  $0.�
,      ',       }  $0.�                  K)      O)       s�                    K)      �+       V
,      ',       V                    K)      �+       s��
,      ',       s��                  l)      �)       q 
���                    �*      b+       u ��
,      ,       u ��                    �)      �)       T�)      �)       s�                        �)      �)       | 
����)      �)       P�)      �+       | 
���
,      ',       | 
���                                     *      )*       Q)*      D*       q�D*      `*       q�`*      |*       q	�|*      �*       q��*      �*       P�*      �*       Y�*      +       P+      "+       p�"+      H+       PH+      S+       p�S+      w+       Pw+      y+       r��+      �+       P�+      �+       p��+      �+       p��+      �+       p��+      �+       Q
,      ,       P                    *      �+       T
,      ",       T                       �*      �*       0��*      �*       1��*      �*       R�*      �*       r��*      �*       {��*      �*       R                d+      �+       T                d+      �+       ��G                  d+      �+       0�                d+      �+       T                d+      �+       ��G                  d+      �+       0�                  d+      q+       Pq+      y+       Ry+      �+       P�+      �+       p��+      �+       R�+      �+       P                 t+      �+       Q                   �+      �+       p����+      �+       r���                   �+      �+       p ����+      �+       r~���                    U,      �-       \�4      �4       \                        =,      },       P},      �.       ���1      �1       ��2      R5       ��                                =,      �-       V�-      �.       ���.      �.       �U��1      �1       ��2      2       ��2      �4       �U��4      +5       V+5      R5       �U�                                      =,      �-       s���-      �.       �T#���1      �1       �T#��2      �4       �T#���4      �4       s���4      5       ��~#��5      
5       �T#��
5      5       ��~#��5      5       �T#��5      +5       ��~#��+5      R5       �T#��                        t,      },       R},      �.       w �1      �1       w 2      R5       w                           v-      �-       q ���-      �.      	 ������1      �1      	 �����2      �3      	 ������4      +5      	 �����                            �-      �-       q x !������-      .      	 q �����.      .       V.      .       v | �.      �.       V�1      �1       V�4      �4      	 q �����                                                �,      �,       P�,      �,       p��,      �,       p��,      -       p�-      -       p�-      8-       p
�8-      R-       p�R-      l-       p�l-      �-       ]�-      �-       p��-      �-       ]�-      .       P2      (2       ^(2      �2       ]�2      �2      
 q 1$~ "#��2      �2      
 q 1$~ "#��2      �2      
 q 1$~ "#��2      �2       }��2      �2       }��2      �2       }��2      3       }�3      �3       \�3      �3       p��3      4       P4      %4       T%4      c4       \c4      �4       P�4      �4       ]�4      �4       p�&5      +5       ]+5      25       T25      E5       \E5      I5       PI5      R5       T                                 �,      .       Z.      �.       ��~�1      �1       ��~2      2       ��~�4      �4       Z�4      5       S
5      5       S5      &5       S&5      +5       Z                          �-      .       P.      .       U.      ".       S".      /.       P/.      a.       p�a.      �.       U�1      �1       U�1      �1       u
��1      �1       u��1      �1       u��1      �1       u��1      �1       U                      .      ".       Sa.      �.       S�1      �1       S                              .      .       Q.      ".       | 
���A.      �.       Q�.      �.       | 
����1      �1       Q�1      �1       | 
����1      �1       Q                      .      .       r 
���l.      �.       r 
����1      �1       r 
���                      �2      �2       Q�2      �2       q��2      �2       Q                    82      j2       [j2      u3       ��                    �3      �4       R+5      R5       R                    =3      �4       ]+5      R5       ]                   F3      I3       4�I3      �3       P                     �3      =4       QF4      �4       Q+5      R5       Q                 �4      5      
 �tH     �
5      &5      
 �tH     �                         �4      �4       s���4      5       ��~#��5      5       �T#��
5      5       ��~#��5      5       �T#��5      &5       ��~#��                        �4      �4       Z�4      5       S
5      5       S5      &5       S&5      &5       Z                 �4      5       �VJ  
5      &5       �VJ                     �4      �4       0��4      5       P
5      &5       0�                       �4      �4       ]�4      �4       P�4      �4       ]�4      �4       }��4      �4       U�4      �4       ]�4      �4       U5      &5       ]                     �4      5       ^
5      5       ^5      &5       ^                      �4      �4       Q�4      �4       Q�4      �4       u���                     �4      �4       } ����4      �4       u~����4      �4       u~���                      �4      �4      
 �tH     ��4      �4       P�4      �4      
 �tH     �                            �
      �
       U�
      c       Vc      h       �U�h      �       V�      �       �U��      �       V                      �
      �
       T�
      b       S�      �       S�      �       Q                            �
      �
       Q�
      g       ]g      h       �Q�h      �       ]�      �       �Q��      �       ]                            �
      �
       R�
      e       \e      h       �R�h      �       \�      �       �R��      �       \                             �
      8       0�8      <       P<      M       RY      h       Rh      v       0�v      �       R�      �       0�                       �
             0�             P!      4       P�      �       0�                   %      h       1��      �       q  $0.��                              `      �       U�      �       S�      �       s��      �       s��      I	       RI	      �	       s��	      �	       R�	      
       s�
      
       R
      -
       s�                            `      l       Tl      �	       \�	      �	       �T��	      �	       \�	      �	       �T��	      -
       \                            `      �       Q�      �	       V�	      �	       �Q��	      �	       V�	      �	       �Q��	      -
       V                             `      �       0��      �       P�      �	       T�	      �	       T�	      �	       0��	      �	       T 
      
       0�
      -
       T                 �	      �	       8�                     �      �	       ]�	      �	       ]�	      -
       ]                                E	      L	       u �8$y �!
���L	      g	       s��8$y �!
���g	      j	       q ��8$q��!
���j	      m	       r 8$q��!
���m	      }	       q ��8$q��!
���}	      �	      @ t��1z ����s "#��8$t��1z ����s "#��!
���
      
       u ��
      
       q ���
      #
       R#
      (
       t��1z ����s "#���                                 E	      I	       s��8$s��!
���I	      R	       r 8$s��!
���R	      g	       s��8$s��!
���g	      y	       q��8$q��!
���y	      }	       u 8$q��!
���}	      �	      & u 8$t��1z ����s "#��!
����	      �	      @ t��1z ����s "#��8$t��1z ����s "#��!
���
      
       y ��
       
       q��� 
      %
       Q%
      (
       t��1z ����s "#���                      E	      E	       RE	      E	       r�E	      I	       r�I	      g	       s�g	      g	       t��1t�����s "#�g	      g	       t��1t�����s "#�g	      �	       t��1t�����s "#�
      
       R
      
       r�
      
       r�
      
       t��1t�����r "�
      
       t��1t�����r "#�
      
       t��1t�����r "#�
      -
       t��1t�����s "#�                                          U&      >       U>      Z       XZ      o       u�o      �       s��      �      
 q 1$s "#��      �      
 q 1$s "#��      �      
 q 1$s "#�                                      T      &       �T�&      {       T{      �       �T�                                      Q      &       �Q�&      v       Qv      �       V                              A      G       r ��G      K       | ��K      R       u ���R      �       ]�      �       q  } "��      �       } q ��      �       q  } "�                      K      O       | ��O      R       ]R      �       | ��                     K      W       RW      o      
 u ��4%�o            
 s ��4%�                                           0�&      �       0��      �       P�      �       U�      �      
 q 2$u "#��      �       q 2$u "��      �      
 q 2$u "#�                                  q &      v       q v             v                           0
      I
       UI
      R
       �U�R
      l
       Ul
      �
       \�
      �
       �U�                        0
      I
       TI
      R
       �T�R
      o
       To
      �
       �T�                          0
      I
       QI
      R
       �Q�R
      c
       Qc
      �
       S�
      �
       �Q�                     G
      I
       q R
      c
       q c
      s
       s                            G
      I
       t u �I
      R
       �T�U�R
      l
       t u �l
      o
       t | �o
      �
       �T| ��
      �
       �T�U�                                          �             U             u�             u�      �       S�      �       ^�      �       X�      �       x��             S      :       X:      o       So      �       ^�      �       X�      �       x��      �       S�      �       X�      �       S4      �       S                          �      8       T8             _      4       �T�4      F       TF      �       _                        �             Q             \      4       �Q�4      �       \                    �      8       P4      Y       P                               w      �       q ����(x "��      �      	 p (x "��      �       q ����(x "��      6       P6      N       pX�N      �       P�      �       pX��      �       P                          p       v ��4      �       v ��                  �      �       0�                                 ]4      �       ]                   8      Q       8�Q      {       P                        %       8�                    M      Y       ZY      �       ��                                      U      F       _F      G       �U�G      2       _                                      T      D       ^D      G       �T�G      2       ^                                                               *       Q*      2       ��~2      G       �Q�G      �       ��~�      e       �Q�e      }       ��~}      �       �Q��      �       ��~�      �       �Q��      g       ��~g      l       �Q�l             ��~             �Q�      x       ��~x      �       �Q��      3       ��~3      �       �Q��      �       ��~�             �Q�      2       ��~                           *       R*      2       �R�                                             *       X*      2       ]2      G       �X�G      �       ]�      e       �X�e      }       ]}      �       �X��      _       ]_      *       �X�*      3       ]3      2       �X�                                                      .      2       PG      Z       PZ      ^       \^      f       Pf      �       \e      }       \�      �       ���      �       \�      �       S�             0�      %       P�      �       0��      #       \      �       \              P       *       0�*      3       \�      �       \             \             ��*      2       S                                       f      �       P�      �       ~� e      }       P�      �       P�      �       ~� �             P      �       ~� 6      l       P
             P      #       ~� x      �       ~� *      3       ~�                       n      �       V�      �       V*      2       V                 �      �       0�                                    x      }       T�      �       T�      �       �      6       ��~l      �       ��~�      
       ��~      x       ��~*      3       �      �       ��~      2       ��~                     �      �       ���~���      �       P�      �       ���~��                     e      }       (�      �       (*      3       (                     e      }       (#��      �       (#�*      3       (#�                  O      o       0��      �       0�                              o       Vo      �      	 | 0$0&��              V       %      	 | 0$0&�                          2      V       RV      o       z v �o      �       z | 0$0&��             R       %       z | 0$0&�                              �             Y-      o       Qo      �       y } "��      �      	 y } " ��      �       Q�             y } "�       *      	 y } " �                      o      w       Pw      �       pp��      �       P                   �      �       Q�      �      
 q v "#���                  �      �       q ?&��      �       V                  o      w       p w      �       pp                   {      �       Q�      �      
 q v "#���                  {      �       q ?&��      �       V                  �             P                              x      }       V�      6       Vl      �       V�      
       V      x       V*      3       V�      �       V             V                                               x      }       P�      �       P�             p�      A       ~� #�A      �       S�      �       P�             Y      (       P(      .       Y.      J       PJ      q       Tq      �       S�      �       P�      �       P�             U      6       Pl      �       P�      �       T�      �       S�      �       T�      
       S      -       P-      H       YH      ]       P]      x       Y*      3       S�      �       S             S                              x      }       _�      6       _l      �       _�      
       _      x       _*      3       _�      �       _             _                     x      }       (�      �       (*      3       (                     x      }       (�      �       (*      3       (                             �      �       Q�      �       q`��      6       Ql      �       Q�      
       Q      x       Q             Q                        �      �       q ���             p ���      �      
 ~� ���*      3      
 ~� ���                  �      �       0�             0�                                  �      �       [�      �       ��~�      6      	 ��~���l      �      	 ��~����      
      	 ��~���      x      	 ��~���*      3       [�      �       ��~            	 ��~���                            A      6       ��~l      �       ��~�      
       ��~      x       ��~*      3       ��~�      �       ��~             ��~                                �              0�       M       UM      �       q�      �       qp�      6       0�l      �       U�      
       q      C       0�C      x       U                                    �      +       0�+      A       TA      �       q�      �       qt�      6       0�l      w       0�w      �       T�      �       q�      
       q      s       0�s      x       T                   m      �       ]�      �       ]                 �      A       V                 �      A       �gZ                   �      A       0�                 �      A       V                 �      A       �gZ                   �      A       0�                            �      �       p��      �       S�             p�             p�             S             ~� #�      -       S-      -       s�-      0       s�0      3       p s "#�3      <       s�<      A       S                    �      <       Q<      ?       q�?      A       Q                                      p���             s p "#���      0       s���0      3       p s "#���3      A       s���                                      p���      -       ~� #���-      0       s ���0      3       p s "���3      <       s ���<      A       ~� #���                          �      y       R�      6       Rl      �       R�      �       R      x       R                             �      e       V�      �       V6      l       V
             Vx      �       V3      �       V�             V                                                             �      �       P�      �       p��      	       S	             Y      D       SD      J       PJ      Y       SY      e       P�      �       p��      �       S�      �       P6      M       p�M      l       S
      X       SX      [       q s "�[      x       Sx      {       q s "�{      �       S�      �       P�      U       \U      l       Pl      �       \�      �       Y�      �       \�      �       Y�      �       \�      ^       \^      �       Y�      �       \�      �       Y�      �       \�      �       Y�             \             Yx      �       S3      �       \�             \      
       Q
             \                             �      e       _�      �       _6      l       _
             _x      �       _3      �       _�             _                        �      �       (�      �       (6      l       (
      #       (x      �       (                          �      e       } ���      �       } ��6      l       } ��
      '       } ��x      �       } ��                              �      �       0��      �       [�      �       0�6      R       0�R      l       [
      #       0�x      �       [�      �       ��~                              �      �       0��      �       P�      e       ��~�      �       0��      �       S�      �       ��~6      l       0�
      #       0�x      �       ��~                     �      �       0�&      6       q�6      J       Q�      �       0�                           �      �       p ���      �       { ���      �       ~� #����      �      	 { ��~�"�
      #       0�x      �      	 { ��~�"��      �       ��~���~�"�                     �      �       0�D      G       s ���G      J       T#      #       0��      �       0�                      �      �       0��             R      e       R#      #       0��      �       0�                  -      �       V      
       V                  -      �       ��\        
       ��\                    -      �       0�      
       0�                  -      �       V      
       V                  -      �       ��\        
       ��\                    -      �       0�      
       0�                         -      <       S<      T       s�T      T       s�T      e       Qe      u       Su      u       s�u      x       s�x      {       q s "#�{      �       s��      �       S      
       q�                     ?      �       P�      �       p��      �       P      
       P                           T      X       s���X      [       q s "#���[      u       s���u      x       s���x      {       q s "#���{      �       s����      �       s���                           T      X       s���X      [       q s "#���[      u       s���u      x       s ���x      {       q s "���{      �       s ����      �       s���                       �             _3      �       _�             _
             _                       �      l       qp�t             qp�             Q8      =       ���P             qp�                              �      �       x ���      �       p ���      �       |���.      R       |���l      �       |����      �       |���3      =       |���                              �      �       T�      �       p ��.      8       T8      =       p ��=      �       T�      �       p ��3      =       T                             �      �       0��             T.      8       0�8      =       
+�=      �       0�P             T3      =       0�                         �      _       U_      l       3�t             U8      =       3�j      l       0��      �       0�P             U                              �      >       R>      L       PL      l       Rt      �       R�             P             R8      =       0�P             R                            �      �       z ���      �       p ���      �       y����      �       z ���      �       p ���      �       y���                      �      �       | �8$8&��      �       y�8$8&�             | �8$8&�             y�8$8&�                 �      �       _                      �      B       ���B      F       QF      G       ����      �       ���                  �      G       _�      �       _                 �      �       (                   G      G       P�      �       P                     =      �       _�             _
             _                     =      �       ����             ���
             ���                     =      �       ����             ���
             ���                     =      �       ����             ���
             ���                    =      ]       (�      �       (�      �       (                     =      ]       (#`��      �       (#`��             (#`�                     �      �       0��      �       P�      �       8�
      
       P                  r      �       Q                r      �       P                    �      �       P�      �       ��~                    �      �       U�      �       �U�                    �      �       T�      �       �T�                        �      �       U�      '       S'      1       �U�1      E       S                      �      �       T�      1       �T�1      E       T                      �      �       Q�      1       �Q�1      E       Q                        �      �       R�      .       ].      1       �R�1      E       R                        �      �       X�      ,       \,      1       �X�1      E       X                       �      �       U�      '       S'      1       �U�1      E       S                       �      �       u���      '       s��'      1       �U#��1      E       s��                       �      	       @<$�	             P      0       ^1      E       @<$�                     �             @<$�      )       P1      E       @<$�                    �      *       V1      E       V                      �      �       T�      �       T�      �       �T1�                 �      �       U                 �      �       6��      �       0�                 �      �       u��                             �       A       0�A      E       PE      J       p�J      Y       PY      \       0�\      j       Qj      �       0��      �       P�      �       Q�      �       P                        �       9       Y9      U       0�U      {       Y{      �       0��      �       Y                         �       �        0��       J       PJ      Y       p�Y      �       P�      �       P                           �       �        u�              R      9       XY      \       Rj      p       Rp      {       X                                           Q      %       X%      )       R)      4       Q4      9       XY      \       Xj      p       X                                             q ����4$z "�      %       x ����4$z "�%      )       r ����4$z "�)      4       q ����4$z "�4      9       x ����4$z "�A      G       p ����4$u "�G      N      	 q 4$u "�N      Y       p����4$u "�Y      \       x ����4$z "�j      p       x ����4$z "�                   p       v        0�v       �        X                          s       �        Q�       �        R�       �        Q�       �        Q�       �        R                           �       �        p ����4$y "��       �        r ����4$y "��       �        q ����4$y "��       �        p ����4$y "��       �        r ����4$y "��       �        r ����4$y "��       �        r ����4$y "�                              �       �        P�       �        R�       �        Q�       �        P�       �        R�       �        R�       �        R                                    T       V        �T�                           P        0�P       V        8�                                   P       V        u                         3        1�                 P      �       U                 P      �       u� �                      m      �       R�      �       {��      �       R                     m      �       0��      �       Q�      �       Q                    �      �       X�      �       X                    �      �       Y�      �       Y                                          U      :       S:      <       �U�<      \       S\      ^       �U�^      t       S                                  T      t       �T�                                  Q      t       �Q�                                          R      ;       V;      <       �R�<      ]       V]      ^       �R�^      t       V                                        U      :       S:      <       �U�<      \       S\      ^       �U�^      t       S                                        u��      :       s��:      <       �U#��<      \       s��\      ^       �U#��^      t       s��                      *      3       �T�<      ^       �T�m      t       �T�                      *      3       �Q�<      ^       �Q�m      t       �Q�                        *      3       V<      ]       V]      ^       �R�m      t       V                        *      3       S<      \       S\      ^       �U�m      t       S                       �      �       U�      �       S�      �       S�      �       U                       �      �       u� ��      �       s� ��      �       s� ��      �       u� �                  �      �       P                 �      �       s� �0$0&�                        `&      �&       U�&      �'       S�'      �'       �U��'      (       U                       `&      �&       U�&      �'       S�'      �'       �U��'      (       U                      r&      �&       U�&      �'       S�'      �'       �U�                  �&      �'       ]                 �&      �'       V                   �&      �&       u���&      �'       s��                    �'      �'       T�'      �'       0��'      �'       \�'      �'       T                  �'      �'       \                    �      �       U�      �       �U�                        �      �       T�             _             �T�      �       _                       �      �       T�             _             �T�      �       _                       �      �       t���             ��             �T#��      �       ��                       �      �       t���             ��             �T#��      �       ��                       �      �       t���             ��             �T#��      �       ��                      �      �       ]�      �       ]             ]                                            �      �       P�      �       P�      �       P�      �       P�             P!      0       PM      c       Pt      �       P�      �       P�      �       P�      �       P�      �       P�      �       P�      �       P                     �      �       ^�      �       ^             ^                                  �      +       ^5      g       ^)             \      �       ^�      �       QU      X       QX      �       ���      �       ^�      �       Q                      �      �       S�      �       S      �       S                        �      �       ��      �       ���      �       P�      �       ��                           �      �       0��      �       ���      �       0�             0�             ��0      �       ��                           �      �       0��      �       ���      �       0�             0�      +       ��0      �       ��                         5       0�5             V                              �      �       P�      w       ��w      �       Y�      �       ^�      �       P�      �       R�      �       P                           �      	 z �()��      0      	 ���()��      �      	 z �()�                            `      o       Uo      �       V�             �U�      4	       V4	      =	       �U�=	      I
       V                            `      �       T�      �       S�      �       U�      (
       �T�(
      4
       S4
      I
       �T�                           `      �       T�      �       S�      �       U�      (
       �T�(
      4
       S4
      I
       �T�                            �       P�      �       w (
      4
       w                                   �             [�      �       [�      �       z �      �       {�X	      p	       [p	      �	       ��(
      ,
       [,
      /
       s /
      4
       {�4
      I
       [                        �      �       P�      �       _�      �       ��(
      4
       _                              �      �       0��      �       ��      �       ���      9       P9      v       ��v      (
       ��(
      4
       0�4
      I
       ��                                           �      �       0��      �       ]      t       ]t      �       Q�      �       ]�      �       R�      �       ]�      �       P�      i       ]i      �       Q�      8	       ]=	      (
       ](
      4
       0�4
      I
       ]                              �      �       [|      �       [�      �       {��      �       [�      �       {��      9       [9      `       ��v      �       [
       
       [                                         �      �       0��      0       ^0      3       P3      �       ^      	       ^=	      S	       ^S	      X	       p�X	      �	       ^�	      �	       | 1&��	      �	       \�	       
       ^(
      4
       0�4
      I
       ^                               �      �       0��      �       ���      �       ���      `       ��=	      �	       ���	      
       \
       
       ��(
      4
       0�4
      I
       ��                               �      �       0��      �       _�      �       0�      .	       _.	      =	       0�=	      �	       _�	      �	       P�	      (
       _(
      4
       0�4
      I
       _                                 �      �       0��      �       ���      �       ���      �       0��      `       ��	      "	       ��=	      �	       ���	      
       1�
       
       ��(
      4
       0�4
      <
       ��<
      I
       1�                                 �      �       0��      �       S�      �       S      6       1�6      �       2��      �       0��      �       1��      	       1�=	       
       S(
      4
       0�4
      I
       S                      �      �       \      	       \
       
       \                          3       P3      e       ^                                 0��      �       0�                      �      �       Q�      �       q}��      	       Q                     �      �       v�#��      �       T�      �       tp��      	       v�#�                                                     "       U"      t       Vt      �       �U��             V      �       ���      �       V�             �U�      N       VN      W       �U�W      j       Vj      s       �U�s      �       V�      c       ��c      u       �U�u      �       ��                                           $       T$      �       ^�      �       �T��             ^             �T�      T       ^T      W       �T�W      p       ^p      s       ����s      �       ^                                          $       T$      �       ^�      �       �T��             ^             �T�      T       ^T      W       �T�W      p       ^p      s       ����s      �       ^                                                 (      ]       _�             _!      ^       V^      ~       ]~      �       V�             _W      r       _s      �       _�      �       V�      �       ]�      �       V�      =       ]=      [       Vc      u       _u      �       V�      �       ]�      �       _�      �       ]                                    t       S�      �       S�      �       w �      �       S      M       SW      i       Ss      �       S                                 t       ]�      �       ]�             ]      R       ]W      n       ]s      �       ]                               �             v��      �       ��#��W      j       v��j      s       �U#��s      �       v���      c       ��#��c      u       �U#��u      �       ��#��                     �      �       P�      �       \s      �       
 �                                  �      �       0��      �       S�      �       T�      �       s��      �       S�      !       0�!      �       w �      0       w 8      c       w u      �       w                        �      �       ~��W      p       ~��p      s       ��s      �       ~��                            �      �       R�      �       w W      h       w h      s       ��s      �       R�      �       w                    �      �       0�s      s       0�s      �       1�                 �      �      
 �1H     �                        N      k       \�      �       w �      �       R�      �       \                    
             P      =       V                            P
      b
       Ub
      �
       S�
      �
       �U��
      �
       S�
      �
       �U��
      o       S                          P
      [
       T[
      �
       V�
      �
       �T��
      �
       V�
      o       �T�                          T
      [
       T[
      �
       V�
      �
       �T��
      �
       V�
      o       �T�                            _
      b
       u��b
      �
       s���
      �
       �U#���
      �
       s���
      �
       �U#���
      o       s��                           _
      b
       u��b
      �
       s���
      �
       �U#���
      �
       s���
      �
       �U#���
      o       s��                    v
      �
       q ��
             q �                    l
      ~
       P�
      �
       P                                  U             �U�                                 U             �U�                              ,       U,      K       SK      L       �U�L      a       U                             ,       U,      K       SK      L       �U�L      a       U                            9       PL      W       PW      a       u                           9       PL      W       PW      a       u                           :       0�:      L       PL      a       0�                      @      Q       UQ      �       S�      �       �U�                      @      U       TU      �       \�      �       �T�                     @      Q       UQ      �       S�      �       �U�                  M      �       V                  e      �       P                      �      �       U�      �       S�      �       �U�                      �      �       T�      �       \�      �       �T�                     �      �       U�      �       S�      �       �U�                  �      �       V                  �      �       P                      p      �       U�      �       S�      �       �U�                     p      �       U�      �       S�      �       �U�                 p      q       u                  p      q       u                       �      �       P�      �       V�      �       P                          �      �       U�      �       S�      �       �U��      �       S�      �       �U�                         �      �       U�      �       S�      �       �U��      �       S�      �       �U�                    �      �       P�      �       P                        �      �       U�             S      �       �U��      �       U                       �      �       U�             S      �       �U��      �       U                     �      �       u���             s��      �       �U#��                     �      �       u���             s��      �       �U#��                  �      �       V                          2       U2      %       �U�                                                              B       TB      �       S�      K       �T�K      �       S�      e       �T�e      �       S�      �       ��z�      �       �T��      �       S�              �T�       �        ��z�       !       �T�!      "       ��z"      �#       �T��#      �#       ��z�#      X$       �T�X$      �$       S�$      �$       ��z�$      �$       �T��$      %       ��z                          K       QK      %       ��y                          $       R$      O       ��z                        $       X$      T       ��y                                                             B       TB      �       S�      K       �T�K      �       S�      e       �T�e      �       S�      �       ��z�      �       �T��      �       S�              �T�       �        ��z�       !       �T�!      "       ��z"      �#       �T��#      �#       ��z�#      X$       �T�X$      �$       S�$      �$       ��z�$      �$       �T��$      %       ��z                                    E      6       ^      �       ^�      �       P�      �       P�             0�      &       \&      S       0�S      e       ^�      �       P�              0�
$      !$       ^                   c      q       Pq      %       ��y                                         �      �       P�      �       ]K      �       ]e      s       Ps      �       ]�      �       ��z�      �       ]       �        ��z!      "       ��z�#      �#       ��zX$      �$       ]�$      �$       ��z�$      %       ��z                                                             B       TB      �       S�      K       �T�K      �       S�      e       �T�e      �       S�      �       ��z�      �       �T��      �       S�              �T�       �        ��z�       !       �T�!      "       ��z"      �#       �T��#      �#       ��z�#      X$       �T�X$      �$       S�$      �$       ��z�$      �$       �T��$      %       ��z                                                             B       t��B      �       s���      K       �T#��K      �       s���      e       �T#��e      �       s���      �       ��z#���      �       �T#���      �       s���              �T#��       �        ��z#���       !       �T#��!      "       ��z#��"      �#       �T#���#      �#       ��z#���#      X$       �T#��X$      �$       s���$      �$       ��z#���$      �$       �T#���$      %       ��z#��                                                             B       t��B      �       s���      K       �T#��K      �       s���      e       �T#��e      �       s���      �       ��z#���      �       �T#���      �       s���              �T#��       �        ��z#���       !       �T#��!      "       ��z#��"      �#       �T#���#      �#       ��z#���#      X$       �T#��X$      �$       s���$      �$       ��z#���$      �$       �T#���$      %       ��z#��                 =      X       U                    c      q       Pq      %       ��y                          �      (       T(      ,       t�,      .       TS      S       TS      `       t�`      e       T
$      !$       T                     �      .       QS      e       Q
$      !$       Q                    �      S       ]�              ]                       �      
       0�
             U&      Q       0�Q      S       U�      �       0��              U               0�               U                                                   �      �       S�      E       �T�K      �       S�             �T�s      �       S�      �       ��z�      �       S       �        ��z�       !       �T�!      "       ��z"      �#       �T��#      �#       ��z�#      
$       �T�!$      X$       �T�X$      �$       S�$      �$       ��z�$      �$       �T��$      %       ��z                             �      6       VK      e       Vs      �!       V�!      �!       U�!      �$       V�$      �$       U�$      %       V                                                     �      �       s���      6       �T#��K      �       s���      e       �T#��s      �       s���      �       ��z#���      �       �T#���      �       s���              �T#��       �        ��z#���       !       �T#��!      "       ��z#��"      �#       �T#���#      �#       ��z#���#      X$       �T#��X$      �$       s���$      �$       ��z#���$      �$       �T#���$      %       ��z#��                          �      �       ^K      �       ^s      �       ^�      �       ^X$      �$       ^                                     �      �       ]K      �       ]s      �       ]�      �       ��z�      �       ]       �        ��z!      "       ��z�#      �#       ��zX$      �$       ]�$      �$       ��z�$      %       ��z                                                     �      �       S�      6       �T�K      �       S�      e       �T�s      �       S�      �       ��z�      �       �T��      �       S�              �T�       �        ��z�       !       �T�!      "       ��z"      �#       �T��#      �#       ��z�#      X$       �T�X$      �$       S�$      �$       ��z�$      �$       �T��$      %       ��z                  �      �       U�      �       V                   �      @       V�             V                   �      @       V�             V                   (      @       V�             V                   (      6       ��{�      �       ��{                                   k      �       ]s      �       ]�      �       ��z�      �       ]       �        ��z!      "       ��z�#      �#       ��zX$      �$       ]�$      �$       ��z�$      %       ��z                       k      |       R|      �       ^s      v       ^�      �       ^X$      �$       ^                     k      �       _s      v       _�      �       _X$      �$       _                     k      �       Vs      v       V�      �       VX$      �$       V                          [       \X$      �$       \                 v      �       ��|                 v      �       ��|                                v      �       V       �        V!      �!       V�!      �!       U�!      "       V�#      �#       V�$      �$       V�$      �$       U�$      %       V                              v      �       S�      �       ��z       �        ��z�       �        �T�!      "       ��z�#      �#       ��z�$      �$       ��z�$      %       ��z                               v      �       V       �!       V�!      �!       U�!      
$       V!$      X$       V�$      �$       V�$      �$       U�$      %       V                 �      �      
 ��|��|"�                	       v      �       D�       
$       D�!$      X$       D��$      %       D�                                     �      �       ]�             ^3      �       ]       7        ]7       E        ^s       �        P!      C!       ^C!      "       ��z�#      �#       ��z�$      �$       ��z�$      %       ��z                                       _!      "       _�#      �#       _�$      �$       _�$      %       _                        E!      "       S�#      �#       S�$      �$       S�$      %       S                                     E!      K!       s  $ &0�wH     "�K!      [!       s $ &0�wH     "�[!      �!       s  $ &0�wH     "��!      �!       r 0�wH     "��!      "       s  $ &0�wH     "��#      �#       s $ &0�wH     "��$      �$       r 0�wH     "��$      �$       s  $ &0�wH     "��$      �$       r 0�wH     "��$      �$       s  $ &0�wH     "��$      %       r 0�wH     "�                           E!      K!       s  $ &0�wH     "K!      [!       s $ &0�wH     "[!      "       s  $ &0�wH     "�#      �#       s $ &0�wH     "�$      �$       s  $ &0�wH     "�$      %       s  $ &0�wH     "                            �!      �!       r 0�wH     "��!       "       s  $ &0�wH     "��$      �$       r 0�wH     "��$      �$       s  $ &0�wH     "��$      �$       r 0�wH     "��$      �$       s  $ &0�wH     "��$      %       r 0�wH     "�                          �!      �!       V�!      �!       U�!       "       V�$      �$       V�$      �$       U�$      %       V                    �!       "       ��z�$      �$       ��z�$      %       ��z                      "       "       P�$      �$       P�$      �$       P                         �!      �!       ��z��!      �!       Q�!       "       ��z��$      �$       Q�$      �$       ��z�                     �!      "       0��$      �$       0��$      %       0�                  7       �        ^                                �"      #       0�#      2#       ��z2#      w#       _w#      ~#       p�~#      �#       ��z�1��#      
$       ��z�1�!$      2$       ��z�$      �$       0�                        b#      ~#       0�~#      �#       ��#      �#       _�#      $       �                        �"      �#       0��#      
$       0�!$      X$       0��$      �$       0�                          �"      #       0�#      �#       ��z�#      
$       ��z!$      2$       ��z�$      �$       0�                      ~#      �#       S�#      �#       S�#      
$       S                        #      2#       \U#      �#       \�#      
$       \!$      2$       \                    p      u       Uu      z       �U�                    p      y       Ty      z       �T�                            �      �       U�      A       ^A      D       �U�D      V       ^V      Y       �U�Y      \       U                            �      �       T�      ?       ]?      D       �T�D      T       ]T      Y       �T�Y      \       T                   �      �       0�Y      \       0�                               T                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       Q�      �       P�      �       �Q�                      �      �       R�      �       Q�      �       �R�                 �      �       U                      �      �       U�      �       V�      �       �U�                      �      �       T�      �       ]�      �       �T�                      �      �       Q�      �       �Q��      �       _                      �      �       R�      �       \�      �       �R�                  �      �       P                     �      �       U�      �       V�      �       �U�                     �      �       T�      �       ]�      �       �T�                 �      �       t                   �      �       ^                 �      �       S                 �      �       ]                 �      �       \                 �      �       V                      �      �       U�             S             �U�                     �      �       U�             S             �U�                 �      �       u                  �      �       u                   �      �       P                  �             S                    0      5       U5      :       �U�                    0      9       T9      :       �T�                 `       �        u�                          P      ;       U;      �       V�      �       �U��      -       U-      �       V                    P      _       T_      �       �T�                        P      �       Q�      �       Q�      �       Q�      -       Q                          P      v       Rv      }       S}      �       �R��      -       R-      �       �R�                            _      �       T�      1       �T�      �       T�      �       �T�             T      -       �T                      w      �       \�      �       \      �       \                 �      �       3�                          �      �       P�      �       p��             p��      �       s } "��      �       p��      �       p�-      e       s } "�e      �       Q                    �      �       4�      -       6�                         g      ;       u��;      �       v���      �       �U#���      -       u��-      �       v��                          �      �       P      �       ]�      �       ](      -       P-      �       ]                      �      v       y 
��
 )��      �       y 
��
 )�      -       y 
��
 )�                    �      �       U-      A       U                      �      �       ^-      �       ^�      �       ~�                  e      �       X                   q      y       Xy      �       R                  q      �       U                                    U      J       SJ      L       �U�                                  T      L       �T�                               U                        K       v�                        �      �       U�             w              ��}             w                         �      �       T�             _             �T�             _                                                  �      �       Q�             V             �Q�      O       VO      	       �Q�	      d	       Vd	      �
       �Q��
      *       V*      P       �Q�P      ;       V;      K       �Q�K      X       ��}X      d       �Q�d      �       V�      B       ��}B      P       VP      �       ��}�      �       V�             ��}                    �      �       R�             �R�                    �      �       X�             �X�                       �      �       T�             _             �T�             _                                      �             ]      O       ]	      d	       ]�
      *       ]P      ;       ]K      X       ��}d      �       ]�      B       ��}B      P       ]P      �       ��}�      �       ]�             ��}                              �      �       ^�             �QO&�Q'�QO&
���      �	       ^�	      �
       �QO&�Q'�QO&
����
      :       ^:      P       �QO&�Q'�QO&
���P             ^                 �      �       U                       D      �       _t      �       _�	      �
       _:      P       _                       D      �       St      �       S�	      �
       S:      P       S                      �	      �	       Q�	      �
       V:      P       V                   �      �       V�	      �	       V                              ^                                           �      �       Q�             V      O       VO      d       �Q�	      d	       Vd	      �	       �Q��
      *       V*      *       �Q�P      ;       V;      ;       �Q�K      X       ��}X      d       �Q�d      �       V�      B       ��}B      P       VP      �       ��}�      �       V�             ��}                               �             \      d       \	      �	       \�
      �
       \�
      �
       U�
      %       \%      )       U)      *       \P      ;       \K      �       \�             \                                    �             ]      O       ]	      d	       ]�
      *       ]P      ;       ]K      X       ��}d      �       ]�      B       ��}B      P       ]P      �       ��}�      �       ]�             ��}                	                 �             S             ^      O       SO      d       ^	      d	       Sd	      �	       ^�
      �
       S�
      *       ^P      �       S�      ;       ^K      �       ^�             ^                 �
      �
       ��}�
����}�
��" $ &�                        �
      �
       P�
      *       ��}d      �       ��}B      P       ��}�      �       ��}                     �
      *       0�d      q       0�q      �       ��}B      P       ��}�      �       ��}                    �
      *       0�d      v       0�v      �       ��}                         �
      �
       P�
             S       )       P)      *       Sd      m       S                    �
             Pd      u       P                          K      X       ��}�      �       P�      B       ��}P      �       ��}�             ��}                        �      �       P�      B       ��}P      d       ��}�             ��}                        R      �       S�      B       sp�P      Y       sp��             sp�                                  �      �       0��      4       SK      X       ��}�      �       S�      �       S�      �       0��      B       ��}P      _       ��}d      �       ��}�             ��}                      �      B       ]P      d       ]�             ]                      �      B       VP      Y       V�             V                 �             _                 �             _                 �             _                  �             S                       0       M        0�M       R        PR       \        0�\       _        P                       0       J        0�J       O        QO       R        RR       \        0�\       _        R                          8       E        QE       M        PM       O        p�R       \        P\       ^        q u��                            #        T#       .        T                         -        0�                                  u                     
               P                u #�                      �      �       U�      '       S'      ,       �U�                 �      �       u�                 �      �       u�                  �             V      '       0�                      @      �       U�      �       �U��      �       U                      @      �       T�      �       �T��      �       T                    F      �       X�      �       X                   F      �       x�#��      �       x�#�                   F      �       x� �      �       x�                         s      y       Qy      }       q`�}      �       Q�      �       Q                    �      �       T�      �       �T�                    �      �       U�      �       �U�                                �      �       U�              S              �U�      �       S�      �       q�~��      �       �U��      �       S�      �       �U�                                �      �       T�             V             �T�      �       V�      �       U�      �       �T��      �       V�      �       �T�                      �      �       P             P      !       P                               �      �       u��              s�              �U#�      �       s��      �       q�~��      �       �U#��      �       s��      �       �U#�                   -      i       p 
��
 )��      �       p 
��
 )�                    7      Y       v��      �       ��                      Y      �       V�      �       U�      �       �T�                      Y      �       S�      �       q�~��      �       �U�                  j      �       P                               9       U9      Z       SZ      \       �U�\      a       U                              9       U9      Z       SZ      \       �U�\      a       U                      *      9       U9      Z       SZ      \       �U�                  5      [       V                                                                        0      \       U\      h       Vh      �       �U��      6       V6      �       �U��      �       V�      "       �U�"      �       V�      �       �U��             V             U             V      �       ��~�      �       �U��      �       V�      Q        �U�Q       U        UU       [        V[       �        �U��       �        V�       !       �U�!      (!       V(!      �!       �U��!      �!       ��~�!      �!       �U��!      �!       ��~�!      "       �U�"      "       V                                                            0      S       TS      h       Sh      �       �T��      �       S�      '       ��~'      6       S6      �       �T��      �       S�      "       �T�"      �       S�      �       �T��             ��~      �       �T��      �       S�      �       �T��      �       S�      �        �T��       �        ��~�       !       �T�!      !       S!      "       �T�"      "       S                                        0      \       Q\      h       \h      �       �Q��      �       \�      "       �Q�"      �       \�      �       �Q��      �       \�      !       �Q�!      !       \!      "       �Q�"      "       \                                                           0      S       TS      h       Sh      �       �T��      �       S�      '       ��~'      6       S6      �       �T��      �       S�      "       �T�"      �       S�      �       �T��             ��~      �       �T��      �       S�      �       �T��      �       S�      �        �T��       �        ��~�       !       �T�!      !       S!      "       �T�"      "       S                 h      n       3�                    X      \       P\      "       ��~                  �      �       0�                                 �      �       P�      �       P�             P'      4       Po      z       P�      �       P�      
        P�       �        PB!      T!       P                           @      c       Pc      o       V        Q        V[       �        V�       !       V(!      |!       V                                     @      �       0��             ��~        Q        0�[       t        0�t       �        ��~�       �        0��       �        ��~�       !       0�(!      B!       ��~B!      l!       0�l!      |!       ��~                                  @      �       0��      �       
��        Q        0�[       }        0�}       �        P�       �        X�       !       0�(!      B!       PB!      l!       0�l!      |!       
��                      o      �       P�      �       V�!      �!       V                     �      �       S�      �       Sj      q       S                             �      �       Sj      q       S�      Q        S[       �        S�       !       S(!      |!       S�!      �!       S                    �      b       \j      q       \                        �              P=      L       Pw      �       P�      �       P                      �      b       Vb      �       \�      �       \                         �      (       ](      6       T6      B       ]o      �       V�      �       V                    b      �       P�      �       P                  g      �       T                  �      �       0�                            X      h       S�      �       S"      [       Sh      �       S�      �       S!      !       S"      "       S                              X      \       U\      h       V�      �       V"      [       Vh      �       V�      �       V!      !       V"      "       V                            X      h       s���      �       s��"      [       s��h      �       s���      �       s��!      !       s��"      "       s��                             $      7       P7      �       ]"      [       ]h      �       ]�      �       P!      !       ]"      "       ]                              X      \       P\      h       ��~�      �       ��~"      [       ��~h      �       ��~�      �       ��~!      !       ��~"      "       ��~                                           $      7       0�7      R       _R      [       Q[      v       _"      3       Q3      F       0�F      �       ��~�      �       P�             0�             R      <       P<      A       Rh      �       ��~�      �       0�"      "       0�                      �      Q       Q!      !       Q"      "       Q                    V      w       X�      A       X                       V      �       [�      �       1��      A       [h      �       [                        �      �       [���      �       [�T�U���      �       p �T�U���      �       p �p�U��                                         �      �       S�      '       ��~'      6       S6      P       �T��      �       S�             ��~      �       �T��      �       S�      �       �T�Q       [        �T��       �        ��~!      (!       �T��!      "       �T�                                               �      6       V6      P       �U��      �       V�             V             U             V      �       ��~�      �       VQ       U        UU       [        V�       �        V!      (!       V�!      �!       ��~�!      �!       �U��!      �!       ��~�!      "       �U�                                           �      �       0��      �       P�      '       _'      6       0�6      A       _A      P       0��      �       0��      �       _�      �       P�      �       ]�      �       _Q       [        _�       �        _!      (!       _�!      "       _                               �      6       0��      �       0��      �       0��             P�      �       0�Q       [        0��       �        0�!      (!       0�                                  �      �       R�      �       ^�      '       ��~�      �       ��~�      �       ��~Q       [        ��~�       �        ��~!      (!       ��~�!      "       ��~                              C      /       ��~�      �       P�             ��~�      �       ��~Q       [        ��~�       �        ��~!      (!       ��~                                      �      �       0��      "       S�      �       S�             0�      �       S�      �       0��       �        4p ��       �        T�       �       	 4��~3��!      �!       S�!      �!       S�!      �!       S                                �      P       \�      �       \�      �       \�      �       \Q       [        \�       �        \!      (!       \�!      "       \                                     r       Pr      {       Q{      �       ^�      �       ��~V       [        P!      (!       P�!      "       ��~                                     �      6       0�6      L       ]L      P       0��      �       0��      �       0��      �       P�      �       ]�      �       0�Q       [        0��       �        0�!      (!       0��!      "       ]                  �             Q                    j      �       
 ��      �       
 �                    j      �       Q�      �       Q                    j      �       T�      �       T                   j      �       0��      �       P                   �      j       S�             S�      �       S                       �      j       V�             V�      �       V�      �       U�      �       V                    �      j       \�             \�      �       \                       �      �       0��      j       ^�      �       0��             ^�      �       0�                  �      �       ]                          Z      �       R�      �       P�      �       R�      �       R�      �       P                       x      q       Sq      �       ��~�      �       S�      �       ��~                                             x      �       V�      �       U�      s       Vs      |       U|      �       V�      �       U�      �       V�      �       U�      �       V�      �       V�      �       U�      q       Vq      u       Uu      {       V|!      �!       V                        �      i       \i      �       ��~�      �       \�      �       ��~                             �      E       0�E      I       PI      �       ^�      �       0��      m       ^m      q       0�q      {       ^|!      �!       ^                              �       ]�      q       ]q      {       ]|!      �!       ]                          �      �       ��~�      �       P�      q       ��~q      {       ��~|!      �!       ��~                                  Q      s       0�s      �       S�      �       S�             4s �             5s �             4s �      $       0�$      V       Pq      {       4s �|!      �!       4s �                     �      �       0��      �       0��      �       0�                      }      �       S�      R       ��~�      ]       ��~{      �       S                                  }      �       V�      �       U�             V             U      K       VK      O       UO      e       V�      ]       V{             U      �       V                       �      �       P�      e       ��~�      ]       ��~{      �       ��~                         �      �       P�      e       ��~�      ]       ��~�      �       P�      �       ��~                           e       ^�      ]       ^�      �       ^                                     P      �       ��~�      �       P�      �       ��~                         !      %       P%      e       ��~�      ]       ��~�      �       P�      �       ��~                         �      �       Q�      �       R�      �       ]�      e       ��~�      ]       ��~                            A       PP      R       P�              P                       �      R       ��~�      �       ��~              P      ]       ��~                          R       _�             _                       �      &       ]&      *       Q*      4       }�4      R       ]�      ]       ]                            �      �       0��      �       P�      R       \R      a       ��~a      e       0��      G       \G      ]       P{      �       0�                        `
      �
       U�
      �
       V�
      �
       �U��
      #       V                        `
      x
       Tx
      �
       S�
      �
       �T��
      #       S                      `
      
       Q
      �
       R�
      #       �Q�                        #       P                       `
      x
       t��x
      �
       s���
      �
       �T#���
      #       s��                          �      �       U�      �       �U��      �       U�             �U�      &       U                        �      �       T�      �       S�             �T�      &       T                          �      �       Q�      �       �Q��      �       Q�             �Q�      &       Q                          �      �       R�      �       �R��      �       R�             �R�      &       R                              �      �       X�      �       �X��      �       X�      �       �h�      �       �X��             �h      &       X                                �      �       Y�      �       �Y��      �       Y�      �       w �      �       �Y��             w              �`      &       Y                             �      �       3��      �       P�      �       3��      �       P�             P             3�      &       P                     �      �       0��      �       T      &       0�                    0      5       U5      :       �U�                    0      9       T9      :       �T�                  �      �       R�      �       �R�                    p	      �	       U�	      �	       �U�                      p	      {	       T{	      �	       P�	      �	       �T�                          p	      �	       Q�	      �	       S�	      �	       �Q��	      �	       S�	      �	       �Q�                    �	      �	       P�	      �	       Q                          @      W       UW      b       Sb      k       �U�k      �       U�      }       S                            @      �       T�      k       �T�k      �       T�      �       �T��      �       T�      }       �T�                      @      w       Qk      k       Qk      �       q��      �       Q                                  @      �       R�      }       \}      k       �R�k      �       R�      �       \�      �       �R��      �       \�      �       R�      }       �R�                          K      j       ^k      �       ^�      �       ^�      �       t �      }       ^                        m      b       ]k      �       ]�      �       ]�      }       ]                           K      �       0��      �       P�      �       P�             Pk      �       0��      B       P                         K      W       u��W      b       s��b      k       �U#��k      �       u���      }       s��                        ~      b       V�      �       V�      �       V�      }       V                        �      )       \)      -       |��      P       \P      S       |�                          )       \)      -       |�                            C       PC      W       p|�W      \       P                  ;      \       Q                    �      #       \#      ;       |�                      �      �       T�      #       t�#      ;       T                                      �      �       Q�      �       R�              t���              R             Q             t��1%Ut��1$�!�             Q             R            > t��1%Ut��1$�!2%3t��1%Ut��1$�!2$�!�              r q !�       2       Q                    B      P       \P      S       |�                      B      k       Pk      q       p~�q      x       P                  c      }       Q                        @      �       U�             V             �U�      1       U                      @      �       T�             �T�      1       T                              L      �       S�      �       u �      �       S�      �       u �             S      /       S/      1       u                              L      �       s� �      �       u #@�      �       s� �      �       u #@�      �       s�       /       s� /      1       u #@                        y             Q      �       q`��      �       Q      1       Q                �      �       0�                �      �       V                 �             s��                          "      /"       U/"      ~"       \~"      �"       U�"      �"       ^�#      $       \&$      U$       \                                "      /"       T/"      �#       S�#      �#       �T��#      �#       S�#      �#       �T��#      $       S$      &$       �T�&$      U$       S                        "      /"       Q/"      �#       V�#      �#       ]�#      U$       �Q�                    "      /"       R/"      U$       �R�                    "      /"       X/"      U$       �X�                                '"      /"       T/"      �#       S�#      �#       �T��#      �#       S�#      �#       �T��#      $       S$      &$       �T�&$      U$       S                              0"      K"       P_"      g"       P�"      �"       P�"      �#       0��#      �#       0��#      �#       P�#      $       P&$      B$       P                      W"      g"       P�#      �#       PC$      K$       P                  �#      $       P                      �"      �"       P�"      �#       s��#      �#       s�                  �"      4#       X                    �"      p#       0�p#      �#       1��#      �#       0�                 �"      #       P                 4"      L"       S                       4"      �"       S�#      $       S$      &$       �T�&$      U$       S                 �#      �#       S                 �#      �#       S                   $      $       S$      &$       �T�                   $      $       S$      &$       �T�                    �       �        U�       �       �U�                   �       �        U�       �       �U�                  �       �       X                     �       �        0��       )       UL      �       U                         �       �        S�       �        [�               Rl      r       [r      �       R                          �              R             P              Rl      r       Rr      �       P                          �              	 y �����       5       0�5      H       ZH      L       u L      Z       0�Z      �      	 y �����                         �       <       0�<      L       PL      k       0�k      l       Pl      �       0�                          �       �        q �              u { "1%4$x "             q               u { "1%4$x "l      r       q                     @       L        UL       �        �U�                   @       L        UL       �        �U�                  D       �        X                   D       L        0�L       �        U                        H       k        Yk       �        R�       �        Y�       �        R                          X       w        Rw       �        P�       �        R�       �        R�       �        P                     D       �        0��       �        P�       �        0�                          b       k        q k       �        u y "1%4$x "�       �        q �       �        u y "1%4$x "�       �        q                          1        U                                 U                                   P               u                       �      �       U�      <       S<      >       �U�                    �             T      >       �T�                  �      =       v��                          @      ^       U^      �       S�      �       u�~��      �       S�      �       �U�                    T      �       ]�      �       ]                        �      �       0��      �       V�      �       v��      �       V                    �      �       \�      �       \                      �      �       U�      �       �U��      �       U                     �      �       U�      �       �U��      �       U                             	      	       Q	      B	       \B	      G	       �Q�G	      `	       \`	      e	       �Q�e	      h	       Q                        	      	       T	      D	       ]G	      b	       ]e	      h	       T                    	      G	       0�G	      e	       1�e	      h	       0�                       	      	       0�3	      =	       s�G	      X	       s�e	      h	       0�                        �	      �	       U�	      �	       �U��	      
       U
      Z
       �U�                        �	      �	       T�	      �	       �T��	      

       T

      Z
       �T�                            �	      �	       Q�	      �	       S�	      �	       �Q��	      
       Q
      Y
       SY
      Z
       �Q�                   �	      �	       0��	      N
       0�N
      Z
       P                    �	      �	       T�	      �	      " `�H     ��H     �T4 $0.( �                    �	      

       T

      Z
       �T�                      �	      
       Q
      Y
       SY
      Z
       �Q�                    �	      
       U
      Z
       �U�                  
      Z
       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    P      W       UW             �U�                      P      �       T�      �       �T��             T                                        P      �       Q�      �       S�      �       �Q��      �       S�      �       �Q��      �       S�      �       �Q��      �       S�      �       �Q��      �       S�      �       �Q��             Q                                �      �       P�      �       Q�      �       P�      �       Q�      �       P�      �       Q�      �       P�      �       Q                      W      �       T�      �       �T��             T                    W      �       U�             U                            �      J       UJ      �       S�             �U�      '       S'      <       U<      \       S                        �      )       T)      '       �T�'      <       T<      \       �T�                      �      �       Q'      7       Q7      <       P                        �      �       R�      '       �R�'      <       R<      \       �R�                    �      	       ^      \       ^                   �      	       ^      \       ^                           �      J       u��J      �       s���             �U#��      '       s��'      <       u��<      \       s��                                        !       �]�Q�p�� !      %       �]�Q�p�\��%      1       �]�Q�p�\��V��1      @       �]�Q�P�\��V��@      J       �]�Q�s��\��V��J      �       �]��\��V���      �       �\��V��      '       �]��\��V��<      \       �]��\��V��                   �      J       ~�#�"�
���'      <       ~�#�"�
���                      p      |       U|      �       S�      �       �U�                    p      �       T�      �       �T�                  �      �       V                                       9       U9      B       ^B      T       ��~T      ~       ^~      M       ��~M      e       ^e      !'       ��~!'      4'       ^                                                                   T       B       SB      T       �T�T      ~       S~             ��~      �       �T��      M       ��~M      e       Se      w       �T�w      #       ��~#      D!       �T�D!      x!       ��~x!      �#       �T��#      �#       ��~�#      �%       �T��%      �%       ��~�%      !'       �T�!'      4'       S                           9       Q9      4'       ��~                           9       R9      4'       �R�                           9       X9      4'       �X�                  �&      �&       P                                      5      B       _B      I       w I      T       ��}T      �       _�      �       w �      T       VT      M       w M      e       Ve      !'       w !'      *'       V*'      4'       w                                           5      B       0�T      e       0�w      5       0�5      7       87      x       0�x      D!       VD!      x!       0�x!      �#       V�#      �#       0��#      U%       VU%      a%       0�a%      �%       V�%      �%       0��%      	&       V�&      '       V!'      4'       0�                                         �             0�             P:      ]       P             PJ      ^       P�      �       P�      �       P(       5        P"      "       P�"       #       0�I$      W$       P�$      �$       P�$      �$       0�                             �      r        \�!      "       \�#      "$       \:$      �$       \�$      U%       \a%      �%       \�&      '       \                                       �              0�       �        ]�!      "       0� #      �#       ]�#      "$       ]:$      I$       ]I$      �$       0��$      %       0�%      :%       ]:%      U%       0�a%      �%       0��%      !'       ]                                   �      R        0��!      "       0��#      �#       0��#      �#       
��:$      �$       0��$      &%       0�&%      :%       Q:%      U%       0�a%      �%       0��&      �&       
���&      '       Q                                 �              Q5       R        P�#      �#       PD$      I$       P[$      `$       Q%      5%       P�&      �&       P�&      �&       q��~��&      '       P                 �            
 ��H     �                 �             V                 /      J      
 Z�H     �                 /      J       V                 s      �      
 K�H     �                 s      �       V                 �      �      
 �H     �                 �      �       V                        (       
 $�H     �                        (        V                    r       �        \ #      "#       \                   �       �        0��       �        Q                        "#      0#       P0#      G#       \�%      �&       \'      !'       \                    1#      G#       P�%      �%       P                        #      �#       0��%      �&       0��&      �&       1�'      !'       0�                   &      �&       V'      !'       V                  #      "#      
 1�H     �                  #      "#       V                 "#      1#      
 B�H     �                 "#      1#       V                     �            
 ~�H     ��"       #      
 ~�H     ��$      �$      
 ~�H     �                     �             V�"       #       V�$      �$       V                       :      
 �H     �                       :       V                       u      O       S�       &!       Sx!      �!       S1"      �"       S                                 }      &!       Sx!      "       S1"      �"       S #      �#       S�#      "$       S:$      �$       S�$      U%       Sa%      �%       S�%      !'       S                      �      �       ]x!      �!       ]1"      �"       ]                 �      �       s�                                �      �       P             P/      >       PV      e       Px!      �!       P1"      <"       P�"      �"       P�"      �"       P                      m      �       \�      O       ]�       &!       ]                         m      �       ^�      �       T�      �       ^      O       ^�       &!       ^                 �      �      
 �H     �                 �      �       s�                 �            
 �H     �                        /      
 �H     �e      g      
 �H     �                  >      V      
 �H     �e      g      
 �H     �                   �             U>      O       U                  �      #       T                  �       !       0�                            �      Y       ��  w      �       ��  D!      x!       ��  �#      �#       ��  U%      a%       ��  �%      �%       ��  !'      4'       ��                                    �      �       ��~��      �       P�      1       � 1      Y       ��~�w      �       ��~�D!      x!       ��~��#      �#       ��~�U%      a%       ��~��%      �%       ��~�!'      4'       ��~�                                    �      �       U�      T       VT      M       w M      Y       Vw      �       w D!      x!       w �#      �#       w U%      a%       w �%      �%       w !'      *'       V*'      4'       w                                 �      ~       ^~      M       ��~M      Y       ^w      �       ��~D!      x!       ��~�#      �#       ��~U%      a%       ��~�%      �%       ��~!'      4'       ^                            �      Y       0�w      �       0�D!      x!       0��#      �#       0�U%      a%       0��%      �%       0�!'      4'       0�                                          �      �       0��      �       P�      ~       _~             ��~      �       ��~H@ ��      M       ��~M      Y       _w      #       ��~#      x       ��~H@ ��      �       0�D!      x!       ��~�#      �#       ��~U%      a%       ��~H@ ��%      �%       ��~!'      4'       _                                   �      �       U�      �       V�      7       0�7      g       v��"�      M       0�M      Y       Vw      Q       0�b      x       w �      �       w D!      x!       0��#      �#       0��%      �%       0�!'      *'       V*'      4'       w                               V                              Q                                 !      
 �pC     ��      M      
 �pC     �w      #      
 �pC     �D!      x!      
 �pC     ��#      �#      
 �pC     ��%      �%      
 �pC     �                                 !       ��  �      M       ��  w      #       ��  D!      x!       ��  �#      �#       ��  �%      �%       ��                                       ~       _~             ��~      !       ��~H@ ��      M       ��~w      #       ��~D!      x!       ��~�#      �#       ��~�%      �%       ��~                                   ~       ^~      !       ��~�      M       ��~w      #       ��~D!      x!       ��~�#      �#       ��~�%      �%       ��~                   `      m       1�m      v       ��~~      �       ��~      %       ��~                             (      m       
 �m             ��}�      M       ��}w      �       ��}�      #       ��}D!      x!       ��}�#      �#       ��}�%      �%       ��}                            m      m       1�~      �       1��             0��      M       0�w      #       0�D!      x!       0��#      �#       0��%      �%       0�                                        Y            	 s 8$8&��      �       Y�      �       ��~�      #      	 s 8$8&��#      �#       S                m      m       
 �m      �       V                 m      ~       0�                  m      ~       0�s!      x!       0�                               �      �       T�      �       ^�             T             ~��      �       T�      #       ~�D!      U!       P�#      �#       P                             m      ~       0��      �       0��              ]�      M       0�w      �       ]�      #       0�D!      s!       0��#      �#       0��%      �%       0�                  m      ~       0�s!      x!       0�                                                  5       0�5      <       P<      ~       [~      �       _�              P              _             [      !       0��      M       _w      �       P�      #       _D!      x!       _�#      �#       _�%      �%       _�%      �%       [                                    1       U1      !       ��~�      M       ��~w      #       ��~D!      x!       ��~�#      �#       ��~�%      �%       ��~                    �              Sw      �       S                 Q      ]       8                                       U       �       S�      �       �U��      �       U                                      U       �       S�      �       �U��      �       U                        �       V                         )       U                    �      �       U�      D       �U�                   �      �       U�      D       �U�                  �      D       X                     �      �       0��      �       U      D       U                         �      �       S�      �       [�      �       R/      5       [5      D       R                          �      �       R�      �       P�      �       R/      5       R5      D       P                     �      �       0��             u�#�             0�      /       q�#�/      D       0�                          �      �      	 y ������      �       0��             Z             u              0�      D      	 y �����                          �      �       q �      �       u { "1%4$x "�      �       q �      �       u { "1%4$x "/      5       q                                   U      y       �U�                                 U      y       �U�                        y       X                                0�      y       U                              +       Y+      P       Rc      i       Yi      y       R                                7       R7      K       PK      P       Rc      i       Ri      y       P                           R       0�S      S       0�S      c       q�#�c      y       0�                          "      +       q +      A       u y "1%4$x "A      K       q K      P       u y "1%4$x "c      i       q                  �      �       U                 �      �       U                    �      �       P�      �       u                     �,      �,       U�,      �,       P                                                        �,      �,       T�,      -       Q-      -       qy�-      #-       Q:-      e-       Qe-      ;.       �T�;.      �.       Q�.      �.       R�.      /       �T�/      j/       Qj/      s/       Rs/      �/       �T��/      P0       QP0      W0       RW0      �1       �T��1      �1       qy��1      
2       Q
2      2       R2      �2       �T��2      �2       Q�2      G5       �T�                    �,      �,       Q�,      G5       �Q�                                        �,      �,       R�,      &-       \&-      :-       �R�:-      .       \.      ;.       �R�;.      E0       \E0      �1       �R��1      �3       \�3      �3       �R��3      4       \4      w4       �R�w4      �4       \�4      G5       �R�                        �,      �,       X�,      5-       ]5-      :-       �X�:-      G5       ]                                       �,      �,       R�,      &-       \&-      :-       �R�:-      .       \.      ;.       �R�;.      E0       \E0      �1       �R��1      �3       \�3      �3       �R��3      4       \4      w4       �R�w4      �4       \�4      G5       �R�                        �-      �-       0��-      �-       P�-      ;.       ~��]�4      m4       ~��]�                           -      -       p�-      #-       T{0      �0       P�0      <1       \�1      �1       p��1      �1       T                              �,      �,       0��,      &-       V:-      N-       VN-      �-       }��-      ;.       _;.      �0       V�1      4       V4      m4       _w4      �4       V                      &-      &-       P/      /       6��3      �3       	���3      �3       3�m4      w4       6�B5      G5       S                    .      ;.       V4      m4       V                    .      ;.       \4      m4       \                    �4      �4       P�4      �4       P                  �.      �.       U                  �/      �/       U                 �/      �/       U                 �0      71       }�                      �0      �1       �Q�m4      w4       �Q��4      G5       �Q�                   �0      �1       Vm4      m4       V�4      B5       V                  <1      �1       \�4      B5       \                  (1      71       Q                              �0      r1       0�r1      �1       P�1      �1       S�1      �1       0�m4      m4       6��4      �4       P�4      85       S85      A5       PA5      B5       S                 (1      01       Q                 (1      01       ��}�                  32      A2       U                 J2      Z2       U                 c2      s2       U                     (      ;(       U;(      L(       \                         (      B(       TB(      �(       V�(      )       �T�)      �,       V                     (      u(       Qu(      �,       �Q�                                             (      ,(       R,(      �(       ^�(      )       �R�)      �*       ^�*      @+       �R�@+      U+       ^U+      �+       �R��+      �+       ^�+      I,       �R�I,      S,       ^S,      ],       �R�],      h,       ^h,      m,       �R�m,      y,       ^y,      �,       �R�                                             (      �(       X�(       )       ] )      )       �X�)      �)       X�)      �)       ]�)      �)       X�)      E*       ]E*      �*       X�*      �+       ]�+      �+       X�+      I,       ]I,      S,       XS,      ],       ]],      �,       X                                            '(      ,(       R,(      �(       ^�(      )       �R�)      �*       ^�*      @+       �R�@+      U+       ^U+      �+       �R��+      �+       ^�+      I,       �R�I,      S,       ^S,      ],       �R�],      h,       ^h,      m,       �R�m,      y,       ^y,      �,       �R�                                           '(      �(       X�(       )       ] )      )       �X�)      �)       X�)      �)       ]�)      �)       X�)      E*       ]E*      �*       X�*      �+       ]�+      �+       X�+      I,       ]I,      S,       XS,      ],       ]],      �,       X                              b)      �)       \Q*      b*       \b*      g*       Sg*      +       \+      8+       [U+      ],       \],      m,       Sm,      �,       \                        b)      g)       |�g)      �)       Q*+      8+       Pg+      �+       S7,      I,       S                                           (      �(       0�)      �)       0��)      �)       P�)      �)       0��)      �)       P�)      ,*       0�,*      @*       P@*      +       0�+      +       P+      ;+       S;+      D+       PU+      �+       0��+      �+       P�+      �,       0�                  �(      �(      
 e�H     �                  �(      �(       U                   �(      �(      
 q�H     �@*      E*      
 q�H     �                       �(      �(       P�(      �(       U�(      �(       P@*      E*       U                        Q*      �*       _U+      �+       _�+      D,       _I,      �,       _                        Q*      �*       �  U+      �+       �  �+      D,       �  I,      �,       �                          Q*      �*       �  U+      �+       �  �+      D,       �  I,      �,       �                          Q*      �*       VU+      �+       V�+      D,       VI,      �,       V                                Q*      b*       \b*      g*       Sg*      �*       \U+      �+       \�+      D,       \I,      ],       \],      m,       Sm,      �,       \                      �*      �*       	���+      �+       	���+      �+       ^],      ],       	��m,      y,       	��                                     Q*      b*       \b*      g*       Sg*      �*       \U+      [+       \[+      �+       S�+      �+       \�+      �+       S�+      �+       P�+      2,       S7,      D,       SI,      S,       \S,      m,       Sm,      �,       \                                 Q*      b*       \b*      �*       SU+      _+       S_+      �+       T�+      �+       S�+      7,       T7,      D,       t�I,      S,       \S,      ],       T],      �,       S                   �*      �*       Rb,      m,       0�                   �*      �*       _�+      �+       _b,      b,       _y,      �,       _                   �*      �*       \�+      �+       \b,      b,       Sy,      �,       \                    �*      �*       P�+      �+       P                    P5      m5       Um5      z5       S                                P5      p5       Tp5      �6       ^7      7       ^7      '7       QG7      �7       ^�7      �7       Q�7      
9       ^9      �B       ^                        P5      �5       Q�5      7       �Q�7      7       Q7      �B       �Q�                    P5      W5       RW5      �B       �R�                        P5      6       X6      >7       V>7      G7       �X�G7      �B       V                        ]<      <      	 r 8$8&��<      �<      	 r 8$8&�\?      `?      	 r 8$8&�uA      |A      	 r 8$8&�                    �<      �<       r 
��v8#�"�
��7��?      �?       r 
��v8#�"�
��7�                        7      '7       T�7      �7       T:      :       P:      b:       S                        L<      �<       T�<      �<       t��<      +=       T\?      �?       TuA      �A       T                             L<      <       0�<      �<       Y�<      �<       q��<      �<       Q�<      �<       Y\?      `?       QuA      �A       0�                        A<      O<       x 1$�O<      +=       U\?      �?       UuA      �A       U                       �5      6       X6      >7       V>7      G7       �X�G7      �B       V                                   �8      �8       _t:      ;       _�;      �;       P8<      @?       _\?      }@       _�@      A       QA      .A       _hA      �A       _�A      aB       _sB      �B       _                               �5      �6       ]7      67       ]G7      �7       ]�7      
9       ]9      �9       ]�9      �9       v8t:      @?       ]T?      �B       ]                    �5      @7       \G7      �B       \                        B      .B       P.B      aB       sB      wB       PwB      �B                           #@      V@       R!A      .A       R                  *6      @6       U                   s>      �>       U�A      �A       U                  �:      ;       U                  �=      �=       U                    P>      f>       U�A      �A       U                             J       UJ      �       S�      �       �U�                             *       T*      �       ]�      �       �T�                               C       QC      �       V�      �       |��      �       �Q�                  �      �       R                  J      f       U                 �      �       U                 �      �       T                        �       1       U1      7       u�7      �       U�      �       u��      �       U                         �              0�      4       P7      a       Pk      �       P�      �       
��                       �       �        0��       b       Xk      �       X�      �       0��      �       1�                                d        Ud       h        u�h       �        U�       �        u��       �        U                           "       K        0�K       `        Ph       �        P�       �        q ��       �        P�       �       
 ��������                              "        0�"       �        Y�       �        Y�       �        0��       �        1�                        `      �       U�      �       S�      �       �U��      �       U                      `      �       T�      �       �T��      �       T                   y      �       Q�      �       Q                          �      �       V�      �      
 q 1%q "#��      �       V�      �       V�      �      
 q 1%q "#�                   �      �       �����      �       ����                     �      �       u�      �       s�      �       u                        �             U             S             �U�             U                    �             P             P                      �      �       U�             u�      9       U                       �      �       0��             P      7       P8      9       0�                      @      u       Uu      �       u��      �       U                       @      b       0�b      x       P�      �       P�      �       0�                      �      &       U&      '       �U�'      K       U                      �      "       T"      '       �T�'      K       T                    �      &       X'      K       X                   �      &       x� '      K       x�                    �      &       x�'      K       x�                        �      �       Q�      �       q`��      &       Q'      K       Q                           "       T"      '       �T�                           &       U&      '       �U�                      P      j       Uj      �
       V�
              �U�                  
      �
       \                                        �      �       0��      	       \	      	       |�	       	       \?	      A	       0�A	      S	       ]S	      r	       }�r	      �	       ]�	      �	       0��	      �	       ]�	      �	       }��	      �	       ]�	      
       0�
      
       ]
      2
       }�2
      K
       ]
      �
       0��
      �
       ]                             ?	      W	       \W	      {	       |H�{	      �	       \�	      �	       |H��	      
       \
      ;
       |H�;
      K
       \                  d      �
       S                            �      e       Ue      �       \�      �       �U��      �       \�      �       �U��             \                    �      p       Tp             �T�                          �      A       QA      �       V�      �       �Q��      �       V�             �Q�                      �      L       RL      �       ^�             �R�                      Y      �       ^�      �       �R��      �       �R��             �R�                          Y      �       V�      �       �Q��      �       �Q��      �       �Q��      �       V�             �Q�                      Y      p       Tp      �       �T��      �       �T��             �T�                      Y      e       Ue      �       \�      �       \�             \                       �      D       0��      �       0��      �       0��      �       0�                         n      p       0�p      �       _�      �       U�      �       _�      �       _�             _                                      n      p       Tp      �       t��      �       T�      �       t��      �       T�             V(      D       S�      �       S�      �       V�      ]       S]      �       V�      �       S�      �       S�      �       V             S                                       �      �       V�      D       S�      �       S�      �       V�             S      ]       V]      �       S�      �       V�      �       S�      �       S�      �       V             S                    �      �       ^�      �       ^�             ^                            �      P       0�P      Y       PY      �       0��      l       0�l      �       P�      �       0��             0�                                       U      7       S7      <       �U�<      C       SC      D       �U�                                   T      "       U"      D       �T�                    #      +       P<      B       P                                      8       U8      \       S\      �       �U��      �       S�             �U�             S      7       �U�7      �       S                                        .       T.      z       V�      9       V�      �       V-      A       V      .       V.      7       �T�7      �       V�      �       V                                  D       QD      �       \�      �       �Q��      0       \0      7       �Q�7      �       \                       �       �+^  �                                    E      M       P�      �       P�      �       P�      �       _      H       PH             _7      Y       P}      �       P�      �       _�      �       _                  �             P                               \      z       S�      �       ^�             S_      u      
 s�Hq "��             ^      -       S�      �       ^�      �       ^                      5      �       ]�      2       ]7      �       ]                               \                 �      �       \                  7      c       1��      �       1�                  7      c       S�      �       S                  7      c       V�      �       V                    L      _       [_      �       ���      �       s��"#S�                   (      <       Z<      �       w                    M      c       _�      �       _                      ['      �'       Y�'      �'       y��'      �'       Y                     w'      �'       Q�'      �'       q��'      �'       Q                  ['      �'       P                  l'      w'       X                        P�      �       U�      /�       S/�      5�       U5�      F�       �U�F�      {�       S                          P�      �       T�      /�       �T�/�      5�       T5�      u�       �T�u�      ��       T��      {�       �T�                                P�      ��       Q��      �       ]�      /�       �Q�/�      5�       Q5�      u�       �Q�u�      ��       Q��      ��       ]��      2�       �Q�2�      {�       ]                            P�      �       R�      /�       �R�/�      5�       R5�      u�       �R�u�      ��       R��      ��       ^��      {�       �R�                                  P�      �       X�      %�       \%�      /�       �X�/�      5�       X5�      F�       �X�F�      u�       \u�      ��       X��      ��       �X���      "�       \"�      {�       �X�                              P�      �       Y�      /�       �Y�/�      5�       Y5�      u�       �Y�u�      ��       Y��      ��       _��      2�       �Y�2�      {�       _                                    P�      5�       0�5�      5�       2�F�      ��       0���      ��       P��      �       V�      ��       P��      ��       V��      �       0��      �       2��      2�       0�2�      =�       P=�      {�       V                u�      x�       �                    u�      u�       Tu�      ��       t 2$s�
"��������      ��       �T2$s�
"������                u�      x�       S                u�      x�       ��~�                      u�      ��       ����      ؠ       Pؠ      x�       Vx�      x�       0�                    u�      ��       s���      ̠       \̠      x�       ��~                   ?�      ?�       T?�      J�       t�J�      J�       t�J�      V�       t�V�      Z�       t.�Z�      x�       | 1$| "4$s�	"#6�                    ȡ      ��       \2�      {�       \                	��      ��       Y                
��      ��       r @B$ $0.�                     ��      %�       � F�      u�       � ��      2�       �                          ��      �       X�      %�       \F�      u�       \��      "�       \"�      2�       �X�                     ��      ��       Q��      �       ]��      %�       ]                     ��      ��       T��      О       QО      �       t 2$u�
"������                       ��      �       U�      %�       SF�      u�       S��      2�       S                    ��      О      H q2$u�	"��H$q2$u�	"#��@$!q2$u�	"#��8$!q2$u�	"#��!�О      �      � t 2$u�
"�����#2$u�	"��H$t 2$u�
"�����#2$u�	"#��@$!t 2$u�
"�����#2$u�	"#��8$!t 2$u�
"�����#2$u�	"#��!�                      1�      ��       ]F�      u�       ]��      "�       ]                  <�      ��       V                        ğ      �       PF�      r�       P��      �       P�      "�       P                        ��      �       0��      �       5��~����      %�       5��~��F�      k�       5��~����      �       5��~��                                      �      �       P�      �       V�      *�       P*�      <�       V��      ��       P��      ��       V��      ��       P��      %�       VF�      u�       V��      ��       V��      �       2��      �       V                   ��      ��      
 q2$u�	"���      О       q2$u�	"#�О      �       t 2$u�
"�����#2$u�	"#�                                      @R      bS       UbS      �S       V�S      �S       �U��S      �S       U�S      <T       V<T      �T       U�T      W       VW      *W       U*W      XX       VXX      ]X       U]X      hY       V                                        @R      rR       TrR      �S       S�S      �S       �T��S      �S       S�S      �S       �T��S      �S       T�S      �U       S�U      �V       �T��V      *W       S*W      �W       �T��W      4X       S4X      hY       �T�                              @R      �R       Q�R      �S       ]�S      �S       �Q��S      �S       ]�S      �S       �Q��S      �S       Q�S      hY       ]                              @R      �R       R�R      �S       ^�S      �S       �R��S      �S       ^�S      �S       �R��S      �S       R�S      hY       ^                          @R      uS       XuS      �S       \�S      �S       �X��S      �S       X�S      hY       \                                    @R      �S       Y�S      �S       �Y��S      7T       Y7T      �T       �Y��T      �U       Y�U      �V       �Y��V      �V       Y�V      �W       �Y��W      $X       Y$X      hY       �Y�                   HR      TR       u� �S      �S       u�                        HR      TR       u� �R      �R       T�R      �R       t��R      S       T�S      �S       u�                                   �R      �R       [�R      �R       { 
����R      �S       [�S      �S       [�S      &T       [�T      [U       [�U      �U       [�V      *W       [�W      �W       [                       �R      �R       p 8$z��!
����R      �R       z��8$z��!
����R      �R       q 8$p��!
����R      S       r 8$p��!
���S      S       p��8$p��!
���                          US      �S       q 
����S      T       q 
����T      �T       q 
����U      �U       q 
����V      �V       q 
���                                        qS      �S       z �8$u �!
����S      "T       z �8$u �!
���"T      7T       z �8$����!
���7T      �T       ����8$����!
����T      U       z �8$u �!
���U      �U       z �8$����!
����U      �U       z �8$u �!
����V      �V       z �8$u �!
����V      �V       z �8$����!
����V      *W       ����8$����!
����W      $X       z �8$����!
���$X      4X       ����8$����!
���                                 HR      �S       0��S      �S       Q�S      �U       0��U      �U       QV      V       Q�V      "W       0�"W      *W       Q�W      
X       0�
X      $X       Q$X      /X       0�                                    HR      �S       0��S      �S       R�S      �U       0��U      �U       RV      V       RV      	V       r q �	V      xV       S�V      %W       0�%W      *W       R�W      X       0�X      $X       R$X      /X       0�                        %S      1S       P1S      GS      / ��4�H0H%�$!0)( 8/��������S      �S       P�S      �S      / ��4�H0H%�$!0)( 8/�������                      -U      [U       0�[U      �U       P�W      �W       0�                            ?U      CU       q ��8$p��!
���CU      GU       u 8$p��!
���GU      JU       u 8$��1��!
���JU      [U       q ��8$��1��!
����U      �U       U�W      �W       q ��8$��1��!
���                      bT      �T       0��T      �T       Q$X      ,X       Q                    YT      �T       T$X      4X       T                             �T      �T       p 8$q��!
����T      �T       q��8$q��!
����T      �T       ��2��8$��1��!
����T      �T       { ��8${��!
����T      �T       p 8${��!
����T      �T       { ��8${��!
���$X      4X       { ��8${��!
���                     V      �V       ��*W      �W       ��4X      hY       ��                     V      �V       \*W      �W       \4X      hY       \                     V      �V       ^*W      �W       ^4X      hY       ^                     V      �V       ]*W      �W       ]4X      hY       ]                   V      	V       r q �	V      xV       S                         V      �V       V*W      �W       V4X      XX       VXX      ]X       U]X      hY       V                               5V      LV       PMV      `V       P;W      ?W       P?W      IW       ��pW      �W       0��W      �W       PPX      ]X       PY      Y       0�                	       V      4V       v4V      �V       _*W      �W       _4X      hY       _                     �V      �V       S*W      �W       S4X      hY       S                        fW      yW       ZzX      �X       Z�X      Y       ��Y      hY       Z                      �W      �W       P�W      �W       qy��W      �W       v#�
���                 �W      �W       R                         �W      �W      
 p r #3%��W      �W      
 qyr #3%��W      �W       v#�
��r #3%��W      �W       P�W      �W       v#�
��r #3%�                  �W      �W       Q                   zX      �X       YY      hY       Y                  zX      Y       VY      hY       V                      zX      �X       0��X      Y       PY      Y       0�Y      hY       0�                                      �X      �X       P�X      �X       P�X      �X       qY       Y       P Y      1Y       q1Y      4Y       P4Y      FY       qFY      IY       PIY      ^Y       q^Y      cY       PcY      hY       q                        �X      �X       t 
����X      �X      
 v�
����X      �X      	 q �
���Y      hY      	 q �
���                     zX      �X       v�X      �X       QY      hY       Q                  �X      �X       T                        pY      Z       UZ      �Z       S�Z      �Z       �U��Z      �Z       S                      pY      �Y       T�Y      Z       _Z      *Z       �*Z      MZ       ~�MZ      MZ       �MZ      gZ       _�Z      �Z       _                    pY      �Y       Q�Y      �Z       �Q�                        pY      Z       RZ      �Z       \�Z      �Z       �R��Z      �Z       R                        pY      �Y       X�Y      �Z       ]�Z      �Z       �X��Z      �Z       ]                        pY      Z       YZ      ZZ       v�ZZ      �Z       �Y��Z      �Z       Y                       pY      RZ       0�RZ      VZ       PZZ      �Z       P�Z      �Z       0�                    �Y      Z       X�Z      �Z       X                    �Y      Z       0��Z      �Z       0�                 pY      rY       u#                 pY      rY       u#                 pY      rY       u#                 pY      rY       u#
                 pY      rY       u#                	 pY      rY       u#                  MZ      QZ       T                 MZ      QZ                               �#      q$       Uq$      �%       �U��%      &       U&      F&       �U�                            �#      4%       T4%      ^%       T�%      �%       T�%       &       T &      *&       t�*&      /&       T/&      7&       t�7&      F&       T                          �#      �#       Q�#      e$       Se$      �%       ���%      &       S&      F&       ��                                �#      \$       R\$      `$       [`$      �$       �R��$      �$       R�$      �$       Z�$      �%       _�%      �%       _�%      &       R&      F&       _                        �#      l$       Xl$      �%       �X��%      &       X&      F&       �X�                    �#      �#       Y�#      F&       �Y�                             �#      �$       y�$      �%       [�%      �%       [�%      �%       S�%      �%       [�%      &       y&      F&       [                         �#      �$       y�$      �%       ���%      �%       ���%      &       y&      F&       ��                        �#      "$       Q"$      q$       u#�
���q$      �$       �U##�
����%      &       Q                                 �#      	$      	 p �
���	$      q$      
 u�
���q$      �$        
����$      �$       } 
����$      �%      	 w �
����%      �%      	 w �
����%      &      	 p �
���&      &      
 u�
���&      F&      	 w �
���                       �#      "$       u"��q �"$      q$       u"��u#�
���q$      �$       �U#"���U##�
����%      &       u"��q �                         �$      �$       } 
����$      �%       ]�%      �%       }��%      �%       ]�%      �%       ]&      F&       ]                              �$      �$       0��$      0%       X0%      [%       R[%      �%       X�%      �%       X�%      �%       X&      #&       X#&      /&       _/&      F&       X                   �#      �$       y �%      &       y                       �#      $       Z$      �$       y�%      &       Z                    �#      �$       Y�%      &       Y                                �$      �$       0��$      �$       P�$      �$       Q	%      D%       PD%      F%       UJ%      �%       P�%      �%       Y�%      �%       P�%      �%       P&      F&       P                               �$      �$       [�$      0%       S0%      <%       Q<%      >%       q�>%      [%       Q�%      �%       [�%      �%       S&      >&       [>&      F&       S                          %      %      	 ~ ����Q%      [%       v 3$z "��%      �%       ^�%      �%       Z>&      F&      	 ~ ����                            �!      �!       U�!      �"       �U��"      �"       U�"      �#       �U��#      �#       U�#      �#       �U�                          �!      d"       Td"      |"       T�"      �#       T�#      �#       Z�#      �#       T                            �!      -"       Q-"      �"       �Q��"      �"       Q�"      �#       �Q��#      �#       Q�#      �#       �Q�                              �!      "       R"      "       r 7�"      G"       RG"      �"       �R7��"      �"       R�"      �#       X�#      �#       R�#      �#       �R7�                            �!      "       X"      �"       �X��"      �"       X�"      �#       �X��#      �#       X�#      �#       �X�                    �!      �!       Y�!      �#       �Y�                             �!      �!       z"      �"       Y�"      �#       Y�#      �#       Q�#      �#       Y�#      �#       z�#      �#       P                   �!      �!       z�#      �#       z                      �!      "       Y�"      �"       Y�#      �#       Y                     �!      �!      	 p �
����#      �#      	 p �
����#      �#      
 u�
���                   �!      �!       u"��y ��#      �#       u"��y �                              G"      �"       [�"      �"       {��"      �"       [�"      c#       [c#      j#       {�j#      �#       [�#      �#       [                   �!      �!       z �#      �#       z                       �!      �!       [�"      �"       [�#      �#       [                      �!      >"       Z�"      �"       Z�#      �#       Z                      G"      `"       Y`"      �"       P�#      �#       P                  `"      y"       y 3$p 3$s "�                         �"      �"       Y�"      "#       QW#      c#       q�p#      �#       Y�#      �#       Q                  �"      *#       S                                    �"      �"       0��"      #       U#      
#       P
#      #       U#      #       P#      *#       UF#      W#       UW#      Z#       u 8$�Z#      _#       Up#      �#       0��#      �#       U                      �       8!       Q8!      Z!       �Q�Z!      �!       Q                      �       &!       P&!      .!       Y.!      K!       p�K!      P!       t #�P!      y!       Y                 �       �!       u                        �E      F       UF      @F       S@F      JF       �U�JF      �H       S                        �E      �E       T�E      �E       TJF      �F       TG      BG       T                            �E      �E       Q�E      AF       VAF      JF       �Q�JF      #G       V#G      BG       QBG      �H       V                      dF      �F       QBG      �G       Q�H      �H       Q                       �F      �F       qBG      qG       q�G      �G       q�H      �H       q                          �F      �F       ZBG      gG       ZgG      qG       q�G      �G       Z�H      �H       Z                         �E      F       u�F      F       UF      8F       ]�G      �G       ]�G      �G       U                  �G      �H       ^                    �G      �G       P�G      �H       _                 �G      �H       s��                 �G      �H        
���                          F      ,F       P,F      0F       \0F      8F       P�G      �G       P�G      �H       \                		 �E      �E      
 t2$u�	"��E      �E       t2$u�	"#�                    �H      �H       U�H      �H       �U�                    �H      �H       T�H      �H       �T�                      �H      �H       Q�H      �H       R�H      �H       �Q�                      �(      �(       U�(      �(       S�(      �(       �U�                 �(      �(       u�                        �H      I       UI      uI       SuI      I       �U�I      �L       S                          �H      �H       T�H      I       QI      vI       VvI      I       �T�I      �L       V                                                   I      *I       P*I      2I       0�I      �I       0��I      �I       P=J      bJ       PcJ      xJ       P}J      �J       P�J      �J       P�J      �J       0��J      �J       P�J      �J       P�J      �J       P�J      'K       0�'K      DK       P�K      L       0�0L      IL       PJL      cL       PdL      oL       P                      �I      �I       P�I      }J       ]K      �L       ]                     BK      BK       QBK      GK       q�GK      IK       | #�IK      �K       | #��L      �L       | #�                      IK      aK      	 p  $ &�aK      �K      , | �H0H%�$!0)( 8/�� $ &��L      �L      , | �H0H%�$!0)( 8/�� $ &�                      SK      �K      	 q ������K      �K      . | #�H0H%�$!0)( 8/��������L      �L      	 q �����                  �K      �K       Q                      �I      �I       P�I      }J       _�L      �L       _                      �I      �I       P�I      �I       \�L      �L       \                      �I      �I       P�I      %J       ^�L      �L       ^                   J      %J       ^)J      }J       ^                         =      X=       UX=      d=       Sd=      j=       �U�j=      (>       S                  =      "=       u�                        =      X=       u��X=      d=       s��d=      j=       �U#��j=      (>       s��                     D=      X=       Pj=      ~=       P�=      >       P                 j=      �=       s��                     �=      �=       0��=      �=       V�=      �=       \�=      �=       V                 �=      (>       s��                                            �~      
       U
             S      $       �U�$      o       So      x       �U�x      (�       S(�      �       ���      Ё       �U�Ё      ق       Sق      ?�       �U�?�      w�       Sw�      ��       �U���      ��       S��      N�       �U�                              �~             V$      o       Vx      ق       V��      �       V?�      w�       V��      ȃ       V*�      9�       V                                               P      #       _#      /       P/      O       _O      o       Po      x       _x      �       P�      �       _Ё      ��       P                      G      o       ^x      �       ^Ё      	�       ^                              @      K       p } "�K      o       | } "�x      0�       | } "�0�      \�       ��} "�Ё      ܁       | } "�ς      ق       | } "�?�      w�       | } "�                       x      0�       | } "�0�      \�       ��} "�ς      ق       | } "�?�      w�       | } "�                           x      Ё       Vς      ق       V��      �       V?�      w�       V��      ȃ       V*�      9�       V                               x      (�       S(�      �       ���      Ё       �U�ς      ق       Sق      ?�       �U�?�      w�       Sw�      ��       �U���      N�       �U�                      �      Ё       ^ς      ��       ^��      N�       ^                        �      �       p 
����      Ё      
 ��~�
���ς      ��      
 ��~�
�����      N�      
 ��~�
���                            a�      m�       0�m�      ��       T��      Ё       ����      �       ��G�      w�       0���      %�       ��*�      I�       ��                           �      �       0��      �       P�      Ё       ��ς      �       ���      ��       0���      ��       ����      N�       ��                                               �             0�      �       P�      Ё       _ς      ق       0�ق      �       ���      ��       0���      �       _�      ?�       ��?�      j�       0�j�      w�       Pw�      ��       ����      Ӄ       _Ӄ      ؃       ��؃      *�       V*�      /�       _/�      9�       ��9�      N�       V                    �      0�       0�?�      w�       0�                  a�      m�       0�G�      w�       0�                    u�      }�       P}�      ��       p�}���      ��       R                              ʀ      �       0��      i�       \��      Ё       \��      �       \��      ΃       \΃      *�       ]9�      N�       ]                              �      �       p ���      �      	 ������      z�       ]��      ��       p ����      ��       } ��ˁ      Ё       ]*�      9�       ]                    ��             s p �      ˁ       ]                  �      �       0�                 w�      ��       s��                 Ё      ܁       | } "�                   Ё      ς       V��      ��       V                   Ё      ς       S��      ��       S                    ܁      ς       ]��      ��       ]                      �      	�       p 
���	�      ς       ^��      ��       ^                         ܁      >�       0�>�      B�       PB�      b�       Rb�      ��       ��~ł      ς       0���      ��       ��~                    s�      ��       0���      ��       P                      ��      ��       P��      ��       r �8$8&���      ��       r p "�8$8&p "���      ��       Q                 ��      ��       s��                        0.      w.       Uw.      ,/       S,/      6/       �U�6/      �0       S                    0.      i.       Ti.      �0       �T�                        0.      p.       Qp.      5/       _5/      6/       �Q�6/      �0       _                        0.      b.       Rb.      1/       ]1/      6/       �R�6/      �0       ]                                0.      �.       X�.      //       \//      6/       �X�6/      a/       \a/      p/       Xp/      0       \0       0       X 0      �0       \                 0.      2.       u�                  �.      �.       P                               �.      �.       R�.      �.       Ta/      z/       Tz/      �/       X�/      �/       ���/       0       T�0      �0       T�0      �0        v 1$#������"�                   �.      �.       U�.      �.       Q                           �.      �.       t q "��.      �.       Qa/      �/       Q�/      0       w 0       0       Q�0      �0       w                         �.      �.       P�.      �.       Va/      ~/       P~/      �0       V                    [.      3/       ^6/      �0       ^                   �.      '/       S6/      a/       S                          �Q      �Q       U�Q      �Q       s�|��Q      R       �U�R      2R       S2R      4R       s�|�                            �Q      �Q       T�Q      �Q       Q�Q      R       VR      R       �T�R      &R       Q&R      4R       V                    �Q      �Q       Q�Q      4R       �Q�                      �Q      �Q       P�Q      R       P'R      4R       P                   �Q      R       S2R      4R       S                   �Q      �Q       u���Q      �Q       S                        �-      �-       U�-      �-       P�-      .       �U�.      %.       P                          �-      �-       T�-      .       V.      .       �T�.      #.       T#.      %.       V                      �-      �-       Q�-      .       �Q�.      %.       Q                      �-      �-       P�-      
.       S
.      .       P                    �-      �-       xtmv��-      �-       T.      %.       xtmh�                    �-      .       \.      %.       \                    �-      .       ].      %.       ]                              @9      e9       Ue9      n9       Vn9      {9       �U�{9      �9       V�9      �9       �U��9      8:       V8:      �:       �U�                              @9      `9       T`9      e9       Qe9      s9       Ss9      {9       �T�{9      �9       S�9      �9       �T��9      �:       S                 �9      �9       8�                      [9      n9       \{9      �9       \�9      F:       \                 8:      F:       0�                  �9      �:       } 
���                     [9      n9       0�{9      8:       0�8:      F:       V                            �L      �L       U�L      �L       S�L      �L       �U��L      M       SM      M       q�x�M      M       �U�                              �L      �L       T�L      �L       Q�L      �L       V�L      �L       �T��L      M       VM      M       UM      M       �T�                  �L      M       P                           �L      �L       u���L      �L       s���L      �L       �U#���L      M       s��M      M       QM      M       �U#��                            �P      �P       U�P      �P       S�P      �P       �U��P      �P       S�P      �P       q�z��P      �P       �U�                              �P      �P       T�P      �P       Q�P      �P       V�P      �P       �T��P      �P       V�P      �P       U�P      �P       �T�                  �P      �P       P                           �P      �P       u���P      �P       s���P      �P       �U#���P      �P       s���P      �P       Q�P      �P       �U#��                      0>      g>       Ug>      7?       \7?      :?       �U�                  O>      5?       V                     O>      g>       u��g>      7?       |��7?      :?       �U#��                     T>      {>       S{>      �>       s`��>      �>       S                  b>      �>       ]                     �>      �>       S�>      �>       sh��>      �>       S                  �>      ?       ]                         M      QM       UQM      fM       ^fM      iM       �U�iM      zP       ^                           M      GM       TGM      QM       QQM      _M       S_M      iM       �T�iM      zP       S                    ;M      bM       \iM      zP       \                      �M      �M       P�M      �N       VO      pP       V                    �M      FO       ]FO      �O        2$#����} "�-P      zP       ]                          �M      �M       P�M      �M       T�M      O       ��O      O       TO      zP       ��                       ;M      QM       u��QM      fM       ~��fM      iM       �U#��iM      zP       ~��                 �O      -P       _                    �O      �O       P�O      -P       w                         +N      GN       _GN      KN       QKN      �N       _-P      zP       _                             +N      GN       YGN      �N       w �N      �N       y��N      �N       Y�N      �N       w �1�-P      nP       w nP      zP       Y                        �P      �P       U�P      �P       S�P      Q       �U�Q      �Q       S                          �P      �P       T�P      �P       Q�P       Q       \ Q      Q       �T�Q      �Q       \                              �P      �P       PQ      Q       PQ      !Q       V!Q      kQ       PkQ      lQ       VlQ      �Q       P�Q      �Q       P                       �P      �P       u���P      �P       s���P      Q       �U#��Q      �Q       s��                    @�      F�       UF�      G�       �U�                    @�      F�       TF�      G�       �T�                    P�      V�       UV�      W�       �U�                    P�      V�       TV�      W�       �T�                        �D      OE       UOE      WE       �U�WE      �E       U�E      �E       �U�                        �D      RE       TRE      WE       �T�WE      �E       T�E      �E       �T�                      �D      �D       Q�D      VE       ZWE      �E       Z                          �D      �D       R�D      VE       QVE      WE       �R�WE      �E       Q�E      �E       �R�                        �D      VE       XVE      WE       �X�WE      �E       X�E      �E       �X�                   HE      OE       u�OE      VE       U                  fE      yE       P                         ;E      HE       YHE      VE       RWE      fE       YtE      �E       Y�E      �E       R                   �D      )E       UfE      yE       U                  �D      )E       T                   �D      
E       PE      )E       P                   E      )E       R                         �      ,�       U,�      i�       ]i�      n�       �U�n�      �       ]                         �      ?�       T?�      d�       Sd�      n�       �T�n�      �       S                        ;�      _�       ^n�      '�       ^�      ��       ^ي      �       ^                      �      '�       0�'�      �       _��      ��       _                                 ;�      _�       0�n�      ��       0���      �       \�      '�       0�'�      Έ       VΈ      ؈       v�؈      ܈       q��      h�       0�h�      ��       \��      ��       Vي      �       0�                                      '�      J�       ^�w �\�P�h�      l�       P��l�      t�       ^��t�      x�       ^�P��x�      �      	 ^�w ���      ��       ^�w �P����      ��       ^�w �\����      �       ^�w �\�P���      ��       ^�w �\�P���      ��       ^�w �\����      ��       ^�w �\�P�                 ��      ��       0�                 ��      �       0�                   �      ��       ���ي      �       ���                   �      ��       �"�  ��      ��       �"�  ي      ي       �"�                     �      ��       S��      ��       Sي      ي       S                 ��      ��       2�                     �      B�       0�B�      ]�       V]�      c�       v�ي      ي       V                   �      B�       0�B�      ��       \ي      ي       \                     �      B�       0�B�      ��       ��~��      L�       1�L�      ��       ��~ي      ي       1�                       �      B�       0�B�      X�       ��~X�      ]�       1�]�      ��       ��~ي      ي       ��~                   �      B�       0�B�      ��       _ي      ي       _                      �      �       P�      ��       w ��      ��       w ي      ي       w                       �(      &)       U&)      +)       �U�+)      6)       U                      �(      #)       T#)      +)       �T�+)      6)       T                      �(      *)       Q*)      +)       �Q�+)      6)       Q                      �(      *)       R*)      +)       �R�+)      6)       R                  )      *)       P                     �(      &)       U&)      +)       �U�+)      6)       U                     �(      &)       U&)      +)       �U�+)      6)       U                    �(      )       T+)      6)       T                   �(      )       P+)      5)       P                    �(      )       X+)      6)       X                      �             T      �        �T��       �        T                      �             Q      �        �Q��       �        Q                           �             0�              ]               P       �        ]�       �        ]�       �        0�                       �      �       S�      �       s��      	        S       �        S�       �        u�
                     �             1�      �        [�       �        1�                             �      �       P�      �       p��             R             r�             r�      J       r�J      c       r�c      �       T�      �       t��      �       T�      �       t��      �       T�              X       �        T�       �        T                    �              V       �        V                              �       R       #        R#       �        tr��       �        R�       �        tr�                  :      �        X                              �       r ��8$r��!
���       #        r ��8$r��!
���#       �        tr��8$ts��!
����       �        r ��8$r��!
����       �        tr��8$ts��!
���                                    %       r��8$r��!
���%      -       x 8$r��!
���-      0       p 8$r��!
���0      �       r��8$r��!
���       #        r��8$r��!
���#       �        tt��8$tu��!
����       �        r��8$r��!
����       �        tt��8$tu��!
���                              �       r��8$r��!
���       #        r��8$r��!
���#       �        tv��8$tw��!
����       �        r��8$r��!
����       �        tv��8$tw��!
���                        c      f       q 
���f             Q�      �       Q       #        Q                                 �       0�       �        0��       �        P�       �        0��       �        P�       �        0�                   #       �        ^�       �        ^                        #       G        QG       x        Y�       �        Q�       �        Y                          /       V        YV       n        Rn       x        Y�       �        Y�       �        R                        8       8        P8       Y        p�[       ^        t p "#�^       ^        P^       x        p��       �        p�                        >       G        Rd       n        Q�       �        R�       �       + p �H0H%�$!0)( 8/�������                  �      �       Q                              �      �      	 p ������      �       P�      �      + r�H0H%�$!0)( 8/��������      �      	 p ������      �       P�      �      + r�H0H%�$!0)( 8/��������       �        P                      `&      �&       U�&      �(       S�(      �(       �U�                            `&      t&       Tt&      �&       Q�&      E'       VE'      g(       �T�g(      u(       Vu(      �(       �T�                      �&      �&       P�&      �&       P�&      �(       Y                              �&      �&       R�&      �&       r��&      '       X'      '       x�'      ,'       x�,'      Y'       x�Y'      '       T'      '       t�'      �'       t��'      �'       t��'      �'       x��'      �'       x��'      �'       ^�'      (       x�(      (       x�(      *(       ^*(      @(       ~�@(      @(       ^@(      Y(       ~�Y(      g(       ^                  �&      �(       U                     �&      Y'       0�Y'      g(       Rg(      w(       0�                    �&      �&       p 
����&      �(       Z                     `&      Y'       0�Y'      g(       Vg(      w(       0�                     `&      Y'       0�Y'      g(       \g(      w(       0�                      �'      �'       p 
����'      �'       P
(      4(       P                    ,'      Y'       p 
����'      �'       p 
���                    0'      Y'       ^�'      �'       ^                 �'      �'       ~ 8%�                       '      Y'       XY'      �'       T�'      �'       X�'      g(       T                     '      Y'       1�Y'      o'       ]v'      g(       ]                    &(      Y(       QY(      ](       q�](      g(       Q                    (      #(       ��������@(      U(       PY(      _(       P                    1(      @(      & ~��@$~ ��H$!~��8$!~��!�F(      U(      & ~��H$~��@$!~��8$!~	��!�                      �      �       U�      �       �U��      �       U                      �      �       T�      �       �T��      �       T                     �      �       U�      �       �U��      �       U                   �      �       u�      �       u                          �Z      �[       U�[      W]       ��~W]      j]       �U�j]      }]       U}]      �]       ��~                          �Z      �Z       P�Z      �[       u��[      j]       ��~j]      }]       u�}]      �]       ��~                          �Z      �[       T�[      i]       w i]      j]       ��~j]      }]       T}]      �]       w                    �Z      �[       u�#j]      }]       u�#                    c\      e\       p q !�e\      �\       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                      0B      BB       UBB      WB       SWB      XB       �U�                 0B      1B       u                  0B      1B       u #�                      P      p       Up      u       Tu      v       �U�                    P      V       TV      v       �T�                  S      u       Y                 S      u       y�                 S      u       y�                    p�      ��       U��      ��       �U�                    p�      ��       T��      ��       �T�                      t�      ��       �h���      ��       Q��      ��       �h�                   p�      ��       T��      ��       �T�                   p�      ��       U��      ��       �U�                                      @4      ^4       U^4      ]5       _]5      6       �U�6      *6       _*6      .6       U.6      /6       �U�/6      @6       _@6      A6       �U�A6      _6       __6      c6       Uc6      �7       �U�                                      @4      J4       TJ4      �4       [�4      �4       Q�4      �4       [�4      6       �T�6      6       Q6      .6       [.6      A6       �T�A6      N6       [N6      c6       Qc6      �7       �T�                      @4      b4       Qb4      �4       T�4      �7       �Q�                                    c4      l4       Pl4      r4       p��4      �4       T�4      �4       t��4      B5       ~�B5      [5       ~�[5      ]5       u~�]5      �5       U�5      �5       u��5      �5       u~��5      6       U6      6       t�A6      N6       ~�d6      �6       U7      K7       UK7      [7       u�[7      p7       u~�p7      �7       U                                           ]5      �5       Y�5      �5       y��5      �5       Y�5      �5       y�d6      z6       Yz6      �6       y��6      �6       Y�6      �6       y��6      �6       Q�6      �6       X�6      �6       x��6      �6       X�6      �6       x��6      7       X%7      .7       T.7      K7       Y�7      �7       Y                    u4      �4      	 } ������4      �4       ]                      |4      �4       U6      6       UA6      U6       U                         �4      ]5       _]5      6       �U�6      6       _A6      N6       _d6      �7       �U�                  �4      �4      & } ��H$}��@$!}��8$!}��!�6      6       0�                        �4      �4      & t ��H$t��@$!t��8$!t��!��4      �4      & ~ ��H$~��@$!~��8$!~��!�6      6      & t ��H$t��@$!t��8$!t��!�A6      N6      & ~ ��H$~��@$!~��8$!~��!�                        B5      �5       Q6      6       Qd6      z6       Q�6      �6       T                         �4      �4       QB5      �5       ]6      6       ]6      6       0�d6      �6       ]�6      7       Y7      �7       ]                          ]5      �5       R�5      6       Rd6      t6       R7      K7       R�7      �7       R                      B5      �5       Z�5      �5       z��5      6       z�d6      �6       Z�6      �6       z��6      �6       z��6      �7       Z                 B5      ]5       1�                      ]5      ]5       1��5      �5       {��5      �5       [d6      �6       [                                     �5      �5       1��5      �5       0��5      6       1�z6      �6       1��6      �6       0��6      �6       1��6      �6       0��6      �6       1��6      �6       0��6      7       1�7      �7       1�                    5      6       Pd6      �7       P                   �4      �4       P�4      �4       p|��4      �4       P6      6       P                  �4      �4      & } ��H$}��@$!}��8$!}��!�6      6      & } ��H$}��@$!}��8$!}��!�                   �4      �4       0��4      �4       Q6      6       0�                            �3      �3       U�3      4       \4      4       �U�4      &4       \&4      '4       �U�'4      54       \                               �3      �3       T�3      �3       t��3      �3       v��3      �3       R�3      �3       r��3      	4       r~�	4      4       R4      $4       v�$4      '4       �T#�'4      54       v�                    �3      �3       Q�3      54       �Q�                            �3      �3       U�3      4       \4      4       �U�4      &4       \&4      '4       �U�'4      54       \                   �3      �3       0�'4      54       0�                    �3      4       P'4      54       P                              �2      �2       U�2      y3       \y3      |3       �U�|3      �3       \�3      �3       �U��3      �3       U�3      �3       \                            �2      �2       T�2      3       V3      03       S03      ;3       s�;3      I3       s�I3      k3       S�3      �3       T�3      �3       t��3      �3       �T#�                        �2      3       Q3      �3       �Q��3      �3       Q�3      �3       �Q�                             �2      �2       U�2      y3       \y3      |3       �U�|3      �3       \�3      �3       �U��3      �3       U�3      �3       \                     3      3      & v ��H$v��@$!v��8$!v��!��3      �3      & t ��H$t��@$!t��8$!t��!��3      �3      0 �T��H$�T#��@$!�T#��8$!�T#��!�                   3      3       RI3      R3      
 s��#��3      �3       0�                        (3      03       P03      ^3       Q^3      a3       q|�a3      k3       Q�3      �3       T                  I3      k3       R                     �2      �2       T�2      �2       t��2      �2       t��2      3       P3      3       p|�3      3       P�3      �3       t�                   �2      �2      & t ��H$t��@$!t��8$!t��!��3      �3      & t ��H$t��@$!t��8$!t��!�                   �2      �2       0��2      3       R�3      �3       0�                        �7      �7       U�7      \8       \\8      c8       �U�c8      �8       \                      �7      �7       T�7      �7       P�7      �8       �T�                                �7      �7       Q�7      &8       ^&8      I8       TI8      `8       ^`8      c8       �Q�c8      8       ^8      �8       T�8      �8       ^                       �7      �7       U�7      \8       \\8      c8       �U�c8      �8       \                    �7      �7       ]�8      �8       ]                           �7      �7       v
��7      �7       S�7      �7       s��7       8       s� 8      8       s|�8      I8       Sc8      �8       S�8      �8       v
�                         �7      �7       _�7      28       ]28      D8       }|�D8      Q8       ]c8      �8       ]�8      �8       _                   �7       8       s ��@$s��8$!s��!� 8      8       su��@$sv��8$!sw��!�                      8      8      	 p �����8      8       U8      8      	 p �����                    8      8      	 q �����8      &8       ��������                            �8      �8       U�8      9       \9      9       �U�9      &9       \&9      '9       �U�'9      59       \                      �8      �8       T�8      �8       Q�8      59       �T�                           �8      �8       U�8      9       \9      9       �U�9      &9       \&9      '9       �U�'9      59       \                      �8      9       V9      $9       V'9      59       V                           �8      �8       s
��8      �8       R�8      �8       r��8       9       rx� 9      9       R9      !9       s
�'9      59       s
�                    �8      9       P'9      59       P                   �8      �8       0�'9      59       0�                    �      �       U�      H       �U�                              �      �       T�             V             �T�      "       V"      .       T.      F       VF      H       T                          �      �       Q�      �       T�      .       �Q�.      4       T4      H       �Q�                    �      �       P�      �       p��      �       p�.      <       p�                    �      �      	 q �����.      <      	 q �����                      �            	 | �����      &      	 | �����.      H      	 | �����                    @      Y       UY      �       �U�                                @      I       TI      �       \�      �       �T��      �       \�      �       U�      �       �T��      �       \�      �       �T�                                @      ]       Q]             V      �       �Q��      �       V�      �       T�      �       �Q��      �       V�      �       T                          @      ]       R]      r       Tr      �       �R��      �       T�      �       �R�                    ^      c       Pc      r       p��      �       p�                    k      r      	 q ������      �      	 q �����                      n      w      	 } ������      �      	 } ������      �      	 } �����                  �      �       U�      <       u�                  �      <      & u ��H$u��@$!u��8$!u��!�                           �      �      & u ��H$u��@$!u��8$!u��!��      �       X�      �       R�             Y             R"      /       Y/      <       X                 �      �       0��      <       Z                          �      �       Y�      �       R�      �       Y�             R"      <       R                          �      �       P�      �       p��      �       P�      �       P�             p�"      ,       p�,      /       P                        �      �      	 q �����             q x !�����            	 q �����"      /      	 q �����                  �      �       U�      �       u�                  �      �      & u ��H$u��@$!u��8$!u��!�                       �      �      & u ��H$u��@$!u��8$!u��!��      )       X)      d       Yg      m       Xm      �       Y                 �      �       0��      �       Z                                6       Y6      _       Q_      d       Yg      m       Ym      �       Q                                     R      9       r�9      >       p u "#�>      >       R>      d       r�g      m       r�                        #      9       PU      X       p x !�X      d       Pg      �       P                  @      L       UL      �       u�                  L      �      & u ��H$u��@$!u��8$!u��!�                           L      L      & u ��H$u��@$!u��8$!u��!�L      �       [�      �       Q�      �       X�      �       Q�      �       X�      �       [                 L      L       0�L      �       Z                          X      �       X�      �       Q�      �       X�      �       Q�      �       Q                          e      e       Qe      z       q�z      �       q��      �       x 2$����u "#��      �       R�      �       r��      �       q 2$����u "#��      �       q 2$����u "#��      �       q 2$����u "#�                      z      �      	 p ������      �      	 p ������      �      	 p �����                    ~      �       q����      �       x 2$����u "#���                         y      Gy       UGy      }       ��}      (}       U(}      2}       ��                         y      Gy       TGy      �|       S�|      �|       �T��|      2}       S                            Gy      Gy       ��#�Gy      jy       ��#�jy      �y       _�y      �y       ��y      z       x�z      &z       |�&z      �z       _�z      C{       ��[|      r|       _�|      �|       _�|      }       _                    jy      �y       T�y      }       ��                 jy      �y       \                  �y      �y       0�                              �y      �y       1��y      �y       ���y      �y       P�y      [z       ��[z      mz       Pmz      �|       ���|      }       ��                        �y      �y       \z      �z       \[|      r|       \}      }       \                        �y      �y       ]&z      iz       ]iz      qz       ^[|      r|       ]                            �y      �y       ��+z      =z       P=z      �{       ��[|      l|       Pl|      r|       ���|      }       ��                               iz      zz       ]zz      �z       ^�z      �z       }��z      �z      
 ~ 2$v "#��z      �z      
 ~2$v "#��z      �z      
 ~ 2$v "#��z      '{      
 ~ 2$v "#�'{      2{      
 ~2$v "#��|      }       ^}      }       ]                        �z      �z       U�z      C{       w �|      �|       U�|      }       w                         �z      �z       0��z      '{       ^'{      ,{       ~�,{      C{       ^�|      }       0�                      iz      �z       0��z      #{       _,{      ;{       _�|      }       0�                    �z      �z       \�z      C{       \                   �z      �z       ~ 2$v "#����z      {       ~ 2$v "#���                          Q{      ^{       ]^{      �{       \�{      �{       |��{      |       |~�|      [|       \r|      �|       \�|      �|       \�|      �|       ]                          ~{      �{       T�{      [|       w r|      �|       w �|      �|       T�|      �|       w                             �{      �{       0��{      [|       ^r|      �|       ^�|      �|       ~��|      �|       ^�|      �|       0�                       Q{      �{       0��{      [|       _r|      �|       _�|      �|       0�                      �{      �{       Q|      0|       Q0|      ?|       ��                   �{      �{       } �8$v �!
���|      [|       } �8$v �!
���                  �      �       T�      �       t�                        p2      �2       U�2      �2       �U��2      �2       U�2      �2       S                          p2      �2       T�2      �2       �T��2      �2       T�2      �2       R�2      �2       V                          p2      �2       Q�2      �2       �Q��2      �2       Q�2      �2       Z�2      �2       �Q�                    y2      �2       P�2      �2       P                        �A      B       UB      B       SB      B       �U�B      !B       U                    �A      B       PB      !B       P                    �      �       p��      �       u#�                    �      �       U�      �       �U�                    �      �       T�      �       t                               �             U      %       V%      +       U+      /       V/      6       �U�6      \       U\      |       V|      �       U                          �      �       T�      /       ]/      6       �T�6      O       TO      �       ]                      �             Q      6       �Q�6      `       Q`      �       �Q�                         �             0�+      /       P6      U       0�U      d      & t��H$t	��@$!t
��8$!t��!�n      |       P�      �       P                          �      �       s��      �       t��      �       T�      �       t��             t�6      O       s�O      |       t�                    �            & s��H$s��@$!s��8$!s��!�6      d      & s��H$s��@$!s��8$!s��!�                     �      �       t �             [6      |       [                      �      �      & t ��H$t��@$!t��8$!t��!��            & t ��H$t��@$!t��8$!t��!�O      d      & t ��H$t��@$!t��8$!t��!�                           �      �       	���      �      & t��H$t��@$!t��8$!t��!��      �       	���            & t��H$t��@$!t��8$!t��!�6      O       	��O      d      & t��H$t��@$!t��8$!t��!�                         �      �      & s��H$s��@$!s��8$!s��!��      �       Y�      �       R�             YO      |       Y                     �      �       0��             ZO      |       Z                          �      �      & s��H$s��@$!s��8$!s��!��      �       R�      �      & s��H$s��@$!s��8$!s��!��             R6      O      & s��H$s��@$!s��8$!s��!�O      |       R                  �             u `      |       Q                        �             U      %       V%      +       U+      /       V`      |       V|      �       U                 �      u       u                      !      0       r�0      5       r|�5      5       R5      @       r�@      m       r�                          !      0      + r �H0H%�$!0)( 8/�������0      5      + rt�H0H%�$!0)( 8/�������@      B      	 p �����B      P       PP      d      + r �H0H%�$!0)( 8/�������                      !      5       PD      P      	 q �����P      m       P                      !      0      , r��H$r	��@$!r
��8$!r��!�����0      5      , r|��H$r}��@$!r~��8$!r��!�����J      d      , r��H$r	��@$!r
��8$!r��!�����                  
      m       T                 
      m       Y                     !      0      & r��H$r	��@$!r
��8$!r��!�0      5      & r|��H$r}��@$!r~��8$!r��!�N      d      & r��H$r	��@$!r
��8$!r��!�                          �w      x       Ux      _x       V_x      �x       �U��x      y       Uy      y       V                          �w      x       Tx      �x       _�x      �x       �T��x      y       Ty      y       _                    x      x       v�x      x       v�x      x       v�x      �x       ]�x      �x       }��x      �x       }x��x      �x       }|��x      �x       ]                      x      7x       P7x      :x       p�:x      Ox      + v�H0H%�$!0)( 8/�������                      x      Ox       ROx      �x       w �x      �x       ��                      Px      _x       0�_x      �x       ^�x      �x       ~��x      �x       ^                    _x      �x       V�x      �x       V                    _x      �x       S�x      �x       S                 �x      �x      , }��H$}	��@$!}
��8$!}��!�����                        Px      _x       0��x      �x       S�x      �x       Q�x      �x       ���x      �x       S                  �      �       T�      �       t�                    �      �       p��      �       u#�                    �      �       U�      �       �U�                    �      �       T�      �       t                               `      �       U�             V             U             V             �U�      3       U3      q       Vq      �       U                          `      �       T�             ]             �T�      /       T/      �       ]                      `      �       Q�             �Q�      U       QU      �       �Q�                        `      �       0�             P      J       0�J      q       P{      �       P                           l      �       s��      �       t��      �       T�      �       t��      �       t�      /       s�/      6       t�6      q       r 1$r "2$����s "#�                    s      �      & s��H$s��@$!s��8$!s��!�      Y      & s��H$s��@$!s��8$!s��!�                     s      �       t �      �       [      q       [                        �      �      & t ��H$t��@$!t��8$!t��!��      �      & t ��H$t��@$!t��8$!t��!�/      6      & t ��H$t��@$!t��8$!t��!�6      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                                   �       	���      �      & t��H$t��@$!t��8$!t��!��      �       	���      �      & t��H$t��@$!t��8$!t��!�      /       	��/      6      & t��H$t��@$!t��8$!t��!�6      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                  >      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                         �      �      & s��H$s��@$!s��8$!s��!��      �       Y�      �       R�      �       Y/      q       Y                     �      �       0��      �       Z/      q       Z                                �      & s��H$s��@$!s��8$!s��!��      �       R�      �      & s��H$s��@$!s��8$!s��!��      �       R      /      & s��H$s��@$!s��8$!s��!�/      q       R                  �      �       u U      q       Q                        �      �       U�             V             U             VU      q       Vq      �       U                   P      d       u 4      =       u                      �      �       Y�      �       y��              y�       )       y|�=      Y       y�                    �      )       X=      Y       X                    �      )       R=      Y       R                    �      )       \=      N       \                         l      �       P�      �       P�      �       Q�             P             Q      4       P=      Y       P                   l      4       [=      Y       [                        �      �       q p "��      �       ]�      �       0��             ]             0�                          pv      �v       U�v      �v       V�v      �w       �U��w      �w       U�w      �w       V                          pv      �v       T�v      �w       ^�w      �w       �T��w      �w       T�w      �w       ^                    �v      �v       v��v      �v       v��v      �v       v��v      [w       \[w      hw       |�hw      tw       |x�tw      ww       ||�ww      �w       \                      �v      �v       P�v      �v       p��v      �v      + v�H0H%�$!0)( 8/�������                      �v      �v       R�v      �w       w �w      �w       ��                    �v      �v       0��v      �w       ]                    �v      [w       _tw      �w       _                      �v      [w      	 v �����ww      �w       X�w      �w       ��                 ww      �w      , |��H$|	��@$!|
��8$!|��!�����                       �v      �v       0�Nw      [w       X[w      �w       Q�w      �w       ��                     !w      )w       v s �)w      <w       T<w      Nw       v  �                  0      4       T4      F       t�                                 p�      )       u#�                    `      q       Uq             �U�                      d      w       Pw      �       yl��             �U#                    �      �       Q�             Q                                         d      �       0��      �      
 y z !
����      �       z 
����      �       0��      �      
 u p !
����      �       p 
����      �       0��      �       P�      �       p 
����      �       p 
����             P             0�             z 
���                             d      d       p�d      w       p�w      y       y|�y      �       Y�      �       R�      �       R�             R             Y             R                              �      �       Z�      �       q u ��      �      � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/����      �      � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/����            � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/���             Z             q u �                           1       T1      S       �T�                    $      A       RA      S       u                 $      R       0�                   $      $       r�$      +       r�+      A       r�A      R       R                    +      A      & r��H$r��@$!r��8$!r��!�A      S      2 u#��H$u#��@$!u#��8$!u#��!�                   +      A      & r��H$r��@$!r��8$!r��!�A      S      2 u#��H$u#��@$!u#��8$!u#��!�                      1      <       T<      A      ) �Tr�H0H%�$!0)( 8/���A      R      , �Tu#�H0H%�$!0)( 8/���                            �u      �u       U�u      v       ]v      v       �U�v      Rv       ]Rv      `v       U`v      jv       ]                            �u      �u       T�u      v       \v      v       �T�v      Rv       \Rv      ]v       T]v      jv       \                         �u      �u       u��u      �u       }��u      �u       }��u      �u       }��u      v       }�v      Rv       SRv      `v       u�`v      jv       }�                      �u      �u       P�u      �u       p��u      �u      + }�H0H%�$!0)( 8/�������                        �u      v       Vv      -v       V-v      1v       v�1v      Rv       V                        v      ,v       s~��8$s��!
���7v      ;v       s~��8$s��!
���;v      >v       p 8$s��!
���>v      Rv       s~��8$s��!
���                                 p�             u#�                             I       UI      �       �U��      �       U                          1       u �      �       u                                   �       0��      �       Q�      �       0��      �       Q�      �       0��      �       Q                               i       Ql      �       Q�      �       Q�      �       Q�      �       t �#�                                          �       0��      �       r x "��      �       P�      �       0��      �       p u ��      �       P�      �       P�      �       0��      �       P�      �       0��      �       P                          I       X�      �       X                                      x�� �      $       x�� �$      I       YI      [       y�[      a       yx�a      f       y|�f      �       Y�      �       x�� ��      �       Y                          1      . x�� ��H$x�� ��@$!x�� ��8$!x�� ��!��      �      . x�� ��H$x�� ��@$!x�� ��8$!x�� ��!�                    l      �      & y��H$y	��@$!y
��8$!y��!��      �      & y��H$y	��@$!y
��8$!y��!�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       R�      �       �U#                       �      �       r�� ��      �       P�      �       p��      �       px��      �       p|��      �       P�      �       P                  �      �      . r�� ��H$r�� ��@$!r�� ��8$!r�� ��!�                     �      �      & p��H$p	��@$!p
��8$!p��!��      �      & p��H$p	��@$!p
��8$!p��!��      �      & p��H$p	��@$!p
��8$!p��!�                               s      (s       U(s      �s       S�s      rt       vt�rt      �t       S�t      �t       vt��t      gu       �U�gu      �u       S                             s      (s       T(s      �t       ]�t      �t       �T��t      gu       ]gu      uu       Tuu      �u       ]                                 s      (s       u�(s      (s       s�(s      Zs       s�Zs      Zs       v�� �Zs      �s       _�s      �s       ��s      �s       x��s      �s       |��s      rt       _rt      �t       s��t      �t       _�t      gu       _gu      �u       s��u      �u       _                          Zs      rt       V�t      �t       V�t      �t       �U#��t      gu       V�u      �u       V                    4s      Gs      & s��H$s��@$!s��8$!s��!�rt      �t      & s��H$s��@$!s��8$!s��!�                    es      �s      . s�� ��H$s�� ��@$!s�� ��8$!s�� ��!��u      �u      . s�� ��H$s�� ��@$!s�� ��8$!s�� ��!�                            ts      �s       0��s      rt       w �t      �t       w �t      �t       P�t      gu       w �u      �u       0�                               t      At       SAt      Ht       QHt      rt       S�t      �t       Su      u       Su      u       Qu      Ku       S                   �s      �s      & ��H$	��@$!
��8$!��!��t      �t      & ��H$	��@$!
��8$!��!�                        t       t       R�t      u       RKu      `u       R`u      gu       ��                          ts      �s       0��s      �s       Q�t      �t       Q�t      �t       ���u      �u       0�                          t      Ht       s @%�Ht      Rt       s @%�Rt      Zt       RZt      rt       s @%��t      �t       s @%�                         t      Ht       s 
���Ht      rt       s 
����t      �t       s 
���u      u       s 
���u      Ku       s 
���                          �s      t       Rt      t       ��t       t       ~ s ��t      u       ~ s �Ku      gu       ~ s �                  d      �       r�                    �      �       U�      X       �U�                         �      �       u�      �       Y�      N       �U#N      R       YR      X       �U#                         �      8       0�8      ;       Q;      K       0�K      N       QN      X       0�                          �      �       Q�      �       t �#��      8       Q;      P       QP      R      # t �#u t �#����u ����*( �R      X       Q                                         �      �       0��             
 z y !
���              y 
���             0�      "      
 u p !
���"      ,       p 
���,      8       0�8      ;       P;      B       p 
���C      K       p 
���K      N       PN      R       0�R      X       y 
���                               �      �       u#��      �       u#��      �       u#
��      �       y
��      �       Z�      8       R;      B       RC      N       RN      R       ZR      X       R                           �      �       u#��8$u#��!
����      �       y��8$y��!
����      :      " �U##��8$�U##��!
���;      M      " �U##��8$�U##��!
���N      R       y��8$y��!
���R      X      " �U##��8$�U##��!
���                           �      �       u#��8$u#	��!
����      �       y��8$y	��!
����      :      " �U##��8$�U##	��!
���;      M      " �U##��8$�U##	��!
���N      R       y��8$y	��!
���R      X      " �U##��8$�U##	��!
���                      �      8       [;      B       [C      X       [                    @      \       T\      �       �T�                    D      w       Rw      �       u                 D      �       0�                   D      D       r�D      D       r�D      w       r
�w      �       R                       D      H       r��8$r��!
���H      K       p 8$r��!
���K      w       r��8$r��!
���w      �       u#��8$u#��!
���                         D      W       r��8$r	��!
���W      b       q 8$r	��!
���b      e       p 8$r	��!
���e      w       r��8$r	��!
���w      �       u#��8$u#	��!
���                  \      r       T                              r      /r       U/r      �r       \�r      �r       sv��r      �r       �U��r      �r       \�r      �r       U�r      �r       \                            r      /r       T/r      �r       V�r      �r       �T��r      �r       V�r      �r       T�r      �r       V                     /r      /r       |�/r      Lr       |�Lr      Lr       |�Lr      �r       |
��r      �r       S�r      �r       |
�                    Lr      rr       p 
���rr      vr       P                    er      �r       ^�r      �r       ^                        �r      �r       s~��8$s��!
����r      �r       s~��8$s��!
����r      �r       p 8$s��!
����r      �r       s~��8$s��!
���                        4       r�                        �      �       U�      �       �U��             U      
       �U�                      �      �       T�      �       t �             t                             �
      �
       U�
      �       ���      �       U�      �       ���             �U�      �       ��                            �
      �
       T�
      �       ���      �       T�      �       ���             �T�      �       ��                        �
      �
       Q�
      �       �Q��      �       Q�      �       �Q�                 �
      �
       u                  �
      �
       u #�u #�"�                  �
      �
      
 | 
��	��                                                       �
             Z<      K       Z�      �       Z      �       Z�             ZW      �       [�      �       { 
����      �       [�             ��R      �       Z�      �       [�      �       ���      N       ZN      �       [�      �       Q�      �       [             ��      !       Z:      d       Zz      �       Z                                                               �
      �
       
����
             [      )       
���)      V       [�      �       
����      �       [      �       [�             [      W       ]W      �       ^�             ^      E       ��E      �       [�      �       
���H      �       [�      �       ^N      �       ^�      �       ^�             ��             ^      !       [!      :       ]N      Y       [Y      d       
���d      z       ]                                             �      �       ��s      w       Vw      �       ���      �       0��             ��W      �       \�      �       z 
����             \�      �       0�H      d       ��d      �       0��      �       \N      �       \�      �       \             \N      d       0�                                               �      �       ��d      o       Vo      �       ���      �       1��             ��W      �       U�      �      	 u 0$0&��             Ud      h       Rh      �       ���      �       ��H      �       ���      �       UN      �       U�      �       U             UN      d       1�                           �
      �
       P�
      D       YD      I       T�      �       P             Y�             TH      d       T                      �
      �
       0��
      I       V�      �       0�      <       V                                                         �
      �
       P�
             T             ��~      q       T�      �       P�      �       T      �       T�             T      �       Y�      �       T�             Y      �       T�      �       Y�      G       XG      :       Y:      d       Td      z       Yz      �       X�      �       Y�      �       X�      �       Y                          �
      �
       P�
      �       ��~�      �       P�      �       ��~      �       ��~                          �
      �
       t �
      �       S�      �       S      C       SH      G       SI      �       S                                                  �
      I       0�K      �       V�      �       p,�      �       V�      �       0��      �       V      �       0��      �       V�      �       0��      �      
 p q !
����      �       p 
����      �      $ s z 1$r "������"#��q !
����      �       V�      �      * s z 1$r "������"#��q !���"
����      �       0��             V             0�      !       p 
���!      �       0��      �       V                                                                                          �
      �
       r��
             P             P      )       t 1$����r "#�)      I       P�      �       r��      �       ^      1       P1      9       t 1$����r "q "#�9      I       PI      d       t 1$����r "q " "#�d      �       ^�             ^      +       ��+      W       VW      j       Pj      �       V�      �       P�      �       v q "��      �       P�      �      	 v q " "��             P      ,       PR      k       Pp      �       R�      �       ���      �       P�      �       s z 1$r "������"��      �       ^�      H       ��H      �       ^�      �       V�      �       P�      �       ���      N       P�      �       P�      �       P�             P      !       s z 1$r "������"�!      N       ��N      d       ^d      z       ��z      �       P�      �       ��                                                                  W       TW      �       x��      �       X�      �       x��             x�      �       X�      �       x��      A       YA      N       UN      �       Z�      �       X�      �       Z�             X             x�!      :       Td      z       Tz      �       Y�      �       u��      �       x��      �       Y�      �       p��      �       x�                        B             ^      �       Z�             ^�      �       Z                           W       ��W      �       P�             ���      �       P                       �             ��N      }       ^}      �       R�      �       ^                                             u 
���              U       -       ^-      }       [}      �       Q�      �       [z      ~       U~      �       ^�      �       ��                  V      �       ���      �       ��                    �             U      |
       �U�                    �             T      |
       ��                            �      �       Q�      c	       _c	      d	       �Q�d	      t	       _t	      u	       �Q�u	      |
       _                 �      �       u                  �      �       u #�u #�"�                    d      Y	       Vu	      |
       V                    \      Y	       [u	      |
       [                       �      )	       t 
���K	      R	       t 
���u	      M
       t 
���b
      |
       t 
���                       �      )	      ( q 1$��"��8$q 1$��"#��!0$0&�K	      R	      ( q 1$��"��8$q 1$��"#��!0$0&�u	      M
      ( q 1$��"��8$q 1$��"#��!0$0&�b
      |
      ( q 1$��"��8$q 1$��"#��!0$0&�                             -      2       0�2      )	       Q)	      C	       q�K	      R	       Qu	      :
       Q:
      M
       q�b
      |
       Q                       �      �       q 1%��      �       P�             q 1%�      (       t 1%�                         �      �       t �      Y	       Rd	      
       R
      u
       Rw
      |
       R                                             �      �       0��      	       P	      R	       0�R	      Y	       Pd	      �	       0��	      �	      
 x } !
����	      �	       x 
����	      �	      " r v 1$| "����z "#��} !
����	      �	       P�	      �	       0��	      �	       P�	      
       0�
      "
       P'
      R
       0�R
      b
       Pb
      |
       0�                  �             ~�      2       ~�                  -      2       U                      �	      �	       P�	      �	       r v 1$| "����z "�
      '
       r v 1$| "����z "�                                     l      %l       U%l      �m       _�m      �p       ��~�p      �p       _�p      �p       �U��p      �p       ��~�p      Bq       _Bq      Pq       UPq      Zq       _Zq      sq       ��~sq      	r       _                                   l      %l       T%l      �m       ^�m      �p       �T��p      �p       ^�p      �p       �T��p      Bq       ^Bq      Mq       TMq      Zq       ^Zq      sq       �T�sq      	r       ^                                                %l      %l       �%l      dl       �dl      dl       �dl      �l       �Cm      [m       R�m      �m       v~��m      An       S]n      kn       Vkn      �n       X�n      o       ��o      Yo       v~�Yo      �o       S�o      9p       ^9p      �p       v~��p      �p       S�p      �p       R�p      �p       |����1$���� "#��p      �p       ��p      �p       ��p      q       �Zq      sq       v~��q      	r       �                                 :l      @l       s 
���@l      Xl       S[l      �m       S�m      �p       ���p      �p       S�p      �p       ���p      Bq       SZq      sq       ��sq      r       S                           m      �m       ��m      �p       ��~#��p      �p       ��p      �p       �U#��p      �p       ��~#��p      �p       �Zq      sq       ��~#�                      m      m       Qm      �p       ��~Zq      sq       ��~                    #m      �m       V�p      �p       V�p      �p       V                      #m      Km       QKm      �p       ��~Zq      sq       ��~                      +m      /m       P/m      �p       ��Zq      sq       ��                      |l      �l       V�l      �l       v 1%�q      &q       V&q      Bq       \                               l      �m       0��m      Ep       ��Jp      �p       ���p      �p       0��p      �p       ���p      Zq       0�Zq      sq       ��sq      	r       0�                            �l      �l       R�l      m       Qsq      �q       Q�q      �q       R�q      �q       ��~�q      �q       Q                     �l      �l       y �8$x �!
����q      �q       y �8$x �!
����q      �q       ��~��8$��~��!
���                    �l      �l       } 
����l      �l      	 } 
��1%��q      �q       } 
����q      �q      	 } 
��1%�                          �m      Zn       ]Zn      ]n       [�n      �p       ]�p      �p       ]Zq      sq       ]                                �m      n        
����n      �n       P�n      o       ��o      5o        
���Yo      ko        
���9p      �p        
����p      �p        
���Zq      cq        
���                           �m      �m       s 
����n      �n       R�n      o       ��o      Yo       s 
���9p      �p       s 
���Zq      sq       s 
���                                   [m      �m       0��m      �m       \�m      �m       Y�m      An       \An      ]n       |�]n      9p       \9p      sp       Ysp      �p       \�p      �p       0��p      �p       \Zq      sq       \                        [m      �m       0�An      Zn       ]Zn      �n       [�n      o       ���p      �p       0�                        [m      �m       0�An      ]n       P]n      �n       Z�n      o       ���p      �p       0�                               �m      An       ��~��8$��~��!0$0&��n      �n       | 1$��~"��8$t �!0$0&��n      �n      ( | 1$��~"��8$| 1$��~"#��!0$0&��n      Ao       ��~��8$��~��!0$0&�Yo      �o       ��~��8$��~��!0$0&�9p      �p       ��~��8$��~��!0$0&��p      �p       ��~��8$��~��!0$0&�Zq      sq       ��~��8$��~��!0$0&�                           [m      �m       ��~�m      ]n       ��~#�]n      ]n       ��~]n      �p       ��~#��p      �p       ��~�p      �p       ��~#�Zq      sq       ��~#�                           [m      �m       ��m      ]n       ��~#�]n      �n       ��~#��n      �p       ��~#��p      �p       ��p      �p       ��~#�Zq      sq       ��~#�                           [m      �m       ��~�m      ]n       ��~#�]n      �n       ��~�n      �p       ��~#��p      �p       ��~�p      �p       ��~#�Zq      sq       ��~#�                             [m      An       VAn      kn       Vkn      �n       X�n      �o       V�o      9p       ��~9p      �p       V�p      �p       VZq      sq       V                  �o      �o       ]                       p      p      
 p r !
���p      p       p 
���p      p       p 
��s "
���p      p       ~��r !
��s "
���                                  @             U      �       _�      �       U�             _      	       �U�	      $       U$      �       _�      �       �U��      �       _                 @      B       u                  @      B       u #�u #�"�                                        �       S�             (      	       �U#($      W       SY      w       Sw      �       (�      �       �U#(�      �       S�      �       S                                       �       � �      �       u� �      �       Q�             �       	       �U#H$      2       Q2      �       � �      �       �U#H�      �       �                               �       T�      �       <�      	       T$      �       T                             �       � �      �       u� �      	       U$      �       U                  �      	       Q                        �      �      
 p r !
����      �       p 
����      �       q��r !
����      	       P                     2      2       Q2      Y       0�j      �       Q�      �       0�                          U       TU      7       T                        7       Y                                        B      ^       Pf      u       Pu      }       t 1$����y "#�}      �       P�      �       t 1$����y "{ "#��      �       P�      �       t 1$����y "r "{ "#��      �       P�      �       r 1$t 1$����"y "{ "#��             P             r 1$t 1$����"y "{ "#�             P      $       r 1$t1$����"y "{ "#�$      /       P/      1       r 1$t 1$����"y "{ "#�                       7       X                        B      ^       q 
����      �       q 
����      �       0��             q 
���      1       q 
���                 �      �       u                  �      �       u #�u #�"�                 �             t�                  �      �       r�                    P      f       Uf      �       �U�                    P      f       Tf      �       Z                  Y      �       Y                         Y      �       0��      �       P�      s       0�s      {       P{      �       0�                     Y      �       0��      �       T�      �       0�                                ]      v       X�      �       X�      �       x���      �       X�      �       X�      �       x��      �       X�      �       
 �T      �       T                        q      �       P�      �       P�      T       P�      �       P                       v      v       Pv      v       p�v      v       p�v      �       p��      7       p�7      �       R�      �       p��      �       R                     v      �       p ��8$p��!
����      T       p ��8$p��!
����      �       p ��8$p��!
���                     v      �       p��8$p��!
����      T       p��8$p��!
����      �       p��8$p��!
���                     v      �       p��8$p��!0$0&��      T       p��8$p��!0$0&��      �       p��8$p��!0$0&�                            �      �      
 q r !
����      �       q 
����             q 
���      T       p��p��8$!
����      �       q 
����      �       p��p��8$!
���                     �      �       x ���             x ���      �       x ��                  �      �       U                      i      l      
 p q !
���l      p       p 
���p      �       r��q !
���                    �      �       U�      C       �U�                      �      �       T�      �       X�      C       �T�                   �      �       u�      �       U                     �      <       0�<      =       P=      C       0�                      �      �       P�              Q=      B       Q                     �      �       Q�      �       q��      �       q��             q�      =       U=      B       q�                          �      )       X)      ,      
 q r !
���,      9       q 
���9      =       u��r !
���=      B       X                         �      �       q ��8$q��!
����      �       t 8$q��!
����      �       u 8$q��!
����              q ��8$q��!
���=      B       q ��8$q��!
���                         �      �       q��8$q��!
����      �       t 8$q��!
����      �       u 8$q��!
����              q��8$q��!
���=      B       q��8$q��!
���                     �              q��8$q��!0$0&�       5       t �8$y �!0$0&�=      B       q��8$q��!0$0&�                    �             R=      B       R                      P      g       Ug      �       u�{��      �       �U�                      P      n       Tn      �       �T��      �       T                     Z      n       t ��n      �       �T���      �       t ��                         Z      j       t 8%�j      x       Rx      �       �T8%��      �       R�      �       t 8%�                        `      q       Qq      �       T�      �       Q�      �       t 8%1$����u "
 �                  g      �       U                   l      �       U�      �       P                                  �i      �i       U�i      �i       ]�i      +j       }�{�+j      :j       ]:j      Bj       }�{�Bj      �k       �U��k      �k       U�k      �k       ]�k      �k       �U�                            �i      �i       T�i      Ak       ^Ak      Dk       �T�Dk      �k       ^�k      �k       T�k      �k       ^                               �i      �i       }��i      �i       }��i      +j       S+j      :j       }�:j      `j       S`j      fj       ]fj      fj       Sfj      fj       s�fj      uj       s�uj      uj       s�uj      ?k       ]Dk      gk       ]gk      �k       V�k      �k       S                        �i      �i       p 
����i      �i       | 
���+j      7j       p 
���7j      :j       | 
���                           �i      �i       0�`j      fj       Pfj      *k       _*k      9k       P9k      Ck       �Dk      �k       _                         �i      �i       0��i      +j       \:j      =k       \Dk      �k       \�k      �k       \                          �i      �i       S�i      +j       }�|�:j      Bj       }�|�Bj      �k       �U#��k      �k       �U#�                   :j      `j       S�k      �k       S                          Nj      Rj       PRj      [j       R[j      �k       ���k      �k       R�k      �k       ��                            �i      �i       V�i      �i       v 3%��i      �i       Pj      +j       V:j      Fj       PFj      `j       v 3%��k      �k       v 3%�                 fj      �j       s ��8$s��!
���                        uj      xj      
 t p !
���xj      �j       p 
����j      &k       v 
���Dk      Vk       v 
���                 uj      �j       s��8$s��!
���                     uj      �j       s��8$s��!0$0&��j      &k       ����8$w ��!0$0&�Dk      gk       ����8$w ��!0$0&�                  �j      
k       T                  Lk      gk       X                        �k      �k      
 p t !
����k      �k       p 
����k      �k       p 
��q "
����k      �k       v��t !
��q "
����k      �k       v��v~��8$!
��q "
���                  $      D       r�                 �      �       u�             u#�                      �      �       X�             R             0�                 �             0�                       �      �       0��      �       P�             0�             P                 �      �       u                            @)      �)       U�)      [*       ][*      `*       �U�`*      +       ]+      Y+       UY+      "-       ]                            @)      w)       Tw)      W*       VW*      `*       �T�`*      +       V+      C+       TC+      "-       V                            @)      �)       Q�)      Y*       \Y*      `*       �Q�`*      +       \+      7+       Q7+      "-       \                           @)      �)       u�
��)      [*       }�
�[*      `*       �U#�
�`*      +       }�
�+      Y+       u�
�Y+      "-       }�
�                      ^)      N*       _`*      p*       _+      �,       _                           ^)      �)       0��)      N*       6�`*      +       6�+      �,       0��,      �,       8��,      �,       6��,      �,       0��,      -       6�-      -       0�-      -       6�-      "-       0�                         �)      �)       }�
#��)      *       Q*      *       q�*      "*       q~�"*      H*       Q`*      +       S�,      "-       S                   �)      �)       }�
`*      g*       P                     �)      �)       r s "#��)      �)      
 s ��"#�*      H*       S                        �)      �)       P�)      H*       ^`*      +       ^�,      "-       ^                       �)      �)       x 8$��#	��!
����)      "*       ��#��8$��#	��!
���"*      ;*       r 
���;*      H*       ��#��8$��#	��!
���                      �)      *       P6*      >*       P`*      g*       P                        *      �*       y 
����*      �*      
 ���
����,      �,       y 
���-      "-       y 
���                  �*      �*      & s ��H$s��@$!s��8$!s��!�                 �*      �*      & s��H$s��@$!s��8$!s	��!�                    U+      Y+       QY+      j,       ��o,      �,       ��                    U+      Y+       UY+      j,       ]o,      �,       ]                 U+      j,       ^o,      �,       ^                     Z+      }+       P~+      �+       Pj,      j,       0��,      �,       8�                  �+      �+       R�+      �+       r��+      �+       r��+      #,       r�#,      @,       Q@,      X,       q|�X,      j,       Q                 �+      ,       r ��8$r��!
���                   �+      �+       y 
����+      j,       T                  �+      ,,       P                 #,      1,       T                #,      j,       U                       1,      <,       q��8$q��!
���<,      @,       p 8$q��!
���@,      C,       p 8$q��!
���C,      ],       q~��8$q��!
���                          @?      q?       Uq?      A       SA      A       �U�A      �A       S�A      �A       U                    ^?      A       VA      �A       V                   ^?      A       \A      �A       \                 @      @       U                   �?      �?       SA      cA       S                     �?      A       s�
�A      A       �U#�
�A      �A       s�
�                 A      5A       s�                 �?      �?       S                 �?      �?       s�                                                          �]      \^       U\^      >_       V>_      D_       TD_      b       �U�b      �b       V�b      Lc       �U�Lc      sc       Vsc      �c       U�c      �c       V�c      !d       U!d      Gd       �U�Gd      �d       V�d      tg       �U�tg      g       Ug      �h       �U��h      �h       V�h      i       �U�i      #i       V#i      Vi       �U�Vi      ci       Uci      ui       V                                        �]      Y^       TY^      b       ]b      b       �T�b      sc       ]sc      �c       T�c      �c       ]�c      !d       T!d      tg       ]tg      g       Tg      Vi       ]Vi      `i       T`i      ui       ]                        �]      ^       Q^      tg       �Q�tg      g       Qg      ui       �Q�                        �]      ^       R^      tg       �R�tg      g       Rg      ui       �R�                        �]      ^       X^      tg       �X�tg      g       Xg      ui       �X�                                 �^      _       P_      �`       _b      "b       P"b      Lc       _!d      �e       _cg      tg       _g      �g       _h      4h       _Uh      #i       _                       O^      q^       1��c      �c       1�i      #i       0�Vi      ui       0�                        O^      �^       0��^      �^       w Lc      Tc       0�Yc      sc       w �c      �c       0�Vi      ui       0�                      c^      q^       p  $0)��c      �c       p  $0)�pi      ui       _                       �]      ^       0�^      8^       \8^      =^       Rtg      g       0�                     �]      ^       0�^      =^       ^tg      g       0�                    �]      �a       Sb      ui       S                   �]      ^       0�tg      g       0�                          �_      �a       ]!d      Gd       ]�d      tg       ]g      h       ]4h      Uh       ]#i      Vi       ]                                    �_      �_       P�_      �`       T!d      Gd       T�d      �d       T�d      �d       0��d      �d       Pg      �g       0��g      �g       p ���g      �g       R�g      �g       p ���g      �g       }��
0$0.��                       �d      
e       0�
e      me       Tme      qe       t�cg      tg       T                     �d      
e       0�
e      �e       [cg      tg       [                    e      �e       Ucg      tg       U                  'e      Ve       X                  'e      Ve       R                   'e      )e      
 `�H     �)e      Ve       P                   'e      �e      
 �H     �cg      tg      
 �H     �                      �e      Yf       ^Yf      cg       ��~4h      Hh       ^                      �e      �e       P�e      cg       w 4h      Hh       P                           �e      �e       V�e      �e       }��e      ef       Vef      cg       ��~4h      Ch       VCh      Hh       }�                       �e      �e       }��e      gf       \gf      cg       ��~4h      Hh       }�                           �e       f       0� f      $f       P$f      7g       ��~7g      Rg       PRg      cg       }�
4h      Hh       0�                      gf      sf       ~�sf      g       ^g      cg       ~�                      gf      �f       ��~�f      g       Pg      cg       ��~                  wf      �f       ��~�����5$| "�                     P`      �`       ]!d      Gd       ]�d      �d       ]                      P`      �`       fylg�!d      Gd       fylg��d      �d       fylg�                   P`      e`       Pe`      �`       Q                      W`      �`       R!d      Gd       R�d      �d       R                  �`      �`       Q                 �`      �`       ]                 �`      �`       2FFC�                   �`      �`       P!d      Gd       P                 �`      �`       R                       �c      �c       T�c      !d       TVi      `i       T`i      ui       ]                      �c      �c       fylg��c      !d       fylg�Vi      ui       fylg�                   �c      �c       R�c      �c       P                          �c      �c       Q�c      !d       QVi      [i       Q[i      `i       t��
��5$t�"�`i      ii       }��
��5$}�"�                    �c      �c       P�c      !d       P                  �c      !d       R                                              `�      ~�       U~�      ��       _��      ��       �U��      s�       �U�s�      ��       _��      `�       �U�`�      ��       }�ۓ      ��       }���      H�       _\�      p�       �U�7�      �       �U��      "�       �U���      
�       _
�      j�       �U���      �       �U��      ��       }�                                    `�      ��       T��      ��       ]��      s�       �T�s�      }�       T}�      ��       ]��      ��       �T���      H�       ]H�      ��       �T���      
�       ]
�      ��       �T�                        `�      ��       Q��      s�       ��~s�      ��       Q��      ��       ��~                        `�      ��       R��      s�       �R�s�      ��       R��      ��       �R�                        `�      ��       X��      s�       �X�s�      ��       X��      ��       �X�                    �      ��       8�]�      j�       :�                        ��      ��       Ss�      ��       S��      H�       S��      
�       S                                               ��      ��       ^��      ��       ��~�      s�       ��~s�      ��       ^��      ��       P��      ��       ^��      �       ��~ۓ      ��       ��~��      H�       ^\�      p�       ��~7�      �       ��~�      y�       ��~��      �       P�      
�       ^
�      j�       ��~��      ��       ��~                            }�      ��       P��      ��       Qۓ      �       P�      ��      	  
��1��      ��       P��      ��      	  
��1�                 ��      ��       }�                    ��      ��       P �      ,�       P                  -�      ;�       P                  �      �       P                        �      9�       \p�      G�       \G�      ��       ��~"�      �       \                    E�      Z�       PZ�      �       _                      c�      }�       R}�      ��       ��~R�      �       R                      ��      ȗ       Pȗ      K�       ^R�      �       ^                      ֗      �       PR�      ј       Yݘ      �       Y                                    )�      9�       0�9�      ��       VH�      W�       Vp�      ��       0���      2�       V2�      ��       ��~�      ��       V��       �       P �      �       V|�      ��       V                      0�      <�       P<�      E�       ��~R�      �       ��~                                ��      �       _�      ۓ       w H�      \�       w p�      7�       w �      �       w "�      E�       _E�      ��       w j�      ��       w                 	                   �      9�       0�9�      D�       _D�      ۓ       0�H�      \�       0�p�      ��       0���      ϔ       Pϔ      O�       _O�      R�       ZR�      ��       ��~�      �       0�"�      ��       0�                
                 �      9�       0�9�      O�       ^O�      ۓ       0�H�      \�       0�p�      ܔ       0�ܔ      ��       P��      7�       ^�      �       0�"�      ��       0�j�      ��       ^                    �      �       pp��      Ε       ��~@�                     �      R�       [R�      r�       \v�      ��       \                      ��      �       Y�      -�       \j�      t�       \                       �      O�       _O�      R�       ZR�      o�       ]o�      v�       }|�v�      ��       ]                      �      R�       0���      �       0��      2�       ]j�      y�       ]                                Ȍ      ��       ]��      �       �T��      s�       �T���      N�       �T�\�      p�       �T�7�      ��       �T��      "�       �T�
�      ]�       �T���      �       �T�                                    Ȍ      T�       _��      �       _�      @�       _��      N�       _\�      p�       _7�      ��       _�      "�       _
�      �       _�      G�       ��~��      ��       ��~Y�      a�       _                                 �      ��       P��      �       ��~�      s�       ��~��      N�       ��~\�      p�       ��~7�      ��       ��~�      "�       ��~
�      ]�       ��~��      �       ��~                        �      �       P�      >�       Q��      Ɏ       Q��      �       Q                         �      �       P�      \�       S��      �       S��      N�       S7�      ��       S                           K�      T�       ]�      ��       ]��      @�       ��~\�      p�       ]�      "�       ]
�      $�       ��~                               K�      T�       _�      @�       _\�      p�       _�      "�       _
�      �       _�      G�       ��~��      ��       ��~Y�      a�       _                            \�      T�       S�      ��       S��      @�       ��~\�      p�       S�      "�       S
�      $�       ��~                                 d�      T�       0�T�      ^�       [_�      y�       0��      	�       0�	�      �       P�      5�       [5�      ��       ��~@�      b�       0�\�      p�       0��      "�       0�                                  d�      T�       0�T�      k�       w k�      y�       0��      D�       0�D�      R�       PR�      @�       w @�      b�       0�\�      p�       0��      "�       0�
�      ]�       w ��      �       w                                   s�      ��       P��      Й       y 2$y "2$#,�Й      �       ��~52$#,��      G�       U��      ��       U��      ��       U��      ۚ       Qۚ      	�       UY�      a�       P                                        d�      :�       0�:�      >�       P>�      y�       V�      *�       0�*�      ��       V��      @�       ��~@�      K�       VK�      b�       0�\�      p�       V�      "�       V
�      $�       ��~2�      `�       P`�      Y�       Va�      �       V                                d�      T�       0�T�      y�       ^�      E�       0�E�      I�       PI�      ^�       ^^�      b�       0�\�      p�       ^�      "�       ^
�      ]�       ^��      �       ^                                   Q�      ��       V��      ��       v���      ��       v���      ��       v���      ��       v���      Ə       v�Ə      ؏       v�؏      ؏       v�؏      �       v��      �       v	��      �       v
��      �       v��      ��       v���      @�       ��~#��      "�       V
�      $�       ��~#�B�      `�       \`�      `�       ]`�      h�       }�h�      s�       }q��      �       ]I�      Y�       ]a�      k�       ]p�      z�       ]                              x�      ٙ       Rٙ      �       ��~�      G�       R��      �       R�      U�       ��~��      ל       PY�      a�       R                                    s�      ��       0���      ��       ]��      ��       }�ΐ      )�       ]x�      �       0�B�      `�       0�`�      Ҝ       ��~ߜ      �       RI�      Y�       ��~Y�      a�       0�a�      �       ��~                
             d�      T�       0��      ��       0���      ��       S��      ��       P��      ��       Sΐ      �       S\�      p�       0��      "�       0�                       `�      ۜ       \ۜ      �       |P�I�      Y�       \a�      �       \                         X�      d�       0�d�      j�       Tj�      o�       Ro�      ��       T�      "�       0�                 ��      ��       ��~�
��4$p �                          X�      d�       Pj�      j�       Pj�      l�       p 1%�l�      o�       P�      �       P�      "�       Q                         ��      Ő       \Ő      ΐ       }3$v "ΐ      @�       \
�      �       }3$v "�      $�       }3$w "                    ��      G�       T��      ��       T                    ��      ��       0���             S                 �      �       u                  �      �       t                   �      �       u #                 �      �       t #                      �A      �A       U�A      �A       S�A      �A       �U�                 �A      �A       u8                              �:      �;       U�;      �;       �U��;      �;       U�;      �;       �U��;      �<       U�<      =       �U�=      =       U                              �:      �;       T�;      �;       �T��;      �;       T�;      �;       �T��;      �<       T�<      =       �T�=      =       T                        �:      �:       Q�:      �;       V�;      �;       �Q��;      =       V                    �:      �;       \�;      =       \                           �:      �;       0��;      �;       P�;      �;       Q�;      �;       0��;      �;       Q�;      =       0�                         �:      �:       0��:      �:       Q�:      �:       q�;      z;       Q<      /<       Q^<      u<       Q                                          �:      �:       Z�:      �;       P�;      �;       z { "��;      �;       S�;      �;       P�;      �;       S�;      <       S<      J<       PJ<      V<       z x "�V<      ^<       S^<      �<       P�<      =       S=      =       P                             �:      z;       	��z;      �;       ���;      �;       [<      /<       	��/<      ^<       ��^<      u<       	��u<      �<       ��=      =       ��                       �:      �:       	���:      �;       ���;      p<       ��u<      =       ��                           �:      �:       	���:      �;       [<      *<       [*<      /<       Q/<      }<       [=      =       [                              �:      �:       	���:      h;       Su;      z;       Qz;      �;       S�;      �;       S<      M<       S^<      �<       S=      =       S                               �:      �:       	���:      �;       X�;      �;       X�;      <       X<      <       Q<      J<       X^<      �<       X=      =       X                	         �:      �:       0��:      �;       ^�;      �;       ^�;      �<       ^=      =       ^                              �;      �;       0��;      �;      
 �C     ��;      �;       ]�;      �;       0��;      <       0�/<      J<       0�J<      ^<      
 ��C     �u<      �<       0��<      =       ]=      =       0�                  �<      =       ^                    �0      �0       U�0      �1       �U�                      �0      �0       T�0      
1       P
1      �1       �T�                     �0      1       0�1      v1       Py1      �1       P                     �0      m1       So1      w1       Sy1      �1       S                    1      71       QH1      ]1       Q                          1      71       0�71      L1       r p �P1      `1       p  r "�`1      e1       r p �y1      �1       0�                      �0      1       V1      e1       To1      x1       V                    �1      �1       U�1      m2       �U�                      �1      �1       T�1      �1       P�1      m2       �T�                     �1      �1       0��1      ^2       Pc2      m2       P                      �1      P2       \Q2      b2       \c2      m2       \                    �1      2       Q*2      <2       Q                          �1      2       0�2      2       u p �/2      ?2       p  u "�?2      D2       u p �c2      m2       0�                      �1      �1       V�1      D2       RQ2      `2       V                    P&      U&       UU&      Z&       �U�                    P&      Y&       TY&      Z&       �T�                            0-      O-       UO-      Y-       SY-      ]-       �U�]-      �-       S�-      �-       �U��-      �-       S                            0-      :-       T:-      \-       \\-      ]-       �T�]-      �-       \�-      �-       �T��-      �-       \                            0-      K-       QK-      Z-       VZ-      ]-       �Q�]-      �-       V�-      �-       �Q��-      �-       V                        P-      o-       Pp-      �-       P�-      �-       6��-      �-       P                    �              U      �       �U�                      �       R       QR      h       �Q�h      �       Q                     �              0�      I       Uh      �       U                                      P             p`�      D       PD      I       p`�h      �       P                          �C      �C       U�C      D       SD      rD       �U�rD      �D       S�D      �D       �U�                        �C      �C       T�C      mD       ]mD      rD       �T�rD      �D       ]                        �C      �C       Q�C      &D       \&D      rD       �Q�rD      �D       \                        �C      �C       R�C      iD       ViD      rD       �R�rD      �D       V                        �C      �C       X�C      qD       _qD      rD       �X�rD      �D       _                          �C      �C       0��C      �C       P�C      ^D       ��rD      �D       ���D      �D       0��D      �D       P�D      �D       ��                       D      &D       ��&D      >D       ^>D      ED       ~�ED      RD       ^�D      �D       ��                   D      ^D       S�D      �D       S                     D      D       PD      &D      	 |�
����D      �D       P                          `B      �B       U�B      �B       S�B      KC       �U�KC      �C       S�C      �C       �U�                        `B      �B       T�B      BC       VBC      KC       �T�KC      �C       V                        `B      �B       Q�B      �B       _�B      KC       �Q�KC      �C       _                        `B      �B       R�B      DC       \DC      KC       �R�KC      �C       \                    `B      �B       X�B      �C       ��                           �B      �B       0��B      �B       P�B      9C       ^KC      YC       ^YC      ]C       T^C      �C       0��C      �C       ^                      �B      �B       ^�B      C       ]C      C       }�C      9C       ]�C      �C       ^                   �B      9C       S�C      �C       S                    �B      �B       Q�C      �C       Q                    �       �        U�       �        q0�                 �       �        U                        ��      �       U�      G�       VG�      V�       �U�V�      j�       U                        ��      �       T�      G�       ]G�      V�       �T�V�      j�       T                       ��      �       U�      G�       VG�      V�       �U�V�      j�       U                   �      G�       Sc�      j�       0�                   ��      �       	��V�      V�       	��V�      j�       P                  *�      :�       P                     �       �       �H� �      )�       Q)�      *�       �H�                 �      *�       S                 �      *�       V                            �        T�       �        �T�                                        P?       @        PG       H        Po       p        P                      @}      j}       Tj}      �}       �T��}      �}       T                  d}      �}       X                  d}      �}       R                  d}      �}       Q                    d}      j}       Tj}      �}       �T�                  d}      �}       U                              �}      �}       U�}      �}       �U��}      �}       U�}      �}       �U��}      �}       U�}      �}       S�}      �}       �U�                              �}      �}       T�}      �}       �T��}      �}       T�}      �}       �T��}      �}       T�}      �}       V�}      �}       �T�                         �}      �}       U�}      �}       �U��}      �}       U�}      �}       S�}      �}       �U�                    �}      �}       V�}      �}       �T�                    �}      �}       S�}      �}       �U�                  �}      �}       P                       ~      ~       U~      ~       �U�~      ?~       U                           ~      ~       T~      ~       �T�~      )~       T)~      >~       V>~      ?~       �T�                      ~      ~       U~      ~       �U�~      ?~       U                    $~      >~       V>~      ?~       �T�                  $~      ?~       U                  9~      <~       P                      @~      W~       UW~      X~       �U�X~      ~       U                          @~      W~       TW~      X~       �T�X~      i~       Ti~      ~~       V~~      ~       �T�                     @~      W~       UW~      X~       �U�X~      ~       U                    d~      ~~       V~~      ~       �T�                  d~      ~       U                  y~      |~       P                          �~      �~       U�~      �~       S�~      �~       �U��~      �~       S�~      �~       �U�                            �~      �~       T�~      �~       Q�~      �~       V�~      �~       �T��~      �~       V�~      �~       �T�                     �~      �~       P�~      �~       P�~      �~       P                    �~      �~       V�~      �~       �T�                    �~      �~       S�~      �~       �U�                  �~      �~       P                                    P�      u�       Uu�      ��       S��      ��       �U���      �       S�      �       �U��      Z�       SZ�      `�       �U�`�      u�       Su�      ��       U��      ��       S                                    P�      y�       Ty�      ��       ]��      ��       �T���      �       ]�      �       �T��      _�       ]_�      `�       �T�`�      u�       ]u�      ��       T��      ��       ]                                    P�      y�       Qy�      ��       V��      ��       �Q���      �       V�      �       �Q��      [�       V[�      `�       �Q�`�      u�       Vu�      ��       Q��      ��       V                    h�      u�       P��      ��       P                                 p�      u�       u��u�      ��       s����      ��       �U#����      �       s���      �       �U#���      Z�       s��Z�      `�       �U#��`�      u�       s����      ��       s��                            ��      ��       P��      ��       P�      �       P�      )�       P`�      g�       P��      ��       P                            a�      ��       \��      �       \�      ]�       \`�      ��       \��      ��       u���      ��       \                   ��      �       s��`�      u�       s��                  ׄ      �       U                   �      J�       s����      ��       s��                      ��      ą       Uą      Ņ       �U�Ņ      օ       U                      ��      ą       Tą      Ņ       �T�Ņ      օ       T                      ��      ą       Qą      Ņ       �Q�Ņ      օ       Q                      ��      ̆       Ŭ      ��       �U���      �       U                      ��      ̆       T̆      ��       �T���      �       T                            ��      Ɔ       QƆ      Ԇ       VԆ      ��       �Q���      ��       V��      ��       �Q���      �       Q                            ��      ̆       R̆      Ԇ       SԆ      ��       �R���      ��       S��      ��       �R���      �       R                 ��      �       ��(	                       ��      ̆       T̆      ��       �T���      �       T                     ��      ̆       Ŭ      ��       �U���      �       U                     Ȇ      ̆       R̆      Ԇ       S��      �       S                     ��      Ɔ       QƆ      Ԇ       V��      �       V                     ��      ̆       T̆      Ԇ       �T���      �       �T�                     ��      ̆       Ŭ      Ԇ       �U���      �       �U�                     І      Ԇ       P��      �       P�      �       \                          ��      	�       U	�      �       S�      �       �U��      ,�       S,�      2�       �U�                            ��      ��       T��      �       V�      �       �T��      -�       V-�      1�       U1�      2�       �T�                      ��      ��       Q��      	�       T	�      2�       �Q�                  
�      1�       P                  �      2�       �Q�                      �      -�       V-�      1�       U1�      2�       �T�                      �      ,�       S,�      1�       q�}�1�      2�       �U�                     �      #�       s��#�      1�       Q1�      2�       �U#��                            `�      �       U�      ��       S��      ��       �U���      J�       SJ�      T�       �U�T�      _�       S                                `�      q�       Tq�      �       Q�      ��       \��      ��       �T���      M�       \M�      S�       US�      T�       �T�T�      _�       \                        ��      ��       P��      ��       P��      ��       VT�      _�       P                        ��      M�       \M�      S�       US�      T�       �T�T�      _�       \                          ��      J�       SJ�      O�       }�{�O�      S�       q�{�S�      T�       �U�T�      _�       S                          ��      ��       P��      �       V�      '�       P(�      S�       PT�      _�       P                        ��      O�       ]O�      S�       QS�      T�       �U#��T�      _�       ]                              ��      ��       U��      �       \�      �       |�}��      �       �U��      /�       \/�      7�       U7�      A�       \                            ��      ��       T��      �       V�      �       �T��      /�       V/�      4�       T4�      A�       V                       ��      ��       |���      �       |��      �       |�}��      �       �U#��      /�       |�                          ӝ       p 
����      ,�       p 
���                  ڝ      �       V                    ڝ      �       \�      �       |�}�                  ߝ      �       S                     ߝ      �       0��      ��      	 s | #���      �      	 s | #��                      �      ��       P��      ��       s�����      �       P                                ��      ��       U��      ��       �U���      ߢ       Uߢ      1�       V1�      T�       UT�      P�       VP�      b�       Ub�      ��       V                      ͢      �       U�      %�       V��      Ĥ       V                  �      �       p ��                   %�      ,�       ]��      Ĥ       P                         1�      T�       UT�      ��       VĤ      P�       VP�      b�       Ub�      ��       V                    G�      ��       ^Ĥ      ��       ^                      N�      ��       SP�      ի       S��      d�       S                        g�      o�       p ����      �       p ���      5�       p ��6�      C�       p ��                         �      0�       0�0�      �       R�      ��       R
�      P�       Rի      ��       R                  x�      ��       0�                                        N�      T�       0��      5�       P5�      ��       \�      �       P�      �       ]��      Ш       _Ш      
�       ]P�      ��       0���      ��       P��      ի       \��      _�       0�_�      d�       Pd�      �       ]                                                       ?�      K�       PK�      p�       Tp�      v�       t�v�      ��       T��      ��       S��      �       P�      >�       S>�      W�       s�W�      a�       Za�      v�       s��      (�       s�(�      X�       SX�      c�       s�c�      ��       S��      ��       s���      Ħ       SĦ      Ϧ       s�Ϧ      �       S�      �       S�      '�       s�'�      1�       S˨      Ш       Se�      e�       Te�      i�       t�i�      m�       ti�x�      ��       P��      ��       T��      ��       t�                      ��      �       \��      Ш       \�      ��       \                      ��      ף       T��      ��       T��      ��       p                 ף      �       p                 K�      ��       R                        Ф      �       \�      ��       \
�      P�       \ի      ��       \                            4�      f�       Qj�      ��       Q��      Ҧ       QҦ      �       P�      ��       Y�      1�       Y                        K�      W�       s�W�      a�       Za�      v�       s��      (�       s�                    K�      j�       P�      (�       P                                             K�      W�       s�W�      ��       Z��      ��       [��      ĥ       {�ĥ      ӥ       [�      �       Z�      �       Y�      �       s��      (�       s�1�      1�       [1�      R�       ZR�      [�       P[�      _�       S_�      n�       Pn�      ��       Z
�      
�       Y
�      P�       Zի      ��       Z                                g�      v�       Tv�      ��       S��      ӥ       Qإ      �       S1�      P�       Sn�      ��       S
�      B�       Sի      ۫       S�      ��       S                        c�      j�       p @%�j�      v�       Pv�      ��       [��      ��       QB�      P�       [                                g�      �       Y�      ��       P��      �       p 
����      �       P1�      D�       Pn�      ��       P
�      ,�       0�B�      P�       Y�      �       P                               �      �       0��      �       s  z "��      �       s  y "�1�      ;�       s  y "�;�      D�       z s �n�      ��       z s �
�      ,�       s  z "��      �       z s �                     "�      �       �[�Ш      
�       �[�d�      �       �[�                      m�      t�       ���x�      ��       U��      ��       u|���      ��       U                       "�      �       �[�Ш      e�       �[���      
�       �[�d�      �       �[�                         "�      �       ���Ш      @�       ���@�      e�       X��      
�       ���d�      �       ���                       "�      �       SШ      ��       S��      
�       Sd�      �       S                       "�      �       ]Ш      e�       ]��      
�       ]d�      �       ]                     "�      �       ]Ш      
�       ]d�      �       ]                            -�      P�       PP�      |�       q �|�      �       ss s  $0-( 4&�Ш      ��       ss s  $0-( 4&���      
�       ss s  $0-( 4&�d�      �       P                                -�      |�       �[�|�      ��       T��      ��       t u "���      
�       T��      ��       T��      ��       R�      �       r p '��      ;�       R;�      L�       PL�      e�       x d�      �       �[�                              -�      |�       �[�|�      ֧       U֧      ٧       u z "�٧      
�       UX�      ��       U��      B�       TB�      D�       t p "�D�      V�       TV�      e�       ��d�      �       �[�                           -�      |�       �[�|�      �       Z�      
�       Z"�      �       Z�      B�       UB�      L�       u p "�L�      e�       Pd�      �       �[�                                -�      |�       �[�|�      ��       [��      ��       P��      ��       t p "���      �       P�      
�       [�      ��       [��      �       S;�      e�       Qd�      �       �[�                     -�      �       ��#�Ш      
�       ��#�d�      �       ��#�                     -�      �       ����Ш      
�       ����d�      �       ����                     -�      �       �J�8�Ш      
�       �J�8�d�      �       �J�8�                     -�      �       ����Ш      
�       ����d�      �       ����                        >�      �       XШ      $�       X��      
�       Xd�      �       X                   >�      |�       Qd�      �       Q                       |�      ��       r ��      ��       P��      ��      
 p ����z���      ��       P��      
�      * rp���#?$��������# %!����z�                       |�      ��       r��      ��       rt��      ��       P��      ʧ      	 p �J�8�ʧ      ӧ       Pӧ      
�      * rt�����z@$��������# %!�J�8�                  |�      ��       r��      �       rx                  	

     |�      ��       r��      �       r|�      �       P�      �      	 p ��#��      ��       P��      
�      * r|�����z># $��������%!��#�                     
�      �       XШ      $�       X��      
�       X                             
�      �       0�Ш      b�       0�b�      l�       Pl�      |�       Q|�      ��       P��      ��      
 p ����z���      ��       P��      
�       0�                             
�      �       0�Ш      ,�       0�,�      6�       P6�      G�       QG�      P�       PP�      V�      	 p �J�8�V�      X�       P��      
�       0�                             
�      �       0�Ш      ��       0���      ��       P��      �       Q�      �       P�      �      
 p ����z��      "�       P��      
�       0�                                 
�      �       0�Ш      Ҩ       0�Ҩ      ٨       Q٨      �       P�      �      	 p ��#��      �       P��      ժ       0�ժ      �       Q�      �       0��      
�       Q                  ��      �       R�      �       r p '�                  �      ��       Q��      ��       T                ��      �       U                  �      !�       S!�      ;�       Q                      x�      x�       u x�      ��       Q��      ��       R��      ��       Q                    ��      ��       P��      ë       [�ë      ի       Q                             �       Q�      �	       �Q��	      �	       Q                           �       R�      �	       �R�                           :       X:      �	       �X�                             b	       Yb	      �	       �Y��	      �	       Y                        m      U	       SU	      _	      & u0�X�R"u �Xu "�Ru0-( | �_	      �	      ( u0�X�R"u �Xu "�Ru0-( u���	      �	       S                  p      �	       Z                            V      �       r p ��      �      	 ��}�p ��      _	      	 ��}�| �_	      �	       ��}�u���	      �	       ��}�u���	      �	      	 ��}�| �                                   0��      �       0��	      �	       0�                         V      m       Sm             u0x u } u0-( �      �       u0�Xr "u } u0-( ��      �       u0�X�R"u } u0-( ��      �	      # u0�X�R"u �Xu "�Ru0-( �                           V      p       Zp      w       ~ u(v { +( �w      �       ~ u(v u8+( ��      �       ~ u(�Xu("�Ru8+( ��      �	      # u8�X�R"u(�Xu("�Ru8+( ��	      �	       ~ u(v u8+( �                     V             X      �       �Xr ��      �	       �X�R�                   �      K	       v�0$0&v�0$0& $ &�K	      U	       v��0$0&v��0$0& $ &�                           	      	       p r "#��@&q "�	      	       v �0$0& r "#��@&q "�	      	       X	      !	       v �0$0& r "#��@&q "�!	      K	      * v �0$0& v �0$0& ?&"#��@&��}"�K	      U	      , v��0$0& v��0$0& ?&"#��@&��}"�                          	      !	       X!	      >	      3 v �0$0& v �0$0& ?&"#��@&p "} "��}"s �>	      B	      ; v �0$0& v �0$0& ?&"#��@&s  $ &��}"p "} "#�B	      K	      9 v �0$0& v �0$0& ?&"#��@&s  $ &��}"p "} "�K	      U	      ; v��0$0& v��0$0& ?&"#��@&s  $ &��}"p "} "�                     	      !	       S!	      >	       P>	      B	       p�                �      	       T                �      	       v �0$0&�                   �      	       P	      	      
 p r "#���                  �      	       p ?&�	      	       R                        g	      r	       Sr	      v	       s�{	      �	       S�	      �	       S                          g	      {	       P	      �	       P�	      �	       s 2$� "
P�	      �	       s2$� "
P�	      �	       P                      g	      {	       R�	      �	       R�	      �	       R                                          �u      �u       U�u      �u       u��u      �u       U�u      �u       u��u      �u       u�v      v       U7v      lv       Ulv      �v       R�v      �v       U�v      �v       u��v      �v       u��v      w       u�-w      ?w       U?w      Jw       u�                      �u      w       Tw      -w       �T�-w      Jw       T                            �u      �u       Q�u      4v       V4v      7v       �Q�7v      *w       V*w      -w       �Q�-w      Jw       V                                  �u      �u       R�u      6v       \6v      7v       �R�7v      �v       \�v      �v       R�v      ,w       \,w      -w       �R�-w      ?w       \?w      Jw       R                 �u      �u       t�                                 �u      �u       Q�u      �u       p O���u      �v       Q�v      �v       p ���v      �v       Q�v      w       Q-w      ?w       Q?w      Bw       p ��Bw      Jw       Q                                           �u      �u       0��u      Sv       XSv      ]v       p ��]v      xv       Xxv      |v       P�v      �v       X�v      �v       p O���v      �v      
 s �O���v      �v      
 s~�O���v      �v       X�v      w       0�w      w       X-w      4w       p ��4w      ?w       X?w      Jw       0�                            �u      �u       Q�u      4v       V4v      7v       �Q�7v      *w       V*w      -w       �Q�-w      Jw       V                     �u      �u       1��v      �v       3��v      �v      
 u  s "x "�?w      Jw       2�                         Yv      cv       2�lv      pv      	 z r u "��v      �v      	 z r u "��v      �v       1��v      �v       0�-w      ?w       3�                                  @I      zI       UzI      4K       ���4K      ;M       �U�;M      �N       ����N      OS       �U�OS      \S       ���\S      ~S       �U�~S      �S       ����S      �T       �U�                    @I      �I       T�I      �T       �T�                    @I      mI       QmI      �T       �Q�                                    @I      wI       RwI      �K       w �K      ;M       �R�;M      \S       w \S      ~S       �R�~S      �S       w �S      �S       �R��S      �S       w �S      T       �R�T      �T       w                           @I      _J       X_J      ~S       �X�~S      �S       X�S      �S       ����S      �T       �X�                     @I      �L       0��L      8M       ^8M      ;M       P;M      �T       0�                        mI      �I       Q�I      �I       ���#�I      _J       | ~S      �S       |                              �I      _J       X_J      �J       �X��J      �J       x 
(!��J      K      
 x 	�
(!�K      K       Q;M      lN       �X�OS      \S       �X�~S      �S       X�S      �S       ���                                �I      �K       w �K      �L       �R�;M      \S       w \S      ~S       �R�~S      �S       w �S      �S       �R��S      �S       w �S      T       �R�T      �T       w                          �I      4K       V;M      fP       VOS      \S       V~S      �S       V�T      �T       V                              �I      4K       ���4K      �L       �U�;M      �N       ����N      OS       �U�OS      \S       ���\S      ~S       �U�~S      �S       ����S      �T       �U�                  �I      �L       ����;M      �T       ����                                    �J      �J       0��J      �J       PK      4K       P4K      �L       ^;M      oM       0�YN      lN       ^lN      wN       PwN      OS       ^TS      \S       ��\S      ~S       ^�S      �S       0��S      �T       ^                      �I      J       RJ      _J       v�~S      �S       v�                      �I       J       P J      _J       v�#P~S      �S       v�#P                  �I      �L       S;M      �T       S                               �I      _J       U_J      eK       ���;M      MQ       ���OS      \S       ���~S      �S       U�S      �S       s��S      �S       ����T      �T       ���                     �I      �I       T�I      �L       ���;M      �T       ���                  �I      �L       \;M      �T       \                           �J      �L       _;M      oM       _YN      lN       0�lN      OS       _TS      \S       Q\S      ~S       _�S      �T       _                   �J      �J        ;M      oM                                �J      kK       ];M      oM       ]lN      �R       ]T      �T       ]                  FJ      _J       ���~S      �S       V                  FJ      _J       ���~S      �S       ���                  FJ      _J       ����~S      �S       ����                    FJ      _J       0�~S      �S       0��S      �S       P�S      �S       0�                   _J      �J       @�oM      YN       @�OS      TS       @�                   _J      �J       ��	  oM      YN       ��	  OS      TS       ��	                     _J      �J       w oM      YN       w OS      TS       w                    _J      �J       �șoM      �M       �ș                            _J      �J       0��J      �J       _oM      �M       _�M      �M       P�M      �M       Q�M      .N       ���TN      YN       0�TS      TS       Q                         _J      �J       @��J      �J       QoM      �M       Q�M      �M       P�M      �M       w �����1$}"�
�?
���                       �J      �J      + q ����3$`�H     "#�����3$ �H     "oM      �M      + q ����3$`�H     "#�����3$ �H     "�M      �M      + p ����3$`�H     "#�����3$ �H     "�M      �M      = w �����1$}"�
�?
��3$`�H     "#�����3$ �H     "                       �J      �J       q ����3$`�H     "oM      �M       q ����3$`�H     "�M      �M       p ����3$`�H     "�M      �M      & w �����1$}"�
�?
��3$`�H     "                    �M      �M       U�M      YN       ���OS      TS       ���                �K      �K                       �K      �K       s� �s� ��                   �K      �K       P�K      �K      
 p t "#���                  �K      �K       p ?&��K      �K       T                �K      �K                          �K      �K       R�K      �K      
 p r "#���                  �K      �K       r ?&��K      �K       P                �L      �L                         �L      �L       P�L      �L       s�                    �L      �L       P�L      �L      
 p q "#���                  �L      �L       p ?&��L      �L       Q                �L      �L                       �L      �L       s�                    �L      �L       Q�L      �L      
 q r "#���                  �L      �L       q ?&��L      �L       R                   �N      =Q       _�T      �T       _                   �N      fP       V�T      �T       V                   �N      =Q       �����T      �T       ����                   �N      8Q       0��T      �T       0�                      �N      �N       P�N      =Q       ����T      �T       ���                     �N      �N       X�N      aO       ����T      �T       ���                 AO      oO        #�����3$ �H     "                      �N      �N       p��N      �P       ���#��T      �T       ���#�                      �N      �N       ����0$p 0$.��N      FP       ��������.��T      �T       ��������.�                      �N      �N       P�N      =Q       �Ș�T      �T       �Ș                      O      DO       PDO      =Q       ����T      �T       ���                  �O      �O       p @$�����                  �O      �O       P                �O      �O       ���#                   �O      �O       p @$��O      �O       P                   �O      �O       P�O      �O      
 p q "#���                  �O      �O       p ?&��O      �O       Q                  fP      yP      	 q �����                  �P      �P       P                  fP      jP       p jP      yP       ���#                  fP      yP       Q                   wP      yP       PyP      yP      
 p q "#���                  wP      yP       p ?&�yP      yP       Q                R      R       �Ț                R      R       s�                   R      R       QR      R      
 p q "#���                  R      R       q ?&�R      R       P                  �R      OS       P                 �R      OS       X                 �R      OS       ]                  �R      OS       U                  �R      OS       T                   |R      OS       �����T      �T       ����                   |R      OS       ����T      �T       ���                        �R      �R       q  $ &X���"X��R      OS       ���� $ &X���"X��T      �T       q  $ &X���"X��T      �T       ���� $ &X���"X�                  �T      �T       T                 �T      �T       ���                 (T      <T       T                (T      <T       ���                 mI      �I       Q                 mI      �I       \                 �I      �I       \                   �I      �I       U�I      �I       ����                 �L      !M       ����                 �      �       U                    �.      �.       U�.      �.       �U�                    �.      �.       T�.      �.       �T�                              pU      ~U       U~U      qV       YqV      wV       �U�wV      �V       Y�V      �V       �U��V      �V       Y�V      �V       �U��V      BW       Y                  pU      �U       T                                                    pU      SV       QSV      WV       SWV      dV       QdV      vV       SvV      wV       �Q�wV      �V       Q�V      �V       S�V      �V       �Q��V      �V       Q�V      �V       S�V      �V       �Q��V      �V       Q�V      �V       S�V      �V       Q�V      �V       S�V      �V       Q�V      4W       S4W      BW       Q                          pU      qV       0�wV      �V       0��V      �V       P�V      �V       0��V      �V       P�V      BW       0�                              tU      ~U       U~U      qV       YqV      wV       �U�wV      �V       Y�V      �V       �U��V      �V       Y�V      �V       �U��V      BW       Y                                 tU      ~U       u~U      UV       yWV      qV       ywV      �V       y�V      �V       y�V      �V       y�V      �V       y�V      �V       y4W      BW       y                                 tU      ~U       u~U      UV       yWV      qV       ywV      �V       y�V      �V       y�V      �V       y�V      �V       y�V      �V       y4W      BW       y                                 tU      ~U       u ~U      UV       y WV      qV       y wV      �V       y �V      �V       y �V      �V       y �V      �V       y �V      �V       y 4W      BW       y                      wV      �V       Q�V      �V       S�V      �V       �Q�                  WV      dV       QdV      qV       S                 WV      qV       y�����3$`�H     "                   �V      �V       S�V      �V       �Q�                   �V      �V       Q�V      �V       S                 �V      �V       S                 �V      4W       y$�                   �V      �V       Q�V      4W       S                  SV      WV       Q                 SV      WV       S                           U      "U       U"U      -U       S-U      /U       �U�/U      WU       SWU      fU       U                             U      "U       T"U      .U       V.U      /U       �T�/U      5U       T5U      WU       VWU      fU       T                           U      "U       Q"U      /U       �Q�/U      9U       Q9U      WU       �Q�WU      fU       Q                       U      (U       0�/U      :U       0�:U      NU       PUU      fU       0�                    p6      �6       U�6      �6       �U�                      p6      �6       T�6      �6       Z�6      �6       �T�                    p6      �6       Q�6      �6       �Q�                      p6      �6       R�6      �6       V�6      �6       �R�                      �6      �6       rp ��6      �6       r p ��6      �6       R                   �6      �6       s p ��6      �6       X                  �6      �6       P                           O       RO      n       t0n      �       R                           g       Pg      n       u�(n      �       P                                  0�      *       q ��*      �       Q                  �      �       Z                 �      �       U                 �      �       T                            @#      �#       U�#      \$       _\$      ^$       [^$      I(       �U�I(      \(       U\(      u(       _                          @#      �#       T�#      ^$       w ^$      I(       �T�I(      \(       T\(      u(       w                         }#      �#       S�#      ^$       ��^$      I(       �T����
�	�U"#H�I(      u(       ��                       }#      %       0�%      +%       P�%      �'       0��'      u(       0�                              �#      �#       S�#      �#       u �#      �#        �#      ^$       ��I(      M(       SM(      \(       u \(      u(       ��                     �#      �#       t ����
�Gv "#P��#      $       w �����
�Gv "#P�I(      \(       t ����
�Gv "#P�                   �#      �#       RI(      \(       R                       �#      �#       0�I(      T(       0�T(      W(       SW(      \(       ��~                     �#      L$       \L$      ^$       SI(      u(       \                      �#      �&       ]�'      	(       ]I(      u(       ]                                     $      L$       \L$      �%       S�%      a&       \a&      q&       Ru&      }&       R}&      �&       P�&      �&       [�&      �'       P�'      	(       S	(      I(       P\(      u(       \                    �#      �#       SI(      \(       u                              $      $       P$      $       U$      /$       P/$      W&       V�'      	(       V\(      d(       Pd(      u(       V                      �#      �'       ^�'      I(       ^\(      u(       ^                      �#      �#       P�#      ^$       ��\(      u(       ��                   m$      �%       0��'      	(       Q                  �$      �$       0�                     �$      �$       Q�$      �$       q���'      	(       Q                      �$      �$       P�'      �'       P�'      	(       u u r  $0-( �                   l%      r%      	 p 0$0&�r%      �%       q �0$0&�                      r%      y%       Py%      �%      
 p r "#����%      �%       P                   r%      y%       p ?&�y%      �%       R                     �%      �%       0��%      &       0�&      C&       Q                  �%      �%       0�                     �%      �%       Q�%      &       q��&      C&       Q                      �%      &       P&      !&       P!&      C&       u u r  $0-( �                 C&      a&       �T����
�	�U"#`                    W&      �'       V	(      I(       V                       W&      a&       �T����
�	�U"#`a&      �&       Q�&      �'       T	(      I(       T                     �&      �&       0��&      �'       Z	(      I(       Z                     �&      �&       0��&      �'       S	(      I(       S                      �&      '       X'      �'       0�(      ;(       X                        �&      Y'       Q�'      �'       Q	(      (       Q-(      ;(       Q                       �&      '       p '      Y'       R�'      �'       p 	(      (       R)(      ;(       U                  '      D'       X                  2'      D'       U                �#       $       S                �#       $       w �����
�Gv "#��                   �#       $       P $       $      
 p q "#���                  �#       $       p ?&� $       $       Q                           �       U�      �       �U�                           �       T�      �       �T�                           �       Q�      �       �Q�                           �       R�      �       �R�                            �       r ����
�	u "#H��      �       �R����
�	u "#H��      �       �R����
�	�U"#H�                  =      �       X                  L      �       Z                      e      q       v 8&�q      �       \�      �      / �U#�(#H�����8&1�U#�(#H�����8&0.( �                    �      �       V�      �       �U#�(#H�����
p;&�                  [      �       ]                     �      �       X�      �       T�      �       X                    �      �       R�      �       P                   �      �      	 u 0$0&��      �      	 u 0$0&�                        �      �       r�0$0&��      �       r��0$0&��             P      �       r�0$0&�                 �      �       t�0$0&��      u       t�0$r�0$+( 0$0&�                 �      �       t�0$0&��      u       t�0$r�0$-( 0$0&�                        �       Y                            (       P(      .       _.      �       r�0$0&u �                  W      �       _                  k      �       P                    9      M       PM      W       r�0$0&u :$} 
 �                        @      j       Uj      |       ��~|      �       �U��              U                        @      C       TC      |       ��~|      �       �T��              T                 @      B       u�(                         @      C       t ����
�	u "#H�C      j       ��~�����
�	u "#H�j      |       ��~�����
�	��~"#H�|      �       �T����
�	�U"#H��              t ����
�	u "#H�                        m      q       Pq      j       u j      |       ��~�              u                             m      �       0��             ��~d             0�             R=      f       0�f      k       ��~k      !       0�}      �       0��      �       ��~�      p       0�p             R              0�                                    m      |       0�|      `       [`      �       _�      �       [�      �       [      [       [f      �       [!      U       [U      h       0�h      �       [�      �       0��      S       [S      �       Q�      �       [p      �       [�              0�                                �      �       P�      �       Q�      ;       u� ;      #       ��~!      ;       P;      �       ��~      �       ��~�              u�                       �      �       P�      |       ��~�              ��~                                     R      |       ��~�      �       R�              ��~                                                     R      |       ��~|      �       ��}�      k       \k      !       ��}!      }       \}      �       ��}�      �       \�             \      �       ��}�             \      �       ��}�      �       R�              ��~                      �      �       P�      |       ��~�              ��~                           )       P)      6       p��6      ;       P                                u,� $ &Pp "�      ;       u,� $ &Pu0"�                       �      �       u0�      �       P�      �       p���              P                 �              u,� $ &Pu0"�                                 �      �       P�      �       ��~�      #       ��}#      �       S�      �       S�             S      �       ��~�      �       Q�      �       P                       �      �       Q�      �       ��~#H�      #       ��}      �       Q�      �       ��~#H                                        �      #       0�#      `       V`      d       0�d             V      �       1��      8       V8      d       1�d             V      =       1�=      k       Vk      U       1�U      h       0�h      �       1��      �       V�      �       V�             V      �       0�                                    �      #       
 }��      �       P.      8       {� #08      d       s0      =       s0k      !       P!      ,       s0h      }       s0}      }       P             P�      �       P      �       
 }�                                    �      #        ���      �       Q.      8       {� #08      d       s0      =       s0k      !       Q!      ,       s0h      }       s0}      }       Q             Q�      �       Q      �        ��                            �      #       
 }�#      �       R.      d       R      =       Rk      �       R      ]       R      �       
 }�                                     �      #        ��#      �       T.      d       Rd      �       T      =       R=      !       T!      }       R}      �       T�      �       T�      ]       T�      �       T      �        ��                            �      #       0�#      �       ^�      �       ^.      �       ^      �       ^�      �       ^�      �       ^      �       0�                                    �      #       0�#      �       ��}�      �       ��}.      d       ^d      �       ��}      =       ^=      !       ��}!      }       ^}      �       ��}�      �       ��}�      �       ��}      �       0�                	                 �      #       
 }�#      �       X8      d       
 }�d      �       X      =       R=      !       X!      >       
 }�h      }       R}      �       X�      L       X      �       
 }�                
                   �      #        ��#      �       U8      d        ��d      �       U      =       R=      !       U!      >        ��h      }       R}      �       U�      ]       U�      �       U      �        ��                                 �      #       0�/      `       ��}d      k       ��}{             ��}�      �       ��}d             ��}=      !       ��}}      �       ��}�             ��}�      (       ��}                            �      #       0�#      =       _T      `       [`      �       _.      �       _�      �       _�             _      �       0�                        �      #       
 }�T      �       P             p } -( ��      �       P      �       
 }�                        �      #        ��T      �       Q�             q { +( ��      �       Q      �        ��                                     �      #       
 }�#      `       ��}d             ��}�      T       ��}T      �       R�      �       ��}d             ��}=      !       ��}}      c       ��}c      �       R�      �       ��}�      �       ��}�      (       ��}      �       
 }�                                     �      #        ��#      `       ��}d             ��}�      T       ��}T      �       T�      �       ��}d             ��}=      !       ��}}      c       ��}c      �       T�      �       ��}�      �       ��}�      (       ��}      �        ��                                     �      #       0�#      `       ��~d             ��~�      T       ��~T      �       ^�      �       ��~d             ��~=      !       ��~}      c       ��~c      �       ^�      �       ��~�      �       ��~�      (       ��~      �       0�                                       �      #       0�#      `       ��~d             ��~�      T       ��~T      ]       _]      �       ��}�      �       ��~d             ��~=      !       ��~}      c       ��~c      �       ��}�      �       ��~�      �       ��~�      (       ��~      �       0�                                     �      #       
 }�#      `       ��~d             ��~�      T       ��~T      �       X�      �       ��~d             ��~=      !       ��~}      c       ��~c      �       X�      �       ��~�      �       ��~�      (       ��~      �       
 }�                      		       		        �      #        ��#      `       ��~d             ��~�      T       ��~T      �       U�      �       ��~d             ��~=      !       ��~}      c       ��~c      �       U�      �       ��~�      �       ��~�      (       ��~      �        ��                            �      �       Y�      7       s0k             s0}      �       s0      K       s0�      �       s0                            �      �       Y�      7       s8k             s8}      �       s8      K       s8�      �       s8                      �      �       ��	  d             ��	  =      f       ��	  �      �       ��	  �             ��	  �      p       ��	                         �      �       ��~d             ��~=      f       ��~�      �       ��~�             ��~�      (       ��~                      �      �       �T����
�	�U"#H�d             �T����
�	�U"#H�=      f       �T����
�	�U"#H��      �       �T����
�	�U"#H��             �T����
�	�U"#H��      p       �T����
�	�U"#H�                              �      �       0��      �       [d             0�             [=      f       0�f      f       [�      �       0��             0��      p       0�p      p       [                        t      �       Q�      �       Q�             Q�      �       Q�      �       ��~��~"#L                             t      �       Q�      �       Z�             ��}�      �       Q�             Z             p q "#��      �       Z�      (       ��}                      t             �����      �       �����             �����             ����                  D      ]       Q                  S      �       X                          ]      �       q� �      �       qp�      �       T�      �       q� �      �       qp                    ]      �       U�      �       U                            ]      h       Rh      �       q� #8�      �       qp#8�      �       R�      �       q� #8�      �       qp#8                      ]      �       P�      �       P�      �       u8                 ]      o       q� #Ho      �       u�                  �      �       q� #H�      �       u�                         �,      -       U-      -       S-      -       U-      -       �U�                        �,      -       T-      -       V-      -       T-      -       �T�                                �(      �(       U�(      �)       S�)      �)       �U��)      e*       Se*      z*       Uz*      �+       S�+       ,       y��~� ,      �,       S                        �(      �(       T�(      e*       �T�e*      z*       Tz*      �,       �T�                                �(      �(       Q�(      �)       ^�)      �)       �Q��)      e*       ^e*      z*       Qz*      �*       ^�*      0,       �Q�0,      �,       ^                        �(      �)       _�)      �*       _0,      �,       _�,      �,       P�,      �,       _                    �(      �)       \�)      �,       \                                     �(      �(       q ����
�Gu "#P��(      �(       q ����
�Gs "#P��(      �)       ~ ����
�Gs "#P��)      �)       �Q����
�G�U"#P��)      e*       ~ ����
�Gs "#P�e*      z*       q ����
�Gu "#P�z*      �*       ~ ����
�Gs "#P��*      �+       �Q����
�Gs "#P��+       ,       �Q����
�Gy "
�I� ,      0,       �Q����
�Gs "#P�0,      �,       ~ ����
�Gs "#P�                              �(      �(       0��(      )       P9)      T)       0�T)      ])       Q])      �)       q��)      �)       Q�)      �)       0�z*      �*       0�D,      ^,       0�                         �(      �)       s����)      e*       s���z*      �+       s����+       ,       y�|� ,      �,       s���                   �(      )       0��)      �)       0��)      �)       p ����Hs "#ȓ�                   *      X*       Q0,      :,       Q                   *      6*       (�6*      9*       P                   =*      X*       P0,      :,       P                  *      X*       R0,      :,       R                     *      #*       P#*      X*       s#�#�
���0,      :,       s#�#�
���                    D,      ^,       T^,      x,       r t +( �x,      �,       T                  �,      �,       T�,      �,       t 	��                  ;,      �,       P                     �,      �,       p  ��,      �,       Q�,      �,       p  �                 �,      �,       T                      �,      �,       T�,      �,      
 q t "#����,      �,       t ?&t "#���                 �,      �,       t ?&�                	�)      �)       _                	 �)      �)       p ����Hs "#���                   �)      �)       P�)      �)      
 p q "#���                  �)      �)       p ?&��)      �)       Q                  h)      �)       R                h)      v)       r                    o)      v)       Pv)      v)      
 p x "#���                  o)      v)       p ?&�v)      v)       X                 �*      �*       ^                     +      +       R+      +       P+      !+       q                    +      !+       P!+      !+      
 p t "#���                  +      !+       p ?&�!+      !+       T                b+      b+       Tb+      b+      
 t  "#���                b+      b+       _                �)      �)       ~ ����
�Gs "#��                   �)      �)       P�)      �)      
 p q "#���                  �)      �)       p ?&��)      �)       Q                        ��      ґ       Uґ      �       V�      ��       �U���      �       V                        ��      ̑       T̑      �       S�      ��       �T���      �       S                        ��      Ǒ       PǑ      ̑       t�̑      ֑       s�֑      �       ��                 �      �       S                 �      �       V                         �      ]�       0�]�      ��       ]��      Ò       1�Ò      ˒       ]�      �       ]                     �      ˒       1�˒      �       ]�      �       1��      �       0�                        H�      ]�       0�]�      ��       w ��      Œ       PŒ      �       w                    ]�      ]�       P]�      �       \                     H�      ��       _��      ��       P��      �       _                H�      ]�       S                 H�      Q�       U                 ]�      ]�       P                   ��      Œ       ^�      �       ^                ��      ��       0�                    ��      ��       �����      ��       R��      ��       ���                ��      ��       \                ��      ��       V                 ��      ��       v�                  ��      ��       ^                ˒      ڒ       \                ˒      ڒ       S                 ˒      ْ       s�                    Є      �       U�      ��       ��w                    Є      �       T�      ��       ��w                           _�      u�       0�u�      .�       ��w�      ��       ��w��      ��       ��w��      Ջ       ��w�#�ڋ      S�       ��w��      ��       ��w                             _�      u�       0�u�      ׇ       ��xׇ      �       ��x�#��      �       P�      .�       ��x�      ��       ��x��      S�       ��x��      ��       ��x                     �      �       ��w#ē�����H��w"#ȓ��      P�       { ����H��w"#ȓ��      �       ��w#ē�����H��w"#ȓ�I�      n�       { ����Hs "#ȓ�                  0�      J�       P                   Є      �       u����      ��      	 ��w#���                                    7�      ��       v��v���v��v��v�����      p�      ; ��w#�#����w#�#���X���w#�#����w#�#���p�      ��      E ��w#�#����w#�#�����w#�#����w#�#����w#�#����      0�      E ��w#�#����w#�#�����w#�#����w#�#����w#�#���0�      ��      ; ��w#�#����w#�#���X���w#�#����w#�#�����      ��      ; ��w#�#����w#�#���X���w#�#����w#�#���ڋ      �      ; ��w#�#����w#�#���X���w#�#����w#�#����      '�       v��v���v��v��v���n�      S�      ; ��w#�#����w#�#���X���w#�#����w#�#�����      ��      ; ��w#�#����w#�#���X���w#�#����w#�#���                
 Є      ҄       u                         �      ��       p��      �       u #�      3�       ��w#3�      J�       S                        �      �       P�      �       ��w!�      #�       P#�      ��       ��w                    /�      3�       P3�      ��       ��x                       8�      ?�       P?�      ��       w ��      ��       ��w��      ��       w                                       _�      u�       Su�      ��       [��      ƅ       Pƅ      ��       [��      �       ��w�      �       [�      ��       ��w��      '�       ��w'�      ��       [n�      S�       ��w��      ��       ��w                     �      �       ��w#ē�����H��w"#ȓ��      P�       { ����H��w"#ȓ��      �       ��w#ē�����H��w"#ȓ�I�      n�       { ����Hs "#ȓ�                     �      �       ��w#ē�����H��w"#����      P�       { ����H��w"#����      �       ��w#ē�����H��w"#���I�      n�       { ����Hs "#���                                   _�      u�       0�u�      p�       S��      �       S�      .�       \0�      }�       S}�      �       ��w��      ڋ       S��      �       ��w�      '�       S'�      n�       \                                   _�      u�       0�u�      p�       ]��      �       ]�      .�       V0�      u�       ]u�      �       ��w��      ڋ       ]��      
�       ��w�      '�       ]'�      n�       V                 �      /�       T                             ��      �       0��      ��       0��      ��       0���      Ջ       0�ڋ      '�       0�n�      S�       0���      ��       0�                                      Q�      ��       	����      ��       Z��      �       R�      ��       P��      �       R�      �       Z�      G�       RG�      V�       PV�      p�       Z0�      9�       Zڋ      �       Z�      '�       	��n�      �       Z                                Q�      ��       0���      p�       ��w0�      ��       ��w��      ��       ��wڋ      �       ��w�      '�       0�n�      S�       ��w��      ��       ��w                                  Q�      ��       0���      �       ��w�      p�       ��w0�      ��       ��w��      ��       ��wڋ      �       ��w�      '�       0�n�      S�       ��w��      ��       ��w                           ��      �       ��w��      ��       ��w�      ��       ��w��      '�       ��wn�      S�       ��w��      ��       ��w                             ��      ��       0���      ��       ��w��      ��       ��w�      ��       ��w��      '�       ��wn�      S�       ��w��      ��       ��w                               ��      ��       0��      p�       \��      ��       \0�      ��       \��      :�       ��w��      ڋ       \��      �       ��w�      '�       \                                    Q�      ��       0���      �       U�      �       p  $ &4$x "#�      G�       UG�      V�       p  $ &4$x "#V�      ��       U�      ��       U��      ��       Uڋ      �       U�      '�       0�n�      S�       U��      Ȑ       U                                 �      p�       0�p�      ��       P�      0�       P0�      ��       0���      ��       1���      ��       0�ڋ      '�       0�n�      S�       0���      ��       0�                    Q�      ��       0��      '�       0�                        Q�      ��       0���      p�       [0�      ��       [�      '�       0�                      ��      p�       T0�      @�       T@�      ��       {�                   ��      �       Z�      V�       Z                                    ��      ̆       P̆      І       p�І      Ԇ       �چ      �       P�      ��       p���      ��       ��      ,�       P,�      0�       p�0�      4�       �:�      V�       P                                r�      ��       Q��      �       ]�      9�       ��wڋ      ��       ��w��      �       ]�      �       ��wn�      �       ��w�      �       z  $ &4$x "                                       {�      ��       T��      ��       R��      ��       T��      �       R�      �       [�      ,�       t v  $t  $-( �,�      A�       t��w�v  $t  $-( ���      �       R�      �       [��      ��       P��      ��       p���      ӎ       P                                   {�      ��       T��      A�       ZA�      P�       TP�      [�       [[�      ڊ       Tڊ      �       {��w�  ${  $+( �ڋ      �       T�      �       {}   ${  $+( ��      ��       {��w�  ${  $+( ���      �       Z                                 r�      ��       T��      ��       R��      �       T�      5�       R5�      9�       ��w9�      ��       R��      ��       Rڋ      ��       ��w��      �       Tn�      �       ��w                                     r�      ��       T��      A�       ZA�      P�       TP�      ��       [��      ��       T��      ��       Tڋ      ��       [��      �       Zn�      ގ       Tގ      �       V�      S�       ��x��      ��       ��x                                                {�      ��       R��      �       S�      ��       R��      �       S�      A�       ��wA�      ��       R��      ��       T��      Պ       RՊ      ��       ��w��      ��       ��wڋ      ��       R��      ��       ��w��      �       S�      �       ��wn�      S�       ��w��      U�       ��w_�      c�       ��w                                                {�      ��       R��      ��       \��      ��       R��      �       \�      A�       ��wA�      ��       \��      ��       T��      ڊ       \ڊ      ��       ��w��      ��       ��wڋ      ��       \��      ��       ��w��      �       \�      �       ��wn�      S�       ��w��      J�       ��w_�      h�       ��w                                                          ��      ��      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&���      Ɖ       PƉ      Љ       { 4$x "#u y 'y �Љ      �      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&��      ,�      x t v  $t  $-(  $ &4$x "#u t v  $t  $-(  $ &4$x "#u ?&'t v  $t  $-(  $ &4$x "#u ?&�,�      A�      � t��w�v  $t  $-(  $ &4$x "#u t��w�v  $t  $-(  $ &4$x "#u ?&'t��w�v  $t  $-(  $ &4$x "#u ?&�A�      P�       yu yu ?&'yu ?&�w�      ��       P��      �       yu yu ?&'yu ?&��      �       t  $ &4$x "x q "��      9�       t  $ &4$x "r  $ &4$x "�ڋ      ��       yu yu ?&'yu ?&���      �      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&�n�      ��       t  $ &4$x "r  $ &4$x "���      ގ      " t  $ &4$x "��w� $ &4$x "�ގ      ��      " v  $ &4$x "��w� $ &4$x "�;�      ��       P��      ��      0  4$x "#y  4$x "#y ?&' 4$x "#y ?&�(�      C�       P��      ��       P��      ��      0  4$x "#y  4$x "#y ?&' 4$x "#y ?&���      ��      6  4$x "#��w 4$x "#��w?&' 4$x "#��w?&�                          �      9�       _n�      z�       _z�      S�       ��w��      ��       ��w��      ��        ��w#H�������Q %3%�����                               ��      ގ       Tގ      �       V�      ��       ]��      ʏ       Vʏ      �       ](�      C�       ]C�      S�       V��      ؐ       ]ؐ      ��       ��w                                 ��      ގ       Tގ      ��       V��      �       P�      S�       V��      ��       V��      L�       TL�      _�       V_�      ��       T��      ��       V                                 ��      �       0��      ��       1���      ��       P��      ʏ       0�ʏ       �       1� �      (�       P(�      C�       1�C�      S�       0���      ��       1�                              ʏ       	��:�      C�       VG�      S�       V��      ��       Q                             ʏ       	��(�      S�       V��      .�       Z.�      _�       V_�      ��       Z                 ��      Ɏ       ��x                     {�      ��       s { +���      А       s { +�А      ��        4$x "{ +�                             ��      ��       p 4$x "#��w���      L�       t 4$x "#��w�L�      _�       v 4$x "#��w�_�      q�       t 4$x "#��w�q�      ��       v 4$x "#��w���      ��       t 4$x "#��w���      ��       v 4$x "#��w�                �      �       ��	                  �      �       0�                �      �       \                �      �       w                 �      �       ��w                �      �       ��w#@                 �      �       T                 ^�      ��       { ����H��w"#ȓ                 ^�      ��       { ����H��w"#��                 ^�      p�       r q +�                      '�      H�       1�H�      ��       U��      ��       u�                 k�      w�       u ����u����3$p "                      ��      Ό       1�Ό      ��       X��      ��       x�                 �      �       x ����x����3$p "                      \�      z�       R��      ��       P��      ��       R                  j�      n�       p���      ��       P                        ��      ��       1���      ��       [��      �       {��      �       ]                  ��      ��       [                    È      �       U��      �       U                    ˈ      �       T��      �       T                 8�      8�       P                .�      C�       w                 .�      C�       ��w                 .�      B�       ��w#�                        p�      ��       U��      p�       Vp�      y�       �U�y�      ʄ       V                        p�      ��       T��      �       ^�      ��       �T���      ȃ       ^ȃ      ʄ       �T�                      T�      ��       Pق      �       P��      �       P                    �      0�       0�0�      ��       _��      ȃ       0���      ʄ       _                           �      ��       S��      ��       s�ȃ      �       0��      b�       1�b�      y�       2�y�      ��       0���      ��       1���      ʄ       S                 ʁ      ʄ       ���}�                	   ʁ      ́       Ṕ      ݁       v                 
   ʁ      ́       p�����3$ �H     "́      ݁       v #�����3$ �H     "                    �      �       P�      �       \��      ȃ       \                       ف      *�       S*�      C�       PC�      c�       S��      ȃ       S                ,�      0�       0�                ,�      0�       \                ,�      0�       V                ,�      0�       v�                  0�      0�       _                   �      ��       s  $ &
�Gv "#P���      ʄ       s  $ &
�Gv "#P�                   �      ��       s  $ &
�	� "
X����      ʄ       s  $ &
�	� "
X��                    �      ��       P��      ʄ       P                        '�      ��       U��      ��       |� � $ &54$|� "���      ��       |�l� $ &54$|�l"���      ʄ       U                          D�      `�       Q`�      d�       p d�      s�       pP��      ��       Q��      ʄ       p                   ��      ʄ       Q                       ȃ      �       v� ��      p�       v���p�      y�       �U#���y�      ��       v� ���      ��       v���                          �      )�       R)�      -�       v�-�      f�       R��      ��       R��      ��       v�                ف      �       ^                 ف      ݁       X                 �      �       P                5�      D�       \��      ȃ       \                5�      D�       ^��      ȃ       ^                  5�      C�       ~���      ǃ       ~�                   ��      ��       ]��      ʄ       ]                 ��      Ԃ       P                  ��      ʁ       X                    ��      ��       ���|���      ʁ       ]                    g      g       Ug      g       �U�                    g      g       Tg      g       �T�                    g      g       Qg      g       �Q�                    g      g       Rg      g       �R�                    �      �       T�      �       �T�                    0#      1#       U1#      2#       �U�                    0#      1#       T1#      2#       �T�                         �      #�       U#�      F�       VF�      I�       �U�I�      l�       V                         �      �       T�      C�       SC�      I�       �T�I�      l�       S                    �      H�       \I�      l�       \                          �?      l@       Ul@      �@       �U��@      �@       U�@      C       �U�C      @C       U                          �?      l@       Tl@      �@       ���@      �@       T�@      C       ��C      @C       T                        @      l@       X�@      �@       XC      ,C       P,C      @C       X                      @      l@       Z�@      �@       ZC      @C       Z                         @      l@       Yt@      SA       Y3B      AB       Y C      C       YC      @C       Y                    !@      �@       _�@      @C       _                              Q@      \@       8�\@      �@       ]�@      �@       4��@      /A       ]FA      C       ]C      ,C       8�,C      @C       4�                                                                  )@      5@       X5@      @@       P@@      L@       p��L@      _@       P_@      l@       ^�@      �@       X�@      �@       x���@      �@       X�@      �@       P�@      �@       p���@      �@       P�@      A       ^A      &A       S&A      8A       X8A      <A       x��<A      FA       XFA      SA       SSA      uA       PuA      �A       p� ��A      �A       V�A      �A       T�A      �A       VAB      GB       p� ��B      �B       P�B      �B       p� �C      ,C       P,C      @C       X                      c@      �@       \�@      /A       \FA      C       \                          c@      l@       ^�@      A       ^A      A       SA      &A       ^FA      �B       ^C      C       ^                        uA      �A       P�A      �A       ��AB      rB       P�B      �B       PC      C       P                   GB      �B       VC      C       V                   GB      rB       PC      C       P                   GB      �B       v��C      C       v��                 �A      �A       S                   �A      �A       P�A      �A       ��                 �A      �A       \                  �A      AB       S                  �A      B       P                    �A      B       TB      AB       s��                  �A      AB       ^                   �B      �B       S�B      �B       s��                 �B      C       \                 �B      �B       ^                            �B      �B       ^�B      �B       ~���B      �B       ^�B      �B       S�B      �B       s���B      C       S                    �B      �B       p s8��B      C       P                    @      �       U�      �        �U�                        @      �       T�      �       ^�      �       �T��      �        ^                 @      D       u0                 @      D       u,� $ &Pu0"�                       @      �       t ����
�	u "#H��      �       ~ ����
�	�U"#H��      �       �T����
�	�U"#H��      �        ~ ����
�	�U"#H�                    ^      �       V�      �        V                  y      �       X                      �      �       ]�      �       	�0�T $0)( 	�#��      �        ]                    �      �       S�      �        S                               �      �       V�      Y       x���      �       V�              x��       ?        Z?       D        y 3$v "�D       U        Zk       �        Z�       �        x��                                    �      v       \�      �       P�      �       P�      �       \�      �       P�      �       \�      �       P�      �        \�       �        P�       �        \                        �      )       P�      �       P�      �       P�              P�       �        P                     �      v       \�      �       \�      �        \                        �      �       t | ��      s       | x��0$0&��      �       t | ��      �        | x��0$0&��       �        | x��0$0&�                             Y       0��              0�       �        U�       �        0�                                   Y       q X��              q X�       )        [)       U        Tk       q        [q       �        T�       �        q X�                                 7        T7       P        PP       U        Tk       q        Tq       �        P                       "       ;        YD       H        z �0$0&�H       U        Yk       �        Y                            -       0�-      P       U�       �        0�                      ^      s       [�       �        [�       �        ��                 s             P                 s      v       | u 0$0&�                         �       P�      �      
 p t "#���                        �       p ?&��      �       T                                �	      c
       Uc
      o       So      �       ���      X       SX      k       �U�k      �       ���      �       �U��      =       S                                    �	      c
       Tc
      h       ^h      �       ���      �       T�      P       ^P      k       �T�k      �       ���      �       �T��             T      =       ^                       �
      o       s0o      �       ��=      X       _k      �       ��                         <
      X
       u8X
      c
       u(�      �       s8�      �       s(�      �       s8�             s(             s8                                             <
      U
       PU
      X
       t �0$0&�X
      n
       Q�      �       P�      �       p}��      �       ~ �0$0&��      �       _�             Q      "       R"      =       _�      �       P�      �       t �0$0&��             Q             P      -       Q                       �	      X       \X      o       s�      X       \�      =       \                       �	      U       ]U      o       s�      X       ]�      =       ]                              
      
       P
      c
       uc
      ]       ���      �       s�      X       ���             s      =       ��                              
      
       P
      c
       u c
      �       ���      �       s �      �       ���             s       =       ��                     
      @       V�      I       V�      =       V                                      3      o       s0o      �       P=      X       _k      �       P#      s       Ss      �       R�      �       R�             Q#      �       P�      �       p���      �       P�             _A      �       _�      �       S                                  >       R>      �       w =      X       Rk      �       w       A       w �      �       w                                   p#��
���      o       s�(##��
���=      X       s�(##��
���                          3      H       PH      �       ��=      E       PE      X       ��k      �       ��                     3      �       [=      X       [k             [                     3      �       Y=      X       Yk             Y                         3      M       x M      h       ~h      o       ��#=      X       x �      �       q 1$s "                           3      �       U=      S       US      X       z 2$z "4$ "�k      �       U�      �       T�      �       U                             3      o       Uo      �       T�      �       t� �      �       T=      S       US      X       z 2$z "4$ "�k      �       P�      �       U�      �       T                       3      o       0�o      �       _=      X       0�k      �       _                 ~      �       p�0$0&t�0$0& $ &�                 ~      �       p�0$0&t�0$0& $ &�                               R            
 r s "#���                               r ?&�             S                  .      5       Q5      5      
 q r "#���                  .      5       q ?&�5      5       R                        A      X       Q�      �       Q�      �       qx��             Q                              S      X       P�      �       P�      �       U�             R             _      A       _�      �       _                      S      X       X�      �       X�      �       x~��             X                      S      X       0��      �       0��      �       P�             P                                   \      A       \�      �       \                                  ^      A       ^�      �       ^                                  _      A       _�      �       _                      #      �       S�             R      A       R�      �       S                     �      �       R�             Q      A       Q                            '      s       Rs      �       T�      �       R�      �       T�      �       R�      �       s�                       �      �       R�      �       P�             P      A       P                                                  9      H       s�0$0&u  $ &�H      M       PM      s       s�0$0&u  $ &�s      s        s�0$0&s� #�0$0& $ &�s      �       u t�0$0& $ &��      �       P�      �       u t�0$0& $ &��      �        s�0$0&s� #�0$0& $ &��      �       0��      �       Y             y u "�      t       Yt      �       z ��      �       0�      &       Y&      +       z �+      <       Y<      A       T�      �       s�0$0&u  $ &��      �        s�0$0&s� #�0$0& $ &�                                             9      Y       s�0$0&x  $ &�Y      c       Qc      s       s�0$0&x  $ &�s      s        s�0$0&s� #�0$0& $ &�s      �       x t�0$0& $ &��      �       Q�      �       x t�0$0& $ &��      �        s�0$0&s� #�0$0& $ &��      �       0��             T�      �       0��             T              T       +       t �+      3       T�      �       s�0$0&x  $ &��      �        s�0$0&s� #�0$0& $ &�                       _             T              T       +       t �+      3       T                          _      t       Yt      �       z �      &       Y&      +       z �+      <       Y<      A       T                    �      �       T       +       T                          &       Y&      +       z �                   �      �       Y      +       	��                     k      �       s {�0$0& $ &��      �       p�0$0&{�0$0& $ &��      �       pH�0$0&{�0$0& $ &�                   k      �       p�0$0&{�0$0& $ &��      �       pJ�0$0&{�0$0& $ &�                     k      �       z�0$0&s  $ &��      �       z�0$0&p�0$0& $ &��      �       z�0$0&pH�0$0& $ &�                   k      �       z�0$0&p�0$0& $ &��      �       z�0$0&pJ�0$0& $ &�                  k      �       Z                 k      �       [                  c      �       ]                  ~      �       ^                       -      M-       UM-      ;.       S;.      B.       �U�                      =-      �-       0��-      �-       1��-      ;.       2�                   =-      M-       u� �M-      �-       s� ��-      ;.       s��                                       ?       U?      �       \�      �       �U��      �       \�      )       U)      �       \�      �       U�      8       \                               ?       T?      �       S�      �       �T��      8       S                                       ?       Q?      �       ]�      �       �Q��      �       ]�             Q      �       ]�      �       Q�      8       ]                                       ?       R?      �       V�      �       �R��      �       V�      9       R9      �       V�      �       R�      8       V                                           3       X3      �       �X��             X             �X�      6       X6      e       Ue      �       �X��      �       X�      �       U�      8       �X�                                           6       Y6      �       ^�      �       �Y��      �       ^�             Y             ^      Y       YY      �       ^�      �       Y�      8       ^                       &      N       0�N      y       Qy      �       q� ��      �       Q�      8       0�                 ?      U       |                               e       Q�      �       Q�      �       u�      �       Q�      �       |                                   1       Q1      �       _�      �       Q�      �       u�      �       _�      �       p q "#��      8       _                         �       ]t��      8       ]t�                          P.      h.       Uh.      �.       V�.      �.       T�.      �.       �U��.      �.       U                    h.      �.       \�.      �.       U                 z.      �.       s `�H     "                 z.      �.      # s `�H     "#�����3$ �H     "                         F      F       UF      MF       VMF      VF       �U�VF      ?I       V                         F      0F       T0F      KF       w KF      VF       ��VF      ?I       w                            F      (F       Q(F      @F       \@F      VF       �Q�VF      
G       \
G      ?I       �Q�                  F      F       u�                          F      8F       0�8F      <F       P<F      UF       _UF      VF       r VF      ?I       _                �F      0I       _                   �F      G       P�H      0I       0�                  �F      �F        �F      0I       V                     �F      �F       P�F      �F       v��F      0I       ��                  �F      �H       S�H      0I       ��                      &G      4G       |�]G      �H       \�H      �H       |�                     �F      �F       0��H      �H       \�H      �H       |�                 �F      &G       	��                 ]G      pG       P                 ]G      pG       p�����3$ �H     "                        hG      �G       ^�G      H       XH      !H       ���H      �H       X                           pG      G       XG      �G       ���G      �G       X�G      �G       X�G      �G       P�G      �G       X                           H      H       TH      hH       ^hH      lH       TlH      uH       ^uH      yH       PyH      �H       ^                  �H      �H       P                  �H      �H       0�                 �      �       U                 �      �       T                        �0      1       U1      D2       �U�D2      [2       U[2      �2       �U�                              �0      
1       T
1      ?2       ]?2      D2       �T�D2      [2       T[2      �2       ]�2      �2       �T��2      �2       ]                            �0      �0       Q�0      C2       _C2      D2       �Q�D2      �2       _�2      �2       �Q��2      �2       _                              �0      1       R1      �1       ^�1      D2       �R�D2      [2       R[2      |2       ^|2      �2       �R��2      �2       ^                        �0      1       X1      D2       �X�D2      [2       X[2      �2       �X�                           1      1       | v �1      1       R1      ;2       | v �[2      �2       | v ��2      �2       | v �                      1      1       P1      D2       Q[2      �2       Q                         1      �1       | v "2~ "��1      ;2       | v "2�R"�[2      |2       | v "2~ "�|2      �2       | v "2�R"��2      �2       | v "2~ "�                              >1      2       R2      "2       rr�"2      "2        | v "?%v "| "1&q ?%q "1&�R"�"2      -2       p r "�[2      �2       R�2      �2        | v "?%v "| "1&q ?%q "1&�R"��2      �2       p r "��2      �2       R�2      �2       | v "?%v "| "1&q ?%q "1&~ "�                                  B1      �1       T�1      2       q r "�2      "2       q r ">�"2      ;2      # | v "?%v "| "1&q ?%q "1&q "�R"�[2      |2       T|2      �2       q r "��2      �2      # | v "?%v "| "1&q ?%q "1&q "�R"��2      �2       T�2      �2      " | v "?%v "| "1&q ?%q "1&q "~ "�                                 B1      N1       r ?�N1      �1       P�1      �1       r ?��1      �1       s x ��1      2       ^[2      b2       Pb2      |2       r ?��2      �2       P�2      �2       r ?��2      �2      " | v "?%v "| "1&q ?%q "1&~ "?�                                 K1      i1      	 @r ?�i1      �1       X�1      2       P[2      q2       Xq2      |2      	 @r ?��2      �2      	 @r ?��2      �2       X�2      �2      	 @r ?��2      �2      % @| v "?%v "| "1&q ?%q "1&~ "?�                        K1      �1       U�1      2       [[2      |2       U�2      �2       U                           K1      �1       @u ��1      �1       Z�1      �1       @u ��1      2       T[2      |2       @u ��2      �2       @u �                               K1      2       0�2      2       P"2      D2       P[2      w2       0�w2      �2       P�2      �2       P�2      �2       0��2      �2       P                     �1      �1       q ?��1      �1       Z�2      �2       q ?�                         �0      �0       @��0      :2       SD2      [2       @�[2      �2       S�2      �2       S                             =       U=      �       �U��      �       U�      �       �U�                             =       T=      �       �T��      �       T�      �       �T�                         =       0��      �       0�                           =       b�=      �       Y�      �       b�                             =       Q=      [       P^             P�      �       Q                        o      x       Rx      �       r/��      �       R�      �       rQ�                  C      �       T                     C      O       q t �O      k       Rk      �       u q t q t 0-( �                      p      �       T�             u�(             T                       �      �       Q�      �       t0�             u�(#0             Q                       �      �       R�      �       r 4!��      �       R�             Q             R                         �      �       0��      �       p ���      �       P�             u�(             P                 p             U                 p      �       T                    �      �       U�      n       �U�                    �      `       T`      n       �T�                    �             Q      n       �Q�                     �      �       q ����
�	u "#H��             q ����
�	�U"#H�      n       �Q����
�	�U"#H�                  �      n       Y                                 S      n       ��                         `       �Q����
88t "#P�`      n       �Q����
88�T"#P�                         `       �Q����
88t "#P`             �Q����
88�T"#P                      <      I       PI      x       Qx      n       ��                        �       0�                          �       0��      T       _                            �       ���      ;       ]>      T       ]                   �      B       PB      T       pH�                   �      �      
 q 2 $0.��      >       p0�2 $0.�                 �      >      ' y�8$8& $�Q����
�	�U"#h� $)�                     
             t { �             Q3      >       Q                        >       [                              Q                         $       Q$      $      
 q r "#���                        $       q ?&�$      $       R                      )       �Q����
88t "#P�                      )       t� ��-(�-� �                   '      )       P)      )      
 p q "#���                  '      )       p ?&�)      )       Q                        �"      #       U#      #       S#      "#       U"#      ##       �U�                        �"      #       T#      #       V#      "#       T"#      ##       �T�                         !      {!       U{!      �"       �U��"      �"       U�"      �"       �U�                         !      {!       T{!      �"       �T��"      �"       T�"      �"       �T�                     !      B!       QB!      �"       �Q�                    $!      �"       _�"      �"       _                    $!      �"       ]�"      �"       ]                         $!      B!       q ����
88u "#P�B!      {!       �Q����
88u "#P�{!      �"       �Q����
88�U"#P��"      �"       �Q����
88u "#P��"      �"       �Q����
88�U"#P�                     c!      {!       0�{!      �"       \�"      �"       \                       {!      �!      ! | ����8�Q����
88"�U"#���!      �!      ! |����8�Q����
88"�U"#���!      �"      ! | ����8�Q����
88"�U"#���"      �"      ! | ����8�Q����
88"�U"#��                   �!      "       p q "#��@& $ &�"      )"        s �r  $ &v q "#��@& $ &�                      ."      4"       p q �4"      �"       R�"      �"       R                                       ."      4"       p q �4"      N"       RN"      ^"       Q^"      r"       Pr"      r"       Rr"      {"       q p �{"      ~"       Q~"      �"       sp ��"      �"       P�"      �"       P�"      �"       p 	���"      �"       P�"      �"       p �                6"      ?"       _r"      �"       _                 6"      ?"       Rr"      {"       q p �                      ="      ?"       P?"      ?"      
 p q "#����"      �"       Q�"      �"      
 p q "#���                    ="      ?"       p ?&�?"      ?"       Q�"      �"       q ?&��"      �"       P                 �!      �!       _                 �!      �!       P                   �!      �!       Q�!      �!      
 q r "#���                  �!      �!       q ?&��!      �!       R                �!      �!       _                �!      �!       R                  �!      �!       Q�!      �!      
 q t "#���                  �!      �!       q ?&��!      �!       T                �!      �!       _                  �!      �!       P�!      �!      
 p q "#���                  �!      �!       p ?&��!      �!       Q                        ��      ��       U��      ˀ       Vˀ      ΀       �U�΀      ��       V                        ��      ��       T��      Ȁ       SȀ      ΀       �T�΀      ��       S                    ��      ̀       \΀      ��       \                        �z      �z       U�z      �|       ^�|       }       �U� }      �       ^                    �z      �z       T�z      �       ��x                         E{      E{       0�E{      �|       ��x�|      �|       ��x�#��|      �|       P�|      �|       ��x }      �       ��x                       E{      E{       0�E{      �|       ��x }             ��x             ��x�#�      �       ��x                               E{      E{       1�E{      �{       \�{      �|       ��x�|      �|       \ }       }       \ }      }       0�}      z}       ��xz}             \      �       \                     L~      W~       ��x#������8��x"#��W~      �~       { ����8��x"#��      -       ��x#������8��x"#��u      �       { ����8u "#��                  �{      �{       P                      E{      E{       PE{      �|       ��x }      �       ��x                                �{      �{       q��q���q���q����{      �{       u�#��u�#���Y��T���{      �{      & ��x#�#����x#�#���Y��T���{      �|      0 ��x#�#����x#�#���Y����x#�#����|      �|      : ��x#�#����x#�#�����x#�#�����x#�#���}      z}      0 ��x#�#����x#�#���Y����x#�#���            : ��x#�#����x#�#�����x#�#�����x#�#����      �       q��q���q���q���                 �z      �z       u                     �z      �z       p�z      {       S                      �z      �z       s 3$��H     "��z      �|       V }      �       V                     �z      �z       P�z      �|       _ }      �       _                            {      �{       S�{      �{       P�{      �|       S }      �}       S             S�      �       S                     L~      W~       ��x#������8��x"#��W~      �~       { ����8��x"#��      -       ��x#������8��x"#��u      �       { ����8u "#��                     L~      W~       ��x#������8��x"#��W~      �~       { ����8��x"#��      -       ��x#������8��x"#��u      �       { ����8u "#��                 �{      �{       T                        �{      �{       0��{      �|       R}      z}       R�      �       0�                                �{      �{       	���{      >|       QA|      n|       Qq|      �|       Q}      7}       Q:}      g}       Qj}      z}       Q�      �       	��                    �{      �{       0��      �       0�                        �{      �{       0��{      (|       P}      }       P�      �       0�                        �{      |       T|      L|       u�]|      �|       u�}      z}       T                            (|      L|       P]|      |       P}      :}       P:}      >}       p�P}      j}       Pj}      n}       p�                �{      �{       0�                �{      �{       _                �{      �{       ^                �{      �{       ~�                  �{      �{       T                 �~      �~       { ����8��x"#�                 �~      �~       { ����8��x"#�                 �~      �~       p r -�                      z}      �}       1��}      �}       X�}      �}       x�                 �}      �}       x ����x����3$p "                      �}      ~       1�~      ;~       U;~      ?~       u�                 +~      /~       u ����u����3$p "                 �z      �z       P                �|      �|       _                �|      �|       ��x                 �|      �|       ��x#�                        Pw      �w       U�w      Pz       VPz      Yz       �U�Yz      �z       V                        Pw      �w       T�w      �x       ^�x      �y       �T��y      �y       ^�y      �z       �T�                      4x      dx       P�x      �x       P�x      �x       P                    �w      x       0�x      �y       _�y      �y       0�kz      �z       _                           �x      �y       S�y      �y       s��y      �y       0��y      Bz       1�Bz      Yz       2�Yz      bz       0�bz      kz       1�kz      �z       S                 �w      �z       ���~�                	   �w      �w       P�w      �w       v                 
   �w      �w       p�����3$ �H     "�w      �w       v #�����3$ �H     "                    �w      �w       P�w      �x       \�y      �y       \                       �w      
x       S
x      #x       P#x      Cx       S�y      �y       S                x      x       0�                x      x       \                x      x       V                x      x       v�                  x      x       _                   �x      �y       s  $ &
88v "#P�kz      �z       s  $ &
88v "#P�                   �x      �y       s  $ &
�	� "
8��kz      �z       s  $ &
�	� "
8��                    �x      iy       Pkz      �z       P                        y      `y       U`y      wy       |� � $ &54$|� "�wy      ~y       |�l� $ &54$|�l"�kz      �z       U                          $y      @y       Q@y      Dy       p Dy      Sy       pPkz      oz       Qoz      �z       p                   xz      �z       Q                       �y      �y       v� ��y      Pz       v�� �Pz      Yz       �U#�q�Yz      bz       v� �bz      kz       v�� �                          �y      	z       R	z      z       v�z      Fz       Rbz      iz       Riz      kz       v�                �w      �w       ^                 �w      �w       X                 �w      �w       P                x      $x       \�y      �y       \                x      $x       ^�y      �y       ^                  x      #x       ~��y      �y       ~�                   �x      �y       ]kz      �z       ]                 �x      �x       P                  uw      �w       X                    uw      �w       ���}��w      �w       ]                              9        U9       �       ���      �       U                                  9        Q9       l       ^l      ~       �Q�~      �       ^�      �       Q                                9        1��       �        1��      �       y��      �       U�      �       1�                  �       �        V�      �       V                            �       �        0��              V0      5       U5      =       V=      F       PF      P       p�P      l       P~      �       V                    �       l       \~      �       \                    �       �        0��              P~      �       0�                      M       S       	 �Y�p�h       |        �Y�U�|       �       	 �Y�p�                                    �.      /       Q/      _/       �Q�_/      �/       Q�/      �/       �Q��/      �/       Q�/      �/       �Q��/      �/       Q�/      "0       �Q�"0      =0       Q=0      �0       �Q�                              �.      �.       R�.      _/       �R�_/      c/       Rc/      n/       r �n/      �/       �R��/      �/       R�/      �0       �R�                 �.      �0       ���  �                 �.      �0       ���  �                             �.      P/       T_/      �/       T�/      �/       u����/      �/       T�/      0       T"0      =0       Tg0      �0       T                                     �.      /       q ����
88t "#P�/      P/       �Q����
88t "#P�_/      �/       q ����
88t "#P��/      �/       �Q����
88t "#P��/      �/       �Q����
88u "
P8��/      �/       q ����
88t "#P��/      �/       �Q����
88t "#P��/      �/       q ����
88t "#P��/      0       �Q����
88t "#P�"0      =0       q ����
88t "#P�g0      �0       �Q����
88t "#P�                                                                     �.      P/       RP/      ^/       P^/      _/       q �_/      �/       R�/      �/       Q�/      �/       P�/      �/       R�/      �/       Q�/      �/       P�/      �/       Q�/      �/       P�/      �/       R�/      �/       P�/      �/       p 	���/      
0       R
0      0       P0      0       Q0      "0       P"0      =0       R=0      D0       PD0      H0       pp�H0      ^0       P^0      b0       Qb0      g0       Pg0      g0       Rg0      }0       P}0      �0       �Q����
88t "#p�0      �0       R�0      �0       rJ�                           �.      �.       0��.      _/       [_/      c/       0�c/      i/       1�i/      �/       [�/      �/       0��/      �0       [                                   �.      /      
 q  $@L$)�/      _/       �Q $@L$)�_/      �/      
 q  $@L$)��/      �/       �Q $@L$)��/      �/      
 q  $@L$)��/      �/       �Q $@L$)��/      �/      
 q  $@L$)��/      "0       �Q $@L$)�"0      =0      
 q  $@L$)�=0      �0       �Q $@L$)�                      �/      0       Q�0      �0       Q�0      �0       q*�                  3      Q3       T                  3      Q3       U                 3      Q3       Q                 3      Q3       R                                    `3      �3       Q�3      �3       P�3      Z4       �Q�Z4      d4       Qd4      w4       Pw4      �4       �Q��4      �4       Q�4      �4       P�4      �4       Q�4      l6       �Q�                                                  `3      =4       R=4      Z4       �R�Z4      w4       Rw4      �4       �R��4      �4       R�4      �4       �R��4      �4       R�4      5       �R�5      "5       R"5      |5       �R�|5      �5       R�5      �5       �R��5      �5       R�5      �5       �R��5      6       R6      16       �R�16      S6       RS6      l6       �R�                                          `3      =4       X=4      Z4       �X�Z4      w4       Xw4      �4       �X��4      �4       X�4      5       �X�5      "5       X"5      |5       �X�|5      #6       X#6      16       �X�16      F6       XF6      [6       �X�[6      l6       X                                `3      �3       Y�3      Z4       �Y�Z4      w4       Yw4      �4       �Y��4      �4       Y�4      �4       �Y��4      �4       Y�4      l6       �Y�                           `3      H4       TZ4      s4       T�4      �4       T�4      �4       u��~�5      "5       T|5      l6       T                                       `3      �3       q ����
�Gt "#P��3      �3       p ����
�Gt "#P��3      H4       �Q����
�Gt "#P�Z4      d4       q ����
�Gt "#P�d4      s4       p ����
�Gt "#P��4      �4       q ����
�Gt "#P��4      �4       p ����
�Gt "#P��4      �4       q ����
�Gt "#P��4      �4       �Q����
�Gt "#P��4      �4       �Q����
�Gu "
�G�5      "5       �Q����
�Gt "#P�|5      l6       �Q����
�Gt "#P�                                                   `3      �3       R�3      �3       SH4      V4       RV4      Y4       p �Z4      d4       Rx4      �4       P�4      �4       R�4      5       P5      5       R5      "5       S"5      C5       PC5      Z5       Rn5      w5       Pw5      |5       R�5      �5       R�5      �5       P)6      ,6       s x "�,6      16       SS6      V6       s x �V6      [6       S                       `3      �3       0��3      �3       1��3      R4       VZ4      d4       0�d4      l6       V                                   `3      �3       q  $@L$)���3      �3       p  $@L$)���3      Z4       �Q $@L$)��Z4      d4       q  $@L$)��d4      w4       p  $@L$)��w4      �4       �Q $@L$)���4      �4       q  $@L$)���4      �4       p  $@L$)���4      �4       q  $@L$)���4      l6       �Q $@L$)��                                  �3      �3       q p ��3      =4       Q|5      �5       Q�5      �5       P�5      6       Q6      ,6      6 u s �Q����
�Gt "#ps �Q����
�Gt "#p0-( �16      66       Q66      V6      6 u s �Q����
�Gt "#ps �Q����
�Gt "#p0-( �[6      l6       P                           
4      =4       0��5      #6       0�#6      )6       Q)6      )6       X)6      16       x �16      S6       0�S6      S6       QS6      [6       X                         +4      =4       P�5      6       P6      16       t#�#�
���16      I6       PI6      S6       t#�#�
���                     C5      I5       r q �I5      L5       r s �L5      n5       P                    �6      �6       U�6      7       �U�                          �6      �6       T�6      �6       S�6      �6       �T��6      	7       S	7      7       �T�                          �6      �6       Q�6      �6       V�6      �6       �Q��6      
7       V
7      7       �Q�                    �6      �6       P�6      7       �\                  �6      7       �U�                    �6      
7       V
7      7       �Q�                    �6      	7       S	7      7       �T�                        7      C7       UC7      A:       _A:      B:       �U�B:      �>       _                        7      $7       T$7      57       P57      �9       \�9      �>       �T�                    �7      3:       0�B:      �>       0�                    7      57       P57      �7       \                   7      C7       UC7      �7       _                               7      57       p ����
�	u "#H�57      C7       | ����
�	u "#H�C7      �9       | ����
�	 "#H��9      A:       �T����
�	 "#H�A:      B:       �T����
�	�U"#H�B:      :;       | ����
�	 "#H�:;      V>       �T����
�	 "#H�V>      �>       | ����
�	 "#H�                  <7      _7       S                    ?7      O7       v  $ &Ps "�O7      _7      	 p Ps "�                  D7      O7       P                  Z7      �7       S                    g7      �7       Q�7      �7       q� �7      �7       Q                  k7      �7       Y                    q7      �7      	 r 3
����7      �7       R                    �7      �7      	 u 3
����7      �7       R                         �7      �9       \�9      3:       �T�B:      :;       \:;      V>       �T�V>      �>       \                   �7      3:       _B:      �>       _                       �7      �9       \B:      �:       \V>      q>       \�>      �>       \                       �7      �9       _B:      �:       _V>      q>       _�>      �>       _                         �7      �9       | ����
�	 "#H��9      3:       �T����
�	 "#H�B:      :;       | ����
�	 "#H�:;      V>       �T����
�	 "#H�V>      �>       | ����
�	 "#H�                   �7      �7       | ����
�	 "#PB:      Q:       | ����
�	 "#P                   �7      �7      0 | ����
�	 "#H� $ &P| ����
�	 "#P"�B:      Q:      0 | ����
�	 "#H� $ &P| ����
�	 "#P"�                   �7      �7       | ����
�	 "#hB:      Q:       | ����
�	 "#h                          8      9       Q9      �9       RQ:      �:       SV>      q>       R�>      �>       R                          88      9       Rb9      �9       Q\:      �:       QV>      q>       Q�>      �>       Q                   �7      �7       �(#H�����8&�B:      Q:       �(#H�����8&�                          �7      �7       T�7      �9       PQ:      �:       PV>      q>       P�>      �>       P                    W8      Z8       x t  $ &�Z8      �8      	 x  $ &�                 `8      `8       q�0$0&�`8      �8       q�0$r�0$+( 0$0&�                 `8      `8       q�0$0&�`8      �8       q�0$r�0$-( 0$0&�                  �8      �8       T                          9      -9       X19      �9       XQ:      �:       XV>      q>       X�>      �>       X                      �9      �9       UV>      q>       U�>      �>       U                    �9      �9       TV>      q>       T                      �9      �9       [�9      �9       [V>      q>       [                       �9      3:       �T��:      :;       \:;      V>       �T�q>      �>       \                     �9      3:       _�:      V>       _q>      �>       _                      �:      �:       S�:      :;       ��q>      �>       ��                       �9      3:       0��:      �=       0��=      �=       Pq>      �>       0�                          �:      �:       S�:      ,;        ,;      :;       ��q>      �>        �>      �>       ��                     �:      !;       | ����
88r "#P�!;      ,;       | ����
88�("#P�q>      �>       | ����
88r "#P�                    �:      :;       Sq>      �>       S                        �:      �:       U�:      :;       ��q>      �>       U�>      �>       ��                                �9      1:       R;      �<       S�<      �<       T�<      �<       T�<      �<       R�<      �<       S�<      �=       R�=      V>       S�>      �>       S                    �:      ,;       T�>      �>       T                                 �9      3:       ^
;      ;       p q "#��@& $ &�;      ;       ~  $ &u q "#��@& $ &�;      V>       ^�>      �>       ~  $ &u q "#��@& $ &��>      �>       ~  $ &��q "#��@& $ &��>      �>      + ~  $ &��~  $ &��?&"#��@& $ &��>      �>       P�>      �>       ^                  �<      �<       P                    �9      1:       V�<      �=       V                       �9      1:       P�<      �<       P�<      �<       Q�<      �=       P                     �9      1:       X�<      �<       0��<      �=       X                     �9      1:       [�<      �<       0��<      �=       [                    =      =       1�y=      �=       0�                      =      V=       Q�=      �=       Q�=      �=       Q                    =      V=       T�=      �=       T�=      �=       T                    =      E=       Y�=      �=       Y                  @=      E=       U                 �:      
;       T                 �:      
;       ^                   ;      
;       P
;      
;      
 p q "#���                  ;      
;       p ?&�
;      
;       Q                      :;      x;       0�x;      /<       Q3<      e<       Q                      :;      x;       
���x;      �;       U�;      e<       U                  :;      x;       0�                   x;      �;       T�;      6<       T                    x;      �;       R�;      A<       R                    x;      �;       [�;      A<       [                    �;      �;       Z�;      A<       Y                     �;      �;       0��;      <       P%<      A<       P                      �;      �;       y <      <       Z<      %<       y                    ,>      2>      	 p 0$0&�2>      E>       q �0$0&�                      2>      9>       P9>      A>      
 p r "#���A>      E>       P                   2>      9>       p ?&�9>      E>       R                          �>      ?       U?      (?       S(?      s?       �U�s?      �?       S�?      �?       �U�                          �>      d?       Td?      l?       \l?      s?       �T�s?      {?       T{?      �?       \                    �>      ?       Q?      ?       R                        �>       ?       R ?      ?       P?      (?       Qs?      �?       Q                           !?      7?       S7?      ;?       s��;?      [?       S[?      _?       s��_?      i?       S�?      �?       S                                (?      @?       PD?      S?       PS?      W?       s8W?      d?       P�?      �?       Q�?      �?       Q�?      �?       s8�?      �?       Q                 ?      ?       r8                   ?      (?       q8s?      �?       q8                    ?      p?       ^s?      �?       ^                      ?      d?       Us?      ~?       U~?      �?       q0                    ?      r?       _s?      �?       _                      ?      d?       Rs?      �?       R�?      �?       ��                  �?      �?       P                   �?      �?       q v ��?      �?       Q                   �?      �?       Q�?      �?      
 q t "#���                  �?      �?       q ?&��?      �?       T                          @C      hC       RhC      �C       \�C      �D       �R��D      �D       \�D       F       �R�                        [C      D       V�D      �D       V�D      �D       V8E      bE       V                    dC      �C      ' s 
��@$����@>$����+( ������D      �D      ' s 
��@$����@>$����+( �����                      lC      nC       PnC      �D       ]�D       F       ]                   �C      �C       | @$������C      �C       �R@$�����                      �C      �C       U�C      �C       U8E      bE       U                        �C      BD       T�D      �D       T]E      bE       T}E      �E       T                          �D      �D       U�D      �D       U3E      8E       UxE      }E       P�E       F       U                      �C      �C       r t #��C      �C       R8E      CE       R                          ~C      6D       P�D      �D       P�D      �D       P8E      bE       P}E      �E       P                              �C      BD       X�D      �D       X�D      �D       v(�D      �D       X8E      bE       X}E      �E       X�E       F       ��                       �C      D       v,�D      �D       v,�D      �D       v,8E      bE       v,                       �C      D       v0�D      �D       v0�D      �D       v08E      bE       v0                       �C      D       v4�D      �D       v4�D      �D       v48E      bE       v4                       �C      D       v8�D      �D       v8�D      �D       v88E      bE       v8                          �C      ED       _�D      �D       _�D      E       _8E      bE       _}E      �E       _                       �C      D       v� �D      �D       v� �D      �D       v� 8E      bE       v�                  �C      �C       ]                     �C      �C       | @$��C      �C       \�C      �C       �R@$�                      �C      �C       \�C      �C      
 r | "#����C      �C       R                     �C      �C       | ?&��C      �C       R�C      �C       | ?&�                  ED      �D       _                  MD      \D       | p �                    �D      �D       Q�D      8E       ��                  �D      E       | p �                8E      NE       S                8E      NE       U                   GE      NE       RNE      NE      
 r t "#���                  GE      NE       r ?&�NE      NE       T                    �E      �E       Q�E       F       ��                  �E      �E       | p �                            PW      lW       UlW      �W       V�W      �W       �U��W      OX       VOX      VX       �U�VX      �Z       V                  PW      sW       T                                PW      ^W       Q^W      �W       \�W      �W       �Q��W      QX       \QX      VX       �Q�VX      �X       \�X      �Y       �Q��Y      �Z       \                    PW      cW       RcW      �Z       �R�                            gW      lW       UlW      �W       V�W      �W       �U��W      OX       VOX      VX       �U�VX      �Z       V                    �W      �W       q��W      �W       Q                   �W      �W       P�W      �W       P                   ?X      QX       \QX      VX       �Q�                            �W      ?X       QVX      tX       Q�X      �X       Q�Y      ,Z       QLZ      `Z       QiZ      pZ       Q                        �W      ?X       \VX      �X       \�X      �Y       �Q��Y      �Z       \                                            �W      :X       P:X      ?X       �T�VX      }X       P}X      �X       �T��X      �X       P�X      �Y       �T��Y      Z       PZ      %Z       �T�%Z      3Z       P3Z      LZ       �T�LZ      `Z       P`Z      iZ       �T�iZ      wZ       PwZ      �Z       �T�                    �W      ?X       VVX      �Z       V                    �X      �X       P�X      �X       S                   :Y      ?Y       ~d�?Y      �Y       \                  CY      �Y       Q                   CY      �Y       |�Y      �Y       Z                  HY      �Y       P                   HY      �Y       |�Y      �Y       Y                   HY      �Y       |�Y      �Y       R                   HY      �Y       |�Y      �Y       X                   HY      �Y       |�Y      �Y       T                 HY      �Y       |                  �X      ?Y       \                 5X      ?X       \                 mX      �X       \                 Z      %Z       \                   %Z      LZ       \`Z      iZ       \                    4Z      LZ       P`Z      iZ       P                 iZ      �Z       \                  xZ      �Z       P                            �Z      ~\       U~\      m]       Sm]      u]       Uu]      �]       �U��]      �]       S�]      H^       U                          �Z      �\       T�\      �]       ���]      �]       �T��]      �]       ���]      H^       T                            �Z      �Z       Q�Z      k\       Sk\      �]       ���]      �]       �Q��]      �]       ���]      H^       S                        �Z      �Z       R�Z      �\       ���\      �]       �R��]      H^       ��                         �Z      �\       t� ��\      �]       ��#H��]      �]       �T#H��]      �]       ��#H��]      H^       t� �                     �Z      [       Q[      �\       t0�]      H^       t0                    �Z      �]       \�]      H^       \                  �Z      �[       P                 �Z      [       1�                     �Z      �Z       Y�Z      �\       t,�]      H^       t,                      �Z      �\       ^�\      �]       ���]      H^       ^                          �Z      [       R[      �\       R�\      �]       ���]      �]       ���]      H^       R                            �Z      [       R[      [       V[      �\       V�\      �]       ���]      �]       ���]      H^       V                      �\      �\       _,]      _]       _�]      �]       _                    �\      �\       ^�\      ,]       ~ :��]      �]       ^                            �Z      �Z       Q�Z      ]       w ]      ]       ��]      �]       w �]      �]       ���]      H^       w                     [      2[       Q2[      5[       x��0$0&�                 /[      s[       \                 /[      s[       R                          A[      Q[       QQ[      Y[      
 q y "#���Y[      `[       [`[      h[       q ?&q "#���h[      s[      # |  $ &��|  $ &��?&"#���                       A[      Q[       q ?&�Q[      \[       Y\[      h[       q ?&�h[      s[       |  $ &��?&�                �[      �[       \                �[      �[       V                 �[      �[       @��[      �[       8�^      0^       @�0^      H^       8�                  �\      ,]       T                         �\      ]       q p r "#��@&�]      ]       q t  $ &��r "#��@&�]      ]      ( q t  $ &��t  $ &��?&"#��@&�]      ]       Q]      ,]      ( v t  $ &��t  $ &��?&"#��@&�                     �\      �\       s �\      �\       s  s� "��\      ,]       V,]      A]       s A]      W]       s  s� "�W]      _]       T�]      �]       V                         �\      �\       s�\      ,]       ],]      W]       sW]      _]       ]�]      �]       ]                �\      �\       T                �\      �\       ��                   �\      �\       P�\      �\      
 p r "#���                  �\      �\       p ?&��\      �\       R                  d]      �]       R                  h]      �]       T                    h]      r]       r | �r]      z]       Pz]      �]       U                h]      �]       ��                   ~]      �]       P�]      �]      
 p q "#���                  ~]      �]       p ?&��]      �]       Q                �]      �]       U                �]      �]       ��                  �]      �]       P�]      �]      
 p q "#���                  �]      �]       p ?&��]      �]       Q                    P^      ]^       U]^      g       �U�                            P^      X^       TX^      �^       _�^      �_       �T��_      �_       _�_      �_       �T��_      @`       _@`      g       �T�                    P^      x^       Qx^      g       ��}                    P^      j^       Rj^      t^       ��}                          }^      �^       P�^      �^       ��}�_      �_       ��}�_      �_       P`      .`       P                      �^      �_       �U��_      `       �U�6`      g       �U�                      �^      �_       ��}�_      `       ��}6`      g       ��}                      �^      �_       ��}�_      `       ��}6`      g       ��}                          �^      �^       _�^      �_       �T��_      `       _6`      @`       _@`      g       �T�                        �^      �^       0��_      �_       0��_      `       P6`      @`       0�                                  �^      �^       Z�^      �^       \�^      �^       \�^      _       0��b      �b       \}c      �c       |��c      �c       2��c      td       0�>e      fe       0�                          �^      (_       \(_      �_       ��~@`      �`       ��~�b      �b       \>e      fe       \(f      ;f       ��~                                           �^      (_       [(_      �_       ^@`      �`       ^�`      �a       _�a      b       [b      �b       _�b      �b       [�d      �d       _�d      �d       [�d      e       _e      9e       [>e      f       [f      (f       _(f      ;f       ^;f      lf       _lf      g       [                    �^      _       | ����
�	{ "#H��b      �b       | ����
�	{ "#H�>e      fe       | ����
�	{ "#H�                               �^      (_       S(_      �_       ��~@`      �b       ��~�b      �b       S�d      �d       ��~�d      9e       ��~>e      fe       Sfe      f       ��~f      g       ��~                                       _      �_       V@`      n`       Vn`      pa       \pa      nb       Vnb      zb       \zb      �b       V�b      �b       V�d      �d       V�d      e       \e      9e       V>e      f       Vf      g       V                 >e      fe       p X�                                        _      �_       S@`      U`       S�`      Ta       STa      Ya       ��~Ya      �a       S�a      b       Pb      �b       S�b      �b       S�d      �d       S�d      *e       S>e      �e       S�e      �e       ��~�e      �e       Sf      lf       S                                 _      (_       0�(_      �_       _@`      ``       _``      >a       ��~>a      Ta       STa      �a       ��~nb      zb       ��~�b      �b       0��d      9e       ��~>e      fe       0�(f      ;f       _                               _      �_       0�@`      �`       0��`      �a       ��~nb      zb       ��~�b      �b       0��d      9e       ��~>e      fe       0�(f      ;f       0��f      g       Q                                   _      �_       0�@`      �`       0��`      �a       ��~�a      �a       Y�a      �a       y��a      b       Ynb      ub       ��~�b      �b       0��d      9e       ��~>e      fe       0��e      �e       Y(f      ;f       0�                                _      �_       0�@`      �`       0��`      Ga       VYa      Ya       1�Ya      ka       Vnb      zb       V�b      �b       0��d      �d       Ve      e       1�>e      fe       0�(f      ;f       0�                                           _      �_       0�@`      �`       0��`      �`       Z�`      �`       ��~�`      8a       Z8a      Ya       ��~Ya      �a       Znb      zb       Z�b      �b       0��d      �d       Z�d      �d       ��~�d      �d       Z�d      e       ��~e      e       Pe      9e       Z>e      fe       0�(f      ;f       0�                     (_      C_       Rn_      �_       R�_      �_       P                       (_      N_       Sn_      �_       0��_      �_       Q(f      ;f       S                          (_      N_       Qr_      �_       Q�_      �_       S�_      �_       \(f      6f       Q6f      ;f       s0                 �_      �_       Q                 �_      �_       \                �_      �_       ��~                �_      �_       ^                   �_      �_       |q��_      �_       R                 �_      �_       P                        �`      �`       ]�`      ba       ]nb      zb       ]�d      e       ]                 �`      �`       ]                 �`      �`       S                �`      �`       ��~                �`      �`       _                   �`      �`       s}��`      �`       R                  �`      �`       P                 �d      e       ]                 �d      e       S                �d      e       ��~                �d      e       _                   �d      �d       s}��d      �d       R                   e      e       P                    }e      �e       R�e      �e       ��~lf      �f       R                        �e      �e       U�e      �e       Ulf      �f       U�f      g       U                      �e      �e       X�e      �e       Xlf      g       X                        �e      �e       Q�e      �e       p r�lf      tf       p r�tf      �f       ur�                   �e      �e       Zlf      g       Z                       �e      �e       q z ��e      �e       Qlf      �f       Q�f      �f       } uz ruz r0-( �                �a      �a       [                �a      �a       T                �a      �a       P                          &b      *b       S*b      nb       Pzb      �b       Pf      f       P;f      Jf       P                        Db      nb       Rzb      �b       Rf      (f       R;f      _f       R                 \b      nb       _                 \b      nb       P                 \b      nb       S                 �b      �b       _                 �b      �b       R                 �b      �b       S                       �b      ]c       \�c      �c       \�d      �d       \9e      >e       \f      f       \                       �b      ]c       [�c      �c       [�d      �d       [9e      >e       [f      f       [                    �b      �b       | ����
�	{ "#H��d      �d       | ����
�	{ "#H�9e      >e       | ����
�	{ "#H�f      f       | ����
�	{ "#H�                      �b      �b       S�d      �d       S9e      >e       | ����
�	{ "#`f      f       | ����
�	{ "#`                        �b      ]c       V�c      �c       V�d      �d       V9e      >e      0 | ����
�	{ "#X� $ &X| ����
�	{ "#`"�f      f      0 | ����
�	{ "#X� $ &X| ����
�	{ "#`"�                   �b      ]c       S�c      �c       S                 �b      �b       U                    �b      ]c       P�c      �c       P                  c      Tc       R                  c      Tc       Q                    �c      �c       Q�c      �c       Q                 3d      td       0�                 3d      td       [                  3d      td       X                  3d      Cd       ��~                   3d      Cd       QCd      td       {0                  >d      td       T                     >d      Qd       QQd      od       q��od      td       Q                  Cd      Qd       q�0$0&�Qd      \d       qH�0$0&�                   Ud      \d       P\d      \d      
 p r "#���                  Ud      \d       p ?&�\d      \d       R                       g      5g       U5g      ng       Sng      ]u       �U�                                               g      (g       T(g      h       _h      &i       ]&i      j       _j      j       �T�j      �m       _�m      �n       ]�n      �n       _�n      ?o       ]?o      Lr       _Lr      �r       ]�r      �s       _�s      �s       ]�s      Nu       _Nu      ]u       ]                                   g      Jg       QJg      vg       ��~vg      j       �Q�j      *l       ��~*l      `m       �Q�`m      �m       ��~�m      Xt       �Q�Xt      �t       ��~�t      ]u       �Q�                                   g      Jg       RJg      vg       ��}vg      j       �R�j      *l       ��}*l      `m       �R�`m      �m       ��}�m      Xt       �R�Xt      �t       ��}�t      ]u       �R�                            Og      ^g       P^g      vg       ��}j      "j       ��}(j      *l       ��}`m      �m       ��}Xt      �t       ��}                        Wg      vg       ��}j      *l       ��}`m      �m       ��}Xt      �t       ��}                        Wg      vg       ��~j      *l       ��~`m      �m       ��~Xt      �t       ��~                                          Wg      h       _h      &i       ]&i      �i       _j      �m       _�m      �n       ]�n      �n       _�n      ?o       ]?o      Lr       _Lr      �r       ]�r      �s       _�s      �s       ]�s      Nu       _Nu      ]u       ]                            Wg      ng       Sng      �i       �U�j      �j       S�j      `m       �U�`m      �m       S�m      ]u       �U�                       fg      ng       0�(j      tj       0�tj      |j       Pm      �m       P�m      �m       0�                                        qg      �g       ^�g      �g       ~��g      �g       ^�g      �g       0��i      �i       ~��i      �i       2�*l      `m       ^�n      �n       ^?o      Ho       0��r      �r       ^�s      �s       ^�t      u       0�                      j      "j       ��}#P�(j      *l      	 ��}#���`m      �m       ��}#P�Xt      �t      	 ��}#���                   �j      *l       ��}Xt      �t       ��}                   �j      *l       _Xt      �t       _                   �j      *l       ��Xt      �t       ��                    �j      *l       UXt      �t       U                      �j      �j       P�j      *l       ��}Xt      �t       ��}                   �j      *l      	 ��}#���Xt      �t      	 ��}#���                   �j      �j       V�j      k       ��}#��                 k      =k       0�                     k      =k       0�=k      *l       \Xt      rt       \                       k      =k       0�=k      �k       ]�k      l       ]l      *l       YXt      rt       ]                      =k      �k       [�k      l       [l      *l       PXt      rt       [                       =k      Dk       RDk      Mk       r��Mk      *l       RXt      rt       r��                  ^k      *l       Z                  ek      *l       Y                 ek      *l       u�8$8& $�� $)�                                    �k      �k       t x ��k      �k       Q�k      �k       ~ t x t x 0-( ��k      �k       x t t x t x 0-( ��k      �k       Q�k      �k       t p ��k      �k       T�k       l      $ q u �0$0&p u �0$0&p 0-( � l      l      & q u �0$0&ru �0$0&r0-( �l      *l       P                   �k      �k       t x -��k      *l       u �0$0&x -�                    �k      �k       T�k       l      $ q u �0$0&p u �0$0&p 0-( � l      l      & q u �0$0&ru �0$0&r0-( �                   �k      l       Tl      l      
 p t "#���                  �k      l       t ?&�l      l       P                    �k      �k       Q�k      �k       ~ t x t x 0-( ��k      �k       x t t x t x 0-( �                   �k      �k       Q�k      �k      
 q ~ "#���                  �k      �k       q ?&��k      �k       ^                            �g      �g       0�Pl      `m       1��n      �n       1�?o      Ho       0��r      �r       1��s      �s       1�                                                �g      h       _h      &i       ]&i      Ai       _Pl      `m       _�m      �n       ]�n      �n       _�n      ?o       ]?o      9p       _�p      Lr       _Lr      �r       ]�r      �r       _�r      �s       _�s      �s       ]�s      Xt       _u      (u       _Nu      ]u       ]                          �g      �g       � �Pl      `m       ���n      �n       ��?o      Ho       � ��r      �r       ���s      �s       ��                      �g      �g       Uil      �l       T?o      Ho       U                                        �g      h       ]h      Ai       ��~|l      `m       ]�m      �n       ��~�n      �n       ]�n      ?o       ��~?o      Ho       ]Lr      �r       ��~�r      �r       ]�s      �s       ��~�s      �s       ]Nu      ]u       ��~                             0i      Ai       ��~X�Ho      �o       ��~X��r      �r       ��~X��r      s       p X�s      �s       ��~X�7t      Xt       p X�u      Nu       ��~X�                
                                      �g      �g       Uh      Ai       S�l      �l       T�l      `m       S�m      ?o       S?o      Ho       Uuo      �o       ��~�o      �o       Q�o      9p       s���p      �p       q� ��p      ,q       Q,q      �q       s���q      Lr       QLr      �r       S�r      �r       s���r      �r       S�s      �s       ��~�s      �s       S�s      7t       s��Nu      ]u       S                                                         �g      �g       0�h      i       _i      Ai       [|l      �l       0��l      `m       \�m      �n       _�n      �n       S�n      �n       \�n      ?o       _?o      Ho       0�uo      9p       [�p      �p       [�p      �p       Q�p      Lr       [Lr      �r       _�r      �r       [�r      �r       \�s      �s       [�s      �s       _�s      �s       \�s      t       [t      7t       ��~Nu      ]u       _                                        �g      h       0�h      Ai       ��~|l      `m       0��m      en       ��~jn      �n       ��~�n      �n       0��n      ?o       ��~?o      Ho       0�Lr      �r       ��~�r      �r       0��s      �s       ��~�s      �s       0�Nu      ]u       ��~                 |l      �l       �(                 |l      �l       �(#�����3$ �H     "                      �g      �g       0�|l      �l       0��l      �l       P?o      Ho       0�                            #h      �h       V�m      �n       V�n      ?o       VLr      �r       V�s      �s       VNu      ]u       V                   �h      �h       ~ "��m      �m       ~ "�                     �h      �h       vs��m      On       vs��n      6o       vs�                   �h      �h       ��~1&~ ""��m      �m       z 1&~ ""�                          �m      n       Rn      $n       q 	��$n      2n       z 1&~ "# 	��2n      Xn       T�n      ?o       X                    o      2o       Y2o      ?o       z ~ "# 	�p �                            n      n       q u �n      n       q t �n      Xn       U o      o       t u �o      o       t { �o      ?o       T                            n      $n       q r �$n      .n       Q.n      ?n       x z 1&r ~ "z 1&r ~ "0-( �o      o       r { �o      "o       r q �"o      ?o       R                    �m      n       Tn      9n        &p A-( �                    �m      n       Xn      9n        Jp A-( �                     jn      �n       vs�Lr      �r       vs�Nu      ]u       vs�                  cr      �r       ^                      kr      �r       R�r      �r       ~ 	���r      �r       Q                      qr      zr       ~ t �zr      �r       ~ q ��r      �r       T                    �r      �r       ~ r ��r      �r       ^                     zn      �n       &�Zr      tr       QNu      ]u       &�                     zn      �n       J�Zr      �r       UNu      ]u       J�                         �l      �l       Q5m      >m       0�Cm      Km       P�n      �n       Q�n      �n       s(�s      �s       s(                                 �l      �l       0��l      �l       S�l       m       Q$m      Cm       0�Cm      [m       V[m      `m       S�n      �n       0��n      �n       S�s      �s       0�                          �l      m       V,m      Cm       VCm      `m       S�n      �n       V�s      �s       V                       �l      �l       p 8��n      �n       p 8��s      �s       p 8��s      �s       s�8�                        �l      �l       r 8��l      �l       v�8��n      �n       r 8��s      �s       r 8�                   s      bs       U7t      Xt       ��~                      s      �s       XLt      Xt       Xu      (u       X                      &s      �s       TSt      Xt       Tu      (u       T                      8s      As       PAs      Ws       r u�Ws      bs       xu�                     8s      �s       S�s      �s       tx�u      (u       S                       8s      As       p s �As      Ss       PSs      Ws       y r s ur s u0-( �Ws      bs       y xs uxs u0-( �                    es      �s       Ru      (u       R                     �o      �o       
���o      �o       p u ��o      �o       P                 �o      �o       _                 �o      �o       R                 �o      �o       Q                      �p      Aq       P�q      3r       P�s      �s       P                   �q      r       q� �r      +r       R                    Ai      �i       ��}9p      cp       ��}�r      �r       0�(u      Nu       ��}                    Ai      �i       _9p      �p       _�r      �r       _(u      Nu       _                   Ai      bi       ��}�����
�	 "#H�9p      cp       ��}�����
�	 "#H��r      �r       � �(u      Nu       ��}�����
�	 "#H�                        Si      gi       PKp      lp       P�r      �r       P:u      Nu       P                        bi      �i       RZp      �p       R�r      �r       RIu      Nu       R                   bi      �i       Pcp      �p       P                      ti      �i       U�i      �i       p�i      �i       p@                 �i      �i       Q                    }i      �i       Q�i      �i       p�                   �i      �i       T                      tp      �p       U�p      �p       p�p      �p       p@                 �p      �p       Q                    }p      �p       Q�p      �p       p�                   �p      �p       T                   j      "j       0�`m      m       0�                   j      "j       ��}#h�`m      m       ��}#h�                   j      "j       V`m      m       V                     j      j       Uj      "j       _`m      m       _                    j      "j       P`m      em       Pm      m       P                 `m      m       0�                 `m      m       ��}#h�                 `m      m       V                 `m      m       _                 m      m       P                 Cj      tj       1�                 Cj      tj      	 ��}#���                 Cj      tj       V                   Cj      Gj       UGj      tj       _                  Hj      fj       Ptj      tj       P                 Lj      tj       1�                 Lj      tj      	 ��}#���                 Lj      tj       V                 Lj      tj       _                 tj      tj       P                 �t      u       0�                 �t      u       _                  �t      u       X                  �t      �t       ��~                   �t      �t       Q�t      u       0                  �t      u       T                     �t      �t       Q�t      �t       q���t      u       Q                  �t      �t       q�0$0&��t      �t       qH�0$0&�                   �t      �t       P�t      �t      
 p r "#���                  �t      �t       p ?&��t      �t       R                  `u      `u       R`u      cu       �R�                    pu      {u       U{u      �u       �U�                   pu      {u       u�{u      �u       �U#�                  �u      �u       P                    �u      �u       U�u      �u       �U�                    �u      �u       T�u      �u       �T�                   �u      �u       u��u      �u       U                        �      �       U�      �       V�      ��       �U���      ��       V                         �      �       0��      S�       ]S�      _�       1�_�      ��       ]��      ��       ]                         �      f�       1�f�      ~�       S~�      �       v8�      ��       �U#8��      ��       1���      ��       0�                          �      �       0��      S�       ^S�      a�       Pa�      ��       ^��      ��       ^                     �      �       P�      ��       \��      ��       \                       �       �       S �      &�       P&�      f�       S��      ��       S                 �      �       U                 �      �       P                   ?�      a�       _��      ��       _                "�      ?�       0�                    "�      /�       ���/�      >�       R>�      ?�       ���                "�      ?�       \                "�      ?�       V                 "�      >�       v�                  *�      ?�       _                f�      v�       \                 f�      u�       ��                    �      �       U�      *�       �U�                    �      �       T�      *�       �T�                    �      
�       Q
�      *�       �Q�                    �      �       R�      *�       �R�                      �      �       X�      (�       S(�      *�       �X�                 �      �       u�                     ��      )�       V)�      *�       P                      �      �       U�      b       w b      m       ��}                    �      �       T�      m       ��}                     �      �       Q�      �       ]�      [       ^                      �      �       R�      [       V[      m       �R�                     �      �       0��      �       _�      �       _                   �      �       Q�      [       ]                       �      �       0��      �       |��      �       \�             |�                     0      D       ��}�D      N       RN      O       ��}�                 0      O       ^                 0      O       ��}                 0      O       w                  �      �       2�                 �      �       U                 �      �       u�                 �      �       u� �                      0      D       UD      �       V�      �       �U�                      0      H       TH      �       \�      �       �T�                      0      H       QH      �       S�      �       �Q�                 c      }       W                 c      }       1�                 c      }       \                 c      }       V                 p      �       1�                 p      �       U                 ~      �       u�                 �      �       u� �                                        }       U}      �       ]�      �       �U��      �       U�             ]             �U�      O       UO      �       ]�      �       U                                    7       T7      �       V�             V      +       T+      �       V�      �       T�      �       V                                    7       Q7      �       \�             \      +       Q+      �       \�      �       Q�      �       \                                          G       RG      }       [}      �       �R��      �       [�             �R�      +       R+      a       [a      �       ���      �       R�      �       [                                        K       XK      �       ^�      �       �X��             ^             �X�      +       X+      �       ^�      �       X�      �       ^                           �       0��      �       P�      �       0��             P      �       0�                                     7       0�7      }       Z�      �       Z             0�      +       1�+      a       Za      �       ���      �       1��      �       3��      �       Z                   �      �       U�             U                       K      Z       0�Z      }       S�      �       S�      �       0�                                G      }       R�      �       R�      �       �+      =       R=      O       u O      a       } a      �       ��      �       R                           K      Z       XZ      }       Q�      �       Q�      �       P�      �       } �����32$x "<��      �       X                u      �       �M�
  �      �       �M�
                    u      �       [�      �       [�      �       ��                  u      }       u��      �       }�                  u      �       0��      �       0��      �       P                    y      �       P�      �       P                  �      �       �
  +      �       �
                        �      �       [�      �       �R�+      a       [a      �       ��                      �      �       U�      �       ]+      O       UO      �       ]                  �      �       0�+      �       0�                    �      �       R�      �       _+      �       _                    �      �       0��      �       P+      �       0�                   +      O       UO      �       ]                   +      a       [a      �       ��                 +      �       _                 +      a       P                   +      T       _T      a       Ra      �       ��                                    �:      �:       U�:      �:       V�:      �:       p��:      �:       �U��:      ;       V;      �;       p��;      �;       �U��;      �;       V�;      �;       p��;      �;       �U�                              �:      �:       T�:      �:       ]�:      �:       �T��:      K;       ]K;      �;       �T��;      �;       ]�;      �;       �T�                              �:      �:       Q�:      �:       \�:      �:       �Q��:      �;       \�;      �;       �Q��;      �;       \�;      �;       �Q�                              �:      �:       R�:      �:       S�:      �:       �R��:      T;       ST;      �;       �R��;      �;       S�;      �;       �R�                    �:      �:       X�:      �;       �X�                              �:      �:       Y�:      �:       ^�:      �:       �Y��:      �;       ^�;      �;       �Y��;      �;       ^�;      �;       �Y�                    �:      �:       P�:      ;       P                    �:      �:       Y�:      �:       ^                   �:      �:       X�:      �:       �X�                   �:      �:       U�:      �:       V                                   �:      �:       U�:      �:       V�:      �:       p��:      �:       �U��:      ;       V;      �;       p��;      �;       �U��;      �;       V�;      �;       p��;      �;       �U�                                   �:      �:       U�:      �:       V�:      �:       p��:      �:       �U��:      ;       V;      �;       p��;      �;       �U��;      �;       V�;      �;       p��;      �;       �U�                  �:      �:       X                   �:      �:       P�:      �:       u                   �:      �:       p ����Hu"H��:      �:       u�����Hu"H�                       �:      �;       ^�;      �;       �Y��;      �;       ^�;      �;       �Y�                         �:      �;       S�;      �;       s��;      �;       S�;      �;       S�;      �;       �R�                       �:      �;       \�;      �;       �Q��;      �;       \�;      �;       �Q�                       �:      K;       ]K;      �;       �T��;      �;       ]�;      �;       �T�                       �:      �;       _�;      �;       �U#��;      �;       _�;      �;       �U#�                   ;      ;       0�*;      �;       P�;      �;       P                     ;      �;       V�;      �;       V�;      �;       ��                 �:      ;       ���
  �;      �;       ���
                   �:      ;       ^�;      �;       ^                 �:      ;       _�;      �;       _                   �:      ;       0��;      �;       0��;      �;       P                       ;      ;       P;      ;       v;      ;        �;      �;       P                  K;      �;       ]                    K;      t;       U|;      �;       ���;      �;       U                 K;      �;       T                       K;      T;       ��T;      �;       R�;      �;       r 1&��;      �;       R�;      �;       ���;      �;       R                          [;      f;       r  q �f;      i;       q x �i;      k;       r  q �k;      r;       r  t ���r;      �;       Q                          �      
       U
      �       ^�      �       �U��      N       ^N      Q       U                      �      
       T
      N       ��N      Q       T                                �      �       Z�      �       ]�      �       Z�      �       Z�      �       }��      �       ]�      �       Z�      N       }�N      Q       Z                              .       ].      �       U�              U�      �       U                     .      �       ^�      �       �U��      N       ^                  .      u       U�      �       U                  .      u       Z�      �       Z                  .      u       { | "#��      �       { | "#�                  .      u       Q�      �       Q                     .      T       { | "# T      q       T�      �       { | "#                    =      u       P�      �       P                  =      u       { | "#�      �       { | "#                  =      u       q �      �       q                       =      d       Rd      l       r�l      u       R�      �       R                   �      �       ^�      N       ^                  �      �       ���      N       ��                     �      �       Z�      P       _�      N       _                   �      �       U�      �       P                    �      �       0��      �       0��             P                 �      �       p ����H{ "�                      �              X�      �       X�      N       ��                 �      �       p ����H{ "                      �              Y�      �       Y�      N       ��                    P      i       Ui      �       _                                      y 3%�             Y      #       p  y "�#      *       y p �*      3       p  y "�      N       Z                                   T      #       t p "#�#      *       t p "�*      3       t p "#�                          #       q p "#�#      *       q p "�*      3       q p "#�                       @       Z                  3      @       q p "�                      u      z       �Y��z      ~      
 �Y�R��~      �       ��������                        �             U      5       S5      ;       �U�;      |       S                          �             T      ;       �T�;      Q       TQ      d       Ud      |       �T�                        �             Q      :       ]:      ;       �Q�;      |       ]                                   R      6       V;      |       V                     �      ,       0�,      ;       P;      |       0�                     �             0�      ;       Q;      |       0�                 G      |       S                  G      d       Ud      z       �T�                G      z       V                 G      d       Q                G      ]       V]      z       \                      P      w       Uw      �       ]�      �       �U�                      P      w       Tw      �       V�      �       �T�                    c      n       Pn      w       u                      g      �       S�      �       sh��      �       S                 w      �       V                   w      �       S�      �       sh�                          �      �       U�      �       V�      �       �U��      �       U�             V                        �      �       T�      �       S�      �       �T��             S                          �      �       Q�      �       �Q��      �       Q�      �       R�             �Q�                    �      �       0��      �       0��             P                  �      �       P                    �             U      �       Q                  �      �       X                        �       T                       ,       X                       ,       T                 ,      M       q��                 M      �       q��                 �      �       q��                      �9      �9       U�9      �:       S�:      �:       �U�                 :      �:       V                 :      N:       V                 (:      N:       V                 N:      {:       V                 N:      {:       s� �                 _:      {:       V                 _:      {:       s� �                    p      �       U�      7       [                      p      �       T�      �       u��      7       �T�                          p      �       Q�      �       S�      �       �Q��      �       S�      7       �Q�                    p      �       R�      7       �R�                          p      �       X�      �       V�      �       �X��      �       V�      7       �X�                   u      �       u��      �       {��      7       {��                      �      �       V�      �       V�      7       �X�                      �      �       S�      �       S�      7       �Q�                        �      �       U�      �       {���      �       U�      7       {��                   �      �       Q�      �       u                            z      �       0�g      �       R�      �       R�      �       0��      �       P�             0�                       �      �       0��      �       {���      �       0��      7       {��                             n       Qn      q       q�q      �       Q�      �       {��      7       {�                  #      4       SP      ]       S                  #      4       QP      ]       Q                       -      4       P4      4      
 p r "#���V      Y       PY      ]       R                      -      4       p ?&�4      4       RV      Y       p ?&�Y      ]       r ?&�]      ]       R                        �      �       P�      [       pP�[      �       P�      �       P                �      �       S                  �      �       p�      �       pX                   �      �       Q�      �      
 q | "#���                  �      �       q ?&��      �       \                �      �       S                   �      �       Q�      �      
 q | "#���                  �      �       q ?&��      �       \                      %       S                        %       \%      %      
 | } "#���                        %       | ?&�%      %       ]                %      ,       S                  %      ,       Q,      ,      
 q ~ "#���                  %      ,       q ?&�,      ,       ^                            �       R�             R      ,       rP�,      7       R                   @      �       u��      �       ^                               P�             P                 @      �       u                   �             {���             {��                          �       U�      7       U                          P      P       PP      Z       p �Z      �       y u� $ &��      �       P�      �       p ��      �       y ~ � $ &��      �       y u� $ &�                P      j       �Q��      �       �Q�                    P      Z       p �Z      j      	 y u���      �       p ��      �      	 y ~ ��                      c      j       Pj      j      
 p ~ "#����      �       P�      �      
 p  "#���                    c      j       p ?&�j      j       ^�      �       p ?&��      �       _                              5       U5             ]      ,       | ,      �       �U�                            $       T$      �       V�      �       �T�                            1       Q1      �       S�      �       �Q�                             9       0�9      =       P=      �       \�      �       �Q                  n      }       U�      �       U                        n      �       P�      �       p~��      �       P�      �       P�      �       p~��             P                 P      �       |��                   P      `       |��`      �       Q�      �       qh��      �       Q                 �      �       |�                   �      �       |��      �       Q�      �       qh��             Q                  +      4       P                    S      �       1��      �       T�      �       T�      �       T      *       T                    X      o       1�o      �       T                   X      �       ���      �       Z                 X      �       X                   X      o       0�o      �       Q                     o      r       r �q ����1$��"��r      �       r �u 1$��"���      �       r|�u 1$��"��                 �      �       T                 �      �       _                 �      �       X                   �      �       0��      �       Q                     �      �       r �q ����1$ "���      �       r �u 1$ "���      �       r|�u 1$ "��                 �      �       T                 �      �       ^                 �      �       X                   �      �       0��      �       Q                     �      �       r �q ����1$~ "���      �       r �u 1$~ "���      �       r|�u 1$~ "��                 �             T                 �             ]                 �             X                   �      �       0��             Q                     �             r �q ����1$} "��             r �u 1$} "��             r|�u 1$} "��                        0      k       Uk      �       �U��      �       U�             �U�                                      0      v       Tv      �       �T��      �       X�      �       X�      �       x��             Y      2       Y2      7       y�7      B       ZB      ]       T]      c       Zc      v       z��      �       T�             z�                        0      v       Qv      �       �Q��      �       Q�             �Q�                          0      f       Rf      �       ]�      �       �R��      �       R�             ]                          0      i       Xi      �       ^�      �       �X��      �       X�             ^                        0      v       Yv      �       S�      �       �Y��             S                      0      �       � �      �       P�             �                     T      [       u���      �       U                  �      �       u��                  �      B       Z                    �      �       T�             T                        �      �       pP��      �       P�      �       pP��      �       p0�                    �      �       [�      �       [                        �             pP�      "       P"      2       pP�2      7       p0�                  �             [                       7      =       1�=      B       {�B      R       {~�X      ]       {��      �       {~�                    c      �       Q�             Q                              �       Y�      �       Y�      �       r<�      �       r                           �       X�      �       y q ��      �       X                         =      B       RX      �       R�      �       rP��      �       R�      �       rP��      �       R�             R                    �              U      b       �U�                    �       �        T�       b       �T�                     �       �        t ����
�u "#��              �T����
�u "#�      b       �T����
��U"#�                     �       �        t ����
�u "#��              �T����
�u "#�      b       �T����
��U"#�                  �       �        P�       �        p�                       �       �        �T����
�u "#��       L       QL      \       qh�\      a       Q                   �              �T����
�u "#�      b       �T����
��U"#�                 �       �        �T����
�u "#�                                   qp3      T       PT      a       qp                                  T3      <       p r �<      a       T                      %       q                          %       P%      %      
 p t "#���                        %       p ?&�%      %       T                �       �        x                    �       �        Q�       �       
 q r "#���                  �       �        q ?&��       �        R                                �      �       U�             S             �U�      �        S�       �        U�       �        S�       �        �U��       �"       S                                �      �       T�             \             �T�      �        \�       �        T�       �        \�       �        �T��       �"       \                                            �      v       Qv             ��      �        Q�       �        ���       �        Q�       4!       ��4!      ]!       Q]!      p!       ��p!      !       Q!      �!       ���!      �!       Q�!      �!       ���!      %"       Q%"      �"       ��                                �      �       R�             ]             �R�      �        ]�       �        R�       �        ]�       �        �R��       �"       ]                                                     �      �       q  $ &
�t "#��      v       q  $ &
�| "#�v             ��� $ &
�| "#�             ��� $ &
��T"#�      �        q  $ &
�| "#��       �        ��� $ &
�| "#��       �        q  $ &
�t "#��       �        q  $ &
�| "#��       �        ��� $ &
�| "#��       �        ��� $ &
��T"#��       4!       ��� $ &
�| "#�4!      ]!       q  $ &
�| "#�]!      p!       ��� $ &
�| "#�p!      !       q  $ &
�| "#�!      �!       ��� $ &
�| "#��!      �!       q  $ &
�| "#��!      �!       ��� $ &
�| "#��!      %"       q  $ &
�| "#�%"      �"       ��� $ &
�| "#�                   �      �       q  $ &
�t "#��       �        q  $ &
�t "#�                   �      �       q  $ &
�t "#��       �        q  $ &
�t "#�                                                               R      �       ���      �       R�      �       s�      �       R      �        ���       �        ���       '!       R'!      /!       s/!      4!       R4!      �!       ���!      �!       R�!      G"       ��G"      L"       QL"      �"       ���"      �"       ���"      �"       ��                                             )             VA      �       V�      �       Q�      �       s�      �       T�      �       s      �        V�       �        V�       �        r t "#��@& $ &��       '!       @�4!      �!       V�!      �!       @��!      �!       @��!      6"       VG"      L"       @�L"      �"       V                              M      Y       1�=      I       1�I      �        ���       �        0�4!      I!       0�p!      �!       ���!      %"       ��                        M             V=      �        V�       �        V4!      �!       V�!      6"       VL"      �"       V                                              Q      Q       0���Q      b       0���0��0��b      �       0��������            	 �����A      A       0���A      �       0���0��0���      }        Y�����0��}       �        Y�����T��       �        0����       �        0���0��0���       4!      	 �����<!      <!       0���<!      I!       0���0��0��I!      p!       0�������p!      �!       Y�����T��!      �!      	 ������!      �!       0���0��0���!      �!       1���0��0���!      �!       1���U�0���!      "       Y�����0��"       "       Y�����0�� "      %"       Y�����T�%"      �"       0�������                     f      �       _I!      p!       _%"      �"       _                 v      �       �1& �" $ &�                       v      �      
 1&"��      �       Q�      �       R�      �      
 1&"�                 v             ���1&x " $ &�                 �      �       t ~ "#��@& $ &�                 v             ���1&�1&x " ��                   �      �       ^�      �      
 t ~ "#���                  �      �       ~ ?&��      �       T                   b"      �"       ~ 	���"      �"      
 ��# 	��                    w"      �"       R�"      �"       ��v "# 	��                   w"      z"       q ~ �z"      �"       U                     w"      �"       r t ��"      �"       ^�"      �"       T                   �      A       0��"      �"       0�                               �      �       V�             Q              V       -       v 	��-      A       R�"      �"       V�"      �"       v`��"      �"       V�"      �"       R�"      �"       V                   �      A       ��� $ &
�| "#��"      �"       ��� $ &
�| "#�                          �      �       v q ��              R       A       Q�"      �"       R�"      �"       Q                 A      �       V                 A      �       ��                      ^      k       r ���k             T      �       r ���                    n      �       Q�      �       ��v "# 	�v ���                     �      �       | t "#��      �       u 
�| "#���      �       ��
�| "#��                   �      �       R�      �       X                   �      �       R�      �      
 r u "#���                  �      �       r ?&��      �       U                              ��
�| "#��                                R             ��                                R            
 r t "#���                               r ?&�             T                      a      �        �
  p!      �!       �
  �!      %"       �
                        a      �        Xp!      �!       X�!      %"       X                          a      �       R�      �       	 x ���"�p!      �!      	 x ���"��!      �!       R�!      %"      	 x ���"�                      a      �        |��p!      �!       |���!      %"       |��                       n      �       |���      �        |��p!      �!       |���!      �!       |���!      %"       |��                       n      �       Y�      �       R�      ;        Z;       S        |�                              �      �      	 u  $ &��      �       r |�� $ &��      �       r t� $ &��      �      	 u  $ &�        G       	 r  $ &�G       S        u�x  $ &�S       ^        u�x  $ &�^       r       	 r  $ &�                         n      
        T
       �        Up!      �!       U�!      �!       T�!      %"       U                        n      }       U}      �        ��p!      �!       ���!      %"       ��                            Q        TQ       �        �T�                             
        t ����0u"�
       &       
 t 0u"�z       �        �T����0u"�                    .       Q        SQ       g        Q�       �        Q                 .       Q        X                   T       g        T�       �        T                  V       g        T�       �        T                      �      �       U�      K       SK      M       �U�                      �      �       T�      L       VL      M       �T�                      �      �       U�      	       �U�	      #	       U                         �      9       0�9      E       T�      �       T�      �       0��      �       ��	      #	       0�                      �      9       0��      �       q ����      �       Y	      #	       0�                     �      �       Q�      �       q��      �       Q	      #	       Q                          9       0�	      #	       0�                   �      7       T	      #	       T                         �      9       0�9      h       Vh      n       v�n      	       V	      	       �U#	      #	       0�                     �      �       U�      	       �U�	      #	       U                     �      �       U�      	       �U�	      #	       U                 �      �       [                       �             P             pP�             P	      #	       P                  Q      r       Z                 [      r       0�                      �      �       1��      �       z��      	       z�"	      #	       1�                 �      �       Z                  �      	       T                  �      	       Q                    �      �       u�      	       �U#"	      #	       u                      0	      �	       Q�	      1
       Q1
      4
       q��4
      �       Q                    0	      �	       R�      �       R                 0	      �       T                 0	      �       U                                   �	      �	       0��	      �	       [�	      �	       0�D
      O
       [O
      �
       q!�8$8&��
      �
       [�
             q!�8$8&�k      �       q!�8$8&��      �       [�      �       q!�8$8&�                             �	      �	       P�	      �	       q0�	      �	       qh�	      �	       q0�	      9
       PD
      �       P�      �       P                      D
      O
       0��
      �
       0��      �       0�                       �	      �	       w D
             w k      �       w �      �       w                        �	      �	       �DD
             �Dk      �       �D�      �       �D                    S
      �
       Vk      �       V                      Z
      ]
       ~ s �]
      �
       ^k      �       ^                    �
      �
       S�
      �
       S                    �
             V�      �       V                      �
      �
       ~ s ��
             _�      �       _                 �	      �	       0�                    �	      	
       V
      9
       V                      �	      	
       ^
      
       ~ s �
      9
       ^                        %       0�                    %      5       V8      k       V                      %      5       _F      L       ~ s �L      k       _                            �      �       U�      
       S
             �U�      �       S�      �       �U��      �       S                            �      �       R�             ^             �R�             ^      �       �R��      �       ^                            �      �       X�             \             �X�             \      �       �X��      �       \                 �      �       ��q  �                            �      �       T�             V      �       V�      �       s �      �       V�      �       P�      �       V�      �       P�      �       ~                        �      �       Q�      �       qP��             Q�      �       Q                       �      �       R�      �       rt��             R�      �       R                      �      |       _�      �       _�      �       _                           j       _j      |       h��      �       h�                        f       S                                      0�      $       V$      (       P1      5       V5      :       0�:      L       ��                                 0�5      :       } ���:      L       Q                         5       ]5      C       }�C      f       ]                                    0�      V       \V      ]       T]      a       |�a      f       \                       f       ^                          x      |       0��      �       \�      �       T�      �       |��      �       \                            �      �       U�      �       S�      �       �U��             S             �U�      !       U                              �      �       T�      �       V�      �       �T��      �       T�             V             �T�      !       T                            �      �       T�      �       V�      �       �T��      �       T�             V             �T�                          �      �       U�      �       S�      �       �U��             S             �U�                      �      �       P�      �       P             P                   �      �       u �      �       s                  �      �       s                    �      �       T�      �       V                 �      �       s�                     �      �       s��             s� �             �U#H�                     �      �       s��             s� �             �U#H�                 �      �       T                   �      �       P�      �       s(                   �      �       p ����Hs0"H��      �       s(�����Hs0"H�                 �             V                 �             s� �                   �             s� �             �U#H�                   �             s� �             �U#H�                  �      �       V                   �      �       P�      �       s�                    �      �       p ����Hs� "H��      �       s� �����Hs� "H�                      0      5       Q5      9       qy�9      �       �Q�                          0      W       RW      `       �R�`      |       R|      �       P�      �       �R�                      R      W       X`      l       Xl      �       Q                         R      W       Q`      i       Qi      o       sy�o      u       �Q#3%�u      �       S�      �       �Q#3%#	��                          �      �       U�             \             �U�      -       \-      0       �U�                    �      �       T�      �       t ����1����-( ��      0       �T����1����-( �                  �      �       Q                      �      �       R�             S      *       S                        �             ]            " �T1�T $0)( ����34$�U"#�      /       ]/      0      " �T1�T $0)( ����34$�U"#�                        0       P                 �             |                         p      {       U{      �       T�      �       �U��      �       T                      x      {       U{      �       T�      �       �U�                  {      �       U                            `      �       U�      �       S�      �       u���      �       �U��      �       S�      �       �U�                          `      �       T�      �       V�      �       �T��      �       V�      �       �T�                  c      w       P                          p      �       T�      �       V�      �       �T��      �       V�      �       �T�                            p      �       U�      �       S�      �       u���      �       �U��      �       S�      �       �U�                    �      �       P�      �       P                      z      �       \�      �       T�      �       \                           z      �       u��      �       s��      �       u���      �       �U#��      �       s��      �       �U#�                 z      �       \                   z      �       T�      �       V                   z      �       u��      �       s�                             z      �       u��      �       s��      �       s� ��      �       u`��      �       �U#H��      �       s��      �       �U#�                             z      �       u��      �       s��      �       s� ��      �       u`��      �       �U#H��      �       s��      �       �U#�                 z      �       T                   z      �       P�      �       u(                   ~      �       p ����Hu0"H��      �       u(�����Hu0"H�                   �      �       \�      �       T                   �      �       V�      �       �T�                     �      �       s� ��      �       u`��      �       �U#H�                     �      �       s� ��      �       u`��      �       �U#H�                     �      �       s� ��      �       u`��      �       �U#H�                  �      �       V                   �      �       P�      �       s�                    �      �       p ����Hs� "H��      �       s� �����Hs� "H�                        �      
       U
      �       ]�      �       �U��      /       ]                      �      �       T�      �       t��      
       �T�                    �      �       Q�      /       Q                    �      �       V�      /       V                          �      �       S�      �       x �      �       S�      �       P�      /       S                   �      
       1�1      �       0��      /       0�                �      �       �H^  �                      "      :       q�0$0&��      �       q �0$0&��      �       q�0$0&�&      /       q �0$0&�                    1      �       U�      /       U                            1      :       S:      F       PF      M       p�M      �       P�      �       Z�      �       V             P                    1      :       T�      �       T&      /       T                  1      �       T�      /       T                       
      :       0��      �       0��      �       1��      �       0�&      /       1�                        &       P                                              �"      �"       U�"      D#       ��|D#      �#       �U��#      *       ��|*      �,       �U��,      �,       ��|�,      $.       �U�$.      O.       ��|O.      q3       �U�q3      �3       ��|�3      �4       �U��4      �4       ��|�4      7       �U�7      a7       ��|a7      �7       �U�                                  �"      #       T#      D#       _D#      �#       �T��#      4'       _4'      �4       �T��4      �4       _�4      7       �T�7      a7       _a7      �7       �T�                    �"      #       Q#      �7       ��|                                              �"      #       R#      D#       ��|D#      �#       �R��#      *       ��|*      �,       �R��,      �,       ��|�,      $.       �R�$.      O.       ��|O.      q3       �R�q3      �3       ��|�3      �4       �R��4      �4       ��|�4      7       �R�7      a7       ��|a7      �7       �R�                         )      -)       P-)      q3       ��{�3      �4       ��{�4      7       ��{a7      �7       ��{                                   *      *       0�*      Y*       ��|Y*      �*       [�*      �,       ��|�,      $.       ��|O.      K3       ��|K3      l3       ��|�#��3      �4       ��|�4      7       ��|a7      �7       ��|                          �"      #       Q#      D#       ��|�#      )       ��|q3      �3       ��|�4      �4       ��|7      a7       ��|                          �"      �"       U�"      D#       ��|�#      )       ��|q3      �3       ��|�4      �4       ��|7      a7       ��|                            �"      #       T#      D#       _�#      4'       _4'      )       �T�q3      �3       �T��4      �4       _7      a7       _                            �"      �"       ��}��"      
#       U
#      D#       ��}��#      )       ��}�q3      �3       ��}��4      �4       ��}�7      a7       ��}�                                +#      D#       S�#      $       S$      *       ��|�,      �,       ��|$.      O.       ��|q3      �3       ��|�4      �4       ��|7      a7       ��|                     $      $       0�$$      2$       T2$      @$       R�$      �$       T                      $      2$       T8$      �$       T�4      �4       T                 $      $       0�                           $      �$       \�$      �$       S�$      #'       ��|�4      �4       \7      7       S7      a7       ��|                   $      �$       P�4      �4       P                          $      '$       Q'$      .$       px<$      j$       Qj$      v$       p�4      �4       Q                     L$      v$       Zv$      �$       Q�$      �$       R�4      �4       Z                         �$      �$       \�$      �$       S�$      #'       ��|7      7       S7      a7       ��|                     �$      �$       \�$      4'       S7      a7       S                          �$      �$       P�$      #'       \7      
7       P
7      7       7      a7       \                       �$      �$       0��$      #'       V7      7       0�7      a7       V                            �$      �$       Q�$      �%       s ��|3&9��8��%      &       Q&      <&       s ��|3&9��8�]&      �&       s ��|3&9��8�7      a7       s ��|3&9��8�                              �$      E%       PE%      �%       s��|3&9��8��%      &       P&      <&       s��|3&9��8�]&      �&       s��|3&9��8��&      �&       P7      a7       s��|3&9��8�                        %      �%       U&      <&       U]&      �&       U7      a7       U                       %      �%       T&      <&       T]&      �&       T7      a7       T                        R%      �%       Q&      <&       Q]&      �&       Q7      a7       Q                        U%      �%       R&      <&       R]&      �&       R7      a7       R                  %      ;%       T�&      �&       T                  %      ;%       U�&      �&       U                       #%      ;%       X;%      ;%       u ?&u 'u ?&��&      �&       X�&      �&       u ?&u 'u ?&�                  #%      ;%       R�&      �&       R                   %      ;%       4��&      �&       4�                    U%      �%       R&      &       R]&      v&       R7      7       R@7      @7       R                    U%      �%       Q&      &       Q]&      v&       Q7      7       Q@7      @7       Q                       l%      �%       Y&      &       q ?&q 'q ?&�]&      d&       Yd&      v&       q ?&q 'q ?&�7      7       Y@7      @7       q ?&q 'q ?&�                     u%      �%       P&      &       P]&      v&       P7      7       P@7      @7       P                   U%      �%       4�]&      v&       4�                      �&      �4       0��4      7       0�7      7       0�a7      �7       0�                          �&      5+       ��}�5+      9+       R9+      �4       ��}��4      7       ��}�7      7       ��}�a7      �7       ��}�                      �&      �&       Q�&      '       qp�'      #'       Q7      7                              �&      '       P'      '       p��'      #'       P7      7       ��}                  �&      �&       R7      7       0�                          #'      4'       0�4'      ='       ��|A'      N'       PN'      �(       ��|q3      �3       ��|                    g'      �'       Y�'      �'       S                             g'      �'       Y�'      �'       V�'      (       V(      �(       ��|�(      �(       S�(      �(       ��|q3      }3       ��|}3      �3       ^                                g'      j'       Yj'      �'       S�'      (       ��|(      &(       S&(      >(       ^A(      �(       ^�(      �(       S�(      �(       V�(      �(       Sq3      �3       S                      �'      �'       \�'      �'       V�'      �'       \                           (      &(       S&(      A(       VA(      E(       ^E(      �(       V�(      �(       Sq3      �3       V                           �'      �'       V�'      (       ��{(      &(       T&(      �(       ]�(      �(       ]�(      �(       T                      �'      (       ^(      �(       ��|�(      �(       \q3      �3       ��|                                  �'      �'       ]�'      �'       ]�'      (       \(      &(       T&(      A(       _](      �(       _�(      �(       ]�(      �(       Tq3      �3       ]                              �'      �'       _�'      (       _(      &(       ��|&(      A(       Sj(      �(       S�(      �(       \q3      �3       \                     �'      (       P(      �(       ��|�(      �(       P                      &(      8(       P�(      �(       Pq3      �3       P                       N'      &(       0�&(      �(       \�(      �(       _q3      �3       _                D#      �#       ��}�                 L#      �#       S                      ()      �)       s��,      �,       s�$.      O.       s�                     ()      �)       s���,      �,       s��$.      O.       s��                            S)      �)       ^�)      �)       T�,      �,       ^$.      +.       T+.      J.       ^J.      O.       T                               S)      �)       U�)      �)       ��|�)      �)       P�)      �)       U�)      �)       Q�,      �,       U$.      '.       P'.      O.       U                                   S)      *       ^*      �,       ��|�,      �,       ^�,      $.       ��|$.      +.       T+.      O.       ^O.      q3       ��|�3      �4       ��|�4      7       ��|a7      �7       ��|                             S)      �)       U�)      �,       ��|�,      �,       U�,      q3       ��|�3      �4       ��|�4      7       ��|a7      �7       ��|                      d)      *       V�,      �,       V$.      O.       V                          h)      l)       t 	��l)      �)       T�)      *       \�,      �,       T$.      O.       \                                 S)      ~)       0�~)      �)       1��)      �,       ��|�,      �,       0��,      $.       ��|$.      O.       1�O.      q3       ��|�3      �4       ��|�4      7       ��|a7      �7       ��|                S)      U)       U                S)      U)       ��|#�                
  S)      U)       PU)      U)      
 p q "#���                  S)      U)       p ?&�U)      U)       Q                    �5      _6       Po6      7       Q                         �5      �5       Q�5      6       x�b6      f6       Pf6      �6       [�6      �6       x�                  �5      7       U                  �5      7       T                    �5      6       R6      X6       R                    �6      �6       R�6      7       R                               *      Y*       ��|Y*      �*       [�*      �,       ��|�,      $.       ��|O.      l3       ��|�3      �4       ��|�4      7       ��|a7      �7       ��|                               *      5+       ��}�5+      9+       R9+      �,       ��}��,      $.       ��}�O.      q3       ��}��3      �4       ��}��4      7       ��}�a7      �7       ��}�                            7*      d*       Qd*      p*       qp�p*      �*       Q�*      �*       qp��*      �*       Q�4      �4       Q                             7*      Y*       ZY*      l*       Pl*      p*       p��p*      �*       P�*      �*       p���*      �*       P�4      �4       Z                   7*      Y*       Y�4      �4       Y                                �*      �*       0��*      �*       [�*      �*       [U,      �,       [�,      -       [�4      �4       [�4      �4       [�4      �4       0�                     �*      �*       v U,      �,       v �,      �,       \                      �,      �,       \�,      �,       U�,      �,       Q�,      �,       U                  a,      �,       P                   �,      �,       U�,      �,       Q                        �*      �*       Q�,      -       Q�4      �4       Q�4      �4       Q                       �*      �*       Q�,      �,       Q�,      -       P�4      �4       P                         �*      �*       Q�,      -       Q�4      �4       Q�4      �4       P�4      �4       P                             +      +       U+      U,       ��|-      $.       ��|O.      Q3       ��|�3      �4       ��|�4      7       ��|a7      �7       ��|                      +      5+       ��}�5+      9+       R9+      G+       ��}�                  +      G+       ��|                  +      +       ��~                       +      -+       V-+      9+       U9+      :+       vP�:+      G+       V                   +      +       P+      +       u                      G+      U,       ��|-      f-       ��|,4      |4       ��|                     G+      U,       ��}�-      f-       ��}�,4      |4       ��}�                     G+      U,       ��|-      f-       ��|,4      |4       ��|                        Y+      �+       \�+      U,       V-      &-       \,4      14       V                  \+      �+       _                          \+      �+       0��+      �+       R�+      �+       \�+      ,       Q-      &-       0�,4      14       \                                          j+      �+       ]�+      U,       ��|-      &-       ]&-      $.       ��|�#�O.      �0       ��|�#��0      l3       ��|�#��3      4       ��|�#�4      ,4       ��|�#�,4      14       ��|14      �4       ��|�#��4      7       ��|�#�a7      �7       ��|�#��7      �7       ��|�#�                   j+      q+       p  $ &
���~"#�q+      }+       } $ &
���~"#�                   j+      q+       p  $ &
�s "#�q+      }+       } $ &
�s "#�                            ~+      �+       P�+      �+       P�+      U,       ��|-      &-       P&-      f-       ��|,4      |4       ��|                      �+      �+       \,      U,       \,4      14       \                  ,      K,       ^                  ,      S,       S                 &-      B-       ��}                   &-      B-       ��}B-      f-       P                 14      K4       ��}                 14      K4       ��}                      �-      $.       S�3      �3       S|4      �4       S                          �-      �-       R�-      .       R.      $.       s(�3      �3       R|4      �4       R                              �-      �-       U�-      .       s0r � $ &�.      $.       s0s(� $ &��3      �3       U�3      �3       s0q ��3      �3       s0r � $ &�|4      �4       U                  �-      �-       u q ��-      .       U                   .      .       Q.      .      
 q r "#���                  .      .       q ?&�.      .       R                 �3      �3       U                   �3      �3       U�3      �3      
 q u "#���                  �3      �3       u ?&��3      �3       Q                      O.      E0       ��|�3      4       ��|�4      o5       ��|a7      �7       ��|                      O.      E0       ��}��3      4       ��}��4      o5       ��}�a7      �7       ��}�                      X.      �.       ��|� $ &
�t "#��4      5       ��|� $ &
�t "#�5      5       ��|� $ &
���~"#�                        q.      x.       t p "#�x.      �.       ��|
�t "#��4      5       ��|
�t "#�5      5       ��|
���~"#�                   q.      �.       ��}�4      5       ��}                            q.      �.       0��.      E0       V�3      4       V�4      5       0�5      )5       P)5      o5       Va7      �7       V                             q.      �.       0��.      �.       R�.      �.       0��.      E0       ^�3      4       ^�4      5       R)5      o5       ^a7      �7       ^                   q.      9/       S�4      )5       S                       �.      E0       \�3      4       \�4      o5       \a7      �7       \                                   �.      �.       S�.      �.       P�.      �.       S�.      /       R/      !/       p !/      9/       R9/      E0       S�3      4       S�4      5       P)5      o5       Sa7      �7       S                  �.      &/       P                    �/      0       r ����3$v ")5      .5       r ����3$v "e5      o5       r ����3$v "                 �3      �3       v                                �/      �/       0��/      �/       Q�/      �/       R�/      �/       Q�/      �/       ^�/      	0       P�3      �3       0�)5      .5       Pe5      o5       P                       0      ,0       UX5      e5       Ua7      k7       Uk7      |7       s0                   �3      �3       u p ��3      �3       U                   �3      �3       U�3      �3      
 p u "#���                  �3      �3       u ?&��3      �3       P                  .5      15       u z �15      =5       U                   ;5      =5       P=5      =5      
 p q "#���                  ;5      =5       p ?&�=5      =5       Q                     ^0       1       ��|�1      73       ��|�7      �7       ��|                     ^0       1       ��}��1      73       ��}��7      �7       ��}�                 ^0      �0       ��|� $ &
���~"#�                 ^0      �0       ��|� $ &
���~"#�                      w0      �0       Y�2      �2       Y�2      73       Y                     w0       1       _�1      73       _�7      �7       _                  ~0      �0       P                      �0      �0       Q�2      �2       Q�2      73                                �0      �0       0��0      �0       S�0      �0       R�2      �2       V�2      73       S                              �0      �0       T�0      �0       R�0      �0       R�1      �1       R�1      �2       V�2      73       T�7      �7       V                         �0      �0       Q�0      �0       P2      �2       R�2      �2       P�2      73       Q                     �0      �0       0��0      �0       R�2      �2       R                      �1      �1       X�1      2       ��|�2      �2       T�7      �7       T                            �1      �1       T�1      �1       T�1      2       ^�2      �2       x t ��2      �2       X�7      �7       X�7      �7       ^                    �1      �1       [�1      �1       [�1      2       ��|                          �1      �1       Q�1      �1       U�1      2       ��|�2      �2       Q�7      �7       Q                     2      P2       r0U2      �2       r0�2      �2       r0                            2      (2       Q(2      P2       r0t �\2      d2       Qd2      �2       r0t ��2      �2       Q�2      �2       r0t �                    H2      U2       Q�2      �2       Q                      �1      �1       @<$��1      2       P�2      �2       @<$��7      �7       @<$�                   %2      (2       q ~ �(2      /2       Q                   /2      62       Q62      62      
 q { "#���                  /2      62       q ?&�62      62       [                 �2      �2       Q                  h2      o2       Qo2      o2      
 q { "#���                  h2      o2       q ?&�o2      o2       [                  a2      h2       Qh2      h2       r0�t �                 h2      h2       Q                h2      h2       q ?&�                �2      �2       s0                   �2      �2       P�2      �2      
 p r "#���                  �2      �2       p ?&��2      �2       R                3      3       q0                   3      3       P3      3      
 p r "#���                  3      3       p ?&�3      3       R                    1      /1       ��|/1      �1       [                  1      �1       ��}�                   $1      /1       0�/1      �1       P                  1      �1       Q                   1      �1       Y                  $1      �1       Z                    �7      �7       U�7      �7       �U�                    �7      �7       T�7      �7       �T�                    �7      �7       Q�7      �7       �Q�                    �7      �7       R�7      �7       �R�                          �7      8       U8      �9       S�9      �9       �U��9      �9       U�9      �9       S                            �7      8       T8      }9       �T�}9      �9       T�9      �9       �T��9      �9       T�9      �9       �T�                            �7      8       Q8      }9       �Q�}9      �9       Q�9      �9       �Q��9      �9       Q�9      �9       �Q�                      �7      8       Q8      �8       _}9      �9       Q                          �7      �7       T�7      8       t ����1����-( �8      }9       �T����1����-( �}9      �9       t ����1����-( ��9      �9       �T����1����-( ��9      �9       �T����1����-( �                        �7      8       U8      �9       S�9      �9       �U��9      �9       S                     O8      `8       P�9      �9       P�9      �9       P                             �7      8      ' t ����1����-( ����0u "#�8      8      ( �T����1����-( ����0u "#�8      }9      ( �T����1����-( ����0s "#�}9      �9      ' t ����1����-( ����0s "#��9      �9      ( �T����1����-( ����0s "#��9      �9      ) �T����1����-( ����0�U"#��9      �9      ( �T����1����-( ����0s "#�                   �7      8       u }9      �9       s                      |8      }9       ^�9      �9       ^�9      �9       ^                     |8      }9       \�9      �9       \�9      �9       \                     |8      }9       V�9      �9       V�9      �9       V                     |8      }9      ( �T����1����-( ����0s "#��9      �9      ( �T����1����-( ����0s "#��9      �9      ( �T����1����-( ����0s "#�                                |8      Q9       0�Q9      U9       PU9      h9       0�h9      l9       Pl9      }9       0��9      �9       0��9      �9       P�9      �9       0��9      �9       P                    �8      �8       P�8      �8      	 s ��"#8                   �8      59       ���9      �9       ��                 �8      �8       V                 �8      �8       V                  9      59       ��                  9      9       \                 9      9       \                 9      59       ��                 9      9       ^                 9      9       ^                          �;      �;       U�;      <       �U�<      *<       U*<      \<       S\<      d<       �U�                        �;      �;       T�;      <       �T�<      0<       T0<      d<       �T�                          �;      �;       Q�;      <       �Q�<      &<       Q&<      ]<       V]<      d<       �Q�                          �;      �;       Q�;      <       �Q�<      &<       Q&<      ]<       V]<      d<       �Q�                        �;      �;       T�;      <       �T�<      0<       T0<      d<       �T�                          �;      �;       U�;      <       �U�<      *<       U*<      \<       S\<      d<       �U�                    8<      S<       PT<      d<       P                         �;      �;       u��;      <       �U#�<      *<       u�*<      \<       s�\<      d<       �U#�                 �;      �;       u                     �;      <       \<      _<       \                    �;      <       ]<      a<       ]                          p<      �<       U�<      �<       �U��<      �<       U�<      �<       S�<      �<       �U�                          p<      �<       T�<      �<       �T��<      �<       T�<      �<       V�<      �<       �T�                        p<      �<       Q�<      �<       �Q��<      �<       Q�<      �<       �Q�                          p<      �<       R�<      �<       �R��<      �<       R�<      �<       ]�<      �<       �R�                          w<      �<       R�<      �<       �R��<      �<       R�<      �<       ]�<      �<       �R�                        w<      �<       Q�<      �<       �Q��<      �<       Q�<      �<       �Q�                          w<      �<       T�<      �<       �T��<      �<       T�<      �<       V�<      �<       �T�                          w<      �<       U�<      �<       �U��<      �<       U�<      �<       S�<      �<       �U�                    �<      �<       P�<      �<       P                         w<      �<       u��<      �<       �U#��<      �<       u��<      �<       s��<      �<       �U#�                 w<      y<       u                     �<      �<       P�<      �<       P                    �<      �<       \�<      �<       \                                �'      
(       U
(      B(       �U�B(      i(       Ui(      H)       VH)      a)       �U�a)      �)       V�)      �)       �U��)      �)       U�)      �)       V                        �'      
(       T
(      8(       S8(      ?(       ~�~�?(      B(       �T�B(      �)       S                          �'      
(       Q
(      B(       �Q�B(      i(       Qi(      �)       �Q��)      �)       Q�)      �)       �Q�                          �'      
(       R
(      B(       �R�B(      i(       Ri(      �)       �R��)      �)       R�)      �)       ��~                     �'      ?(       ^?(      B(       �T#��B(      �)       ^                       �'      
(       t��
(      8(       s��8(      ?(       ~P�?(      B(       �T#��B(      �)       s��                   �'      A(       _B(      �)       _                         �'      (       0�(      0(       \B(      �(       0��(      �)       \�)      �)       0�                         �'      (       0�(      0(       ]B(      �(       0��(      �)       ]�)      �)       0�                    �'      �'       U�'      �'       �U�                      �'      �'       T�'      �'       u�~��'      �'       �T�                    �'      �'       Q�'      �'       �Q�                      �      �       U�      �       P�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                      p      }       U}      �       P�      �       �U�                         $      ;$       U;$      3%       �U�3%      >%       U>%      R'       �U�                         $      �$       T�$      3%       �T�3%      >%       T>%      R'       �T�                      $$      �%       Q�%      �&       �T#'      R'       �T#                           $$      �$       t �$      (%       X(%      3%       �T3%      >%       t >%      �&       X'      R'       X                   �$      (%       R>%      X%       R                    �$      (%       P>%      q%       P                     �%      
'       W
'      '       w��~�'      R'       W                    �&      �&       P'      '       P                   �%      �%       p 
 �+'      R'       p 
 �                   �%      �%       W+'      R'       W                      �      �       U�      �       T�      �       �U�                   �      �       u �      �       U                      `'      �'       U�'      �'       V�'      �'       �U�                      `'      x'       Tx'      �'       S�'      �'       �T�                   `'      �'       0��'      �'       P                                            �      �       U�      �       ^�      �       �U��      �       ^�      �       �U��      �       ^�      �       U�             ^      #       U#      �       ^�      �       U�      �#       ^�#      �#       �U��#      $       ^                    �      �       T�      $       ��~                      F      H       QH      �       U�#      $       U                        O      n       Qn      �       r��      �       q��#      $       Q                         S      
       ��~�8$8&��      �       ��~�8$8&��      �       ��~�8$8&�i      �       ��~�8$8&�z#      �#       ��~�8$8&��#      �#       ��~�8$8&�                                   S      
       ^�      �       ^�      �       ^�      �       U�             ^      #       U#      �       ^�      �       Ui      �       ^z#      �#       ^�#      �#       ^                               f      w       0�w      
       ���      �       ���      �       ���      �       ���#�c      �       ��z#      �#       ���#      �#       ��                       f      w       0�w      �       S"      �       Sc      �       S                   `      �       ~�c      �       ~�                    �      �       T�      �       T                          �      
       ��~�8$8&��      �       ��~�8$8&��      x       ��~�8$8&��      �#       ��~�8$8&�$      $       ��~�8$8&�                      �      =       ��1$~�"=      �       U�      �       U                                          �      
       ^�      �       ^�      �       ^�      �       U�             ^      #       U#      �       ^�      �       U�      x       ^�      �#       ^�#      �#       �U��#      �#       ^$      $       ^                                         T��             T�Q�      !       R�Q�!      j       T�Q�j      m       �Q��      �       T�Q�                                           !      d       V�\�d      g       �\�/      2       T��2      ?       T�Q�?      B       P�Q�B      �       T�Q��      �       S�V��             T�Q��      �       V�\��      �       V���      �       S�V��      �       S�Z��      �       S��z#      �#       T�Q�                                              �      �       V���             V�\�             R�\�             R�V�      !       \�V�!      d       V�\�d      g       �\�~      �       V���      �       V�\��      �      
 ������      
      
 �������      �       V�\��      �       T�Q��      �      
 ������z#      �#      
 �������#      �#      
 ������                      �      �       P�      �       ~��      �       ~�                             !      �       P�      �       _      
       _�      �       P�      �       _z#      �#       _�#      �#       _                            �      Q       ]Q      
       \�      �       ]�      �       \z#      �#       ]�#      �#       ]                                          +      �       S�             V             S      A       VA      �       s��             S      S       VS      �       ]�      
       V�      �       S�      �       ]z#      �#       V�#      �#       s��#      �#       s�                                     C      U      	 r 8$8&��      �       q 38$8&��      �       v �38$8&�      �       v �38$8&�      S       v �38$8&�S      e      	 p 8$8&��            	 p 8$8&�z#      �#       v �38$8&��#      �#       s�38$8&��#      �#       v �38$8&��#      �#       s�38$8&�                      �      �       T�      �       P�      �       T                  �      �       Q                        f      �       T�      �       Y�      �       T�#      �#       T                    i      �       Q�#      �#       Q                          r      �       Z�      �       Y�      �       X�      �       Z�#      �#       Z                        u      �       X�      �       Z�      �       X�#      �#       X                      �      �       Y�      �       R�      �       Y                  �      �       P                          S      �       S�      �       S�      �       R�      
       S�      �       S                        S      �       V�      �       V�             Z�      �       V                                 �             ^      #       U#      c       ^�      �       U�      �       ^�      z#       ^�#      �#       ^�#      �#       �U�$      $       ^                                �             \      !       |�!      c       \�      x       \�      7       \�"      �"       \�#      �#       \$      $       \                            �      c       S�      x       S�      7       S�"      �"       S�#      �#       S$      $       S                     �      �       s(�      �       TN      c       T                             �      #       ]N      c       Q�      i       ]�      7       ]�"      �"       ]�#      �#       ]$      $       ]                        �      �       U�      i       ^�      z#       ^�#      �#       ^$      $       ^                                   	      7       ��7      C        VC       !       _!      !       v��!      ""       V""      0"       v�0"      D"       �D"      �"       _�"      �"       V�"      #       V#      Z#       V                              �!       \""      �"       \Z#      z#       \                         	      7       0�7      *        ��*       I        PI       �"       ��#      z#       ��                                                        �      Z       QZ      i       U�      �       U�             PM      ]       P]      l       Tl      �       P�      �       T�      �       P"!      )!       Q)!      8!       U8!      x!       Qx!      �!       p �!      �!       Q�!      �!       U�!      �!       Q�!      ""       P�"      �"       P�"      �"       Q#      Z#       PZ#      z#       Q�#      �#       U$      $       P                                                 i       U�      �       U]      l       Tt      �       T)!      8!       UA!      �!       U�!      �!       U�!      �!       U�!      ""       T�"      �"       T�"      �"       U#      Z#       TZ#      z#       U�#      �#       U                    R       !       S""      �"       S                    W       !       ]""      �"       ]                    	      <       R�"      �"       R                            i       T�      �       T�"      �"       T�#      �#       T                         M       h        0�h       �        V�       �        PD"      ["       P�"      �"       V                        s       �        Q�       �        T�       �        Q�"      �"       Q                    w       �        R�"      �"       R                      �       �        x  $ &q ��       �        ~� $ &q ��"      �"       x  $ &q �                       �       �        r t "1x  $ &��       �        r x "1x  $ &��       �        ~� $ &r "1~� $ &��"      �"       r x "1x  $ &�                	 �      �       ���                 �      �       ���                 �      �       ���                   (      Z       Q�"      �"       Q                     (      Z       ����"      �"       ����"      �"       R                           (      <       ���<      F       RF      J       ���J      Z       R�"      �"       ����"      �"       R                       (      <       ��<      S       P�"      �"       ���"      �"       r                    (      Z       0��"      �"       0�                   �!      �!       QZ#      j#       Q                     �!      �!       ���Z#      e#       ���e#      j#       P                         �!      �!       ����!      �!       p��!      �!       ����!      �!       p�Z#      e#       ���e#      j#       P                            �!      �!       P�!      �!       T�!      �!       P�!      �!       TZ#      e#       Pe#      j#       p                      v      �       P�"      �"       PI#      Z#       P                       v      �       ����"      �"       ���I#      U#       ���U#      Z#       Q                           v      �       ����      �       q��      �       ����      �       q��"      �"       q�I#      U#       ���U#      Z#       Q                              {      �       Q�      �       R�      �       Q�      �       R�"      �"       RI#      U#       QU#      Z#       q                    �      �       P#      1#       P                     �      �       ���#      %#       ���%#      1#       U                           �      �       ����      �       U�      �       ����      �       U#      %#       ���%#      1#       U                    �      �       Q#      1#       Q                   �      �       R#      1#       R                   �!      ""       P1#      I#       P                     �!      ""       ���1#      =#       ���=#      I#       U                           �!      �!       ����!      	"       U	"      "       ���"      ""       U1#      =#       ���=#      I#       U                    �!      ""       Q1#      I#       Q                   �!      ""       p 1#      I#       p                    C!      {!       Qj#      z#       Q                     C!      �!       ���j#      u#       ���u#      z#       P                         C!      W!       ���W!      c!       p�c!      c!       ���c!      u!       p�j#      u#       ���u#      z#       P                            H!      W!       PW!      c!       Tc!      g!       Pg!      u!       Tj#      u#       Pu#      z#       p                  �"      �"       s�7
���                             p       Tp      �       �T��      4       T                                     H       QH      �       �Q��             Q      �       �Q��      �       Q�      �       �Q��      4       Q                                     H       RH      �       �R��      '       R'      �       �R��      �       R�      �       �R��      4       R                                       H       XH      �       �X��      �       X�      �       �X��      �       X�      �       �X��      #       X#      4       �X�                                       H       YH      �       �Y��      �       Y�      �       �Y��      �       Y�      �       �Y��             Y      4       �Y�                               >      H       ZP      �       P�      �       Z�      B       ZB      �       [�      �       Z�      �       [�      4       Z                                A      H       [H      �       u� $ &�R��      ?       [?      B       QB      �       u� $ &�R��      �       [�      �       u� $ &�R��      4       [                           A      M       Z�             Z      I       X�      �       Z�      �       X�      4       Z                       c      p       t 3&0$0&u� "�p      �       �T3&0$0&u� "��      �       PP      f       t 3&0$0&u� "�f      �       Q                    �      �       XP      T       �q 70$0&&�T      �       �t 70$0&&�                             �      �       x�7
����      �       �X#�7
����      �      	 | 7
����      �       �X#�7
����            	 | 7
���      #       x�7
���#      4       �X#�7
���                    �      �       T�             �T�                    �      �       Q�             �Q�                        �      �       R�      �       �R��      �       R�             �R�                    �      �       X�             �X�                    �      �       Y�             �Y�                      �      �       Q�      �       Q�            % u� $ &�Q"1u� $ &u ��&�                         �      �       p r ��      �       P�      �       P�      �       x  $ &�R��             u� $ &�R�                  �             R                   �      �       t 3&0$0&u� "��             �T3&0$0&u� "�                                P                                �      �       T�             �T�      Y       TY      �       �T��      �       T�             �T�      V       TV      g       �T�                              �      �       Q�             �Q�      g       Qg      �       �Q��      �       Q�             �Q�      g       Q                              �      �       R�             �R�      �       R�      �       �R��      �       R�             �R�      g       R                                �      �       X�             �X�      Y       XY      �       �X��      �       X�             �X�      R       XR      g       �X�                                   �      �       Z�      �       R�      �       P�      
       Z      �       Z�      �       [�      �       Q�             Z             [      g       Z                                �      �       [�      
       u� $ &�R�      �       [�      �       Q�      �       u� $ &�R��              [              u� $ &�R�      g       [                           �      �       Z      ~       Z~      �       T�      �       Z�             T      g       Z                         �      �       r 3&��      �       p 3&��      
       z 3&��      �       { 3&��      �       q 3&��      �       Q                   �      
       z 7��      �       { 7��      �       q 7�                                   Y       x�7
���Y      �       �X#�7
����      �      	 v 7
����             �X#�7
���      I      	 v 7
���I      R       x�7
���R      g       �X#�7
���                      �      T       UT      y       �U�y      �       U                  �      �       T�      �       �T�                    �      �       Q�      �       �Q�                    �      �       R�      �       Z                    �      �       X�      �       �X�                    �      �       Y�      �       �Y�                            �      �       P�             R             Y      D      Q u� $ &�Q"1u� $ &u ��&0u� $ &�Q"1u� $ &u ��&0*( �y      �       P�      �      Q u� $ &�Q"1u� $ &u ��&0u� $ &�Q"1u� $ &u ��&0*( �                        �      �       P�             Q             P�      �       Q                     7      W       RW      o       P�      �       R                       �      �       x�7
����      �      	 x 7
����      D       �X#�7
���y      �       �X#�7
���                          y       Y�      �       Y                        ,       P                           A       X�      �       X                    7      y       T�      �       T                    0      :       Q:      r       �Q�                      :      <       Q<      g       Rg      r       u�� $ &�                      �
      �
       U�
      �
       R�
      !       U                      �
      �
       U�
      �
       R             R      !       R                    �
      �
       Q�
      �
       P�
      !       Q                    �
             P      !       P                              `      �       U�      �	       S�	      �	       v�}��	      �	       �U��	      o
       So
      p
       v�}�p
      u
       �U�                    `      �       T�      u
       �T�                    `      �       Q�      u
       �Q�                    `      �       R�      u
       �R�                    `      �       X�      u
       �X�                    `      �       Y�      u
       �Y�                       �      N	       s� #8�	      �	       s� #8�	      
       s� #8

      ;
       s� #8                       �      N	       s� #(�	      �	       s� #(�	      
       s� #(

      ;
       s� #(                       �      N	       s� #�	      �	       s� #�	      
       s� #

      ;
       s� #                       �      N	       s� #�	      �	       s� #�	      
       s� #

      ;
       s� #                       �      N	       s� �	      �	       s� �	      
       s� 

      ;
       s�                       �      	       R�	      �	       R�	      

       R                      �      	       T�	      �	       T�	      
       T                      �      !	       Q�	      �	       Q�	      %
       Q                      �      N	       X�	      �	       X�	      ;
       X                    	      <	       1�

      ;
       2�                    <	      m	       Ym	      w	       Q                              p      �       U�      �       S�      �       |�}��      �       �U��      O       SO      R       |�}�R      U       �U�                    p      �       T�      U       �T�                    p      �       Q�      U       �Q�                    p      �       R�      U       �R�                    p      �       X�      U       �X�                       �      �       s� #(      T       s� #(�      �       s� #(�             s� #(                       �      �       s� #      T       s� #�      �       s� #�             s� #                       �      �       s� #      T       s� #�      �       s� #�             s� #                       �      �       s�       T       s� �      �       s� �             s�                      �      �       s� #(              s� #�             s� #(                     �      �       s� #              s� #(�             s� #                           B       2��             1�                    B      s       Ys      }       Q                            �      �       U�      ,       S,      2       �U�2      r       Sr      x       �U�x      �       S                                        �      �       T�      /       \/      2       �U#h2      >       T>      u       \u      x       �T�x      �       T�      �       \�             T      ?       \?      ^       T^      �       \                                      �      �       Q�      -       V-      2       �U#p2      s       Vs      x       �Q�x      �       Q�      �       V�             Q      ?       V?      G       QG      �       V                     �      �       u��      �       Y�      �       y �                   �      �       u� �      �       p �                �             V                �             \                 �      �       u�                    �      �       u� �      �       T                  �      �       U�             S                 �             P                 �             ]                             4       U4      ^       V^      a       �U�                           >       T>      a       �T�                           >       Q>      a       �Q�                               &       R&      )       P)      >       p �>      a       �R�                             :       X:      >       r �>      a       �X�                        ]       S                  ?      a       P                  1      `       \                            �      %       U%      8       S8      B       �U�B      �       S�      �       �U��              S                    �             T              �T�                            �             Q      A       _A      B       �Q�B      �       _�      �       �Q��              _                            �      -       R-      E       PE      B       �R�B      S       PS      Y       VY              �R�                        �      E       XE      B       �X�B      K       XK              �X�                                N       Q�      �       ZB      y       Q�      �       Z�              Q                                     5       ^5      N       |�      �       P�      �       u�      �       PB      v       |�      �       u�      �       |                        E      N       PN             VV      �       P�      �       V�              P                      5             ^B      �       ^�              ^                       <      Z       PB      S       PS      V       VV      �       P�              P                                �      �       \�      �       U�      �       ���             U      &       \B      �       \�      �       U�      �       U�              \                                   �       T�      �       ���      �       T�             t�      v       Tv      v       Rv      �       r��      �       T�      �       t��      �       T�              R                                �      <       U<      �       \�      �       �U��      �       \�      �       U�      >       \>      E       �U�E      �       \                                �      <       T<      �       V�      �       V�      �       T�      �       X�             ��      <       VE      �       V                                  �      <       Q<      F       SF      �       �Q��      �       S�      �       Q�      ;       S;      E       �Q�E      �       S�      �       �Q�                            �      (       R(      <       Z<      �       �R��      �       R�      !       ��!      �       �R�                            �             X      �       ^�      �       �X��      B       ^B      E       �X�E      �       ^                          �      <       Y<      �       �Y��      �       Y�             ]      �       �Y�                                 �             r t �      <       [<      >       �R�T�>      C       1�C      �       P�      �       �R�T��      �       [�      !       ��!      y       �R�T�y      �       	���      �       P                          �      �       _�      �       �X�Q��      D       _D      E       �X�Q�E      �       _                          4      7       P7      �       ]�      �       }��      �       ]�      �       ]      !       ]                        T      T       UT      �       Y�      �       ���      �       U�      �       Y                     <      �       P�      �       P      !       0�                     T      �       R�      �       ���      �       R                          �      "       Y"      N       ��N      \       Y!      Z       YZ      �       ���      �       Y                        0      5       P5      �       Uk      p       Pp      �       U                    >      �       Qy      �       Q                      N      k       Rk      n       r q "�n      �       R�      �       R                   N      �       X�      �       X                              G      [       P[      f       uf      �       Q�      �       u �      �       P�      �       u�      �       Q                  Q      m       Tm      }       u� �      �       T                       6      ;       R;      Q       u�      �       R�      �       u�      �       R                      6      V       QV      }       u �      �       Q�      �       u(                            �      �       P�      �       Q�      �       u0�      �       P�      	       Q	             u8                          �      �       R�      �       u�      �       P�      �       u             P             u                         �      �       T      =       T=      F       p F      V       QV      a       T                  �      u       Y                                  �      �       p��      �       z��      �       r��      �       R�      �       P�      �       R�      �       p��      �       P      ,       RV      a       R                    =      F       p O      V       Q                             '       T'      �       �T��      �       T                                    	 p q8�             r 8�      Y      	 p q8��      �       r 8�                 >      h       Q                     *      '*       U'*      S*       �U�                     *      **       T**      K*       SK*      S*       �T�                     *      .*       Q.*      S*       �Q�                     *      .*       R.*      K*       VK*      S*       �R�                 7*      K*       �U�                 7*      K*       �Q�                 7*      K*       V                 7*      K*       S                 K*      K*       0�                           
       U
             �U�                           
       T
             �T�                           
       Q
             �Q�                           
       R
             �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                    �      �       R�      �       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       Q�      �       Q�      �       �Q0�Q $@L$.( �                    �      �       R�      �       �R�                                    �      �       U�      &       Z&      E       �U�E      d       Zd      �       �U��      �       Z�      �       �U��      �       Z�             ��~      �       �U�                                        �      &       T&      E       �T�E      d       Sd      �       �T��      �       S�      �       �T��      v       Sv      �       �T��      �       S�      ;       ��~;      P       �T�P      �       S                                              �      &       Q&      E       �Q�E      d       Qd      �       �Q��      �       Q�      �       ^�      �       �Q��      �       ^�      �       Q�      <       ^<      �       �Q��      �       ^�             �Q�      6       ^6      �       �Q�                                        �      &       R&      E       �R�E      d       Rd      �       �R��      �       R�      h       _h      �       �R��      �       _�      �       �R��      �       R�             _      �       �R�                                �      &       X&      E       �X�E      d       Xd      �       �X��      �       X�      �       �X��      �       X�      �       �X�                                       �      &       ]&      E       �T#��E      d       ]d      �       �T#���      �       ]�      �       �T#���      v       ]v      �       �T#���      {       ]{      ;       ��~;      P       �T#��P      �       ]                                       �      &       t��&      E       �T#��E      d       s��d      �       �T#���      �       s���      �       �T#���      v       s��v      �       �T#���      �       s���      ;       ��~#��;      P       �T#��P      �       s��                                     P      :       w :      E       ��~E      �       w                                                &       0�&      <       VE      `       0�`      �       V�      C       0�C      �       V�             0�      �       V�             vk�      �       V�      �       vk��      �       vV��      �       V�      ;       ��~P      �       V                                               &       0�&      >       \E      `       0�`      d       Vd      �       \�      C       0�C      Y       RY      �       \�             0�      �       \�      �       |��      �       \�      ;       ��~P      `       |�`      j       |*�j      �       \                                                   &       q  $HM$)��&      E       �Q $HM$)��E      d       q  $HM$)��d      �       �Q $HM$)���      �       q  $HM$)���      �       ~  $HM$)���      �       �Q $HM$)���      �       ~  $HM$)���      �       q  $HM$)���      <       ~  $HM$)��<      �       �Q $HM$)���      �       ~  $HM$)���             �Q $HM$)��      6       ~  $HM$)��6      �       �Q $HM$)��                                                   &       q  $@N$)��&      E       �Q $@N$)��E      d       q  $@N$)��d      �       �Q $@N$)���      �       q  $@N$)���      �       ~  $@N$)���      �       �Q $@N$)���      �       ~  $@N$)���      �       q  $@N$)���      <       ~  $@N$)��<      �       �Q $@N$)���      �       ~  $@N$)���             �Q $@N$)��      6       ~  $@N$)��6      �       �Q $@N$)��                  �             U                         0      v       0��             0��      O       0�O      [       P[      G       ^G      P       0�                        W      �       0��             \             |�      1       \                   �      �       0��      �       P                          @      F       PF      d       s�d      v       ��~�             ��~�      P       ��~                              J      L       PL      P       s�P      d       Rd      v       ��~�      �       ��~�             ��~�      P       ��~                       J      v       ^�             ^�      O       ^O      P       ��~                    6      �       ^P      �       ^                    �      �       U�      �       �U�                      �      �       T�      �       u�~��      �       �T�                    �      �       Q�      �       �Q�                      P       W        UW       [        P[       b        �U�                    P       a        Ta       b        �T�                    P       a        Qa       b        �Q�                              -        U-       1        P1       A        �U�                      p       v        Uv       z        Tz       {        �U�                   p       v        u v       z        U                      �      �       U�      �       V�      �       �U�                      �      �       T�      �       S�      �       �T�                   �      �       0��      �       P                        P      n       Un      �       �U��      �       U�      �       �U�                                  P             T      �       S�      �       T�             S             �T�             T      (       �T�(      �       T�      �       S                               P      �       t�             U�      �       U�      �       t�      �       U             U(      �       U�      �       t                     P      �       t �      �       t �      �       t                                  �      �       0����      �      
 0��0����      �       0��0��Y���      �       0��0��Y�X��      �       Z�U�Y�X��      �       Z��Y�X��      �       Z���      �       Z�U���      �       Z�U�Y���      �       Z�U�Y�X�                      �      �       U�      5       _5      K       �U�                    �             Q      �       u�                    �      �       u� �      K       ���~                                   R      �       u� �      K       ���~                       �       T                               %       U�%      0       R]      u       Qu      �       |�4�-�-��������@�-%�4� 4%��      5      ! w #�4�-�-��������@�-%�4� 4%�                     y      �       ���~�      �       P�      K       ���~                     �      �       ]�      �       V�      �       v��      5       V                          �      �       S�      �       s 1&��      �       S�             | ~ 1&�       ]       S0      5       S                      �             PH      ]       P0      5       P                 L             _                  P             \                    p      �       S�             S                     p      z       � �      �       T�      �       T                     p      z       0��      �       ^�             ^                     �      �       ~ s���      �       R�      
       R                    `      v       Uv      �       �X                        �       �        U�       �        �U��       )       U)      �       �U�                        �       �        T�       �        �T��              T      �       �T�                            �       �        Q�       �        Z�       �        �Q��              Q             Z      �       �Q�                                �       �        R�       �        Y�       �        P�               Y       L       Pk      s       Pu      {       P}      �       P                        �       �        X�       �        �X��       �       X�      �       �X�                                  )      @       T@      F       t�F      L       UL      R       PR      X       UX      ^       Q^      d       Pd      k       Uk      �       T�      �       U                       )      L       Pk      s       Pu      {       P}      �       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                      �      �       R�      �       P�      �       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       Q�      �       P�      �       �Q�                          !       U!      9       �U�                                   T      1       P1      9       �T�                    @      Q       UQ      �       �U�                        @      `       T`      o       Uo      �       \�      �       �T�                      Y      �       V�      �       |��      �       �T#�                      ]      �       S�      �       |��      �       �T#�                                    `      �       U�      �	       ]�	      D
       SD
      K
       ]K
      b
       Ub
      �
       ]�
      �
       �U��
      j       ]j      ]       S]             ]                    `      �       T�             ��~                    `      �       Q�             ��                            	      	       R	      w	       _�
      �
       ��~q ��
      j       _]      �       _�      �       ��~q ��      �       _                          	      s	       U�
      �
       ��p ��
             U]      i       U�      �       ��p ��      �       U                                          �      �	       S�	      	
       ^
      
       Q
      K
       ^
      �
       S�
      ^       S^      j       ��j      �       ^�      �       
 ��             ^
             Z      6       ^6      S       r�~�X      ]       0�]      �       S�             ��                                               	      �	       [�	      �	       V
      
       
 �
      I
       VI
      K
       _�
      �
       _�
      L       [L      j       0�j      �       V�      �       Q�      �       V
             0�      P       VX      ]       Q]      v       [v      �       ���      �       _�      �       [�      �       { ��             
 �                        
      
       Q�
      �
       ��~��� $ &8$��
      �
       Ru      �       0��             Z       ]       
 �                           
      
       0��
      �
       Q�
      �
       ��x �      j       
 ��      �       Q�             
 �>      ]       Q�             0�                                          �      �       Q�      �	       Y�	      K
       \x
      �
       U�
             Y      �       \�      �       |��      0       \0      X       |�X      ]       \]      r       Yr      v       Tv      �       ���      �       U�      �       Y�      �       _                             �      	       Z	      K
       ��x
      �
       [�
      �
       ���
      �       ���      �       [�             ��                                            �      �	       T�	      �	       ]�	      
       }�
      =
       ]K
      �
       T�
             T      '       V'      L       v�L      c       Vj      �       ]�      
       }�
      ]       ]]      f       Tf      �       \�      �       T�      �       S�      �       s��      �       S                                �      �       Q�      �
       ���
      �
       ��8&��
             ��             V      m       ��m      �       V�             ��                          5	      �	       ^�	      �	       _
      :
       _j      �       _�      �       _�             Q              _       ]       U                    N	      K
       ��j      ]       ��                    o	      K
       ��j      ]       ��                            �             U      &       S&      '       �U�'      @       S@      A       �U�A      _       S                        �      �       T�             TA      T       TT      _       �h                        �             Q      A       �Q�A      T       QT      _       �l                    �      X       UX      Y       �U�                      �      �       Q�      �       p��      C       QM      X       Q                      �      '       P'      =       T=      X       P                      �      ,       R,      =       u� =      X       R                            �       U�      9       ��y9      n       Un      �       �U�                         9      �       ��y��      �       S�             sP�      �       S�             sP�      9       S9      n       ��y�                        �      �       Y�             ~ | �      #       ~ | �#      9       Y                        �      �       P�      �       z v �      -       z v �#      9       P                            �             Y      ?       ]?      �       y ?&y 'y ?&��             ~ | ?&~ | '~ | ?&�      #       ~ | ?&~ | '~ | ?&�#      9       ]                            �             P      <       [<      �       p ?&p 'p ?&��      �       z v ?&z v 'z v ?&�      -       z v ?&z v 'z v ?&�#      9       [                     X      \       U\      �       _�      �       r | �                      ~      �       U�      �       ]�      �       t | �                    �      �       U�      �       q v �                  (      L       U                         �      �       } p u y ��      �       z v } u y ��      �       z v } ~ | u ��      �       t | z v ~ | u ��      �       t | z v q v ~ | �                  X      �       [                         �       S�             sP�                                V      |       P|      �       s�      �       P�      �       s �      �       P�      �       sh�      	       P	             sx                   g      �       U�      �       R�      �       T�             Q             X                    E      g       s�      �       s�      �       sh                    E      �       s �      �       s(�             sx                          �      �       U�      �       V�      �       �U��      �       V�      �       U                              �      �       W�      �       S�      �       ]�      b       Sb      s       ]�      �       S�      �       s ��      �       W�      �       ��{�                     P      S       p t 3${ "�S      W       w t 3${ "��      �       P                 P      d       x q 3$y "�                            �      �       1��      �       \�      s       \s      w       |�w      �       \�      �       \�      �       |��      �       \                      �      �       1��      �       Rb      r       R�      �       1�                 �      b       S                      �      �       Y      D       PD      r       Y                      �             s0      K       sK      N       QN      b       s                           '       U'      S       �U�                           *       T*      K       SK      S       �T�                           .       Q.      S       �Q�                           .       R.      K       VK      S       �R�                 7      K       �U�                 7      K       �Q�                 7      K       V                 7      K       S                 K      K       0�                          �/      0       U0      00       �@00      �0       �U��0      �0       U�0      �0       �U�                          �/      0       T0      00       ��00      �0       �T��0      �0       T�0      �0       �T�                                    �/      00       Q00      o0       So0      q0       �Q�q0      �0       S�0      �0       �Q��0      �0       S�0      �0       �Q��0      �0       S�0      �0       Q�0      �0       S                        �/      00       R00      �0       �R��0      �0       R�0      �0       �R�                        �/      00       X00      �0       �X��0      �0       X�0      �0       �X�                                  10      A0       PD0      P0       PP0      p0       Vq0      }0       P�0      �0       V�0      �0       P�0      �0       V�0      �0       P�0      �0       V                          �,      �,       U�,      8.       S8.      B.       �U�B.      N.       UN.      �/       S                                              �,      �,       T�,      .       V.      B.       �T�B.      N.       TN.      n.       Vn.      r.       Ur.      �.       V�.      �.       �T��.      �.       V�.      �.       U�.      �.       V�.      /       �T�/      /       V/      �/       �T��/      �/       V                  �.      �.       0�	/      /       0�                    �,      =.       ]N.      �/       ]                             �,      2-       0�2-      H-       PH-      3.       \B.      N.       0�N.      �.       \�.      �.       0��.      �/       \�/      �/       0��/      �/       \                       .      .       0�s.      �.       _�.      �.       0��.      /       _/      �/       _                         �.      �.       0��.      �.       P�.      �.       V�.      	/       V	/      /       0�/      �/       V                        �.      �.       P�.      /       ^/      #/       P#/      �/       ^                 /      �/       \                     /      /       |�/      #/       U#/      �/       |�                        �-      .       VN.      n.       Vn.      r.       Ur.      s.       V�.      �.       U�.      �.       V                         �-      .       ^N.      n.       ^n.      r.       Tr.      s.       ^�.      �.       T�.      �.       ^                      �-      .       0�N.      j.       0�j.      r.       Pr.      s.       _�.      �.       P�.      �.       0�                  :-      �-       V�.      �.       V/      /       V                  :-      q-       Sq-      �-       V�.      �.       V/      /       V                    :-      H-       PH-      �-       \�.      �.       \/      /       \                        :-      H-       p�H-      �-       |��-      �-       U�-      �-       |��.      �.       |�/      /       |�                     :-      v-       0�v-      �-       P�-      �-       0��.      �.       P/      /       3�                    �,      �,       U�,      �,       �U�                    �,      �,       T�,      �,       �T�                    �,      �,       Q�,      �,       �Q�                    �,      �,       R�,      �,       �R�                   �,      �,       u�,      �,       U                          p	      �	       U�	      �	       V�	      �	       �U��	      
       V
      
       �U�                  {	      �	       S�	      �	       0�                    	      �	       \�	      
       \                 �	      �	       S                     �	      �	       s��	      �	       U�	      �	       s�                                    P)      �)       U�)      P*       SP*      S*       |�~�S*      U*       }h�U*      V*       �U�V*      �*       S�*      �*       |�~��*      �*       }h��*      �*       �U��*      �*       S                          ])      U*       ]U*      V*       �U#�V*      �*       ]�*      �*       �U#��*      �*       ]                       ])      F*       0�F*      V*       U�V*      �*       0��*      �*       U��*      �*       0�                    �)      �)       P�*      �*       P                        �)      �)       S�)      5*       SV*      �*       S�*      �*       S�*      �*       S                        �)      �)       s��)      5*       s�V*      �*       s��*      �*       s��*      �*       s�                         �)      �)       V�)      5*       VV*      �*       V�*      �*       V�*      �*       V                               �)      �)       P�)      �)       P�)      *       vt �*      *       vv�V*      g*       vv��*      �*       P�*      �*       vt ��*      �*       vv�                        �
      �
       U�
      �
       S�
      �
       �U��
      �       S                  �      �       P                  r      �       t 
���                                 p ��             q ��                    =      A       p ��A      R       q ��                    0
      4
       U4
      5
       �U�                    0
      4
       T4
      5
       �T�                   0
      4
       T4
      5
       �T�                   0
      4
       U4
      5
       �U�                    `
      u
       Uu
      {
       �U�                    `
      l
       Tl
      {
       �T�                    `
      q
       Qq
      {
       �Q�                  `
      q
       Qq
      v
       �Q�                  `
      l
       Tl
      v
       �T�                  `
      u
       Uu
      v
       �U�                    `
      l
       q ����t �����l
      u
       Tu
      v
       �Q�����T�����                  `
      v
       0�v
      v
       P                    0      :       U:      b	       �U�                            0      ^       T^      �       Z�      \       zp�\      �       Z	      %	       Z%	      C	       PR	      b	       T                              0      v       Qv      �       U�      �       ���      	       Q	      	       U	      R	       ��R	      b	       Q                                                        6      �       _�      �       P�      �       ^�      �       ]�      �       \�      �       V�             S             T             ��      0       R0      8       [8      >       Y>      D       XD      J       UJ      P       TP      V       RV      \       Q\      �       _	      a	       _a	      b	       �U
���                                   J      ^       P^      �       ���      �       ��p "��      �       ��p "~ "��      �       ��p "} "~ "��      �       zp��} "��"~ " "��      �       zp��| "~ " "��"} "�\      g       ���      �       ���      �       U	      	       ��%	      R	       RR	      X	       PX	      b	       ��                        p      �       P�      �       p��      �       �D�#�	      	       P                                                                        �      C       UC      
       S
             �U�      )       S)      �       �U��      o       So      y       Uy      �       S�      �       �U��      %       S%      r       �U�r      �       S�      �       �U��      �       S�      �       �U��      �       S�      �       �U��      �       S�              �U�               S       `        �U�`       f        Uf       \"       �U�\"      f"       Uf"      �#       �U��#      �#       S�#      �$       �U��$      �$       S�$      B)       �U�                        �      '       T#      )       	��`       f        T\"      f"       T                                            '      H       	��H      P       Py      �       P�      �       P�      �       P      )       	���      �       	���      �       	���      �       P@      �       	���      �       P�      �       P�      %       	��%      0       P�      �       P�      �       	��-      C       Pi      t       P�      �       	���#      �#       	��                                
       p ��
      @       x ��r      |       x ��|      �       s 1����$      �$       s 1���                                                                                                                     �      �       Q�      �       Z�      �       Q             P      g       0�g      z       Zz      �       0��      �       Z�      	       0�	      )       0�r      w       Qw      z       Z~      �       	���             Z             0�      8       0��      �       Z�      �       0��      �       Z�      X       ��X      [       Z_      �       1��      �       ���             Z.      E       ZE      Q       0�Q      q       0��      �       Z�      -       Z.      b       Pb      �       0��      �       Z�      �       Q�             P�      �       0�'       *        ZC       `        	��f       s        Zs       �        0��       �        Z�       �        Q�       !       Z!      �!       ���"      �"       Z�"      �"       0��"      �"       0�Q#      f#       0��#      $       Z$      $       Z�$      �$       Z�$      �$       	���$      �$       P�$      %       Z%      8%       ��8%      Y%       	���%      �%       Z�%      �%       P�%      &       Z&      2&       ���&      �&       P�&      *'       	��@'      E'       	��w'      �'       	���'      �'       P�'      �'       	���'      �(       ��)      )       	��                                        �      �       S�      �       �U��      �       S�      �       �U��      �       �U��      -       �U��              �U�       `        �U�f       \"       �U�f"      �#       �U��#      �$       �U��$      B)       �U�                    �      �       Z�      �       Z                                                               �      �        7��      �       R�      �       Q�      �       P�      �       |�      S       TS      �       X)      X       ��#      #       0�      *        7�|      �       P�      �       |g      �       R�      �       ��~�       !       |�!      �!       Ps"      �"       X�"      0#       |$      -$       X-$      i$        7��$      �$        7�"%      Y%       	��$&      2&       	��*'      1'       |1'      E'       zE'      R'       |R'      X'       ��~#�'      �'       	���(      )        7�                                                                    �      �       _:      O       _d      q       _z      H       _H      w       0�w      �       _�      �       _�      �       _�             _      �       _�             0��             _�      �       _'       `        _f       �        _�       �        _�       �!       _s"      �"       _�"      �"       P�"      Q#       _$      $       0�$      i$       _�$      �$       _�$      Y%       _�%      �%       _&      2&       _�&      �'       _�'      �(       _�(      )       _                                                                                                            �      �       ]?      O       ]d      q       ]z      �       ]�      �       }x��      �       ]�      �       }��      �       ]�             R             rx�      )       R)      C       ]H      w       0�w      �       ]�             ]      +       R+      .       rx�.      8       R8      k       ]s      �       ]�      �       R�      �       rx��      �       R�      �       r��      I       RI      �       ]�             ]      E       ]E      c       Rc      f       rx�f      q       Rq      �       ]�      �       }��      �       ]�             0��             ]�      �       R'       `        ]f       �        ]�       �        R�       �!       ]s"      �"       ]�"      �"       R�"      �"       rx��"      �"       R�"      �"       ]�"      Q#       ]$      $       0�$      m$       ]m$      �$       }��$      �$       ]�$      �$       }��$      %       R%      Y%       ]�%      �%       ]&      2&       ]�&      �'       ]�'      �(       ]�(      )       ]                                                                                           �      �       V1      �       V�      �       Y�             V             v�      �       V�             V      %       v�%      �       V�             Q      �       V�             V      1       Y1      U       VU      ]       v�]             V�              V'       `        Vf       �        V�       �        Q�       "       Vs"      �"       V�"      �"       v��"      f#       V�#      -$       V-$      L$       YL$      �$       ��~�$      �$       V�$      �$       Y�$      �$       V�$      %       Q%      Y%       V�%      �%       V�%      �%       V�%      2&       V�&      '       V*'      �'       V�'      �(       V�(      )       ��~)      &)       V                                                    �      �       ^5      �       ^�      �       ^�             ^             ^�              ^'       `        ^f       �        ^�       "       ^s"      f#       ^�#      �$       ^�$      Y%       ^�%      �%       ^�%      �%       ^�%      2&       ^�&      �'       ^�'      �(       ^�(      &)       ^                                                                    �      �       [?      �       [�      �       [�      �       [X      �       [      �       [�      �       ��~�      -       [3      �       [�      �       [�             ['       Z        [s       �        [Q#      f#       [�#      �#       [�#      $       P$      $       [-$      L$       [L$      �$       ��~�$      �$       [�$      �$       [�%      �%       [�%      �%       [�%      �%       |� �%      �%       [�%      &       P*'      E'       [�'      �'       |� �'      �'       [�(      )       ��~                               K      O       x�L      P       x��      �       x r ��      �       Xs       �       	 |� �{ ��#      �#       q��$      �$       q { ��%      &       { p �                                                                                       �      �       Z�             	���             Z             0�H      q       Zr      �       P�      �       0��      �       Z�      �       0��             0�      0       Z0      9       0�9      Z       0��      �       Z�      �       0��      �       0�      u       Zv      �       P�      �       0��      �       Z�      -       1�-      b       Zc      �       P�      �       Z�      �       0��      �       0�%      -       Z       '        0�f       s        Z�       �        Z"      &"       0�f"      s"       Pf#      p#       Zp#      �#       P�#      �#       Z�#      �#       	��Y%      �%       P�%      �%       P�%      �%       Z2&      a&       P�&      �&       Z�'      �'       P�(      �(       	���(      �(       P=)      B)       	��                   �             Sf       s        S                   �             \f       s        \                                             H       |�             |!      �       |�             Q�      �       |�      �       Q�             |�%      �%       |g&      p&       |�&      �&       |�&      �&       u�(      �(       u&)      /)       |/)      B)       p                                   H       Qp      �       Q�      �       Q�%      �%       Qg&      �&       Q�&      �&       Q�(      �(       Q&)      B)       Q                                          -      8       P8      C       RC      H       q ���      �       p ���      �       q ����      �       P�      �       R�%      �%       p ���%      �%       |���g&      s&       Ps&      �&       R�&      �&       P�(      �(       P&)      ))       p ��))      B)       q ���                                                     �             _�             _      �       _
             _       -       _       '        _f       s        _�       �        _"      \"       _f"      s"       _f#      �#       _�#      �#       _Y%      �%       _�%      �%       _�%      �%       _2&      �&       _�&      �&       _�'      �'       _�(      �(       _&)      B)       _                                                               �             ]�             ]      %       ](             ]             }x�      H       ]H      R       }x�R      y       ]      �       ]�      �       }x��      �       ]
      �       ]�      �       }x��      �       ]       -       ]       '        ]f       s        ]�       �        ]"      \"       ]f"      s"       ]f#      �#       ]�#      �#       ]Y%      �%       ]�%      �%       ]�%      �%       ]2&      �&       ]�&      �&       ]�'      �'       ]�(      �(       ]&)      B)       ]                                                                   �             V�             V      �       V�             v�      =       V=      L       v�L      �       V�      �       v��      �       V�      �       v��      -       V       '        Vf       s        V�       �        V"      \"       Vf"      s"       Vf#      �#       V�#      �#       VY%      �%       V�%      �%       V�%      �%       V2&      �&       V�&      �&       V�'      �'       V�(      �(       V&)      B)       V                                                   �             ^�             ^      -       ^       '        ^f       s        ^�       �        ^"      \"       ^f"      s"       ^f#      �#       ^�#      �#       ^Y%      �%       ^�%      �%       ^�%      �%       ^2&      �&       ^�&      �&       ^�'      �'       ^�(      �(       ^&)      B)       ^                                                                                 �             [�             [      H       [H      q       R�      �       R�      u       [�      �       U�      '       [-      b       [h      -       [       '        [f       s        [�       �        [�       �        U"      V"       [f"      s"       Uf#      t#       Ut#      }#       x� }#      �#       U�#      �#       [Y%      b%       Ub%      �%       [�%      �%       [�%      �%       x� �%      �%       [2&      ]&       U]&      a&       u� g&      �&       [�&      �&       [�&      �&       R�&      �&       P�'      �'       R�'      �'       U�'      �'       R�(      �(       [�(      �(       U�(      �(       R&)      B)       [                                          �      �       t��      �       t��       �        p�j"      s"       r u �f#      p#       { u ��#      �#       q��#      �#       TY%      b%       r u ��'      �'       q��'      �'       T�'      �'       u r ��(      �(       r u ��(      �(      	 x� �u �                                        �       S�      �       s��      �       S       '        S�       �        Sf"      s"       Sf#      �#       SY%      b%       S�%      �%       S2&      I&       S                                                                             �      �       \�             X             |             \      �       \-      6       \6      9       P9      b       Xb      �       ��~�      -       \       '        \f       s        X�       �        \"       "       \f"      s"       \f#      �#       \�#      �#       \Y%      b%       \b%      �%       ��~�%      �%       \�%      �%       \2&      F&       \g&      �&       \�&      �&       \�&      �&       U�&      �&       \�'      �'       \�(      �(       U�(      �(       \&)      /)       \/)      B)       P                         O       Ss       �        S                       #       |                              K      a       Pa      h      	 r 3$| "�h      s         t 2$��H     "�����3$| "�s"      "       P"      �"      	 r 3$| "��"      �"      (  |�����2$��H     "�����3$| "�$      -$       P                          �"      �"       P�"      0#       |0#      8#       P<#      Q#       PE'      R'       |R'      X'       ��~#                 �"      �"       ��~�"      #        x ����2$��H     "�p ��~�"�                         S      �       Us"      .#       U.#      0#       Q$      -$       UE'      N'       U                   ~      )       S%      "%       S&      $&       S                     ~      �       X�      )       ��%      "%       ��&      $&       ��                           ~      �       Y�      �       ���      )       | �%      %       | �%      "%       ��~# �&      &       | �&      $&       ��~# �                           ~      �       R�      �       ��~�      )       |�%      %       |�%      "%       ��~#�&      &       |�&      $&       ��~#�                        ~      �       P�      '       ��~%      %       ��~&      &       ��~                     �      (       P(      )       ��%       %       P %      "%       	��&      !&       P!&      $&       	��                     �      �       P�      )       ��~%      "%       ��~&      $&       ��~                 �      �       P�&      '       0�                    �      #       S!      �!       S�'      �(       S                      �      #       ��~!      �!       ��~�'      @(       ��~b(      �(       ��~                        �      �       ����      �       Y�      #       ���!      �!       ����'      �(       ���                        �      #       ���!      ^!       ���^!      b!       Yb!      �!       ����'      �(       ���                        �      �       ����      �       P�      #       ���!      �!       ����'      �(       ���                        �      #       ���!      O!       ���O!      b!       Pb!      �!       ����'      �(       ���                    �      #       ��!      �!       ���'      �(       ��                     �      !       ���#�!      �!       ���#��'      �(       ���#�                 !      !       ��~                                    �      �       P�      "       Pc!      �!       P�!      �!       	���!      �!       P�!      �!       ��~�'      1(       P1(      <(       	��N(      O(       PO(      b(       ��~b(      q(       Pq(      x(       	��x(      �(       P                       �      #       ��~)!      O!       PO!      �!       ��~�'      �(       ��~                 T      �       S                  T      Y       ��~                   T      [       R[      �       ��                    T      [       X[      �       ��~                    T      [       Y[      �       ��~                 \      �       P                  E$      �$       9��(      )       9�                	  E$      �$       5��(      )       5�                
  E$      �$      
  �H     ��(      )      
  �H     �                  E$      �$      
  �H     ��(      )      
  �H     �                   E$      �$       S�(      )       S                 E$      �$      
  �H     ��(      �(      
  �H     �                 E$      �$      
  �H     ��(      �(      
  �H     �                 E$      �$       5��(      �(       5�                 E$      �$       9��(      �(       9�                   M$      �$       P�(      �(       P                   E$      �$       S�(      )       S                E$      E$       �V�                  E$      E$       �I�                  E$      E$       �<�                  E$      E$       �/�                          �      �       U�      #       S#      %       �U�%      .       U                   �      �       U�             S                 �             V                        P      �       U�      �       T�      �       �U��      �       U                      �      �       U�      N       SN      P       �U�                      �      �       T�      O       VO      P       �T�                    �      �       Q�      P       �Q�                             V                              s                        �      	       U	      B       SB      L       �U�L      �       S                          �             T      C       VC      L       �T�L      U       TU      �       V                          �      �       Q�      G       ]G      L       PL      U       QU      �       ]                         �             P      ,       ^L      U       Pk      �       Q�      �       0�                      �      $       \$      (       UL      U       \                               �      ,       _,      I       ^I      L       �U#PL      U       _U      `       ^`      �       R�      �       w �      �       R                                  �       U�             �U�      )       U)      �       �U��      �       U                                      �        T�       L       XL      ]       T]      J       XJ      �       P      )       T�      �       X                            t        Qt       �       ��}                            �        R�       �       ��}                            |        X|       �       ��}                            �        Y�       �       ��}                              �       �      )       ��      �       �                            �      �       U�      �       ��}4�      �       ��|�1�             ��|�1�)      ]       ��|�1�]      v       r�                            A      V       PV      [      	 p ��|���      �      	 p ��|���      �       | r �$��|���      �       Pt      �       U�      �       | ��|�{ �$�                                L       0�d      j       ��}j      �       T�      �       ��}�      �       T�      �       ��}                                   R      �       	���      �       Q�      )       Z)      =       Q=      �       Z      �       Q�      �       q��      �       T�      �       Q)      v       Q                                           h       �        T�       �        ?��              T             t�      /       T7      L       	��]      �       T�      �       ��}      &       P&      *       p�J      �       0��      �       S             S)      v       S�      �       T�      �       t��      �       T                                                   �       �        1��       �        P�       �        p��       �        r�)      L       0�L      Y       PY      ]       R�      �       0��             Q      v       Q�              T              R=      o       Uo      �       T�      �       T�      �       t��      �       T}      �       R�      �      
 1��|�1$��      �       R�      �       0�                        �      �       ��|             ��|)      b       ��|f      v       U                           �       �        P�       �        q �              Y      L       0�L      ]       q ]      �       Y�      �       Y                 �      �       1{ $1��      �       1r $1�                 		

                                       ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               W               ��}�               ��}�               ��}�               ��}�               ��}�       h        ��~�h       �        U�       �        P7      L       ��}��      �       ��}��      �       p 2$� "
8��      �       p 2$� "
<��             p 2$� "
8�             p 2$u "�      *      
 p 2$u "#�*      4      
 p2$u "#�R      �       �      >       �a             �             PL      ]       �#�]      �       ��      �       ��}�                         R      �       0��      P       ^      �       ^             ^)      v       ^                                                       �       �0���      �       ���}��      �       �Y����}��             T�Y����}�             T�Y��_�      �       ���}�      #       ���}�#      D       �X����}�D      a       �X��a      �       T�X����}��      �       T�X��V��            
 �X��V�      )       �0��)      L       �X��L      X       T�X��X      ]       T�X��U�]      v       ���}��      �       �0��                              R      �       [�      )       X)      =       [=      �       X      �       [�      �       R�      �       R�             [)      �       [                                    7      L       ��~��      �       ��~��      �       p 2$� "���      �       p 2$� "���             p 2$� "��V      [       ��}4��      �       ��}4��      �       ��}�      �       _�      �       |��      �       _�      �       ��~�                                               p z �      L       S�      �       p q 2$� "
@���      �       P�      �       p 1$��      �       P�      �       p q 2$� "
@���      �       S�      �       p q 2$� "
@���      �       S                            R      �       0��      �       P)      7       P=      =      	 ��}�x �=      [      # ��}�x ������|�����-( �[      o       1u $��      �      # ��}�x ������|�����-( ��      �       1t $�             P)      v       P                     
      $
       U$
      %
       �U�                     
      $
       T$
      %
       �T�                    @
      U
       UU
      [
       �U�                    @
      L
       TL
      [
       �T�                    @
      Q
       QQ
      [
       �Q�                     @
      L
       q ����t �����L
      U
       TU
      [
       �Q�����T�����                   @
      V
       0�V
      [
       P                                   /       U/      %       S%      -       �U�-      �       S�      �       U�      �       S                                     D       TD      �       V-      >       V>      l       T�      �       V�      �       T�      �       V                   �             ]l      v       ]�      �       ]                   �             ^l      v       ^�      �       ^                   �             Sl      v       S�      �       S                     �      �       P�             Vl      v       V�      �       V                                �*      +       U+      f+       Sf+      n+       �U�n+      �+       S�+      �+       �U��+      �+       S�+      �+       �U��+      �,       S                                  �*      +       T+      +       V+      �+       �T��+      �+       T�+      �+       V�+      �+       �T��+      �+       V�+      O,       �T�O,      �,       V                              �*      +       Q+      )+       ])+      �+       �Q��+      �+       Q�+      �+       ]�+      �+       �Q��+      �,       ]                              �*      +       R+      )+       \)+      �+       �R��+      �+       R�+      �+       \�+      �+       �R��+      �,       \                     )+      e+       \e+      n+       0�n+      �+       \�+      �+       \                          )+      I+       ^T+      m+       ^m+      n+       Pn+      |+       ^�+      �+       ^�+      �+       P                  �+      �+       P                    A+      F+       VF+      i+       \n+      �+       V                  �+      �+       SO,      �,       S                 �+      �+       s                     �+      �+       PO,      X,       P                    O,      T,       s�T,      X,       UX,      �,       s�                       �+      ,       V,      ,       0�,      1,       V1,      4,       v q �4,      O,       V                  �+      O,       S                    �+      B,       0�B,      M,       P                    �+      ,       Q,      ,       V,      A,       Q                        �             U             S      $       �U�$      �	       S                          �             T      $       �T�$      �       _�      �       T�      �	       _                          �             Q      $       �Q�$      �       \�      �       Q�      �	       \                                 �             0�             V      $       P$      �       V�      v       0�v      �       1��      �       0��      �	       V�	      �	       1��	      �	       V                                         �      !       ^!      $       �U#L$      H       ^O      O       0�O      n       ^n      �       P�      �       ^�      �       Q�      G	       ^G	      [	       Q[	      o	       ��o	      �	       ^�	      �	       ���	      �	       ^�	      �	       P�	      �	       ^                                   �             ]      $       �U#H$      K       ]O      O       0�O      �       ]�      �       w �      n       ]n      �       P�      B	       ]B	      G	       QG	      �	       ]�	      �	       P�	      �	       ]                                        �      �       P�             w              P      $       ��$      W       w W      �       0��      �       w �      �       P�             
 ��      �       w �      	       Po	      �	       w �	      �	       0��	      �	       P                           $      O       PW      [       P�      �       P�      �       P�      	       P�	      �	       P                                       $      O       P�      �       P�      �       Q�      �       P             Q=      l       Ql      �       ���      	       P2	      B	       ]B	      [	       Q[	      o	       ���	      �	       ���	      �	       P                   �      �       So	      �	       S                    �      �       [�      �       ��o	      �	       [                    �      �       [�      �       ��o	      �	       [                    �      �       Uo	      �	       U                      �             U      T       ST      g       �U�                  �      f       V                 �             U                                  U      �       Q                 p      �       Q                                 h       Uh      �       S�      �       �U��      �       U�      �       �U�                    4      l       Z�      �       Z                   4      X       Q�      �       Q�      �       0�                       4      4       Q4      E       VE      X       @<$�[      �       V�      �       V�      �      
 q 1%q "#�                        p       �        U�       �       S�      �       �U��      �       S                          �       J       VR      e       Re      s       vx�s      �       R�      �       V�      �       9��      �       V                            �       �        u�       �        U�       �        ss      �       T�      �       s�      �       U�      �       s                    M      M       QM      V       q�V      �       X                  O      �       P                   �       >       S�      �       S                    �       >       P�      �       P                          �      �       U�      <       S<      D       �U�D      N       UN      �       S                          �      �       T�      =       V=      D       �T�D      N       TN      �       V                    �      ?       \N      �       \                           �             0�             P      7       ]D      N       0�N      �       ]�      �       0��      �       ]                 N      �       V�      �       V                 N      �       S�      �       S                 N      �       ]�      �       ]                  _      �       ^�      �       ^                    �      �       P�      �       P�      �       ��                    �	      
       U
      �       �U�                        �	      �	       T�	      !
       V!
      ~
       �T�~
             V      �       �T�                        �	      �	       Q�	      y
       ]y
      ~
       �Q�~
      �       ]                            �	      �	       R�	      B
       \B
      ~
       �R�~
      �       \�      �       �R��      �       \                    �	      t
       S~
      �       S                     �	      �	       R�	      l
       \l
      l
       0�~
      �       \�      �       \                       �	      �	       Q�	      y
       ]y
      ~
       �Q�~
      �       ]                       �	      �	       T�	      !
       V!
      ~
       �T�~
             V      �       �T�                   �	      t
       S~
      �       S                          �	      B
       0�B
      Y
       _^
      l
       _~
      �       0��      �       _�      �       _�      �       0�                 �
      �
       0�                   E
      S
       VS
      l
       \�      �       V                 �      �       S                     �      �       s��      �       U�      �       s�                  �      �       P                 �      �       0�                ~
      �
       S                 ~
      �
       s                   �
      �
       P                 �
      �
       s�                                      V       #       v q �#      b       Vb      i       v�`�i      �       V�      �       V�      �       0�                          �       S�      �       S                         �       0��      �       0�                        9       Q                       9      o       
 �o      t       
 �t      �       ^�      �       ^                      O      o       P�      �       P�      �       P                      p      �       U�      �       V�      �       �U�                  x      �       S�      �       0�                   x      �       u8�      �       \                 �      �       S                                              U               S               �U�       G        SG       H        �U�H       b        Sb       c        �U�                             1        P2       F        PH       ]        P                                                        �l      �l       U�l      �q       ^�q      �r       ��~�r      (t       �ط~8�(t      Ct       ^Ct      �z       ��~�z      �z       �ط~8��z      r�       ��~r�      ��       ^��      0�       ��~0�      I�       ^I�      �       ��~�      �       q�~�      O�       ��~O�      [�       q�~[�      c�       ��~c�      ��       �ط~8���      ��       ��~��      ��       �ط~8���      �       ��~                                  �l      �l       T�l      �q       S�q      (t       �T�(t      Ct       SCt      r�       �T�r�      ��       S��      0�       �T�0�      I�       SI�      �       �T�                            �l      m       Qm      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      �       ���~                            �l      *m       R*m      �       �ȷ~�      �       qȷ~�      O�       �ȷ~O�      [�       qȷ~[�      �       �ȷ~                    �l      �n       X�n      �       �X�                  �l      �n       Y                  �l      �n       �                           �l      �       ��      �       q�      O�       �O�      [�       q[�      �       �                                 �l      �r       0��r      �r       ](t      �z       0��z      �z       P�z      �z       0��z      �z       ]�z      V�       0�V�      c�       Pc�      �       0�                                    �l       m       P m      �n       ~��n      �r       ���~(t      �z       ���~�z      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      W�       ���~��      �       ���~                                  bm      �m       T�m      �p       _�p      (t       �ط~(t      Ct       _Ct      �       �ط~�      �       qط~�      O�       �ط~O�      [�       qط~[�      �       �ط~                       bm      �q       \(t      Ct       \r�      ��       \0�      I�       \                           bm      �n       ~8�n      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      �       ���~                       bm      �q       v @$�(t      Ct       v @$�r�      ��       v @$�0�      I�       v @$�                	                                             bm      �q       0��q      �r       ��~(t      Ct       0�Ct      �z       ��~�z      r�       ��~r�      ��       0���      0�       ��~0�      I�       0�I�      �       ��~�      �       q�~�      O�       ��~O�      [�       q�~[�      X�       ��~e�      �       ��~�      �       P�      !�       ��~!�      y�       0�y�      ��       1���      ��       0���      ��       Y��      ��       0���      �       2��      ��       ��~��      ��       0���      ��       ��~��      '�       0�'�      �       ��~                
                                   bm      �q       0��q      �r       ���~(t      Ct       0�Ct      �z       ���~�z      r�       ���~r�      ��       0���      0�       ���~0�      I�       0�I�      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      3�       ���~3�      7�       P7�      ٕ       ���~��      :�       ���~��      T�       ���~T�      [�       0�[�      �       ���~                                           bm      �q       0��q      �r       ���~(t      Ct       0�Ct      �z       ���~�z      G{       ���~G{      C|       1�C|      r�       ���~r�      ��       0���      0�       ���~0�      I�       0�I�      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      �       ���~                                                                bm      �q       0��q      �r       ���~(t      Ct       0�Ct      �z       ���~�z      �       ���~	�      r�       ���~r�      ��       0���      0�       ���~0�      I�       0�I�      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      ��       ���~��      X�       ���~e�      .�       ���~;�      ��       ���~��      �       P�      !�       ���~!�      �       0��      �       ���~��      Ė       0�Ė      ̖       P̖      �       ���~�      ��       0���      -�       ���~��      �       ���~                       bm      �p       ]�p      �p       ��~(t      6t       ]6t      Ct       ��~                                                                                                                                                                                                                       bm      3q       0�3q      �r       _(t      Ct       0�Ct      x       _x       x       U x      �x       _�x      �x       U�x      �z       _�z      �z       _�z      {       U{      l|       _l|      �|       U�|      �|       _�|      �|       U�|      X~       _X~      \~       Q\~             _      4       U4      �       _�      �       U�      X�       _X�      k�       Uk�      ��       _��      ۄ       Uۄ      �       _�      0�       U0�      I�       0�I�      q�       _q�      ��       U��      <�       _<�      ��       U��      ��       _��      ��       U��      �       _�      *�       U*�      ?�       _?�      C�       UC�      �       _�      '�       U'�      ׌       _׌      �       U�      �       _�      a�       Ua�      ��       _��      ȍ       Uȍ      +�       _+�      q�       Uq�      ��       _��      w�       Uw�      ��       _��      ʏ       Uʏ      ֏       _֏      ��       U��      ��       _��      ��       U��      �       _�      �       U�      <�       _<�      ��       U��      ��       _��      �       U�      ϒ       _ϒ      �       U�      �       _�      M�       UM�      i�       _i�      ��       U��      Z�       _Z�      h�       Uh�      ��       _��      ��       U��      �       _�      �       U�      i�       _i�      ��       U��      ��       _��      ݖ       Uݖ      �       _�      �       U�      ��       _��      �       U�      �       _�      >�       U>�      ��       _��      �       U�      ��       _��      ��       U��      ՙ       _ՙ      ޙ       Uޙ      ��       _��      �       U�      �       _�      �       U�      =�       _=�      [�       U[�      j�       _j�      v�       Uv�      �       _�      �       U�      3�       _3�      ?�       U?�      �       _                            �p      (t       �з~Ct      �       �з~�      �       qз~�      O�       �з~O�      [�       qз~[�      �       �з~                                                                                            �q      |r       S�r      �r       S�r      �r       r �r      �r       SCt      �t       S�u      �u       S�v      �v       S�w      x       SGx      jx       S�x      Jy       S"z      Kz       S�z      �z       S{      P{       SC|      _|       S�|      �|       S^}      �}       S
~      .~       S�~      �~       S�      ��       S�      ;�       S;�      ځ       ���~	�      C�       S��      �       SI�      u�       SI�      o�       So�      s�       P��      q�       S��      ��       SQ�      Z�       SZ�      _�       P_�      ��       S��      ̇       SJ�      X�       S�      �       S;�      L�       S�      ��       SD�      V�       Sc�      ��       S                                               bm      �q        -1��q      Br       ���~Br      Gr      	 ���~�1�Gr      �r       ���~(t      Ct        -1�Ct      �z       ���~�z      r�       ���~r�      ��        -1���      0�       ���~0�      I�        -1�I�      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      �       ���~��      	�       ���~��      �       ���~                                       bm      aq       0�aq      �q       P(t      Ct       0�9�      D�      	 �ȹ~p "�D�      L�       PL�      �       w r�      ��       0�9�      A�      	 �ȹ~p "�A�      R�       P��      I�       w 0�      I�       0���      ��       w e�      ��       w                                                      bm      jq       	��jq      �q       0��q      �r       ���~(t      Ct       	��Ct      �z       ���~�z      �{       ���~�{      �{       S�{      �{       p��{      |       PC|      r�       ���~r�      ��       	����      ��       ���~��      ��       P��      <�       ���~I�      0�       ���~0�      I�       	��I�      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      �       ���~��      �       ���~                    �z      {       P{      {       q�                          �z      �z       P<�      A�       PA�      y�       Sy�      $�       ���~?�      J�       ���~                       <�      y�       ��~#`�y�      $�       ~� �$�      ?�       ��~#`�?�      J�       ~� �                       <�      A�       PA�      y�       Sy�      $�       ���~?�      J�       ���~                               <�      ��       U��      ��       _��      ��       U��      �       _�      *�       U*�      1�       _?�      C�       UC�      J�       _                            e�      y�       Vy�      ��       Y��      ��       T��      ވ       Zވ      �       T�      $�       Y                  a�      y�       [                     e�      �       0��      $�       1�?�      J�       0�                   ��      ��       1��      �       1�                    ^�      1�       ]?�      J�       ]                               ^�      ��       U��      ��       _��      ��       U��      �       _�      *�       U*�      ?�       _?�      C�       UC�      J�       _                        ��      ��       S��      ��       s|���      $�       S?�      J�       S                      ��      ��       Pۈ      ވ       x p "�ވ      �       X                  ��      ͈       P                 ��      ψ       s|                   ͈      ψ       Pψ      ψ      
 p q "#���                  ͈      ψ       p ?&�ψ      ψ       Q                   �      �       [?�      J�       [                     �      �       U?�      C�       UC�      J�       _                     �      $�       U?�      C�       UC�      J�       _                       �|      �|       0��|      }       V}      0}       v~�0}      4}       V                    �|      �|       P�|      4}       S                 �|      4}       _                       _|      l|       0�l|      �|       \�|      �|       |��|      �|       \                    \|      l|       Pl|      �|       V                  _|      �|       S                    l|      w|       P�|      �|       P                       L|      l|       _l|      �|       U�|      �|       _�|      �|       U                 M}      ^}       _                        $�      ;�       P;�      �       ]Q�      X�       P��      <�       ]                           $�      ;�       0�;�      B�       VB�      H�       vz�H�      L�       TL�      Ɂ       vz�Ɂ      ځ       VQ�      X�       0�                    Z�      ^�       P^�      ��       Z                    l�      p�       Pp�      ��       [                  x�      ˁ       ^                  ��      ��       X                    ;�      B�       \��      ځ       \                    ;�      B�       S��      ځ       S                     �      �       _Q�      X�       _��      <�       _                 7�      <�       _                      M�      o�       P�      ��       P��      �       P                    s�      x�       Px�      �       Q                      �      �       P�      )�       ���~� $ &#�)�      9�       P                 �      H�       ���~�                 H�      H�       P                  �      )�       ��                  �      )�       Q                    ��      �       w ��      ��       w e�      ��       w                  ��      ��       P                        ��      �       ���~��      ��       S��      ��       ���~e�      j�       Sj�      ��       ���~                        ��      �       P��      ��       P��      ��       Te�      ��       P                ��      2�       w                  ��      �       P                ��      2�       ���~                    �      �       P�      "�       R                      ��      ��       P��      ڌ       [��      ȍ       [                      ��      ��       P��      n�       Z��      ȍ       Z                      ��      ��       P��      �       Y��      ȍ       Y                    ��      ڌ      	 z p { ���            	 z p { �                   ��      �       2���      ȍ       2�                   ��      �       U��      ȍ       U                         Ì      �       U�      ��       _��      a�       Ua�      n�       _��      ȍ       U                    ��      �      	 y z p ���      ��      	 y z p �                   ��       �       4���      ��       4�                   ��       �       U��      ��       U                     ��      a�       Ua�      n�       _��      ��       U                  ��      ��       P                    �      ��       P��       �       T                  Қ      ��       P                    ͚      њ       Pњ      Ԛ       T                  ��      ��       P                            ��      
�       P
�      ��       ]g�      ��       P��      ��       ]B�      O�       PO�      Ԙ       ]                        ��      ��       V�      �       P�      �       V>�      w�       V                      ��      ��       \�      �       P>�      ��       \                       	�      �       R���      �       ���~���      �      	 ���~�R��      ��       ���~����~�                   :�      >�      	 R����~�>�      ��       ���~����~�                      3�      ��       X��      �       X�      >�       X                        ;�      ?�       P?�      ��       \��      �       \�      >�       \                        B�      F�       PF�      ��       V��      �       V�      >�       V                              J�      N�      	 p  $ &�N�      ��       w � $ &���      ��       w � $ &���      җ       ��~� $ &�җ      K�       w � $ &�K�      ��       ��~� $ &���      ��       w � $ &�                          R�      ��      	 s  $ &���      �       S��      �       S�      9�      	 s  $ &�9�      ��       S                      c�      n�      	 p  $ &�n�      S�       ��~� $ &���      ��       ��~� $ &�                    ȕ      �       R�      �       ���~                    ܕ      �       Q�      9�       ���~                    �      *�       T*�      =�       t0�=�      ��       ���~#0�                       ��      B�       ]B�      ��       ���~��      ��       P��      ��       ���~                         ��      5�       �л~�5�      >�       Q>�      s�       �л~�s�      w�       Tw�      ��       �л~�                   ��      ߗ       Uߗ      �       }                 ��      ��       ���~                 ��      ��       �л~�                   ��      ��       Q��      Ƙ       ���~#                  ǔ      �       P                          Ɣ       PƔ      �       T                 ��      �       ���~                  c�      m�       P                  6�      =�       P                    1�      5�       P5�      8�       T                  �      �       P                    �      �       P�      �       T                    �      �       PT�      [�       P                        �      �       P�      �       XO�      S�       PS�      [�       X                    Ι      י       Pי      ޙ       p �                  _�      m�       P                    Z�      ^�       P^�      e�       T                                         �      �       P�      q�       Y��      ��       Yڎ      w�       Y��      Ώ       Y֏      R�       YR�      e�       Q��      ʐ       Y��      �       Yϒ      ��       Y�      �       Y��      �       Y��      '�       Y                                             �      q�       X��      Ď       Xڎ      �       X'�      w�       X��      Ώ       X֏      K�       X��      �       Xϒ      ��       X�      �       Xi�      �       X��      Ė       XĖ      ̖       P̖      �       ���~�      ��       X��      '�       ���~                                                                !�      C�      	 up 8�C�      q�      
 uu8���      ��      	 up 8�ڎ      ��      	 up 8�'�      H�      	 up 8���      ��      	 up 8�֏      �      	 up 8��      �      	 up 8�%�      3�      	 up 8�B�      e�      	 up 8���      �      	 up 8���      ��      	 up 8�      �      	 up 8��      �      
 uu8��      �      
 8�ϒ      �      	 up 8��      ��      	 p 8��      -�      	 up 8�-�      M�      
 uu8�M�      i�      
 8�i�      �      	 up 8��      ��      
 uu8���      ��      
 8���      ��      	 up 8���      ̖      
 uu8�                                                            
�      !�       0�!�      C�       up 8x �C�      q�       uu8x ���      ��       up 8x �ڎ      �       up 8x �'�      H�       up 8x ���      ��       up 8x �֏      �       up 8x ��      �       up 8x �%�      3�       up 8x �B�      K�       up 8x ���      �       up 8x ���      ��       up 8x �      �       up 8x ��      �       uu8x ��      �       8x �ϒ      �       up 8x ��      ��       p 8x ��      �       up 8x �i�      �       up 8x ��      ��       uu8x ���      ��       8x ���      ��       up 8x ���      ̖       uu8x �                 ��      _�       S                    *�      7�       P7�      g�       p�                   �      �       Q�      ϒ       ���~                 �      �       1�                    ��      ��       S�      ��       S                    ʐ      ��       Y�      ��       Y                     �      n�       0�n�      ��       1��      ��       0�                         �      �       1��      '�       ['�      <�       {�@�      ��       [�      ��       [                                �      �       \�      �       V�      �       T�      '�       { ~ "#�'�      <�       { ~ "�@�      ��       T��      ��       V�      ��       T                       �      �       up 8x ��      E�       ZE�      r�       z�r�      ��       Z�      ��       z�                    �      �       P9�      <�       } p "�                 �      -�       V                  �      +�       P                   +�      -�       P-�      -�      
 p q "#���                  +�      -�       p ?&�-�      -�       Q                   E�      n�       Z�      ��       Z                     E�      n�       U�      �       U�      ��       _                       I�      ��       U��      ��       _�      �       U�      ��       _                  f�      ��       P                  R�      ��       Y                  ;�      B�       P                    6�      :�       P:�      =�       T                  �      �       P                    �      �       P�       �       T                  �      �       P                  �      ��       T                �      ��       T                 �      �       P                   �      ��       P��      ��      
 p q "#���                  �      ��       p ?&���      ��       Q                  ��      Ώ       P                  ��      Ώ       T                  L�      w�       T                 '�      H�       ���~#�	                  ��      '�       P                 ڎ      ��       ���~#�	                  Ў      ֎       P                    ˎ      ώ       Pώ      ؎       T                    Ď      Ȏ       PȎ      ڎ       X                    ��      ��       P��      ڎ       Y                    P�      Z�      	 q 
��#�Z�      q�       r�	�
��#�                    P�      W�       QW�      f�       Pf�      f�       p t '�                     Ė      ̖       1�̖      �       T��      '�       T                                                                     !�      q�       Uq�      ��       _��      w�       Uw�      ��       _��      ʏ       Uʏ      ֏       _֏      ��       U��      ��       _��      ��       U��      �       _�      �       U�      <�       _<�      ��       U��      ��       _��      �       U�      ϒ       _ϒ      �       U�      �       _�      M�       UM�      i�       _i�      ��       U��      �       _��      ݖ       Uݖ      �       _�      �       U�      ��       _��      �       U�      '�       _                 ��             U                 �      �       ���~                 �      ��       6�                 #�      >�       ���~�>�      i�       �й~�                 J�      d�       �ط~                 J�      d�       ���~�                 >�      i�       �й~�                  x�      ��       P                  s�      ��       T                  Q�      h�       P                  <�      B�       P                    7�      ;�       P;�      D�       T                    0�      4�       P4�      I�       X                    (�      ,�       P,�      I�       Y                    ��      �      	 q 
��#��      �       r�	�
��#�                    ��      ��       Q��      �       P�      �       p t '�                  7�      =�       P                  2�      G�       T                7�      ?�       T                 7�      =�       P                   =�      ?�       P?�      ?�      
 p q "#���                  =�      ?�       p ?&�?�      ?�       Q                        ��      ��       P��      ��       S��      ��       V��      ƙ       S                  ��      ��       P                    ��      ��       P��      ƙ       P                    ~�      ��       P��      ��       T                    ��      ��       P��      ��       X                    ��      ��       P��      ��       T                    ��      +�       P�      �       P                          �       �       Q �      "�       q�"�      '�      
 uu3&�'�      +�      
 3&��      �       Q                    $�      +�       T�      �       T                     ��      '�       U'�      .�       _�      �       U                            #�      '�       P'�      ^�       X^�      a�       Pa�      ��       X՛      כ       Pכ      ��       X                    *�      7�       P7�      �       T                               *�      ^�       X^�      a�       Pa�      ՛       Q՛      כ       Pכ      ܛ       Xܛ      ޛ       Qޛ      ��       X�      �       Q                   *�      7�       P7�      �       T                   *�      ?�       U?�      �       _                          *�      ��       0��2����      ��       V�S���      Û       x ��Û      Ǜ       x �x�՛      ��       0��2���      �       V�S�                        ��      ��       ]��      Ǜ       PǛ      ՛       ]�      �       ]                              ��      ��       P��      ��       p t ���      ��       P��      ��       }���      Ǜ       PǛ      ɛ       p q "�ɛ      ћ       Pћ      ӛ       p t "�ӛ      ՛       P�      	�       P                      ��      ��       ^��      ��       ~���      ՛       ^�      �       ^                   ;�      ?�       U?�      �       _                   ��      ��       V����      ��       V�S�                  �      ��       ��                    �      ��       P��      ��                         ��      ń       P                 c�      ń       ���~                    Њ      Ԋ       PԊ      �       X                    ׊      ۊ       Pۊ      �       V                        �      )�       P)�      V�       ]��      ��       P��      �       ]                 Q�      �       ���~                 Q�      t�       �л~�                 ��      �       ���~                 ��      ܋       �л~�                Ey      �y       ���~                    Ey      �y       ��}��y      �y       P�y      �y       ��~                    Ey      �y       ��L��y      �y       P�y      �y       �ػ~                Ey      �y       ��~                    Ey      ]y       �л~�]y      py       Upy      �y       �л~�                 �y      �y       �ط~                 �y      �y       U                      �v      w       Vw      �w       \X�      _�       V                       �v      �v       0��v      w       ]w      lw       Slw      �w       sz��w      �w       SX�      _�       0�                    7w      ;w       P;w      �w       Z                    Iw      Mw       PMw      �w       [                  Uw      �w       ^                  aw      �w       X                  pw      �w       ]                  �w      �w       V                   �v      �w       _X�      _�       _                �      �       _                  �u      �v       S                      �u      �u       V�u      �u      	 p 3&��u      �u      
 3&�                       �u      �u       0��u      (v       V(v      dv       v|�dv      �v       V�v      �v       v��v      �v       p�                      �u      Sv       [�v      �v       P�v      �v       [                    v      v       Pv      Sv       Z                  v      �v       \                  ,v      Sv       X                 ,v      �v       \                  ?v      �v       ]                 �u      �v       _                      �t      �t       S�t      �u       S�      �       S                    �t      �t       V�t      �t      	 p 3&�                             �t      �t       0��t      �t       V�t      u       Vu      u       v�u       u       Y u      Nu       VNu      �u       v|��u      �u       V�      �       V                    7u      ;u       P;u      {u       Z                              �t      u       \u      u       ^u      u       Pu      Qu       \Qu      �u       ^�u      �u       ^�      �       ^                  Cu      {u       [                      Qu      �u       \�      ��       \��      �       �                     fu      �u       ]�      �       ]                     fu      �u       \�      ��       \��      �       �                      �t      �t       _�t      �u       _�      �       _                 �      �       _                      �~      �~       R�~      �       ���~�      0�       ���~                    �~      �~       Z�~      �~      	 p 3&�                     �~      �~       0��~             ZW      �       Z�      �       z��      +�       Z+�      0�       z�                    �~      �~       ^      �       ^                        �~      �~       P�~      8       [�      �       [�      0�       [                            �~      �~       R�~             �Է~      8       R�      �       R�      �       �Է~�      0�       �Է~                            W       V�      �       V+�      0�       V                       �~      W       ]�      �       P�      �       ]�      0�       ]                                8       X�      �       X�      �       S�      �       X�      0�       X                            W       S�      �       S�      0�       S                   �t      �t       _a�      r�       _�      �       _                         �~             _      4       U4      �       _�      �       U�      0�       U                 �t      �t       t 8$p !0$0&�                      �t      �t       P�t      �t       T��             T                  �t      �t       P                   I�      V�       p�~�V�      c�       T                       ��      Â       s ��Â      ؂       R؂      ؂       r p "�؂      �       p r "#l�a�      q�       R                       Y�      _�       s ��_�      |�       R|�      ��       	�r ���      ��       TJ�      X�       R                  
�      Q�       T                    ��      ��       R��      �       R                    Æ      ��       T��      ȉ       T                    ܆      �       X��      ��       X                  �      �       P                         �n      �       �ȷ~�      �       qȷ~�      O�       �ȷ~O�      [�       qȷ~[�      �       �ȷ~                    �n      ]o       ~��]o      �o       P�o      {p       ��~                �n      {p       ]                    �n      p       ���~�p      "p       Q"p      {p       ��~                    �n      �o       ���~��o      p       Qp      {p       ��}                    �n      Oo       �й~�Oo      �o       Q�o      {p       ��}                  �n      �n       ~8�n      {p       ���~                �n      {p       ���~                �n      {p       ^                    �n      �n       U�n      �n       ���~��n      {p       T                �o      �o       U                �o      �o       ��}�                �o      �o       ��L                �o      �o       ^                �n      �o       @�                �n      �o       _                �n      �o       \                �n      �o       ��}�                �o      �o       U                �o      �o       ��}�                �o      �o       ��L                �o      �o       ^                �o      �o       ����                �o      �o       U                �o      �o       ��}�                �o      �o       ��L                �o      �o       ^                �o      �o       ���~�                 �m      �m        �                 �m      �m       T                 �m      �m       \                 �m      �m       ���~�                 �m      On       D�                   �m      �m       T�m      On       _                 �m      On       \                 �m      On       �й~�                 On      �n       D�                 On      �n       _                 On      �n       \                 On      �n       ���~�                �n      �n       _                �n      �n       ���~�                                   �p      �p       R�p      �r       ���~(t      Ct       RCt      �z       ���~�z      �       ���~�      �       q��~�      O�       ���~O�      [�       q��~[�      W�       ���~��      �       ���~                 �p      �p       R                 �p      3q       �з~0�      D�       �з~                   �p      �p       _�p      3q       �ط~0�      D�       �ط~                 �p      3q       \0�      D�       \                        �p      �p       0��p      �p       P�p      3q       _0�      9�       _9�      C�       TD�      D�       0�                   3q      Eq       A�r�      ��       A�                       3q      Eq       ���~�r�      ��       ���~���      ��       U��      ��       ���~�                 |r      �r       _                   �r      �r       ]�z      �z       ]                   �r      �r       �ط~�z      �z       �ط~                 �r      0s       ���~�                 �r      0s       ��}�                	 �r      s       ��}                 0s      us       ���~�                 0s      Xs       U                 us      �s       �й~�                 us      �s       U                 �s      �s       ���~�                 �s      �s       U                �s      t       _                 �s      t       S                 Qt      ft       _                   �w      x       _̅      �       _                     Gx      �x       _�x      �x       Uk�      ��       _                   �x      "z       _��      ��       _                 G{      h{       ���~�h{      C|       �й~�                 t{      �{       �ط~                 t{      �{       ���~�                 h{      C|       �й~�                 �{      �{       P                �{      �{       ���~�                 �{      �{       ��                 �{      �{       ���~                   ^}      �}       _��      ̅       _                      ��      �       P�      +�       ���~� $ &�+�      9�       P                 ��      M�       ���~�                 M�      M�       P                  �      +�       ��                  �      +�       R                     L�      �       _D�      V�       _c�      ��       _                       �      ��       ���~�D�      L�       ���~�L�      P�       UP�      V�       ���~�                 ��      �       _                        `Y      �Y       U�Y      �Z       S�Z      �Z       �U��Z      @[       S                        `Y      �Y       T�Y      �Z       ]�Z      �Z       �T��Z      @[       ]                        `Y      �Y       Q�Y      �Z       V�Z      �Z       �Q��Z      @[       V                        `Y      �Y       R�Y      CZ       w CZ      �Z       ��~�Z      @[       w                       `Y      Z       XZ      �Z       �X��Z      @[       X                            `Y      Z       YZ      �Z       �Y��Z      �Z       Y�Z      �Z       �Y��Z      [       Y[      @[       �Y�                             �Y      �Y       0��Y      �Y       T�Y      �Y       ^�Y      -Z       T�Z      [       T[      [       Y[      )[       T                       �Y      ;Z       | �0)��Z      �Z       | �0)��Z      �Z       | �0)��Z      3[       | �0)�                         �Y      �Y        �#	��Y      ;Z       | �0.�#	��Z      �Z       | �0.�#	��Z      �Z       | �0.�#	��Z      3[       | �0.�#	�                   �Y      �Y       0��Y      �Y       p�                     ?Z      hZ       0�hZ      �Z       1��Z      �Z       2�                   )Z      ?Z       y  $x  $+��Z      �Z       y  $x  $+�                   .Z      ?Z       P�Z      �Z       P                   �Z      �Z       S�Z      �Z       �U�                   �Z      �Z       S�Z      �Z       �U�                         W      "X       U"X      �X       S�X      �X       �U��X      VY       S                           W      QW       TQW      `W       R`W      �X       ]�X      �X       �T��X      VY       ]                         W      KW       QKW      `W       X`W      �W       _�W      VY       �Q�                         W      6W       R6W      �W       \�W      �W       Q�W      VY       �R�                       W      =W       X=W      �W       V�W      VY       �X�                         W      \W       Y\W      �X       ^�X      �X       �U#Ȓ�X      VY       ^                         X      X       Z��X      "X       Z�_�"X      �X       �_��X      �X       Z�_��X      �X       ���_��X      VY       �_�                   X      X       \��X      �X       \�V��X      VY       \�V�                     X      X       [��X      "X       [�P��X      �X       [�P��X      �X      
 ������                 �W      �W       V                 �W      �W       \                 �W      �W       _                 �W      �W       ]                          �U      &V       U&V      rV       SrV      �V       �U��V      �V       U�V      W       S                        �U      �U       T�U      �U       \�U      |V       ]|V      W       �T�                        �U      �U       Q�U      �U       V�U      ~V       ^~V      W       �Q�                   V      V       \��V      rV       \�V��V      W       \�V�                  �V      �V       0�                        @T      UT       UUT      �T       S�T      �T       �U��T      �T       S                          @T      UT       TUT      �T       \�T      �T       �T��T      �T       T�T      �T       \                              @T      UT       QUT      �T       V�T      �T       Q�T      �T       s��T      �T       �Q��T      �T       Q�T      �T       V                   @T      UT       U�T      �T       S                              _       T_      �       �T��      �       T�      �       �T�                              f       Qf      �       �Q��      �       Q�      �       �Q�                              9       R9      �       �R��      �       R�      �       �R�                              B       XB      �       �X��      �       X�      �       �X�                          �       � �      �       Z                                        9       S9      �       R�      �       S�      �       R�             r �J      `       R`      m       r ��      �       R�      �       r �                                      B       PB      �       X�      �       P�             X`      c       Xc      y       x ��      �       X�      �       x ��      �       x �                 c      c       �X�                 c      c       �R�                 c      c       Q                �      �       u��                �      �       
3��                 �      �       P                �      �       p ?&�                 �      �       u��                 �      �       Ι}�                  �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       u��                �      �       
�L�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                             u��                             
3��                              P                             p ?&�                 �      �       u��                               P            
 p q "#���                               p ?&�             Q                )      9       u��                )      9       3� �                   7      9       P9      9      
 p q "#���                  7      9       p ?&�9      9       Q                        �T      U       UU      SU       SSU      WU       �U�WU      sU       S                    �T      TU       T�Q�WU      sU       \�V�                             N      _N       U_N      �O       S�O      �O       �U��O      \P       S\P      fP       �U�fP      `S       S                     N      �N       T�N      `S       ��~                             N      [N       Q[N      �O       ]�O      �O       �Q��O      aP       ]aP      fP       �Q�fP      `S       ]                   N      WN       R�X�                     N      |N       Y|N      `S       �Y�                        )N      )N       u���)N      IN       \IN      PN       u���PN      �N       \fP      Q       \                        PN      O       _fP      R       _,R      9R       _GS      [S       _                                      N      �N       0��0���N      �O       V�\��O      �O       �\��O      WP       V�\�fP      �P       0��0���P       Q       V�0�� Q      8Q       V�\�8Q      PQ       V�\�PQ      pQ       V�\�pQ      �Q       V�\��Q      `S       V�\�                            N      O       0��O      �O       0�fP      �Q       0��Q      ,R       1�,R      9R       0�GS      `S       1�                     iN      �N       SfP      ,R       SGS      `S       S                   iN      �N       \fP      Q       \                     iN      �N       _fP      R       _GS      [S       _                     iN      �N       ]fP      ,R       ]GS      `S       ]                     iN      �N       �7�  fP      ,R       �7�  GS      `S       �7�                       iN      �N       �  fP      ,R       �  GS      `S       �                        �N      �N       t p ��N      �N       TfP      �P       T                  �P      	Q       P                �N      �N       Y                 �N      �N       P                   �N      �N       P�N      �N      
 p t "#���                  �N      �N       p ?&��N      �N       T                �N      �N       X                  �N      �N       Q�N      �N      
 q ~ "#���                  �N      �N       q ?&��N      �N       ^                 fP      �P       Y                 fP      rP      
 r v #5&�                   �P      �P       Y�P      �P      
 p y "#���                  �P      �P       y ?&��P      �P       P                  �P      �P       Q�P      �P      
 q x "#���                  �P      �P       q ?&��P      �P       Q                      �P      �P       t x ��P      �P       Q�P      �P       t x �                  �P      �P       P                      �P      �P       Q�P      �P      
 q r "#����P      �P       U                   �P      �P       q ?&��P      �P       R                   �P      Q       RQ      Q       q y �                 �P      	Q       P                      Q      Q       RQ      Q      
 p r "#���Q      Q       P                     Q      Q       r ?&�Q      Q       PQ      Q       r ?&�                        ?      F?       UF?      �@       S�@      �@       �U��@      I       S                                    ?      P?       TP?      @       w @      S@       ��~S@      �@       w �@      �@       ��~�@      (A       w (A      ~A       ��~~A      �G       w �G      �G       T�G      I       w                                     ?      P?       QP?      g?       Vg?      �@       �Q��@      �@       V�@      F       �Q�F      �F       V�F      �G       �Q��G      �G       Q�G      �G       V�G      I       �Q�                        ?      P?       RP?      �G       ��~�G      �G       R�G      I       ��~                        ?      P?       XP?      �G       ��~�G      �G       X�G      I       ��~                        ?      P?       YP?      �G       �Y��G      �G       Y�G      I       �Y�                                       �?      �?       ����?      �?       ]�?      l@       ]�@      �@       ]�@      �A       ]E      WE       ]WE      F       ��~�F      �F       ]8G      JG       ��~JG      �G       ���H      3H       ���3H      I       ��~                            *?      �@       _�@      �A       _�C      ND       _E      �F       _8G      �G       _H      I       _                   �?      �?       w #(JG      qG       w #(                                          �?      �?       0��?      �@       V�@      �@       V�@      �A       VE      F       V�F      �F       V�F      �F       0��F      �F       r��F      �F       R�F      8G       r�8G      JG       VH      3H       0�3H      I       V                                        �?      �?       	���?      �?       \�?      �?       	���?      �@       \�@      �@       \�@      �@       \A      A       	��A      �A       \E      F       \�F      �F       \8G      JG       \H      3H       	��3H      I       \                   JG      `G       ��~�`G      mG       Q                           O@      c@       ��~�c@      l@       UE      3E       U3E      F       ��~�8G      JG       ��~�3H      I       ��~�                         c@      l@       UE      3E       U3E      F       ��~�8G      JG       ��~�3H      I       ��~�                       E      3E       U3E      
F       ��~�8G      JG       ��~�3H      I       ��~�                     E      
F       ��~�8G      JG       ��~�3H      I       ��~�                     E      
F       ��8G      JG       ��3H      I       ��                            E      �E       T�E      �E       �8G      JG       T3H      |H       T�H      �H       T�H      I       �                        �E      �E       PYH      H       P�H      �H       P�H      I       P                             E      �E       0��E      �E       Q8G      JG       0�3H      jH       0�jH      |H       Q�H      �H       0��H      I       Q                        E      �E       0��E      
F       1�8G      JG       0�3H      jH       0�jH      �H       1��H      �H       0��H      I       1�                           E      bE       0�bE      �E       Q8G      JG       Q3H      YH       Q�H      �H       Q�H      �H       Q                     bE      �E       ��~�3H      |H       ��~��H      �H       ��~�                   �E      �E       ��~��H      I       ��~�                 �E      F       ��~�                	  jH      �H       ��~��H      I       ��~�                   �C      D       ��~�D      D       T                 &D      0D       Q                   �F      �F       P)G      8G       P                      �F      G       PG      G       qG      %G       P                 �F      )G       U                 )G      )G       P                  G      G       ��                  G      G       X                   �F      �F       Q)G      8G       Q                �?      �?       ���                        �@      �@       R�@      �@       ~ v("��@      �@      
 ~ �Q#("�F      nF       R                    �@      �@       ��~F      �F       ��~                        FF      XF       0�XF      cF       p ��~ �cF      gF      
 p ��~O�gF      lF       p ��~ �                       �@      �@      
 1r 7$1��@      �@       1~ v(�7$1��@      �@       1�Q#(~ 7$1�F      nF      
 1r 7$1�                      �@      �@       R�@      �@       ~ v("��@      �@      
 ~ �Q#("�F      AF       R                  �@      �@       ��~F      AF       ��~                      �@      �@       R�@      �@       ~ v("��@      �@      
 ~ �Q#("�                  �@      �@       ��~                  �@      �@       B�                  �@      �@       P                     �A      �C       S8D      E       S�F      �F       S�G      H       S                                   �A      �A       0��A      �B       V*C      IC       [IC      TC       TTC      �C       t��C      �C       TDD      ND       0�ND      ]D       V�D      E       V�F      �F       0��G      H       V                    �C      �C       R�C      �C       r�                	   	 	 �A      �A       s�A      �A       P8D      ND       s�F      �F       s                           �A      �A      
 p < $0.��A      �B       v5$s "#�< $0.�ND      UD      
 p < $0.��D      �D       v5$s "#�< $0.��D      �D       v5$s "#�< $0.��G      
H       v5$s "#�< $0.�                           �A      �A       s u "#��A      �A       s u "H��A      �B      
 v5$s "#�ND      ]D      
 v5$s "#��D      E      
 v5$s "#��G      H      
 v5$s "#�                
           �A      �B      
 v5$s "#��B      �B       s u "#(�ND      UD      
 v5$s "#��D      �D      
 v5$s "#��G      �G      
 v5$s "#��G      �G       s u "#(�                            B      NB       XNB      �B       y 
����D      �D       y 
����D      �D       t 
����D      �D       y 
����G      
H       y 
���                            /B      HB       PHB      �B       z 
����D      �D       z 
����D      �D       | 5$s "#<�
����D      �D       | 5$s "#<�
����G      
H       z 
���                           /B      NB       x �NB      �B       y 
����D      �D       y 
����D      �D       t 
����D      �D       y 
����G      
H       y 
���                           /B      HB       p �HB      �B       z 
����D      �D       z 
����D      �D       | 5$s "#<�
����D      �D       | 5$s "#<�
����G      
H       z 
���                           /B      ]B       T]B      �B       @<$y 
��{ y 
�� $0.( ��D      �D       @<$y 
��{ y 
�� $0.( ��D      �D       @<$t 
��{ t 
�� $0.( ��D      �D       @<$y 
��{ y 
�� $0.( ��G      
H       @<$y 
��{ y 
�� $0.( �                              <B      AB       QAB      HB       @<$p { p  $0.( �HB      �B       @<$z 
��{ z 
�� $0.( ��D      �D       @<$z 
��{ z 
�� $0.( ��D      �D      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( ��D      �D      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( ��G      
H       @<$z 
��{ z 
�� $0.( �                          AB      �B       Q�D      �D       Q�D      �D      � @<$y 
��{ y 
�� $0.( @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( @<$y 
��{ y 
�� $0.(  $@<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.(  $,( ��G      �G       Q�G      
H      } @<$y 
��{ y 
�� $0.( @<$z 
��{ z 
�� $0.( @<$y 
��{ y 
�� $0.(  $@<$z 
��{ z 
�� $0.(  $,( �                          QB      �B       X�B      �B       p ��D      �D       X�G      �G       X�G      
H       p �                 �B      �B       X                     QB      �B       
 ���D      E       
 ���G      H       
 ��                     QB      �B       
 ���D      E       
 ���G      H       
 ��                     QB      �B       0��B      �B       q  $p  $-��D      �D       0��G      �G       0�                  �B      �B       s u "#(��G      �G       s u "#(�                  TC      vC       T                 TC      vC       ]                  `C      vC       ��                  `C      vC       P                 �C      �C       0�                 �C      �C       ��~                     �F      �F       Q�F      �F       q`��F      8G       Q                   �G      �G       Q�G      �G       r                    �G      �G       ����G      �G       R                            0      q       Uq             Y      !       U!      �       Y�      �       U�             Y                            0      u       Tu             �T�      !       T!      �       �T��      �       T�             �T�                                      0      �       Q�             �Q�      !       Q!      *       �Q�*             Q      �       �X�      �       �Q��      �       Q�      �       �X�      �       Q�             �Q�                        ]      �       0��      �       P*      ,       0��      �       0�                   5      ]       T      !       T                                     5      �       Q�             �Q�      !       Q!      *       �Q�*             Q      �       �X�      �       �Q��      �       Q�      �       �X�      �       Q�             �Q�                    �      �       P�      �       T                     �      �       r t "#��@&��      �      8 �X#�{�O%�X#�{�"1& $ &y� $ &t "#��@&��      �      g �X#�{�O%�X#�{�"1& $ &y� $ &�X#�{�O%�X#�{�"1& $ &y� $ &?&"#��@&�                �      �       y                �      �       �X#�{�2�                   �      �       R�      �      
 r t "#���                  �      �       r ?&��      �       T                      �             t�             U             u�      D       U                 �             T                        �             t z �             z  t "��      �       | z ��             z  | "�             p�                     �      �       [Y      �       [�      �       [�      �       [                       =      ?       p ����#5$y "#�?      C      
 r5$y "#�C      G      
 r 5$y "#�G      b       p ����#5$y "#�                                       �       T�      �       �T��      �       T�      �       �T��             T             �T�             T      (       �T�                                   :      P       PP      R       RR      u       Pu      �       R�      �       P�      �       Q�      �       P�      �       0�             P      (       u$                   �      �       P�      �      
 p r "#���                  �      �       p ?&��      �       R                 �             u                   �             t r �             �Tr �                 �      �       u                   �      �       T�      �       �T�                      �      �       T�      �      
 p t "#����      �       P                     �      �       t ?&��      �       P�      �       t ?&�                        p-      �-       T�-      �.       �T��.      �.       T�.      �.       �T�                        p-      �-       R�-      .       �R�.      6.       R6.      X.       �R�X.      �.       R                              p-      �-       X�-      .       �X�.      $.       X$.      X.       �X�X.      r.       Xr.      �.       �X��.      �.       X                                          �-      �-       T�-      
.       { p��.      6.       T6.      D.      
 p�p��X.      o.       To.      �.       p�z ��.      �.       T�.      �.       p�z ��.      �.       T�.      �.       { z ��.      �.       T�.      �.       { z ��.      �.       T�.      �.       { z �                       �-      
.       P.      D.       PX.      �.       P�.      �.       P                     �-      �-       Q�-      �-       P�.      �.       Q                  �-      �-       T�.      �.       T                 �-      �-       P                    �-      �-       ���.      �.       ��                    �-      �-       Z�.      �.       Z                 .      .       U                6.      H.       Y                 6.      A.       X                   A.      H.       XH.      H.      
 p x "#���                  A.      H.       x ?&�H.      H.       P                        �,      �,       U�,      �,       V�,      �,       �U��,      m-       V                        �,      �,       T�,      �,       �T��,      %-       T%-      m-       �T�                          �,      �,       Q�,      �,       S�,      �,       �Q��,      %-       Q%-      m-       S                 `-      d-       T                 �,      �,       P                     -      %-       T%-      Y-       �T�`-      `-       �T�                   -      Y-       \`-      `-       \                    &-      D-       0�D-      Y-       T`-      `-       T                   &-      Y-       P`-      `-       P                 -      %-       |�&                                              �      ^�       U^�      ��       _��      ��       �U���      �       _�      V�       �U�V�      x�       Ux�      �       _�      ��       �U���      �       _�      $�       �U�$�      2�       _2�      ��       �U���      ��       U��      �       �U��      *�       _                                              �      ^�       T^�      ��       V��      ��       ����      ��       �T���      ޡ       ��ޡ      V�       �T�V�      u�       Tu�      �       V�      ��       �T���      ˦       ��˦      ڦ       �T�ڦ      �       ���      ��       �T���      ��       T��      *�       �T�                                              �      ^�       Q^�      �       ^�      ��       �Q���      �       ^�      V�       �Q�V�      p�       Qp�      �       ^�      ��       �Q���      �       ^�      $�       �Q�$�      2�       ^2�      ��       �Q���      ��       Q��      �       �Q��      *�       ^                     J�      ^�       u V�      x�       u x�      ��                                  U�      ��       S��      ��       S��      ��       p ��      ��       S��      *�       S                         7�      �       \��      �       \V�      �       \��      �       \��      ��       \                                         t�      ٜ       s�ٜ      ��       _��      ��       �U���      �       _�      ��       �U���      V�       �U��      ��       �U���      �       _�      $�       �U�$�      2�       _2�      ��       �U���      �       �U��      *�       _                      ��      X�       P��      �       P��      �       P                        ��      ��       Y��      �       Y��      �       Y�      *�       Y                       ��      ��       X��      �       X��      �       X�      *�       X                          ��      ]�       0�]�      ��       s��      V�       0��      ��       0���      ��       0���      ʩ       sʩ      *�       0�                     ]�      x�       Qx�      ��       | ��      ʩ       ��~                           ̜      ��       q���      ġ       q�ġ      ޡ       #���      Ǧ       q�Ǧ      ˦       #�ڦ      �       #�                        Ӝ      ��       R��      �       R��      �       R�      *�       R                                         ̜      ٜ       s�ٜ      ��       _��      ��       �U���      �       _�      ��       �U���      V�       �U��      ��       �U���      �       _�      $�       �U�$�      2�       _2�      ��       �U���      �       �U��      *�       _                   ̜      �       �#�  ��      ѡ       �#�                     ̜      �       ��  ��      ѡ       ��                     ̜      �       �����      ѡ       ���                   ̜      �       �����      ѡ       ���                                   j�      ��       _��      ��       �U��      ��       �U���      V�       �U��      ��       �U��      $�       �U�$�      2�       _2�      ��       �U���      �       �U��      *�       _                     n�      ��       ���$�      2�       ����      *�       ���                     n�      ��       T��      ��       s��      *�       T                  ��      ��       P                              ��      ��       ���  �      ]�       ���  ��      V�       ���  �      ��       ���  �      $�       ���  2�      ��       ���  ��      ��       ���  ʩ      �       ���                                ��      ��       ����      ]�       �����      V�       ����      ��       ����      $�       ���2�      ��       �����      ��       ���ʩ      �       ���                                  ��      ��       ����      �       ����      �       T�      ]�       �����      V�       ����      ��       ����      $�       ���2�      ��       �����      ��       ���ʩ      �       ���                              ��      ��       S�      ]�       S��      V�       S�      ��       S�      $�       S2�      ��       S��      ��       Sʩ      �       S                             ��      ��       0��      ��       0���      V�       0��      ��       0��      $�       0�2�      ��       0���      �       0�                    գ      D�       V�      ��       V��      �       0�                               �      ��       ����      ��       �����      V�       ����      ��       ����      $�       ���2�      ��       �����      ��       ���ʩ      �       ���                               �      ��       S�      ��       S��      V�       S�      ��       S�      $�       S2�      ��       S��      ��       Sʩ      �       S                   �      =�       s�t�      ��       s�                            �      �       0��       �       1� �      S�       \S�      Y�       1�Y�      ˞       \˞      Ϟ       1�؞      ؞       1�<�      V�       \t�      ݧ       \�      �       1��      $�       \                     &�      =�       �#�'�t�      �       p�'��      ��       �#�'�                   �      &�       0�&�      =�       �#�'�0.�t�      ��       �#�'�0.�                         �      =�       [|�      ��       [t�      ��       [��      $�       w b�      m�       P                	           �      ߠ       ]<�      V�       ]�      ��       ]t�      $�       ]2�      m�       ]ʩ      �       ]                       
�      �       ^<�      V�       ^�      �       ^t�      $�       ^                            K�      \�       P\�      r�       u�#�
��@$��      C�       V4�      ��       V2�      m�       Vʩ      �       V                   &�      =�       s�t�      ��       s�                 ��      ��       s�                     ��      ��       ��~���      ��       R��      ��       ��~�                     ��      ��       ��~���      ��       T��      ��       ��~�                 ��      ��       s�#                 ��      ��       P                     �      2�       �B$x �ʩ      �       �B$x ��      ��       �B$��~��                    ��      ��       Q��      	�       Q                          ߞ      2�       X�      /�       X/�      4�       s�ʩ      �       X�      ��       ��~                  a�      ��       s��                  a�      ��       Y                  a�      ��       0�                  a�      ��       s��                  a�      ��       Q                  a�      ��       V                  П      �       s��                  П      
�       Y                  П      �       ]                  П      �       s��                  П      ݟ       s�                  П      �       V                           `�      ��       S�      ��       S��      <�       S�      t�       Sm�      ��       S��      ��       S                           `�      ��       s���      ��       s����      <�       s���      t�       s��m�      ��       s����      ��       s��                 `�      ��       V                            ��      ?�       Zs�      v�       q t �v�      ��       Z8�      :�       p r �:�      P�       PP�      _�       p r �_�      h�      	 q��r �                             `�      ��       0���      ��       \�      �       \��      <�       \�      >�       \m�      ��       \��      ��       0�                      y�      �       P��      <�       P�      �       P                     Ϡ      ��       Y�      x�       Y��      ��       Y                       נ      ��       X�      ��       X��      �       x���      ��       X                           ߠ      ��       ]�      ��       ]��      <�       ]�      t�       ]m�      ��       ]��      ��       ]                           �      ��       ^�      ��       ^��      <�       ^�      t�       ^m�      ��       ^��      ��       ^                      Ϡ      ��       v���      �       v����      <�       v����      ��       v��                      נ      ��       v���      �       v����      <�       v����      ��       v��                      ߠ      ��       v���      �       v����      <�       v����      ��       v��                      �      ��       v���      �       v����      <�       v����      ��       v��                               �      ��       0���      ��       R�      �       0�y�      ��       0���      �       [=�      a�       0�a�      ��       R��      <�       [                           �      ��       NB$��      ��       NB$���      <�       NB$��      t�       NB$�m�      ��       NB$���      ��       NB$�                           �      ��       �B$��      ��       �B$���      <�       �B$��      t�       �B$�m�      ��       �B$���      ��       �B$�                 ��      ��       V                 ��      ��       s��                 ��      ��       s��                 ��      ��       s��                ��      Ϡ       ��                  ��      Ϡ       ���                  Ϡ      נ       ��                  Ϡ      נ       ���                  נ      ߠ       �"�                  נ      ߠ       ���                  ߠ      �       �/�                  ߠ      �       ���                            ��      ��       2���      ��       X��      ��       0���      �       Y1�      <�       Y                              ��      ��       ������      �       Y�      ��       U��      ��       Y��      ��       ������      ۤ       Rۤ      �       X�      �       R1�      <�       X                      ͢      ��       R��      �       U��      <�       U                        ܢ      ��       Uˤ      �       X�      1�       Q1�      <�       X                      ��      ��       Q��      �       Q1�      <�       Q                �      [�       T                �      [�       ���|�                   T�      [�       Q[�      [�      
 p q "#���                  T�      [�       q ?&�[�      [�       P                ��      ��       T                  ��      ��       Q��      ��       s�                   ��      ��       P��      ��      
 p q "#���                  ��      ��       p ?&���      ��       Q                   ��      ��       s����      ��       ��~b�      m�       s��                   ��      ��       0�b�      m�       0�                   ��      ��       [b�      m�       P                   ��      ��       s����      ��       Rb�      m�       s��                   ��      ��       Qb�      m�       Q                   ��      ��       Vb�      m�       V                   �      ��       s���      �       s��                 �      ��       P                 D�      ��       s��                 D�      ��       V                 l�      ��       s��                    l�      x�       Qx�      ��       |                    l�      �       R�      ��       s�                 å      �       s�                 å      �       s��                            �]      �]       U�]      �]       \�]      �]       �U��]      �^       \�^      �^       �U��^      �^       \                            �]      �]       T�]      �]       V�]      �]       �T��]      �^       V�^      �^       �T��^      �^       V                     �]      �]       P�]      �]       P�^      �^       P                           �]      �]       U�]      �]       \�]      �]       �U��]      �^       \�^      �^       �U��^      �^       \                   �]      �]       t�]      �]       v                   �]      �]       t �]      �]       v                   �]      �]       0��]      �]       P                 �]      �]       3�                   �]      �]       0��]      6^       0�                   �]      �]       v�]      &^       v                   �]      �]       v�]      "^       v                    �]      �]       P�]      6^       P                  ^      -^       R                 ^      1^       Q                    �]      �]       0�6^      y^       0��^      �^       0�                    �]      �]       v(6^      i^       v(�^      �^       v(                    �]      �]       v 6^      e^       v �^      �^       v                   b^      p^       R                 b^      t^       P                  �]      �]       1�y^      �^       1�                 �]      �]       v8y^      �^       v8                 �]      �]       v0y^      �^       v0                  �^      �^       R                 �^      �^       Q                          �k      l       Ul      Ll       \Ll      Ol       �U�Ol      al       \al      hl       �U�                      �k      l       Tl      .l       V.l      hl       �T�                  l      l       P7l      Ol       P                         �k      l       Ul      Ll       \Ll      Ol       �U�Ol      al       \al      hl       �U�                      l      Il       SOl      ^l       S^l      gl       U                   
l      l       tl      l       Q                   
l      l       t l      l       T                
l      l       S                  
l      l       0�l      l       P                      .l      7l       ]Ol      cl       ]cl      gl       Q                      .l      7l       VOl      _l       V_l      gl       T                      .l      7l       SOl      ^l       S^l      gl       U                    3l      7l       POl      gl       P                     .l      7l       SOl      ^l       S^l      gl       U                 .l      3l       1�                    �<      �<       U�<      �<       �U�                    �<      �<       T�<      �<       �T�                   �<      �<       U�<      �<       �U�                  �<      �<       S                        �              U       $       S$      &       �U�&      I       S                          �             T      %       V%      &       �T�&      4       T4      I       V                    
             q u �             U                   
            
 q u s8"�             U                          0      [       U[      w       Sw      {       �U�{      �       S�      �       �U�                          0      [       T[      {       �T�{      �       T�      �       \�      �       �U#                   S      [       u {      �       s                        S      [       r t �{      �       r t ��      �       st ��      �       s| �                  �      �       ��                  �      �       P                  _      r       @�                  _      r       Q                           =      '=       U'=      �=       V�=      �=       �U��=      �=       U�=      	>       V                         =      '=       T'=      �=       �T��=      �=       T�=      	>       \                         =      '=       Q'=      �=       �Q��=      �=       Q�=      	>       �Q�                          =      '=       U'=      �=       V�=      �=       �U��=      �=       U�=      	>       V                    =      �=       S�=      	>       S                       =      '=       s��'=      �=       Q�=      �=       s���=      	>       Q                   =      '=       s�&�=      �=       s�&                      �=      �=       P�=      �=       Q�=      �=       P                 �=      	>       \                 �=      	>       |�                 Q=      r=       R                Q=      r=       t�                 r=      r=       P                  S=      r=       t�                  S=      r=       R                      �j      �j       U�j      Sk       SSk      Wk       �U�                    �j      �j       T�j      Wk       �T�                    �j      �j       Q�j      Wk       �Q�                      �j      �j       R�j      �j       Z�j      Wk       �R�                    �j      �j       X�j      Wk       �X�                      �j      �j       Y�j      Vk       \Vk      Wk       �U#�                  �j      �j       �                   �j      �j       �                    �j      Tk       VTk      Wk       �U#�                k      -k       Q                k      -k       v�                 -k      -k       P                  k      -k       v�                  k      -k       Q                      P      �       U�      �       S�      �       �U�                  ]      �       V                 ]      �       U                 ]      �       P                          p7      �7       U�7      d8       Sd8      n8       �U�n8      z8       Sz8      �8       �U�                          p7      �7       T�7      i8       ]i8      n8       �T�n8      8       ]8      �8       �T�                      p7      �7       Q�7      �7       ���7      �8       �Q�                          p7      �7       R�7      k8       ^k8      n8       �R�n8      �8       ^�8      �8       �R�                          p7      �7       X�7      g8       \g8      n8       �U#�n8      }8       \}8      �8       �X�                          p7      �7       Y�7      e8       Ve8      n8       �U#�n8      {8       V{8      �8       �Y�                  p7      �7       �                   p7      �7       �                  p7      �7       �                   �7      8       Pn8      y8       P                   �7      �7       t��7      �7       U                    �7      8       Pn8      y8       P                           n       Tn             u�                           =       Q=             �Q�                   K      n       Pn             u�                                      `      u       Tu      �       t��             t�             {�             T      &       t�&      :       RZ      h       Th      y       t�y      �       t��      �       t��      �       [�      �       t�                            Y      �       Q�      �       u��      �       Q�      �       u��      �       Q�             u�                               U                         n      �       u��      �       u�@��      �       u��      M       u�M      h       Xh      �       u��             u� �                               n      �       0��      �       2��      �       0��      �       0��      �       4��      �       0��      �       2��             4�                                       n      �       0��             0�             P      &       0�&      ,      & t��H$t��@$!t��8$!t��!�,      7      & r|��H$r}��@$!r~��8$!r��!�7      :       Ph      �       0��      �       P�      �       0��      �       P�             0�                      �      �       2��      �       4��      �       2��             4�                        �6      �6       U�6      7       S7      `7       �U�`7      f7       U                      �6      �6       T�6      `7       �T�`7      f7       T                       �6      
7       0�
7      7       s�7      B7       SB7      H7       P                      �6      �6       P�6      G7       ]H7      _7       ]                      �6      �6       P`7      e7       Pe7      f7       u�	                  !7      67       U                                 U             �U�                                 T             �T�                              u                               u #�                                  U             �U�                                  T             �T�                               u                                u #�                      �             U             S             �U�                 �      �       u                  �      �       u #�                      �      �       U�      �       T�      �       �U�                    �      �       T�      �       �T�                  �      �       Y                 �      �       y�                 �      �       y�                      P      m       Um      �       �U��      �       U                                 P      s       0�s      �       P�      �       0��      �       X�      �       0��      �       P�      �       X�      �       P�      �       0�                               P      P       t P      Y       t �#�Y      z       Qz      �      ' t �#�U#�t �#�����U#�*( ��      �       Q�      �       R�      �       0��      �       Q�      �       0�                    0      J       TJ      K       �T�                 0      J       0�                    �      �       P�             u                    �      �       p���             u #��                �      �       1�                �      �       U                   �      �       P�      �       u                  �      �       Q                `      �       0�                `      �       U                   c      w       Pw      �       u                  j      �       Q                      Pc      ic       Uic      �c       V�c      �c       �U�                          Pc      ic       Tic      �c       \�c      �c       �T��c      �c       \�c      �c       �T�                         Pc      ic       0�ic      sc       Psc      �c       0��c      �c       P�c      �c       0��c      �c       P                              \c      �c       S�c      �c       | �c      �c       �T�c      �c       S�c      �c       S�c      �c       | �c      �c       P                {c      �c       S                {c      �c       V                  {c      �c       0��c      �c       P                    �      �       T�              �T�                    �      �       Q�              �Q�                 �              ��                   �              T                 �              U                       �      �       u t "��      �       P�      �       u t "��              u �T"�                 �              �                   �              U                    �      �       0��             Y             R                   �      �       q 
����             Q                    �             P             r ���                                X                      �.      �.       U�.      /       �`/      t1       �U�                    �.      1       T1      t1       �T�                    �.      1       Q1      t1       �Q�                   �.      1       q��1      t1       �Q#��                                              d/      h/       0�h/      ~/       P~/      �/       p��/      �/       0��/      �/       P�/      �/       p��/      �/       0��/      �/       P�/      �/       p��/      �/       0��/      0       P0      0       p�c0      g0       0�g0      �0       P�0      �0       p��0      �0       0��0      �0       P�0      �0       p�                            d/      �/       U�/      �/       U�/      �/       U�/      Z0       Uc0      �0       U�0      t1       U                    1      1       Q1      +1       P+1      +1       p q '�                          �1      �1       U�1      t2       St2      v2       �U�v2      C3       SC3      E3       �U�                    �1      �2       Q�2      E3       �Q�                 �1      v2       T                 v2      E3       T                  �      �       P                    �+      �+       U�+      �,       X                 5,      [,       T                 p,      �,       T                        �             U      `       �U�`      f       Uf      �       �U�                      �      Z       PZ      `       �U#(`      �       P                                 U`      n       0�                      6      C       Tn      ~       T~      �       u  $ &4$p"�                    ;      C       Xn      �       X                   ;      C      	 py "1�n      �      	 py "1�                      �3      �3       U�3      ;4       �U�;4      H4       U                      �3      4       S4      G4       SG4      H4       u(                  ,4      44       P                  t      �       P                      �5      �5       U�5      �6       S�6      �6       �U�                    �5      �5       T�5      �6       �T�                      �5      �5       Q�5      %6       \%6      �6       �Q�                      �5      �5       R�5      %6       V%6      �6       �R�                    �5      �5       X�5      �6       �X�                  �5      �5       U                 �5      %6       \                    6      6       P6      %6       |�                           �      �       U�      �       �U��      �       U�      c       �U�c      o       U                      �      #       P#      )       �U#()      o       P                      �      �       R�      �       0�c      o       R                      �             T)      >       T>      Q       r  $ &4$p"�                                   U)      4       U4      Q      	 pz "@�                               	 py "1�)      Q      	 py "1�                          P3      g3       Ug3      �3       �U��3      �3       U�3      �3       �U��3      �3       U                            U3      �3       S�3      �3       S�3      �3       u(�3      �3       S�3      �3       S�3      �3       u(                  �3      �3       P                          �[      �[       U�[      �[       S�[      �[       �U��[      �[       S�[      �[       �U�                          �[      �[       T�[      �[       V�[      �[       �T��[      �[       V�[      �[       �T�                          �[      �[       Q�[      �[       \�[      �[       �Q��[      �[       \�[      �[       �Q�                    �[      �[       P�[      �[       �\                  �[      �[       1�                    �[      �[       U�[      �[       S                    P      �       U�      �       �U�                    P      �       T�      �       �T�                      P      �       Q�      �       \�      �       �Q�                    P      �       R�      �       �R�                      \      s       Vs      z       u(z      �       V                  �      �       ]                   �      �       P�      �       S                      P4      �4       U�4      n5       Sn5      t5       �U�                    P4      �4       T�4      t5       �T�                      P4      �4       Q�4      �4       ]�4      t5       �Q�                      P4      �4       R�4      �4       V�4      t5       �R�                    P4      �4       X�4      t5       �X�                  �4      �4       U                    P#      x#       Ux#      y#       �U�                      P#      [#       T[#      x#       Zx#      y#       �T�                      P#      e#       Qe#      x#       [x#      y#       �Q�                      P#      e#       Re#      x#       Xx#      y#       �R�                 P#      f#       U                                @*      �*       U�*      2+       ^2+      5+       �U�5+      B+       UB+      M+       ^M+      Z+       UZ+      x+       ^x+      �+       U                    @*      _*       T_*      �+       ��                        @*      c*       Qc*      .+       \.+      5+       �Q�5+      �+       \                 @*      d*       U                   k*      #+       \5+      �+       \                   k*      #+       ��5+      �+       ��                           k*      �*       ]�*      �*       T�*      #+       ]5+      Z+       ]Z+      f+       Tf+      �+       ]                             k*      �*       U�*      #+       ^5+      B+       UB+      M+       ^M+      Z+       UZ+      x+       ^x+      �+       U                  d+      f+       S                              p*      �*       0��*      #+       _5+      B+       0�B+      M+       _M+      Z+       0�Z+      v+       _v+      x+       	��x+      �+       0�                        |*      �*       P5+      B+       PM+      Z+       Px+      �+       P                   |*       +       0�5+      �+       0�                     �*      	+       SB+      K+       Sf+      x+       S                    �+      �+       U�+      �+       �U�                      �+      �+       T�+      �+       Y�+      �+       �T�                 �+      �+       U                                @
      �
       U�
      �
       Y�
      �
       �U��
      �
       U�
      Y       YY             U      �       Y�      �       U�      �       Y                    @
      R
       TR
      �       [                            @
      Y
       QY
      �
       V�
      �
       �Q��
      �
       V�
      Y       �Q�Y      c       Vc      �       �Q�                                @
      Y
       RY
      �
       S�
      �
       �R��
      Q       SQ      Y       �R�Y      �       S�      �       �R��      �       S                         _
      �
       Z�
      �
       U�
      C       ZK      Y       UY      v       Z�      �       Z                 @
      Z
       U                         ~
      ~
       V~
      �
       v 1$��
      �
       V�
      C       RY      c       v 1$�c      m       Vm      v       R�      �       R                   ~
      �
       [�
      C       [Y      v       [�      �       [                          ~
      �
       R�
      �
       R�
      �
       u�
      �
       yY      f       Rf      v       u�      �       u                   ~
      �
       �  �
      C       �  Y      v       �  �      �       �                     ~
      �
       Z�
      C       ZY      v       Z�      �       Z                            ~
      �
       0��
      �
       0��
      �
       V�
      �
       U�
      $       V$      3       UY      v       0��      �       0�                      ~
      �
       0��
      �
       0��
      8       ]8      C       }�Y      v       0�                          ~
      �
       1��
      �
       1��
             P	             P             1�      ;       PY      v       1��      �       1�                        �
      �
       t ���
      �
       t ���
      �
       u ����
      ,       T                     
      1
       U1
      2
       �U�                  
      )
       U                            �(      Y)       UY)      �)       _�)      �)       �U��)       *       _ *      -*       U-*      ?*       _                            �(      V)       TV)      �)       S�)      �)       �T��)      -*       S-*      4*       �T�4*      ?*       S                            �(      Q)       QQ)      �)       V�)      �)       �Q��)       *       V *      -*       Q-*      ?*       V                            �(      L)       RL)      �)       \�)      �)       �R��)       *       \ *      -*       R-*      ?*       \                          �(      ])       X])      �)       �X��)       *       �X� *      -*       X-*      ?*       �X�                      �)      �)       ��y��)      �)       S-*      4*       S                           �(      �)       0��)      �)       P�)      �)       0��)      �)       P�)      4*       0�4*      ?*       ��                      |)      �)       ^*       *       ^-*      4*       ^                      �)      �)       ]*       *       ]-*      4*       ]                    �#      �#       U�#      �(       ��~                              �#      �#       T�#      �#       S�#      �'       ��~�'      �'       S�'      &(       ��~&(      =(       S=(      �(       ��~                    �#      �#       Q�#      �(       ��~                        �#      �#       R�#      r$       ]r$      w$       �R�w$      �(       ]                    �#      �#       X�#      �(       �X�                    �#      �#       ^�'      �'       ^&(      �(       ^�(      �(       ~�                                      �#      �#       1�($      Y$       ��~���~�"| �w$      %%       ��~���~�"| �%%      �%       ��~���~�"��~���%      &       ��~���~�"| �&      &       |  ��~�"��~�"�&      ,&       ��~���~�"| �,&      �'       ��~���~�"| ��'      �'       ]�'      &(       ��~���~�"| �&(      �(       1��(      �(       ��~���~�"| �                                   �#      �#       0�($      Y$       \w$      %%       \%%      �%       ��~�%      &       \&      �'       \�'      �'       0��'      �'       1��'      &(       \&(      �(       0��(      �(       1��(      �(       \                 Y$      e$       3�                                 �#      �#       R($      Y$       ��~w$      �%       ��~�%      &       7�&      �'       ��~�'      &(       ��~&(      Z(       RZ(      �(       ��~�(      �(       8��(      �(       ��~                  H(      �(       \                  L(      �(       V                            A$      Y$       Sw$      �$       S�%      &       S,&      �'       S�'      &(       S�(      �(       S                       :&      _&       P�&      �&       P�&      �&       P�'      �'       P                               A$      Y$       0�w$      &       0�,&      M'       0�M'      Q'       PQ'      h'       Ru'      �'       0��'      &(       0��(      �(       0�                    �&      -'       ��~# -'      :'       ��~�'      �'       R                   '      u'       V�'      �'       V                 �%      &       S                  �%      �%       P                      �$      �$       P�$      �%       ��~�(      �(       ��~                       �$      �$       0��$      �$       P�$      �%       V�%      �%       0��(      �(       V�(      �(       0�                    �$      �$       P�(      �(       P                        �$      ,%       0�,%      3%       |�3%      ~%       \~%      �%       |�                    ,%      3%       S<%      �%       S                    _&      �&       U�'      &(       U�(      �(       U                     e&      �&       Q�'      &(       Q�(      �(       Q                     e&      �&       0��'      (       0�(      &(       1��(      �(       0�                              �!      V"       UV"      #       ��#      #       U#      #       ��#      '#       U'#      H#       ��H#      M#       U                        �!      Q"       TQ"      �"       S�"      #       �T�#      M#       S                              �!      V"       QV"      #       ��#      #       Q#      #       ��#      '#       Q'#      H#       ��H#      M#       Q                                �!      V"       RV"      �"       ]�"      #       �R�#      #       R#      #       ]#      '#       R'#      H#       ]H#      M#       R                    �!      	"       X	"      M#       ��                  4#      6#       _                                       "      V"       0�V"      }"       X}"      �"       ^�"      �"       X�"      #       X#      #       0�#      #       X#      '#       0�'#      6#       X6#      F#       ^F#      H#       	��H#      M#       0�                       *"      V"       P#      #       P#      '#       PH#      M#       P                   *"      �"       0�#      M#       0�                     i"      �"       _#      #       _6#      H#       _                             	      H	       UH	      X	       \X	      _	       �U�_	      
       \
      
       �U�
      
       \                             	      D	       TD	      \	       ^\	      _	       �T�_	      

       ^

      
       �T�
      
       ^                       	      H	       QH	      U	       SU	      
       �Q�                             	      H	       RH	      V	       VV	      _	       �R�_	      
       V
      
       �R�
      
       V                      i	      
       ]
      
       �U
      
       ]                      n	      r	       Pr	      �	       |�	      
       ��~                     n	      �	       ^�	      �	       S
      
       ^                      v	      
       _
      
       �Q����33$�T"�
      
       _                        P      �       U�      �       S�      �       �U��      	       S                        P      z       Tz      �       V�      �       �T��      	       V                  �      	       Q                       �      �       \�      �       \�      �       T�      	       \                     �      �       1��      �       ]�      �       }��      	       ]                 v             U                 �      �       S                 �      �       S                                  %       U%      4       V4      5       �U�5      J       VJ      K       �U�K      ?       V                         -      3       S3      4       v 4      5       �U5      =       SK      ?       S                                   -             0�      K       PK      �       0��      �       P�      �       0��      �       P�             0�             P      (       0�(      -       3�-      ?       0�                            �             U      �       S�      �       �U��      �       S�              �U�              S                          �             T      �       Z�      �       �T��              Z              T                  �              Q                           �             0�      R       [R      V       {�V      �       [�      �       [�      �       {��      �       [�             0�                                 �      !       0�!      =       P=      l       0�l      �       P�      �       0��      �       P�      �       0��              P              0�                  �      �       Q                    p      }       U}      �       Y                      p      �       T�      �       X�      �       T                  �      �       Q                   w      �       0��      �       P                          �      �       R�      �       Q�      �       R�      ^       Q^      h       R                         �      �       0��      �       Y�      P       YP      T       y�T      ^       Y^      h       0�                     �      �       3��      �       P�      h       3�                        �             0�             R             r�      7       R                         �      �       r �      �       r �             r              q7      ^       r                           K       Pf      r       P                    D      j       Pj      o       p�                      �             U      D       SD      F       �U�                 �      �       u8                                 C       UC      S       SS      \       �U�\      �       S�      �       �U�                        "       u8                    +      [       \\      �       \�      �       0�                 o      �       \                 o      �       S                  �      �       T                 �      �       P                 �      �       R                            @      g       Ug      �       S�      �       �U��             S             �U�      )       S                      @      O       TO      �       \�      )       �T�                            @      d       Qd      �       V�      �       �Q��             V             �Q�      )       V                                          �      .       U.      7       X7      n       ��n      *       �U�*      M       UM      d       �U�d      �       U�      �       ���      '        �U�'       5        U5       �!       �U��!      �!       ���!      �!       U                                                �      &       T&      I       ^I      n       Tn      *       ^*      E       TE      M       ^M      d       �T�d      �       ^�      �       T�      �       ^�              T       n!       ^n!      u!       Tu!      �!       ^�!      �!       T�!      �!       ^                                �             Q      n       ]v      �       ]�      �       }��      M       ]d      �        ]�       �        }��       @!       ]@!      D!       }�D!      �!       ]�!      �!       } p "��!      �!       ]                      3      7       u �      �       u �              ��n!      �!       ��                                                         �      @       0�@      e       Pe      n       S�      �       S�             R             S      *       R*      M       0�d      �       0��      �       P�      �       S       "        S"       '        p �'       5        0�!      (!       S(!      :!       R:!      V!       SV!      n!       R�!      �!       S�!      �!       S�!      �!       0�                                           �      v       0�v      %       V(      *       V*      M       0�d      �       0��              V'       �        0��       e!       Vl!      �!       V�!      �!       P�!      �!       V�!      �!       0��!      �!       V�!      �!       0�                                           �      v       1�v      �       \�      �       P�      *       \*      M       1�d      �       1��      '        \'       �        1��       !       \!      4!       \7!      �!       \�!      �!       1��!      �!       \�!      �!       1�                           �      &       0�*      *       0�*      M      	 p �-)�d      n      	 p �-)�n      �       _'       *        _�!      �!       _                                       �      `       0�`      n       Y�      *       Y*      M       0�d      �       0��      �       Y               1�'       5        0�!      n!       Y�!      �!       Y�!      �!       Y�!      �!       0�                               �      �       0��      �       T*      M       0�d              0�'       !       0�!      &!       Tn!      �!       0��!      �!       0�                      �       �        Q�       !       Q�!      �!       Q                    �              Pn!      �!       P                          �      �       U�      �       \�      �       �U��             \             �U�                    �      �       S�      �       S�             S                    �      �       P�             P                            0       {        Q{       �        [�       �        Q�       �        [�       �        Q�       �       [                          3       ]        X]       �        Y�       �        X�       �        Y�       �        X�       �       Y                           3       �        0��       �        Z�       �        0��       f       Zi      k       Zk      �       0�                         3       Y        0�Y       y       	 s �-)�y       �        x �-)��       �        0��       �        S�       �        0��       �       S                         3       �        0��       �        \�       �        0��       k       \k      �       0�                      ~       �        P�       �        P�       �       P                   �       �        Q�       �       Q                      �              R             XB      k       R                           d      Sd       USd      0e       S0e      Ee       �U�Ee      h       Sh      h       Uh      �j       S                  d      "d       u                     5d      <e       VEe      �j       V                                   5d      �d       ���d      �d       \�d      0e       \Me      �e       \�e      �f       \�f      �f       ���f      _g       \_g      dg       7�h      h       ���h      �h       0��h      �h       \                    Td      xd       P�d      �d       P                    5d      �d       0�Kg      dg       ��~h      h       0�                 �e      (f       0�                �e      (f       �t.                  �e      (f       S                 (f      �f       A�                      *f      >f       z�>f      Cf       ZCf      Jf       z�                 (f      �f       S                      :f      Cf       PJf      \f       P|f      �f       P                  ]f      of       P                   �d      �d       ���h      �h       0�sj      xj       0�                  �e      �e       P                    �d      �d       Sh      �h       S�h      yi       S                       �d      �d       P�d      �d       ��~h      �h       ��~�h      yi       ��~                    �h      i       Ri      Di       ��~                  Eh      Zh       P                          �d      �d       	��h      8h       	��8h      �h       \�h      �h       |��h      Di       \Di      yi       	��                    h      2h       PDi      \i       P                  �d      �d       �0  h      h       �0                    �d      �d       Sh      h       S                 Di      \i       s                     dg      h       Syi      sj       Sxj      �j       S                       �g      �g       P�g      h       ��~yi      sj       ��~xj      �j       ��~                      �i      j       Rj      Lj       ��~xj      �j       ��~                    �g      �g       P�g      h       P                      �g      �g       	��yi      �i       	���i      Gj       \xj      �j       \                    �g      �g       Pyi      �i       P                �g      �g       �2                  �g      �g       S                            �g      �g       P�g      �g       X�i      j       Xj      Lj       ��~Lj      rj       Xxj      �j       ��~                      j      @j       Pxj      zj       P|j      �j       P                 yi      �i       s                 (g      Kg       �+.                  (g      Kg       S                         )        U                         )        T                         )        R                           %        Q%       )        t �����@$t�����!�                      �      �       U�      �       S�      �       �U�                 �      �       u                       �      �       U�      1       S1      7       �U�                      �      �       T�      2       V2      7       �T�                      �      �       Q�      4       \4      7       �Q�                      �      �       R�      6       ]6      7       �R�                     �      �       0��      �       P�      7       Q                      �8      �8       U�8      9       \9      9       �U�                      �8      �8       T�8      9       ]9      9       �T�                         �8      �8       0��8      �8       p��8      �8       P�8      �8       ^�8      	9       P                      �:      �:       U�:      ;       ^;      ;       �U�;      �;       ^                  �:      �:       T�:      �;       �T�                      �:      �:       Q�:      ;       ];      ;       �Q�;      �;       ]                            �:      �:       \�:      �:       U�:      ;       \;      :;       \:;      >;       U>;      �;       \                     �:      ;       V;      ;       P;      �;       V                                        �:      �:       R�:      �:       �;      ;       R;      :;       �I;      i;       Ri;      n;       �n;      ;       R;      �;       ��;      �;       R�;      �;       ���;      �;       R�;      �;       ��;      �;       R                  �:      �:       sx�,;      :;       sx�                 �;      �;       U                    :      ":       U":      x:       T                    4:      d:       Pi:      x:       P                    S:      d:       Ri:      x:       R                 :      ":       U                        �9      �9       U�9      �9       T�9      �9       U�9      :       T                    �9      �9       P�9      :       P                      �9      �9       Q�9      �9       q����9      :       Q                 �9      �9       U                  d      �       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                  �      �       X                  �      �       U                 �      �       P                                 '       U'      .       U.      3       P3      5       u p '�5      6       P                  S9      ]9       P                  <      �<       U                      $<      9<       QH<      V<       0��<      �<       Q                      o<      |<       R�<      �<       R�<      �<       q  $ &4$u"�                      t<      |<       T�<      �<       T�<      �<      	 uz "@�                   t<      |<      	 uy "1��<      �<      	 uy "1�                    >      2>       U2>      ?       [                      >      5>       T5>      �>       U�>      ?       �T�                    >      9>       X9>      ?       �X�                      p>      u>       S��u>      �>       S�P��>      �>       �P�                   >      9>       X9>      G>       �X�                  >      >       uȑ                   9>      G>       XG>      G>      
 p x "#���                  9>      G>       x ?&�G>      G>       P                G>      S>       Y                G>      S>       {̑                  G>      S>       QS>      S>      
 q r "#���                  G>      S>       q ?&�S>      S>       R                u>      �>       r�                    �>      �>       T�>      �>      
 t u "#���                  �>      �>       t ?&��>      �>       U                �>      �>       P                �>      �>       r�                   �>      �>       Q�>      �>      
 q x "#���                  �>      �>       q ?&��>      �>       X                  �>      �>       S�>      �>      
 q s "#���                  �>      �>       s ?&��>      �>       Q                 �>      �>       P                  �>      �>       R�>      �>      
 r t "#���                  �>      �>       r ?&��>      �>       T                  I      $I       U�                  I      $I       P                 0I      FI       �̎  �                  4I      EI       ��                  4I      EI       P                   J      8J       U                  $J      8J       Q                      @J      |J       T|J      }J       �T�}J      �J       T                 DJ      �J       U                  }J      �J       T                  }J      �J       U                  �J      �J       ��                  �J      �J       Q                      �J      �J       T�J      �J       �T��J      �J       T                 �J      �J       U                  �J      �J       T                  �J      �J       U                  �J      �J       P                        �J      K       UK      4K       S4K      6K       �U�6K      AK       U                       �J      K       UK      4K       S4K      6K       �U�6K      AK       U                      �J      K       UK      4K       S4K      6K       �U�                  K      5K       V                              PK      �K       U�K      �L       V�L      �L       �U��L      �L       V�L      M       UM      M       VM      M       �U�                            PK      �K       T�K      �L       \�L      �L       �T��L      M       TM      M       \M      M       �T�                              PK      �K       Q�K      �L       _�L      �L       �Q��L      �L       _�L      M       QM      M       _M      M       �Q�                              PK      �K       R�K      %L       ��%L      �L       ]�L      �L       �R��L      �L       ���L      M       RM      M       ��                            �K      �K       R�K      %L       ��%L      �L       ]�L      �L       ���L      �L       RM      M       ��                          �K      �K       Q�K      �L       _�L      �L       _M      M       _M      M       �Q�                        �K      �L       \�L      �L       \M      M       \M      M       �T�                  �L      �L       0�M      M       P                       �K      �K       S�K      �K      
 s 2%s "#��K      �L       S�L      �L       SM      M       S                           �K      �K        ~ ��K      �K       Y�K      *L       ���L      �L       ���L      �L       YM      M       ��                   �K      �L       S�L      �L       SM      M       S                   �K      �L       V�L      �L       VM      M       V                      �K      �K       P�K      �L       ���L      �L       ��M      M       ��                    �K      }L       ^}L      �L       0��L      �L       ^M      M       ^                 /L      xL       ^                 /L      xL       V                  KL      lL       U                 KL      xL       P                   KL      oL       ToL      xL       v � $ &3$v("�                           M      \M       Q\M      �M       \�M      �M       �Q��M      �M       Q�M      �M       \                           M      \M       R\M      �M       ]�M      �M       �R��M      �M       R�M      �M       ]                       M      pM       XpM      �M       �X��M      �M       X                         M      >M       Y>M      �M       _�M      �M       �Y��M      �M       _                     kM      �M       S�M      �M       s~��M      �M       S                      FM      pM       YpM      �M       ^�M      �M       Y                    PM      pM       S�M      �M       S                   PM      �M       V�M      �M       V                          M      \M       Q\M      �M       \�M      �M       �Q��M      �M       Q�M      �M       \                          M      \M       Q\M      �M       \�M      �M       �Q��M      �M       Q�M      �M       \                 �M      �M       \                 �M      �M       Q                      `S      �S       T�S      �S       �T��S      �S       T                          `S      �S       Q�S      �S       S�S      �S       �Q��S      �S       Q�S      �S       S                     `S      �S       0��S      �S       P�S      �S       0�                   `S      |S       U�S      �S       U                   `S      |S       u���S      �S       u��                      sS      S       P�S      �S       P�S      �S       u�#h                �S      �S       w                 �S      �S      	 q  $ &�                        �S      �S       U�S      T       ST      T       �U�T      9T       S                    @[      D[       UD[      g[       �U�                    @[      f[       Tf[      g[       �T�                      p[      u[       Uu[      v[       �U�v[      �[       U                      p[      u[       Tu[      v[       �T�v[      �[       T                            �[      \       U\      !\       S!\      %\       �U�%\      2\       S2\      9\       U9\      :\       �U�                            �[      \       T\      "\       V"\      %\       �T�%\      3\       V3\      9\       T9\      :\       �T�                            �[      \       Q\      $\       \$\      %\       �Q�%\      5\       \5\      9\       Q9\      :\       �Q�                          \      $\       \$\      %\       �Q�%\      5\       \5\      9\       Q9\      :\       �Q�                          \      "\       V"\      %\       �T�%\      3\       V3\      9\       T9\      :\       �T�                          \      !\       S!\      %\       �U�%\      2\       S2\      9\       U9\      :\       �U�                  \      9\       P                    @\      f\       Tf\      g\       �T�                    p\      �\       U�\      �\       �U�                    p\      �\       T�\      �\       �T�                    p\      �\       Q�\      �\       �Q�                   p\      �\       Q�\      �\       �Q�                   p\      �\       T�\      �\       �T�                   p\      �\       U�\      �\       �U�                  t\      �\       R                  �\      �\       U                 �\      �\       P                          �\      �\       U�\      A]       SA]      G]       �U�G]      v]       Sv]      �]       U                            �\      �\       T�\      D]       \D]      G]       �T�G]      b]       Tb]      v]       \v]      �]       T                            �\      �\       Q�\      F]       ]F]      G]       �Q�G]      W]       QW]      v]       ]v]      �]       Q                     ]      <]       0�U]      W]       0��]      �]       3�                        �\      �\       U�\      ]       SG]      U]       SW]      v]       Sv]      �]       U                      �\      ]       VG]      U]       VW]      �]       V�]      �]       u(                  l]      v]       P                 ]      <]       ]                 ]      <]       \                 ]      <]       S                    "]      7]       P7]      <]       �L                 ]      <]       S                 ]      "]       1�                    �^      �^       U�^      _       �U�                    �^      _       T_      _       �T�                      _      _       U_      _       �U�_      #_       U                      _      _       T_      _       �T�_      #_       T                      0_      F_       UF_      �_       \�_      �_       �U�                      0_      >_       T>_      h_       Vh_      �_       �T�                      0_      F_       QF_      o_       So_      �_       �Q�                  G_      �_       P                  5_      G_       1�                    5_      F_       UF_      G_       \                   K_      o_       So_      �_       �Q�                   K_      h_       Vh_      �_       �T�                 K_      �_       \                K_      �_       1�                  K_      o_       So_      �_       �Q�                  K_      h_       Vh_      �_       �T�                K_      �_       \                 Y_      �_       T                  w_      �_       U                  z_      �_       R                            �_      �_       U�_      �_       S�_      �_       �U��_      �_       S�_      �_       U�_      �_       �U�                            �_      �_       T�_      �_       V�_      �_       �T��_      �_       V�_      �_       T�_      �_       �T�                            �_      �_       Q�_      �_       \�_      �_       �Q��_      �_       \�_      �_       Q�_      �_       �Q�                          �_      �_       \�_      �_       �Q��_      �_       \�_      �_       Q�_      �_       �Q�                          �_      �_       V�_      �_       �T��_      �_       V�_      �_       T�_      �_       �T�                          �_      �_       S�_      �_       �U��_      �_       S�_      �_       U�_      �_       �U�                  �_      �_       P                        �_      `       U`      2`       �U�2`      I`       UI`      �b       S                        �_      `       T`      2`       �T�2`      K`       TK`      �b       V                        �_      `       Q`      2`       �Q�2`      ;`       Q;`      �b       �Q�                          �_      `       R`      1`       _1`      2`       �R�2`      >`       R>`      �b       _                          �_      `       X`      +`       \+`      2`       �X�2`      O`       XO`      �b       \                        �_      `       Y`      2`       �Y�2`      Z`       YZ`      �b       �Y�                            r`      a       ]a      [a      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&�[a      �a       ]�a      �a      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&��a      ub       ]ub      �b      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&�                        �`      �`       Ra      �a       R�a      �a       Rb      "b       R                                    ~`      �`      	 >u r ��`      �`      + >u O} (  / 0@K$(	 1$#/��O'��`      a      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'�a      [a       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'�[a      ea      	 >u r �ea      oa      + >r Ov (  / 0@K$(	 1$#/��O'�oa      �a      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'��a      �a       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'��a      ub      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'�ub      �b       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'�                            K`      �`       T[a      �a       T�a      �a       p �a      �a       Tb      /b       T/b      Jb       �                             O`      �`       X[a      �a       X�a      �a       p�a      �a       Xb      Jb       XJb      �b       ��                         O`      �`       p�`      �`       � #[a      �a       p�a      �a       � #b      Jb       � #                         O`      �`       p�`      �`       � #[a      �a       p�a      �a       � #b      Jb       � #                         O`      �`       p�`      �`       � #[a      �a       p�a      �a       � #b      Jb       � #                         O`      �`       p�`      �`       � #[a      �a       p�a      �a       � #b      Jb       � #                          Z`      �`       Y[a      �a       Y�a      �a       Yb      Jb       YJb      �b       ��                         Z`      �`       p�`      �`       � #[a      �a       p�a      �a       � #b      Jb       � #                     Z`      a`       Qa`      i`      
 q r "#���i`      r`       ]                   Z`      a`       q ?&�a`      r`       R                    �`      �`       P�`      Aa       ��                    �`      a       } p �a      $a      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                 [a      a       V                 [a      a       ]                      ia      sa       Qsa      {a      
 q r "#���{a      a       R                     ia      sa       q ?&�sa      {a       R{a      a       q ?&�                    �a      �a       Y�a      �a       w                     �a      �a       } p ��a      �a      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                    Fb      Jb       RJb      �b       ��                 Fb      Jb       � #�����                    Kb      ub       } p �ub      �b      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                      �b      �b       U�b      �b       S�b      -c       �U�                    �b      �b       T�b      -c       �T�                 �b      �b       t ����1$u"�
���                       �b      �b       0��b      �b       s��b      c       Sc      #c       s�                      �b      �b       P�b      c       ^c      ,c       ^                 �b      c       U                      0c      <c       U<c      =c       �U�=c      Cc       U                      0c      <c       T<c      =c       �T�=c      Cc       T                    �c      �c       U�c      d       �U�                    �c      �c       T�c      d       Y                  �c      d       X                         �c      �c       0��c      �c       P�c      �c       0��c      �c       0��c      d       P                        `k      �k       U�k      �k       X�k      �k       �U��k      �k       U                        `k      �k       T�k      �k       �T��k      �k       T�k      �k       �T�                      `k      �k       Q�k      �k       �Q��k      �k       Q                  `k      k       Q�k      �k       Q                  `k      k       U�k      �k       U                  �k      �k       Q                  �k      �k       U                  �k      �k       P                    �k      �k       0��k      �k       R                   �k      �k       T�k      �k       T                  �l      �l       ��                  �l      �l       Q                  �l      �l       U                  �l      �l       Q                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  �      �       U                      �       �        U�       y       �U�y      �       U                       �              0�      m       Pt      y       Py      �       0�                          �       �        p��       F       XF      _       0�_      y       Xy      {       p�{      �       t �#�                     �              0�      m       Uy      �       0�                        �              S      9       Y=      B       QB      k       Yy      �       S                        �              Q#      &       R&      Q       Qc      m       Q                      �               Z#      Q       ZQ      c       Qc      t       Z                                 R1      m       R                      @       _        U_       �        �U��       �        U                  D       �        Q                      R       U        q p "�U       �        R�       �        R                  _       �        U                           @       j        0�j       �        X�       �        U�       �        X�       �        U�       �        0�                    j       �        P�       �        P                    �      �       U�      &       ��~                          �      �       T�             S      �       ��~�      �       S�      &       ��~                        �      �       Q�             \      %       �Q�%      &       \                        �      �       R�             w       %       ��~%      &       w                     �      �       X�      &       ��~                        �      �       Y�              ]       %       �Y�%      &       ]                                     0�      �       S%      �       S�      �       0�                   �             V�      &       V                                �       V�      �       vx��      �       V%      �       V�      �       vx��      �       V�      �       vx��      �       V                    q      �       PT      �       P                      .      :       P:      �       _%      �       _                        :      H       ~�H      _       ^_      c       ~�%      O       ^                       i      w       q�w      {       Q{             q��      �       Q                                    U       7        �U�                                   U       7        �U�                         7        T                         7        U                                         P       !       	 q ����!       ,        P,       3       	 q ����3       7        t �����                          p      �       U�      �       �U��      �       U�      �       �U��      �       U                   :      @       4�@      n       u r #�                     6      @       0�@      j       Pp      �       P                      :      n       Rn      p       r�p      y       R                     @      n       r n      y       ry      �       X                    H      M       TM      Q       x��Q      �       T                         �      �       6��             T             t�             T$      /       T                       �      �       0��             P      !       P$      /       P                        �             X             x�      !       X$      /       X                     �             x              x$      /       x                       �      �       R�      �       y���      !       R$      /       R                    w      �       U�      �       T                    �      �       0��      �       T                 �      �       T                   �      �       U�      �       �U�                 �      �       0�                 �      �      
 �I     �                 �      �       T                   �      �       U�      �       �U�                 �      �       0�                 �      �      
 �I     �                          �      �       U�      l       u�p      t       u�t      y       Uy      �       u��      �       U�      n       u�                            �      l       [p      y       [�      �       R�      �       [�      g       Rg      n       [                              �      l       4�p      y       4��      �       4��      �       z����             z~���             x �I     "���      0       z���g      n       4�                         �      �       0��      l       Yp      y       Y�      �       Yg      n       Y                           �      �       4��      '       S'      l       R�      �       R�      �       Sg      n       S                                     �      l      
 �I     �p      t      
 �I     �t      �       Z�      �       z��      �       p��      �       Z�      �      
 �I     ��      �       Z�      �       z��      �       z~��      �       P�      g       Qg      n      
 �I     �                          �      6       R6      g       Qg      l       R�      �       Qg      n       R                                     �             r 1$ $ &�I     "�      6       Z6      X       q 1$ $ &�I     "�X      l       Zp      �       Z�      �       P�      �       Z�             z}�             x �I     "�      :       Z:      I       p �I     "�I      n       Z                                  '      	 x ��'      ^      F s y "1&1$ $ &�I     "�8$
��
��#%!
���I     "���^      g       Pg      l      F s y "1&1$ $ &�I     "�8$
��
��#%!
���I     "����      �       Pg      n      	 x ��                  �      0       q ��8$p��!�0      W       q ��8$q��!�                            :       Z:      I       p �I     "�I      g       Z                    �      �       U�      �       �U�                  �      �       P                            �       �        U�       ^       S^      `       �U�`      r       Sr      t       �U�t      ~       U                        �       �        T�       	       U	      t       �T�t      ~       T                                   P      _       V`      s       V                          0       O        UO       f        �U�f       u        Uu       |        �U�|       �        U                          0       O        TO       f        �T�f       y        Ty       |        �T�|       �        T                              0       O        QO       _        V_       e        Ue       f        �Q�f       r        Qr       |        V|       �        Q                              0       O        RO       Y        SY       e        Qe       f        �R�f       y        Ry       |        S|       �        R                      I       a        \a       e        Rf       |        \                                      U       %        S%       &        �U�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                    �       �        Q�       �        �Q�                    �       �        R�       �        �R�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                      �      �       U�      �       �U��             U                        �      �       T�      �       S�      �       �T��             T                   �      �       u �      �       U                      0      k       Uk      �       S�      �       �U�                  �      �       P                  h      �       W                            0      �       U�      �       �U��      �       U�      �       �U��      �       U�      +       �U�                            0      �       T�      �       S�      �       �T��      �       S�      �       T�      +       S                            0      f       Qf      �       V�      �       �Q��      �       V�      �       Q�      +       V                                0      �       R�      �       �R��      	       R	      �       �R��      �       R�      �       �R��      �       R�      +       �R�                     i      �       u �      �       u �      �       �U                          �      �       \L      �       \�      n       \x      �       \�      +       \                             �      �       v�      �       XL      �       X�      }       X�      n       Xx      �       X�      +       X                       �      �       0��             Q�      �       Q�      �       r q ��      �       P                         �      �       v�      �       p ��      �       q ��      �       } ��             v���      �       v��                      �      �      	 q ������            	 z ������      �      	 z �����                       �      X       [X      c       {�c      n       [x      �       [�             [                       �      �       \�      �       T�      @       t�@      L       T�             \                          �      �       X�      �       Q�      @       qx�@      H       Q�      �       P�      �       p��      �       P�             X                             �      �       q 3%��      �       PL      O       q 7�O      Q       Qx      �       Q�             P             q 3%�                    �      0       P0      3       U                   �      �       R�      �       R                  \      �       ^                   `      �       ]�      �       }��      �       ]                       �      <       [<      G       {�G      N       [�      �       [             [                       �      �       \�      �       U�      !       u�!      ,       U             \                          �      �       X�      �       Q�      !       q|�!      ,       Q�      �       Y�      �       y��      �       Y             X                             �      �       p 2%��      �       Q�      �       p 2%�,      /       p 3�/      5       P�      �       P             Q                    �             P             T                   �      �       Q�      �       Q                     [      �       U�      �       u��      �       U      +       U                         `      x       \x      �       | p "#��      �       | p "��      �       | p "#��      �       | q "�      +       \                         `      x       Xx      �      
 p 1$x "#��      �       p 1$x "��      �      
 p 1$x "#��      �      
 q1$x "#�      +       X                        c      g       p 1%�g      x       Q      #       Q#      +       p 1%�                      �      �       r ���      �       q ���      �       | p "���                         �       Z�      �       z��      �       Z                           '       \'      3      
 t 2$| "#�3      �       t 2$| "��      �      
 t 2$| "#�                           '       X'      3       x t "#�3      �       x t "��      �       x t "#�                        '       P                 3      �       t 2$| "�                    >      �       U�      �       [                                T      X        r r 
|p p 
�"q q 
m6"@%�X      \      4 t 2$| "��t 2$| "��
|p p 
�"q q 
m6"@%�\      `      1 t 2$| "��t 2$| "��
|p 
�"q q 
m6"@%�`      g      I t 2$| "��t 2$| "��
|p 
�"t 2$| "#��t 2$| "#��
m6"@%�g      n      . t 2$| "#��t 2$| "#��
m6p 
�"r "@%�n      u      I t 2$| "#��t 2$| "#��
m6t 2$| "#��t 2$| "#��
�"r "@%�u      }      * t 2$| "#��t 2$| "#��
�q "r "@%�}      �      I t 2$| "#��t 2$| "#��
m6t 2$| "#��t 2$| "#��
�"r "@%�                                                  �       U�      u	       �U�u	      �	       U�	      
       V
      
       U
      W
       VW
      �
       �U��
      �
       V�
      �
       U�
      :       V:      p       Up      �       V�      �       U�      �       V�      ]       �U�                                                �       T�      u	       �T�u	      
       S
      
       T
      �
       S�
      �
       w �
      t       St      �       �T��      �       w �      �       �T��             S      U       ��U      ]       S                                  W       QW      �       �Q��      �       Q�      
       �Q�
      
       Q
      ]       �Q�                                  \       R\      �       �R��      �       R�      
       �R�
      
       R
      ]       �R�                            �      f	       0��	      �	       P�      �       B��      �       0��      �       0��      �       0�                      �      f	       V�      �       V�      �       V                         �      �       T	      	       0�	      &	      	 t q "v �&	      *	       q t "v #�      +       1�+      �       T                         �      �       X�      �       1��      ;	       U�             ~�      �       X                           �      W	       ��~�#��      �       s�      �       ^�      �       ��~�#��      �       s�      �       ^                       �      B	       w G	      W	       U�      �       0��      �       w                                z      �       S�      �       ��~�      
       ��~
      
       S
      �
       ��~�
      �
       P�
      E       ��~E      ]       ��~                                        ~      �       R�      u	       ��~u	      ~	       R~	      
       ��~
      
       R
      �
       ��~�
      �
       R�
      :       ��~:      E       RE      �       ��~�      �       R�      �       R�      ]       ��~                   u	      �	       ����	      �	       Q                     �      �       \      +       u +      �       \                  	      ;	       v t �                                �	      
       ��~
      �
       ��~	      :       ��~b      �       ��~�      �       ��~�      �       ��~�      �       ��~�      ]       ��~                                �	      
       ��~
      �
       ��~	      :       ��~b      �       ��~�      �       ��~�      �       ��~�      �       ��~�      ]       ��~                                          �	      
       S
      �
       S�
      �
       w �
      �
       S	      :       Sb      �       S�      t       St      �       �T��      �       w �      �       �T��             S      U       ��U      ]       S                                      �	      �	       P�	      
       ��~
      �
       ��~	             P      :       ��~b      g       Pg      �       ��~�      �       ��~�      �       ��~�      �       ��~�      ]       ��~                              �	      
       \
      �
       \      :       \p      �       \�      e       \�      �       \�      ]       \                                        *
      0
       ^0
      j
       _�
      �
       ^�
      �
       _/      5       ^5      :       _~      �       _�      �       _�      �       ^�      �       ^�      �       _�      ]       _                    
      0
       4��
      �
       2�      :       1�p      �       8�                         �	      
       ]
      p
       ]�
      �
       ]	      :       ]b      �       ]�      �       ]                            �	      
       P
      �
       P�
      �
       P      :       Pm      �       P�      �       P                                 �	      
       0�
      �
       0�	      :       0�b      �       0��      �       0��      �       P�      �       V�      �       0��      �       V�      ]       V                   G
      �
       | 3$��      �       | 3$�                    _
      x
       Rx
      |
       _                        �
      �
       _�
      �
       U�
      �
       _�      �       _                   �
      �
       ^�      �       ^                     �
      �
       R�
      �
       S�      �       S                   �
      �
       ]�      �       ]                       �
      �
       P�
      �
       v��
      �
       V�      �       V                   �
      �
       _�
      �
       U                            E       ]E      I       TJ      e       ]U      ]       ]                                 7       V7      J       ^J      S       ~ | "�S      Y       UY      _       ~ | "�_      t       ^U      ]       V                         7       s �| ����} "�U      ]       s �| ����} "�                         e        | �U      ]        | �                      �      �       s      -       ]-      1       T2      U       ]                           �      �       U�             V             P      2       S2      6       s | "�6      ?       U?      @       s | "�@      E      	 s | "~ "�                 �      �       s �| ����s"�                 �      U        | �                            0       �        U�       Y       �U�Y      �       U�      �       �U��      �       U�      !       �U�                                  0       �        T�              \      Y       �T�Y      �       T�      �       �T��      �       T�      �       \�      �       T�      !       \                                0       �        Q�              V      Y       �Q�Y      �       Q�      �       �Q��      �       V�      �       Q�      !       V                      �       �        U�      �       U�      �       U                           �       �        S�       �        s ��       �        t���      �       t���      �       |���      �       t���      �       |��                      �       	       ]�      �       ]�      !       ]                        �       X       _Y      �       _�      �       _�      !       _                        �       V       ^Y      �       ^�      �       ^�      !       ^                     �       �        P�       �        p ��       �        v���      �       v��                    �       �        Q�      �       Q                 �       �        v                           $       P$      +       VB      F       V                           7       \7      ;       T?      R       \                          ;       XB      Y       X                                ]@     �@     �@     :@     :@     l@     l@     �@     �@     �@     �@     �@     �@     �@     �@     @     @     �@     �@     t@     t@     �@                     \      b      f      h                      �      �      �      �                                                 (      ?      G      K                                    (      ?      G      K                                    (      ?      G      K                      K      O      [      [      [      n                      K      O      [      n                      w      w      w      w            �      �      �                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �                               #      ,      >      `      c      g      m      w      �      �      �                      �      �      �                   0                      �      �      �            8      B                      �      �      �      �      �      �      	      
	      	      	      !	      %	      )	      ,	                      �      �      �      �      �      �      	      
	      	      	      !	      %	                      �      �      �      �      �      �      
	      
	      	      	      	      	      ,	      4	      7	      ;	      ?	      A	                      �      �      �      �      �      �      
	      
	      	      	      	      	      ,	      4	      7	      ;	                      �      �      �      �      	       	      %	      )	      G	      V	                      �      �      �      �      	       	      %	      )	      G	      S	                      �      	      
	      	      )	      )	      4	      7	      ;	      ?	      V	      d	                      �      	      
	      	      )	      )	      4	      7	      ;	      ?	      V	      b	                      b      e      {      ~      �      �      �      �      �      �      �      �      �      �      �      �                      b      e      {      ~      �      �      �      �      �      �      �      �      �      �      �      �                      b      e      {      ~      �      �      �      �      �      �      �      �      �      �      �      �                      e      i      ~      �      �      �      �      �      �      �      �      �      �      �      �      �                      e      i      ~      �      �      �      �      �      �      �      �      �      �      �      �      �                      e      i      ~      �      �      �      �      �      �      �      �      �      �      �      �      �                      q      u      �      �      �      �      �      �      �      �      �      �      �      �                      q      u      �      �      �      �      �      �      �      �      �      �      �      �                      q      u      �      �      �      �      �      �      �      �      �      �      �      �                      v      z      �      �      �      �      �      �      �      �      �      �            $      .      6      B      F                      v      z      �      �      �      �      �      �      �      �      �      �            $      .      6      B      F                      v      z      �      �      �      �      �      �      �      �      �      �            $      .      6      B      F                      �      �      �      �      �      �      �      �      �      �      �      �      6      ;      J      R      c      g                      �      �      �      �      �      �      �      �      �      �      �      �      6      ;      J      R      c      g                      �      �      �      �      �      �      �      �      �      �      �      �      6      ;      J      R      c      g                      �      �      �      �            	                  $      (      ?      ?      ?      ?                      �      �      �      �            	                  $      (      ?      ?                      �      �      �      �      	            +      .      ;      ?      R      Z      g      k                      �      �      �      �      	            +      .      ;      ?      R      Z      g      k                      �      �      �      �      	            +      .      ;      ?      R      Z      g      k                                  ?      ?      ?      B      F      J      [      c      n      r                                  ?      B      F      J      [      c      n      r                      �      �      �      �      �      �      �      �      �      �      �      �            
                      �      �      �      �      �      �      �      �      �      �      �      �                      �      �      �      �      �      �      �      �                  
                            �      �      �      �      �      �      �      �                                        >      �      �      �      �            0                      E      g      �      �             2      �      �                      n      �      �             6      [      �      �      0      H                      �      �      [      y      �      �      �            K      p                      �            (      I                      P      P      Y      h      l      o      q      s                      a      h      l      o      q      s                      �      �      �                             �      �      �      �                                                                      <      @      H                            "      &      -                      1      <      @      H                            �      �      �                      �      �      �      �                      	      	            L      X      v      z      �      �      �                      r      v      z      �      �      �                      �      �      �      �                      7       A       E       ]       �       �                       <       A       E       ]       �       �                       <       A       J       T                       �       �       �       �                       �!      �!      �!      �!                      �"      �"      �"      �"                      $      B$      p$      �$                      F$      a$      �$      �$      �$      �$      �$      %      %      .%                      [%      �%      �%      K'      U'      )                      `&      �&      @(      p(                      �&      �&      p(      �(      �(      �(                      �&      �&      �&      '      '      '      '      '      '      '      #'      ''                      �&      �&      �&      '      '      '      '      '      '      '      #'      ''                      �&      �&      �&      '      '      '      '      '      '      '      #'      ''                      �&      �&      '      '      '      '      '      '      '      #'      ''      +'                      �&      �&      '      '      '      '      '      '      '      #'      ''      +'                      �&      �&      '      '      '      '      '      '      '      #'      ''      +'                      �'      �'      (      @(                      $)      P)      p)      p)      t)      {)                      �+      �+      �+      �+      �+      �+                      �+      �+      �+      �+                      �+      �+      �+      �+      �+      
,                      �+      �+      �+      �+      �+      ,                      ,      �,      �,      M-                      #,      U,       -      M-                      d,      �,      �,       -                      Z-      m-      r-      w-      �-      �-      �-      �-                      �/      �/      �/      �/                      �0      �0      �0      �0      �0      1      1      1      1       1      (1      C1      P1      �1                      �0      �0      �0      �0      �0      1      (1      C1      P1      g1      p1      1                      (1      ;1      P1      W1                      �1      �1      �1      �1      �1      �1      �1      �1      02      j2      p2      2                      �2      �2      �2      �2      �2      �2      �2       3      3      3                      �2      �2      �2      �2      �2      �2      �2      �2      3      3                      �2      �2      �2      �2                      +3      >3      A3      F3      J3      M3      Q3      S3                      �3      �3      �3      �3      �3      �3                      04      C4      P4      U4      Y4      \4      `4      b4                      �4      �4      �4      �4      �4      �4                      �6      �6      �6      �6      �6      �6                      �6      �6      �6      �6      �6      �6                      �6      �6      �6      7                      97      X7      Y7      `7                      J7      X7      Y7      `7                      }7      }7      �7      �7      �7      �7      �7      �7                      �7      �7      �7      �7      �7      �7                      �7      �7      �7      8      8      
8      8      8                      �7      8      8      
8      8      8                      �8      �8      �8      �8                      69      69      D9      �9      �9      �9                      O9      �9      �9      �9                      p9      t9      y9      �9                      �9      �9      �9      �9                      �;      �;      �;      �;      �;      �;      �;      e<      i<      k<      �<      H=      N=      k=                      <      #<      +<      e<      �<      H=      N=      k=                      �<      �<      �<      �<                      �<      0=      N=      k=                      �<      �<      �<      �<      �<      0=      N=      k=                      �<      �<      �<      �<                      �<      0=      g=      k=                      �<      =      g=      k=                       =      =      	=      =                      J>      e>      j>      �>      J?      V?                      �?      �?      �?      �?                      �@      �@      �@      �A      B      rD      wD      }D      �D      �D      �D      �D      �D      �D      E      .E                      �A      �A      �B      �B      �B      ]C                      �C      VD      �D      �D      E      .E                      �C      <D      @D      @D                      5E      zE      �E      �E                      �E      �E      �E      F      #F      .F      2F      GF      PF      ZF      eF      pF      sF      �F                      yG      �G       K      `K                      �G      �G       K      @K                      �G      �G      @K      `K                      �G      oH      `K      �K      �L      �L                      �G      oH      `K      �K      �L      �L                      �G      �G      �G      FH      `K      `K                      0H      4H      =H      FH                      _H      fH      fH      oH                      K      �K      �K      �K                      �L      �L      �L      �L                      �H      �H      �H      �H      �H      �H                      wI      J      )J      -J                      �I      J      )J      -J                      cJ      K      �K      L                      L      �L      �L      �L                      AM       N      N      N      0N      PN      tN      }N      ~N      �N      �N      �N                      N      N      tN      }N      ~N      �N      �N      �N                      �N      O      PO      VO      ZO      fO      gO      lO      qO      �O                      �Q      �Q      �Q      R      R      5R                      �R      �R      �R      S                      T      T      T      (T                      tT      bV      bV      �V      �V      PW      aW      jW      �W      �W      �W      �W                      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U                      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U                      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U                      �U      �U      �U      �U      �U      �U      �U      �U      �U      �U                      jV      tV      {V      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      jV      tV      {V      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      jV      tV      {V      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      tV      wV      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      tV      wV      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      tV      wV      ~V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V      �V                      �V      �V      �V      �V                      �V      �V      �V      �V                      �V      �V      �V      �V                      8Z      `Z      �Z      �Z                      xZ      �Z      �Z      �Z                      �[      \      X\      X\                      R]      V]      Y]      p]      t]      v]      �]      �]                      �^      �^      �^      �^                      �^      �^      _      _      _      q_      �_      �_      �_      �_       `      `                      _      _      _      _      _      )_      �_      �_      �_      �_      �_      �_       `       `      `      `                      n`      s`      w`      }`                      �b      �b      �b      �b      �e      �e                      �b      �b      �b      �b                      &d      *d      .d      Vd      Pe      Ze      ^e      ce                      Zd      jd      wd      ~d                      �d      �d      �e      �e                      �d      �d      �e      �e                      e      :e      �e      �e                      �g      �g      �h      �h      �h      �h                      �g      �g      �h      �h      �h      �h                       h      5h      hh      h                       h      5h      ph      h                      �i      �i      j      7j      �j      �j      �j       l      6l      �l                       j      7j      l       l      6l      �l                      Gj      Lj      Pj      ^j                      n      *n      /n      3n      �n      �n      �n      �n                      3n      Ln      �n      �n                      Vo      oo      �o      �o                      ip      �p      �p      �p                      @q      @q      Lq      \q      �q      �q      �q      �q                      �u      �u       v      v      v      v                      �v      �v      �v      �v      �v      �v                      �v      �v      �v      �v                      Gy      Ly      Qy      cy                      �z      U{      �{      �{      �{      |                      �{      �{      �{      �{      �{      �{                      J}      U}      �}      �}      �}      �}      �}      ~                      c}      q}      )~      .~                      +      .      2      7                      ր      ��      Ё      Ձ      /�      J�                      ��      ��      ��      ��      /�      6�                      Z�      Z�      a�      i�                      i�      ��      ��      ��      /�      6�                      i�      ��      /�      6�                      ��      ��      ��      ��                      ��      ��      Ё      Ձ      6�      J�                      �      �      �      1�                      $�      -�      4�      ?�      C�      N�      Q�      ]�      a�      z�                      �      ��      ��      Q�                      b�      i�      m�      u�      z�      ��      ��      ��      ��      Ç      ȇ      �      �      �      �      "�      '�      Q�                      ��      È      ƈ      ؈                      �      �      �       �      �      ,�                      I�      I�      S�      ��      ��      T�      h�      v�                      ��      T�      h�      v�                      ��      ��      ��      ��                      ��      ��      ��      ��                      �      %�      ,�      .�      6�      9�      =�      ��      ��      �                      ��      /�      @�      @�      @�      N�                      �      +�      G�      N�                      ��      ��      ��      ��      h�      ��                      Ǐ      �      �      �      @�      O�                      @�      Y�      �      �                      @�      Y�      ��      �                      }�      ��      4�      @�                      ��      ��      4�      @�                      ��      ��      ��      ؕ      8�      u�      ��      ��      ��      ֘      [�      ��                      Œ      T�      ��      ��      ɕ      ؕ      8�      >�      C�      u�      ��      ��      ��      ��      [�      ��                      �      �      "�      "�      ��      ��                      ��      ��      ��      ��      Ǔ      Ǔ      C�      P�      U�      u�                      �      ��      ��      �      �      �                      Y�      t�      ��      ɕ      >�      C�      Ř      ֘                      ��      ��      ��      m�      ؕ       �       �      &�      u�      ��      ��      ��      ֘      [�      ��      ��                      ��      ��      O�      S�      W�      b�      g�      m�      ݕ      �      u�      ��                      p�      ��      ݗ      ��                      ��      ��      ��      ��                      m�      ��       �       �      &�      8�                      y�      Ě      �      �                      �      �      ��      �                      ��      ɛ      ֛      0�                      X�      \�      `�      t�                       �      |�      ��      ��      Н      E�      Ȣ      �                      ՝      �      8�      =�                      ֢      ڢ      ޢ      �                      M�      g�      ՟      ۟      �      V�      V�      ��       �      ��      ��      ��                      V�      }�      ��      ��                      }�      ��      ��      ��                      �      #�      #�      V�      V�      s�       �      )�      M�      ��      ��      ��                      �      �      ��      �                      V�      V�      V�      d�      i�      s�                      ��      ��      ��      ��                      ��      ��      ��      ��                      P�      Y�      n�      s�      {�      ��      ��      ̣      ��      ��                      ��      ��      ��      ģ                      k�      x�      ��      ��                      ��      ��      դ      ڤ      ޤ      �      G�      G�      P�      ��      Ц      0�      0�      H�      ��      ��                      h�      ��      ��      ��      Ц      �      ��      �                      p�      ��      ��      ��      Ц      �      ��      �                      �      L�      �      ��                      &�      L�      �      ��                      Ѥ      դ      ڤ      ޤ                      ��      *�      G�      P�      ��      Ц      0�      0�                      ��      *�      ��      Ц                      v�      z�      ~�      ��      H�      `�                      �      �      ��      ��                      �      �      ;�      ��      ��      ��                      F�      ��      ��      ��                      R�      T�      ��      ��                      �      �      �      �      :�      @�      s�      s�                      �      �       �      %�                      ��      ��      ��      �      %�      �                      �      �      %�      �                      ��      ��      %�      �                      Y�      ]�      a�      |�      ի      ۫      �      �                      ��      ��      ��      ��                      �      �      
�       �      $�      L�                      ��      ��      ��      ��      ج      ��                      ��      ��      Į      ߮                      c       c       g       �                       p      �      �      �                      �      �      �      �                      �      �      �      �                      �      �      (      �      �      �                                                          "      &      *      -      0      4      8      @      H      L                                        "      &      *      -      0      4      8      @      H      O      S                      �      �      �      8                      �      �      �      �      �      �      �      �      �      �                                                           �      �      �      �      �      �      �                                           #                      �!      Z#      b#      p#                      �'      �'      0(      8(      J(      R(      e(      q(      x(      �(      �(      �(      �(      �(      �(      �(                      �(      �(      �(      )                      �*      �*      �*      �*                      +      +      #+      �+                      +      +      #+      ?+                      1      1      1      1      $1      61                      I1      P1      Q1      e1                      �2      �2      �2      �3      y5      �5                      84      T4      \4      _4      h4      �4                      �5      �5      �5      �5      �5      6                      �6      �6      �6      �6                      �6      �6      �6      �6                      �9      r;      �;      R<      j<      H=                      �:      �:      �:       ;                      �:      �:      �:      �:      ;      ;                      �<      �<      �<      �<       =      !=                      \C      �C      �C      �C      �C      �C      �C      �C                      }E      �E      �E      �E                      �E      �E      �E      F                      PF      �F      �F      �F      �F      �G      �G       I                      'I      0I      0I      5I      AI      OI                      �I      �I      �I      J                      MJ      WJ      ZJ      oJ                      pK      uK      zK      �K      �K      �K                      M      �M      �M      �M                      _M      pM      �M      �M                      wP      �P      �P      �P                      �R      �R      PS      bS                      �R      PS      pS      �S                      �R      �R      �R      �R      �R      S      S      	S      S      S      S      S      S      #S      +S      /S                      �R      �R      S      S      	S      S      S      S      S      S      #S      +S      2S      6S                      T      �T      �T      IU      OU      RU      XU      oU                      T      �T       U       U      "U      <U                      vX      X      �X      �\      &]      ha      xa      �a                      vX      X      �X      �X      �`      �`      �`      ha                      �`      �`      �`      �`                      �`      �`      �`      �`                      `Z      cZ      yZ      �Z                      `Z      cZ      �Z      �Z      �Z      �Z      �Z      �Z                      �Z      �Z      �Z      �Z      �Z      �Z                      �Z      �[      &]      �]      >^      �^      �_      M`                      X]      k]      �]      �]                      �[      �[      �[      ,\      �^      _      �_      �_      M`      _`                      Fc      �d      �i      j      -j      �j      �t      �t                      3d      �d      �i      j      j      j      �j      �j      �j      �j      �t      �t      �t      �t                      `d      cd      gd      ~d                      -j      �j      �j      �j                      �f      �f      �f      �f                      �f      �f      �f      �f                      Vi      �i      �j      |l      �l      �t      �t      mu      �u      �w                      ei      li      }i      �i      �l      �l                      �j      |l      �q      �q      �q      r      
r      �t      �t      u      �u      aw      pw      �w                      �j      |l      �u      �v      @w      aw      pw      �w                      �j      �k      �k      �k      �v      �v      pw      �w                      �k      �k      �k      Cl                      �q      r      
r      �r      �r      �t      �t      u      �u      �u      �v      w                      �q      r      
r      rr      �s      �t      �t      u      �v      w                      t      .t      2t      6t                      .t      2t      6t      :t      =t      Pt                      �v      �v      �v      �v      �v      �v      �v      �v      �v      w      w      w                      �v      �v      �v      �v      �v      �v      �v      �v      w      w      w      w      w      w                      "m      �p      aw      pw                      �p      �p      �p      �p                      �p      �p      #q      Aq                      �w      `x      `x      wx      {x      �x      �x      hy                       x      `x      �x      Py      Zy      hy                      rx      rx      �x      �x      �x      �x                      �y      Uz      �z      <{                       z      #z      &z      *z      2z      Iz      Lz      Pz      �z      <{                      �z      �z      �z      �z      �z      �z      �z      �z                      mz      �z      �z      �z      �z      �z                      �|      }      A}      H}                      �}      �}      �}      A~                      w~      �~      (      5      9      ;                      �      �      �      �      �      �      ��      ڀ                      ρ       �      �      8�                      ֆ      ��      ؋      ��                      ��       �      ��      _�                      .�      �      ��       �       �      8�      ��      ��      ��      ͓                      `�      ��      ڏ      �      ��      ��      ��      ��                            K�      \�      `�      ڏ       �                      f�      f�      k�      ��                      ő      q�      ͓      	�                      ��      �      0�      `�                      ��      ��      ��      ��      ��      Ü      Ü      �      �      <�                      ��      %�      )�      8�                      ��      ҝ      ם      ڝ      �      �      �      �                      �      ��      ��      ��      ��      ��                      ��      @�      P�      ݣ      (�      P�      ��      ��      ��      ��                      P�      ݣ      (�      P�      ��      ��      ��      ��                      P�      ݣ      (�      P�      ��      ��      ��      ��                      (�       �      ��      ��                      ^�      d�      i�       �      ��      ��                      �      �      P�      v�      ~�      ~�      ~�      ��      ��      ��      
�      =�                      Q�      ��      ֨      ��                      ��      ��      =�      \�                      Ѥ      դ      ۩      C�      =�      ��                      դ      �      ��      ֨                      ��      ��      ��      ��      q�      ��      ��      ©      T�      =�                      s�      s�      z�      ��      �      =�                      ��      �      �      �      �      �      �      �                      ;�      P�      `�      c�      p�      ~�                      :�      B�      l�      u�      ��      ��                      ߮      �      �      ��                      �      �      ��      ��      ��      ��      ��      ��      ְ      �      ��      ��      `�      ��      ڳ      ��      ��      ��      ��      	�      	�      .�      @�      H�      X�      a�      k�      ��      ��      ��      �      =�      B�      `�      w�      ��      ��      �      !�      ��      ��      h�      q�      ��      ��      ��                      �      �      �      ��      X�      a�      ��       �      ��      ��                      կ      �      ��      ��                      �      ��      ��      ��      ��      d�      (�      =�      ��      0�      ��      ��      n�      ��                      ��      0�      n�      ��                      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      �      �      �      �                      ��      ��      ��      ��      ��      ��      ��      �      �      �      �      �                      ְ      �      e�      ��                      t�      ��       �      ��      0�      a�                      �      0�       �      .�      ��      n�                      ��      ��      ��      ŷ                      ҷ      �      �      ��                      ]�      ��      ��      ��      E�      W�                      ��      ��      ��      ��      ��      ��                      ��      z�      ��      ��      ��      ��      q�      ��                      Ⱥ      ��      ��      ��                      Q�      m�      q�      y�                      һ      ��      ��      ��                      ��      v�      ��      )�                      ��      ƾ      8�      X�                      ƾ      Ͼ      Ӿ      ��      ��      �                      �      ��      �      W�                      ��      .�      W�      ��                      2�      ��      ��      ��                      ��      ��      ��      &�                      ��      �      ��      ��      )�      F�      ��      ��                      �      M�      ��      ��                      ��      ��      ��      ��                      C�      ��      a�      h�                      ��      ��      B�      `�      ��      �      W�      ��                      ��      ��      ��      ��                      ��      ��      ��      ��                      ��      ��      :�      M�                      ��      	�      	�      �      ��      �                      �      ��      ��      ��                      ��      ��      ��      ��                      ��      L�      k�      ��                      ��      ��      w�      ��      ��      ��      ��      ��                      ��      ��      !�      E�                      ��      ��      �      (�                      ��      ^�      M�      ��                      ^�      ��      ��      ��      ��      ��                      ��      ��      ��      ��                      ��      �      ��      ��                      �      �      ��      ��                      �      ��      F�      ��      ��      ��                      @�      ��      c�      j�      ��      ��                      ��      ��      j�      ��      ��      ��                      ��      ��      F�      K�      ��      ��                      ��      ��      K�      c�      ��      ��                      	�       �      ��      ��                      ��      �      ��      ��                      �      ��      ��      ��                      ��      `�      ��      ��      ȳ      ڳ      .�      @�                      �      `�      ��      ��      ȳ      ڳ      .�      @�                      -�      E�      ȳ      ڳ                      �      G�      J�      ~�      ��      ��                      ��      ��      ��      a�                      ��      ��      ��      ��      ��      p�      1�      a�                      ��      ��      ��      }�      @�      V�      1�      a�                      ��      ��      �      !�      *�      V�                      .�      <�      D�      [�      ^�      h�      m�      ��      ��      �      ��      D�      L�      \�                      0�      5�      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      �      �                      <�      C�      [�      ^�      ��      ��      ��      ��      �      }�      1�      ��                      ��      ��      ��      @�                      ��      ��      ��      ��      0�      H�                      3�      3�      7�      R�                      e�      e�      i�      �                      ��      O�      ��      ��      ��      (�      H�      p�      ��      ��      ��      0�                      ��       �      ��      0�                      ��       �      ��      �                      �      O�      ��       �      H�      p�      ��      ��                      1�      ��      H�      p�                      ��      ��      ��       �                      ��      ��      ��      ��      ��      �      �      �                      ��      ��      ��      ��      �      �      �      !�      $�      (�                      4�      R�      T�      Z�                      �      �      �      �                      �      �      �      �                      Z      ^      h      �                      �      �             }                            �      �      �            %      8      k                                                               h      �      0      �      N      k                      ^      @      P      %                            #      '      +                      #      '      1      H                      �      �      P      �                      �      �      �      �                      z      �      �      �                                  �      �      �      �      �      �      �      �                      :       D       P       �       �       !      (!      �$                      �       �       f"      �#      �#      �$                      �"      �#      �#      �#      �#      �$                      �"      �"      �"      �"      �"      �#      �#      �#      �#      �$                      #      �#      �#      �#      �#      �$                      F#      �#      �#      �#      �#      �$                       &      N&      T&      p&                      P'      p)      �*      %+                      �'      `)      �*      �*                      .      �.      �.      �/      (0      -0                      0.      �.      (0      -0                      �2      �2      �2      3      (3      H3                      �3      �3      P6      �6                      �8      �8      �<      �<                      )9      `9      b<      �<                      �<      g=      p=      =                       =      $=      )=      b=      p=      =                      �=      F>      p>      �>                      lB      �B      �B      �B                      �C      �C      CD      �D                      �C      �C      �C      �C      CD      CD      pD      pD                      �F      G      G      EG                      eH      �H      �I      kK      pK      �K                      �I      cK      pK      �K      �K      �K                      rL      yL      �L      �L      �L      �L      �L      �L                      yL      {L      �L      �L      �L      �L      �L      �L      �L      �L      M      �M      �N      O      0O      PO      pO      �O      �O      �O      HW      �W                      �M      iN      O      0O                      !N      1N      =N      iN      O      0O                      P      QS      mV      �V      �V      %W      PX      Y      Y      �Y                      ;P      �R      mV      �V      Y      �Y                      �V      %W      PX      Y                      �S      T      �W      �W                      &U      mV      �V      �V      �W      �W      Y      Y                      5U      bU      jU      �U      �U      mV                      �Y      �Y      �Y      �Y      �Y      �Y                      3Z      1\      �\      `]      �]      �]      �]      8^                      �Z      �Z      8]      `]       ^      ^                      �Z      �Z      8]      `]       ^      ^                      �[      �[      �[      �[      
\      \      �]       ^                      1\      �\      �]      �]      8^      p^                      :\      �\      �]      �]      8^      p^                      b       �       �       �                       �      �      �      �                      �      @      U      i                      -      -      1      g                      �      �      �      �      �      �      �      �      �      �                      0      d      h      k      m      o                             S      h      h      l      r      x      z                      �      �      �      �      8      0                      X      �      �      0                      N      j      �      Q      Q      Y      �      �      �      �            	                      �      �      �                  &      �      �                      e      �      �      �      �      �      �      �      	      �                      v      �      �      �      	      �                      h      n      p      �                      n      n      p      �                      �            (      -      0      _                            �      �      �                      ;      �      �      �                      x      �      �      �                      '      a      e      k      q      �                      �      �      �      �                      8            �      �                            C      `      �                                  �      H      c      �      �      t                       �       �       !      !                      �!      �!      "      �"      �"      �"                      �#      �#      �)      �)                      Y$      ^$      q$      �$      0(      �)      .      X.      `.      }.                      h(      �)      .      X.      `.      }.                      �$       %      %      %      %      %      .%      1%      8%      F%      L%      Q%      W%      `&      �)       *      �-      .                      �&      �&      �&      	'                      p'      �'      �'      0(                      *      F*      K*      ]*                      �*      �*      �*      �*      �*      �*      �*      �*                      D+      M+      R+      `+      e+      i+                      `+      e+      o+      �+                      �+      5,      �,      X-                       -      -      -      -                      /      �/      0      �0                      Z1      i3      s3      ~3                      �1      �1      �1      �1      �1      2                      �1      �1      
2      62      @2      `2                      �1      �1      
2      2      2      12                      e2      e2      l2      t2                      t2      �2      �2      �2                      �3      �3      �3      	4      4      84      H4      ]4                      �4      �4      �4      �4                      �4      �4      �4      �4                      �4      �4      �4      �4                      �5      6      $6      �6      �6      �8      �8      �8      �8      9                      N6      �6      �6      �7      �7      V8      �8      �8                      �6      (7      @7      �7      �7      V8      �8      �8                      �9      `:      �:      ;      ;      ;                      �9      :      :      `:      �:      ;      ;      ;                      �<      �<      �<      �<      �<      �<                      4=      8=      <=      l=      y=      ~=                      &>      �?      �?      �?      @      �@                      �>      �?      @       @                      A      �B      �B      �C      �C      ED                      @A      �A      �A      8B      �C      �C      �C      ED                      @A      �A      �A      8B      �C      ED                      �B      �B      �B      C      C      PC      �C      �C                      }D      �D      �D      �D      �D      �D                      E      9E      =E      BE      PE      XE      \E      gE      mE      oE                      rE      vE      �E      �E      �E      �E      �E      BF      HG      aG                      G      'G       I      I                      �I      �I      �I      �I      �I      �I                       J      J      J       J                      DK      `Q      �Q      �T       U      0Y      0Y      3Y      PY      �o                      uK      |K      �K      N      N      $N      +N      7Q      �Q      �Q       U      HU      �X      Y      PY       [      �^      B_      ]_      �o                      ZN       Q      �_      T`      �j      �o                      aN      �N      �_      �_      �_      �_      �_      T`      �j      �m      n      �o                      �_      T`      �j      �m      n      �o                      P      P      1P      �P      �m      n                      �`      �a      �a      �j                      �`      �`      �`      �a      -c      Yc      �f      Gi      [i      �j                      fg      �h      j      �j                      �a       b      b      -c      Yc      kc      c      �c      �c      �f                      �b      �b      c      -c                      �e      ;f      �f      �f                      �R      �R       [       \                      0S      �S      �S      �T                      YU      �W      �W      �W      F\      �]      �]      �^                      aV      �V      �\      �\      �]      �]      �]      �^      �^      �^                      �]      ^      ^      ^      ^      ^                      ^      �^      �^      �^                      >^      �^      �^      �^                      �V      �V      �V      �V                      W      W      W      W      W      !W      $W      dW                      m\      �\      �\      �\                      z]      �]      �]      �]                      �W      �W      �W      �X      [       [      \      F\      �]      �]                      �X      �X      \      F\      �]      �]                      V      �      �      �      �      �                      �      �      �      �                      �      �      �      �      �      �      �      �                      �      S      V      �      �      �                      `      �      �      �                      �      �      �      �      �      �                      A	      ^             %      0      E                      �	      �	      �	      �	                      �	      �	      
      
                      S
                                         �
      �
      �
      �
                      j                               �                      8      h      �      @      @      F      P                  �$                      8            �      �             @      �             P      �            �$                      8      =      \      h      v      v                      =      D      K      N      h      q      v      �      �            `      �             0      �      �                  ;      E      �      �                      �      �      `      �      ;      E                            �      `      �      �      �      ;      E                      &      �      0      0      �      �      P            �                           )#      X#      g#      y#                      9      =      B      �      P            �                           )#      X#      g#      y#                      9      =      B      P      P      �      P      �      �                           )#      X#      g#      y#                      �      �      �                           )#      X#      g#      y#                      �      �      �                           )#      X#      g#      y#                      �      �      �      �      �      �      �                           )#      X#      g#      y#                      !      �      �                           )#      X#      g#      y#                      ]      �      �                           )#      X#      g#      g#      o#      y#                      �             o#      y#                      �      �      �      `             �            ;      E      b                    X#      ]#                      0      �      ,      ;                      (      �      �      �                      H       )#      ]#      g#      y#      /$      8$      �$                      �       #      ]#      g#      y#      �#      <$      �$      �$      �$                      �       =!      �$      �$                      �!      �!      ]#      g#                      #      �      �             @      h             @      �                            �      �      @      h      �                                   G       P       U                       {       �       �       �                       �       �       �       U      Y      �      �      �                      /      6      B      n      �      �                      �      �      �      �                      �      �      �      	                            "      %      Q                      )	      �	      
      -
                      �      �      �      �                      *      3      @      U      e      i      m      t                      �      h      �      �      @      p            -      -             �      �      3      �      �                            -      -      -      �            
                      �      �      �      �                      �      �      �      �      �             3      �      �            
                            �      �      �             3      �      �            
                            �                        P                             �      G      �      �                      =      �      �      �      �      �      
      
                      ]      �      �      �                      h      �      �      �      �      @      p                   �      �                        %      3      �      �            2                      l      t      x      �      �      �      �      @      p      �      �                   �      �      �                                  �      �      [      �      �      �                      �      �      �      H                      �      �      �      �      �      @      p      �      �                   �                      �      �      �                                        Z      e      �      �                      p      s      w      �                      �      �      �      �                                         �      �      �      �      �                      �      �      �                            D      G      J      N      R      e                      G      J      N      R      k      ~                      �      �      �      �$      %      W&                      /      4      ;      D      H      ]      d      r      w      �      �      �      �      �      �      �      -      �      �$      �$                      �      �      �      �      �      �      �                  �      -      {      �$      �$                      �                  �                      �      �      -      -                      �      -      �      �$      �$      �$      %      W&                      %       �       	#      �$                      �!      �"      �$      �$      %      W&                      "      H"      P"      m"      s"      �"      �$      �$      %      �%      �%      �%      �%      W&                      s"      �"      �$      �$                      r&      r&      v&      �'                      �&      �&      �&      �'      �'      �'                      �'      �'      �'      �'      �'      �'                      #(      %(      )(      2(      O(      f(      n(      w(                      �(       )       ,      
,                      �(      )       ,      ,                      ;)      D)      K)      d+      d+       ,      
,      ',                      �)      �)      �)      d+      d+       ,      
,      ,                      d+      d+      d+      �+                      3,      7,      =,      N,      U,      �.      �1      �1      2      �4      �4      R5                      �-      �.      �1      �1                      �-      .      ".      �.      �1      �1                      3      �4      +5      R5                      �3      64      F4      �4      +5      R5                      �4      �4      �4      5      5      5      &5      &5                      �4      �4      �4      5                      �.      �1      �1      2      2      2                      �.      7/      �1      2                      X0      d0      q0      v0      �0      �0      �0      �0                      �0      1      2      2                      �      �      �            	      5                      �      �      �      �      �      �            	      @	      /
      4
      <
                            e      4
      <
                            Y      �      	                      �      �      �      	                      �      �      �      �      `      d      x      p      �      �                      �      �      �      �                      8      k      �      @      �      �                      �                              S      W      b      i      �                      +      2      =      B      F      K      T      Y      ^      c                      �      �      �      E      P            x      �      �      �              $      2$      %                      �      �      �      �      �      �                      �      @      �                            (      @      �                            [      `      k      �      x      c      k      v      �      �      X$      �$                      v      �              �       &!      "      �$      �$      �$      %                      �      "      3      �              �       &!      "      �$      �$      �$      %                      �            &!      "      �$      �$      �$      %                      +!      "      �$      �$      �$      %                      -!      H!      [!      "      �$      �$      �$      %                      �!      �!      �!      �!      �!      �!      �!      �!      �!       "      �$      �$      �$      %                      �"      $      2$      X$      �$      �$                      �"      �"      �"      $#      2#      $                      �      0      X      h      $      2$                             '      .      3      ;      �                      �      X      �                              �      �      �      �      0      \      h      �                      Y      r      v      �      �      �                      �      �      �      �      �      �      �                   d      	      �	      �
      *      P      ;      X      �      �                            	      y	      �
      *      P      ;      X      �      �                            �
      *      ;      ;      f      �                      �
                              %      f      v      v      �      �      �                      P      ;      X      f      �      �      �                            D      �      x      �      �	      �
      :      P                      �      �      �      L      �	      �	                      �                                        *      *      .      U                      H       J       Q       �       �       �                       �             `      d      h      k      l      �                      8      ?      C      W                      �      �      �      #                      `      g      k      q                       
      N
      N
      T
                      Q      S      X      h      �      �      (      [      p      �      �      �      !      !      "      "                      I      �      p      �                      `      �      p      �                      h      n      z      �      �      �      j      q      �      Q       [       �       �       !      (!      �!                      h      n      @      \              Q       [       �       �       !      (!      �!                      �      �      �      �      j      q                      B      �      �      �                      b      �      �      �                      \      �      �!      �!                      �      P      �      �      �      �      �      �      Q       [       �       �       !      (!      �!      "                      �      �            P      _      �      �!      �!                      j      �      �      �      �      �                      �      j      �            �      �                      x      �      �      �      �      q      q      {                      }      e      �      ]      {      �                      4"      @"      G"      L"                      @"      G"      L"      _"      0$      K$                      �"      �#      �#      �#                      p#      �#      �#      �#                      �#      �#      �#      �#                            
            K      X      y                      �      �                           $      (      .      /      D                      y      �      �      �                      Y      �      �      �      �      �      �                            W      �      �      �                      @      c      �      �                      X      h      r      z      �      Y      �      i      k      �      H!      �!      �#      �#      �%      �%                      �      �      �      �      �                                        �      �      �      �      �      �      �      �                        %      �      P      �      (      H!      �!      �#      �#      �%      �%                      �            �      �      �%      �%                      �      H!      �!      �#      �#      �#      �#      ($      @$      �%      �%      ('                      �            �"       #      �$      �$                      u      O      �       7!      �!      �!      8"      �"                            /      e      e                      >      V      e      e                      �      K      �       7!                      �      >      �       7!                      �      W       �!      "      �#      ($      @$      �$      �$      �%      �&      '                      �      �      �                             #      �#      �#      �#      �%      �&      '      ('                       #      #      #      "#                      #      #      "#      1#                      G#      �#      �#      �#                      �%      �&      '      ('                      �&      �&      '      ('                      �(      �(      @*      H*                      H*      M*      Q*      �*      [+      �+      �+      �,                      �*      �*      �*      �*      �+      �+      b,      b,      p,      y,      y,      �,                      �-      �-      �-      @.                      �/      �/      �/      �/                      �0      1      1      �1      m4      m4      m4      w4      �4      B5                      1      1      1      !1      (1      (1      +1      01                      -2      /2      32      B2                      *6      A6      O6      R6                      �7      �7      �8      �8      e9      p9      �9      �9      ;      ;      s>      �>      n@      p@      �A      �A                      P>      j>      �A      �A                      �?      n@      p@      x@      !A      .A      hA      uA                      �A      jB      sB      �B                                        =      p      �                      Z      �      �      �                      v      �      �      �                      !      &      ,      /      1      4      6      U      ^                  
                  $      1                      b      o      �      �      �      �      �      �      �      �      (      v      w      {      �      �                      b      o      (      Y      d      v      w      {      �      �                      �      �      �      �      �      �                      �      �      �      �                      |      $	      x	      B
      h
      |
                      V      �      �      �      �      �                      �                              �      H      Q      Y      d      �      �      �            !      :      d      �                            �      �      �      �      �                      �      �      �      �      ~      �                      �            N      �                      �      /      Y      �                      F      L      Q      �      �      �                      �      _      g      �                      �            (      <                      �            	                  �      �      �              �                       �      �      	                         �      �              �       �       �                       �      �      �       �                       �      �      �       �                               �       �       �                       (       n       �       �       �       �                       0"      �"      �#      �#                      �"      c#      t#      �#                      T$      Y$      `$      e$      l$      �$      �$      �$      �$      �%      �%       &      &      F&                      '      @'      G'      `'      l'      p(                      �(      �(      �(      )                      �)      �)      �)      C*                      p*      +      �,      "-                      �*       +      �,      "-                       +      0+      7+      P+      U+      j,      p,      �,      �,      �,                      I.      P.      b.      p.                      �.      '/      @/      h/                      �2      �2      �2      3      �3      �3                      �4      6      6       6      *6      06      H6      N6      R6      U6      _6      7      %7      �7                      �4      �4      �4      �4      6      6                      �7      �7      �7      D8      h8      �8                      �?      �?       A      hA                      �?      �?      �?      �?                      @      @      @      @      &@      1@                      �D      �D      �D      E      E      0E                      �E      8F      �G      �H                      PF      G      HG      �G      �H      �H                      �I      rJ      �L      �L                      K      �K      �L      �L                      L      xL      �L      �L                      N      �N      �N      �N      0P      zP                      �O      �O      �O      	P                      �Q      �Q      �Q      �Q      �Q      �Q                      �S      �T      /X      /X                      kT      �T      �T      �T                      �T      �U      �W      /X                      6U      WU      `U      �U      �W      �W      �W      X                      �U      V      V      V      V      UV      lV      qV      uV      �V      *W      �W      9X      hY                      �V      �V      *W      /W      IW      �W      iX      hY                      �W      �W      sX      zX                      zX      Y      Y      hY                      �V      W      W      W      W      %W                      �[      �[      �[      `]      �]      �]                      �[      �[      �\      `]      �]      �]                      ]      M]      �]      �]                      �]      �]      �]      =^                      �_      �a      (d      Gd      �d      tg      g      h      8h      Uh      #i      Vi                      A`      I`      P`      �`                      �`      �`      (d      Gd                      �d      �e      hg      tg      �g      �g                      e      e      e      qe      hg      tg                      e      e      'e      Ve                      �e      hg      8h      Hh                      �e      hg      8h      Hh                      ,f      ?f      Gf      pf      sf      g                      xc      �c      �c      �c                      �i      �i      �i      +j                      fj      &k      Dk      �k                      �j      &k      Dk      Qk      pk      �k                      �l      m      xq      �q                      [m      �p      �p      �p      `q      xq                      �o      �o      �o      @p                      ts      �s      �s      xt      �t      �t      �t      pu                      �s      xt      �t      �t      �t      pu                      �s      �s      �s      xt      �t      �t      �t      pu                      v      v       v      Xv                      �y      �|      �|       }                      �y      �y      �y      �z      �z      �{      �{      �|      �|       }                      dz      �z      �z      6{      �|       }                      �z      �z      �z      #{      '{      ,{                      C{      �{      �{      `|      x|      �|      �|      �|                      �{      �{      �{      `|      x|      �|      �|      �|                      $~      $~      %~      <~                      d~      d~      e~      |~                      �~      �~      �~      �~                      �      ր      ڀ      ߀      �      Ё      Ђ      ��      ؃      N�                      �      a�      ?�      G�                      a�      ��      G�      G�      p�      w�                      ��      ր      ڀ      ߀      �      Ё      G�      p�      ؃      N�                      ڀ      ߀      �      n�      z�      Ё                      ڀ      ߀      �      ��      ��      Ё                      Ё      Ђ      ��      ؃                      |�      ��      ��      ��                      ��      ��      `�      x�                       �      S�      ��      ��                      ��      ��      ��      ��      �      
�                      ��      Ԇ      ��      �                      0�      J�      Z�      ��      ��      ��                      ��      ��      ��      ��      ي      ي      ي      �                      H�      h�      v�      h�      ي      ي                      ��      P�      ي      ي                      �      �      �      +�      -�      2�                      ��      :�      >�      I�      O�      X�      X�      Z�                      ��      ��      ��      ��                      Ȍ      ��      ��      ��      �      x�      ��      N�      `�      t�      @�      ��      �      (�      $�      `�      `�      y�      ��      ��                      ̌      ь      K�      y�      �      b�      `�      t�      �      (�      $�      `�      ��      ��                      ̌      ь      P�      `�      `�      ͜      I�      Y�                      ̌      ь      P�      `�      q�      ��                      Q�      Ϗ      ԏ      ؏      ݏ      �      �      �      �      �      �      �      �      (�                      ��      ��      ��      Ő      ΐ      @�                      ~�      �      �      P�                            ��      ��      ��      @�      ܖ      `�      y�                      ݒ      ��      ��      œ      t�      @�      ��      �      (�       �      y�      ��                      7�      9�      �      �      X�      @�      y�      ��                      ��      0�      f�      x�       �      �      �      8�                      ��       �      8�      {�                      ͢      8�      ��      Ȥ                      8�      ��      Ȥ      ��                      ��      ��      ��      Ш                      ף      ��      ��      ��                      Ȥ      �       �      ��      �      P�      ث       �                      &�      ��       �      ��      �      P�      ث       �                      &�      0�      K�      S�      W�      (�      8�      ��      �      P�      ث       �                      "�       �      Ш      �      d�      ��                      "�       �      Ш      ;�      @�      P�      Z�      ^�      a�      e�      ��      �      d�      ��                      
�       �      Ш      ��      ��      �                      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ©      ĩ      ǩ      ʩ      ̩      Ω      ԩ      �      �      �      �      �      �                      ��      ��      ��      ��      ��      ��      ��      ��      ©      ĩ      ǩ      ʩ      ̩      Ω      ک      �      �      �      �      ��      ��      ��                      ԩ      ک      �      �      ��      ��      ��      �                      �      �      �      �      �      ;�                      P�      ث       �      d�                      �      �                              !      :                      X      e      �      B                      p      p      t      ~      �      �                      �      �      �      �      �      �                      �      �      �      �                      �      �            �                      �      �      $      `                      �      �      �      �                      /      >      B      S      V      �                      �      �      �      	      	      
	      	      	                      U	      �	      �	      �	                      U	      v	      {	      �	      �	      �	                      �
      �      =      \      k      �                      �
      �
      �
      �
            
                  &      )      3      �      k      �                      p      �      �      �      k      �                      �                                                                 .      A                      =      \      �                             	                  �                        A      �      �                      	            �      �      �      �                        A                      _      �      �      �            A                            (      E      �      �      �                      �      �      F      �                      Q      t      |      �                   �      �                      Q      t      �      �      �      �      (      d      d      �      �      �                   �      �                      Q      j      o      t      �      �      h            @      f      �      �                   �      p                      Q      j      o      t      t      �      �      �      �            �      �                   �      Y      `      d                      `      �      �      �                            k      m      �      �      �      �      �      �      8                      �      �      �      �                       �      �      �      �                       �      �            �              �                             Y      �       �                       Y      �      �       �                       s      s      v      �                      �!      �"      �"      �"                      �!      �!      �!      �!      �!      �!                      �!      �!      �!      �!      �!      �!                      �!      �!      �!      �!      �!      �!      �!      "                      "      �"      �"      �"                      6"      K"      x"      x"      {"      �"                      �#      �#      �#      �#      �#      �#      �#      $                      '$      `$      m$      �%      �'      (                      /$      4$      ?$      `$      �$      %      %      �%                      �%      �%      &      &                      H&      �'      (      I(                      �&      �'      �'      �'      (      I(                      �&      ]'      b'      �'      �'      �'      (      @(                      �&      Y'      �'      �'      �'      �'      (       (      )(      @(                      �(      )      �)      P*      0,      �,                      �)      P*      0,      �,                      �)      �)      �)      �)      �)      *      *      	*                      �,      �,      �,      �,      �,      �,                      X)      Z)      ])      �)                      �)      �)      �)      �)                      �*      �*      +      �+       ,      0,                      �*      �*      �+      �+       ,      0,                      +      +      	+      +      +      +      +      )+      7+      ;+                      +      +      ,+      /+      3+      7+      ;+      C+      E+      I+      �+      �+                      )+      ,+      /+      3+      L+      O+      V+      Z+      b+      n+                      [.      [.      \.      �.      �.      �.      �.      �.                      �/      0      �0      �0                      �3      H4      �5      l6                      
4      H4      �5      [6                      4      @4      �5      [6                      h4      �4      �4      5      (5      �5                      7      7      !7      $7      )7      �7                      �7      3:      H:      �>                      �7      �9      H:      �:      `>      x>      �>      �>                      `8      �8      �8      �8                       9      �9      `>      x>      �>      �>                      �9      �9      `>      x>                      �9      �9      �9      �9      `>      x>                      �9      3:      �:      `>      x>      �>                      �9      3:      ~<      �=                      �9      $:      1:      3:      �<      �=                      1:      3:      �<      Z=      c=      �=      �=      �=                      1:      3:      =      V=      ~=      �=      �=      �=                      =      E=      �=      �=                      �:      
;      
;      ;                      ,;      j<      �=      `>                      ,;      E;      �;      �;      �;      6<                      �;      �;      �;      6<                      �;      �;      <      (<                      �?      �?      �?      �?      �?      �?                      \@      p@      �@      &A      PA      /B      AB      �B      C      C                      PA      WA      PB      �B      C      C                      �C      �C      �C      �C                      dF      kF      �F      0I                      BI      FI      �I      �L      @M      �T                       J      'J      FJ      _J      �S      �S                      _J      �J      pM      YN      PS      TS      TS      `S                      xM      �M      �M      YN      PS      TS                      kK      �L      `S      �S      �S       T                      kK      oK      {K      }K      �K      �K      �K      �K                      �K      �K      �K      �K                      �L      �L      �L      �L                      �L      �L      �L      �L      �L      �L      �L      �L                      �N      @Q      �T      �T                      �O      P      P      #P                      �O      �O      �O      �O                      ^P      cP      fP      jP      sP      �P                      @Q      �Q      pT      �T                      �Q      �Q      �Q      �Q      R      R      R      )R                      |R      PS      �T      �T                      ]I      eI      mI      mI      pI      }I      �I      �I                      }I      �I      �I      �I                      �L      M      	M      !M                      �W      �W      �W      �W                      �W      �W      @X      GX                      �W      �W      �W      @X      `X      �Z                      �W      �W      �X      �Y                      %Z      LZ      `Z      iZ                      /[      5[      8[      A[      J[      Y[      \[      `[      p[      s[                      5[      8[      A[      J[      Y[      \[      `[      d[      h[      p[      s[      w[      �[      �[                      �[      \      �]      ^      ^      H^                      �\      ]      ,]      `]      �]      �]                      �\      �\      �\      �\      �\      ]      ]      ]                      h]      h]      r]      �]      �]      �]                      �]      �]      �]      �]      �]      �]                      �^      �^      �^      �_      �_      �_      �_       `      6`      g                      �^      �^      �^      _      0_      �_      E`      �b      �b      �b      �b      �b      �d      �d      �d      9e      >e      f      f      g                      0_      U_      b_      �_      0f      @f                      �_      �_      �_      �_                      K`      P`      X`      n`      w`      �`      �`      Pa      Ta      Ya      pb      �b      �d      e                      �`      �`      �`      �`      �`      �`                      �d      �d      �d      e      e      e                      �a      �a      pe      �e      �e      f      pf      g                      �a      �a      �a      �a      �a      �a      �a      �a                      b      pb      �b      �b      f      0f      @f      pf                      �b      ]c      �c       d      �d      �d      9e      >e      f      f                      �b      Tc      �c       d                      �c      �c      �c       d                      +d      /d      3d      �d                      Hd      Md      Qd      hd                      Wg      �i      j      "j      "j      &j      0j      ]u                      ng      qg      �j      0l      `t      �t                      ng      qg      �j      0l      `t      rt                      ng      qg      Mk      0l                      ng      qg      yk      0l                      ng      qg      �k      0l                      �j      �j      �j      �j      k      k                      �g      �g      �g      Ai      El      Hl      Pl      `m      �m      9p      �p      �r       s      `t      u      (u      Nu      ]u                      h       i      �m      �n      �n      @o      Pr      �r      �s      �s      Nu      ]u                      �h       i      �m      `n      �n      @o      �s      �s                      pn      �n      Pr      �r      Nu      ]u                      �l      m      m      `m      �n      �n      �s      �s                      �l      �l      �n      �n      �s      �s                      �o      �o       s      �s      @t      `t      u      (u                      �o      9p      �p      Pr      �r      �r      �s      @t                      �o      �o       q      Aq      �q      Pr      �s      @t                      Ai      �i      9p      �p      �r       s      (u      Nu                      j      j      j      "j      `m      `m      em      lm      pm      m                      5j      =j      Cj      Lj      Qj      [j      bj      tj                      Lj      Lj      Qj      [j      bj      tj                      �t      �t      �t      u                      �t      �t      �t      �t                      �u      �u      �v      w      ?w      Jw                      @v      fv      lv      �v      0w      ?w                      Rw      Yw      uw      uw      �w      �w      �w      �w      �w      �w                      |w      �w      �w      �w      �w      �w      �w      z      z      Bz      Yz      �z                      |w      �w      �w      �w      �w      �w      �w      �w                      x      $x      �y      �y                      �x      �x      �x      �x                      �x      �y      kz      �z                      y      y      y       y      kz      �z                      �y      z      z      Bz      Yz      kz                      �z      �z      �z      �z      �z      �z                      {      �|       }      �                      X{      �|       }      z}                  �      �                      �{      �{      �{      �{      �{      �|      }      z}                      �{      L|      `|      ||      }      z}                      �      �      �      �      �      �                      �      S�      V�      _�      ��      ��                      r�      y�      ��      ��      ��      ��      ��      ��      Ł      ʁ                      ��      ��      ��      ��      ��      Ł      ʁ      7�      :�      b�      y�      ʄ                      ��      ��      ��      ��            Ł      ف      �                      5�      D�      ��      ȃ                      ��      ��      ��      Ԃ                      �      ��      ��      ʄ                      ,�      4�      7�      @�      ��      ʄ                      ȃ      7�      :�      b�      y�      ��                      �      �      "�      *�      /�      8�                      P�      �       �      ��      ��      X�      ��      ��                      ��      �       �      ��      ��      '�      n�      X�      ��      ��                      �      ��      ��      ��       �      ��      ��      ��      �      '�      n�      X�      ��      ��                      Z�      s�      ��      e�                      m�      p�      ��      �       �      e�                      p�      p�      0�      @�      G�      ��      ��      ��      �      �      n�      X�      ��      ��                      �      @�      n�      X�      ��      ��                      ��      X�      ��      ��                      �      ��      ��       �      (�      X�      ��      ��                      y�      ��      ��       �      X�      ��                      ��      ��      ��       �                      ��      ��      ��      ۈ      �      ��                      X�      z�      ��      ��                      �      �      �      �                      �      (�      0�      7�      H�      H�      M�      R�      Z�      ]�                      f�      ��      ��      Ò      �      �                             "       '       +       .       g       �       �                       >       K       N       Q       V       c                             H      L      \                                        1                      �      �      �      7                      #      @      P      i                      z      z            d      l      �                      �      �      �      �                      �                                                                                          !      %      ?      K                                        !      %      8                      �      �      �      7                      �      �      E      r      u      �                        ,                      �      �      P      P      ]      r      u      y      �      �      �      �                      �      �            ,                      �      �      �      �                      �      	      "	      #	                      P	      S	      a	      �	      �	      -
      1
      4
      H
      �                      �	      �	      H
            p      �                      P
      r
      p      �                      �
      �
      �      �                      �	      -
      1
      4
                      	
      -
      1
      4
                      ~      �      �      �      �      �                      �      s      |      �      �      �                            f      |      �                      x      |      �      �                      @      G      G      e      g      z                      �      �      �      �      �                            �      �      �      �      �                            �      �      �      �                      C      �      �            0      �      �      �                      u      �      �      �      �      �                      �      �      0      �                      �                   %                      �      �            0      0      �      �      �                      �            �      �      �      �      �      P                      �            �      �      �      �      �      P                      �            �      �      �      3      �      P                      �                   @                      p      p      t      �      �      �                      t      w      z      �                      �      �      �      �                            �      �      /                      �      7      7      =                      7      7      =      B      E      �      �      �                                   E      L      P      �      �      �      �      �                      �      �      �      �      �      �      �      �      �      �                      �      �      �      �      �      �      �      �      �                  �       �       �"                      �      �      �      �                      Y      b      M      ]      a      }       �!      ("                      b      �      �      �      P!      z!      ("      �"                      k      �      P!      z!                      v      v      �      �      �      �      �      �                      �      �      �      H      �"      �"                      H      M      Q      �                      �"      �"      �"      �"      �"      �"      �"      �"      #      #      #      D#      �#      )      �3      �3      �4      �4      7      a7                      �#      �#      $      �$      �4      �4                       $      )$      2$      �$      �4      �4                      �$      �&      7      a7                      �$      �%      �%      �&      7      a7                      %      ;%      �&      �&                      U%      �%       &       &      `&      v&      7      7      @7      @7                      �&      �&      �&      #'      7      7                      #'      �(      �3      �3                      8'      8'      N'      �(      �3      �3                       )      �3      �3      �4      �4      7      a7      �7                      ()      -)      4)      ;)      B)      E)      J)      N)      S)      a)                      �)      �)      *      *      �5      7                      �)      �)      *      *      �5      7                      �*      �*      X,      �,      �,       -      �4      �4      �4       5                      �*      �*      X,      �,                      �*      �*      �,       -      �4      �4      �4      �4                      G+      X,       -      f-      14      |4                      �+      �+      �+      �+      �+      X,                      �-      $.      �3      �3      |4      �4                      �-      �-      �-      $.      �3      �3      |4      �4                      �-      �-      �-      $.      �3      �3      |4      �4                      �-      �-      �-      �-      �-      .                      P.      ^0      �3      4       5      r5      a7      �7                      �.      /      /      !/                      &/      @/      �/      00      �3       4      )5      r5      a7      �7                      0      00      X5      r5      a7      �7                      �3      �3      �3      �3                      .5      .5      15      I5                      ^0       1      �1      @3      �7      �7                      �0      �0      �1      @3      �7      �7                      �0      �0      �1      �2      �2      �2      �7      �7                      �0      �0      %2      %2      (2      B2                      2      2      h2      {2      �2      �2                      �2      �2      �2      �2                      �7      �7      �7      �9      �9      �9                      �7      �7      �7      �9      �9      �9                      |8      �9      �9      �9      �9      �9                      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8                      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8                      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8       9      9                      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      �8      9      9                      �8      �8      �8      �8      �8      �8      9      $9                      �8      �8      �8      �8      �8      �8      9      $9                      �9      �9      :      	:      :      �:                      �9      �9      :      <:      F:      N:                      (:      <:      F:      N:                      <:      F:      N:      {:                      �:      �:      �:      �:                       ;      �;      �;      �;                       ;      ;      �;      �;                      .;      9;      <;      �;                      �;      �;      �;      �;      <      [<                      �;      �;      �;      �;      <      X<                      w<      w<      <      �<      �<      �<                      w<      w<      <      �<      �<      �<                                        h                      C      F      F      O                      %      s      �                             	      m	      
      @
                      �      �      �      �                      �      �      �                            �      �            &      *      ?      S            �      �      �      �      x      �      �#      �#      �#      �#                      �            �      �      �      �      h      �      �#      �#      �#      �#                      �      �      �      �      �            �      �      �      �      �#      �#      �#      �#                      �      �      �      �      �      �      �            �      �      �      �      �#      �#      �#      �#                            �      �#      �#                      X      �      �                            �      h      x      �                      �            #      h                      �      x      �      �#      �#      �#                      �      �      �      �                      �      �      �      �                      (      Z      �"      �"                      0      @      �!      �!      `#      p#                      v      �      �"      �"      P#      `#                      �      �       #      %#                      �      �      �!      ("      %#      P#                      C!      {!      p#      �#                      �%      '      '      R'                      �%      �%      +'      R'                            f      p      �                      �      �      �      �                  0      5                      `      �      �                            	      P
      p      `                             �      �             �      K                             �      P      �                             �      �      �      �                            �      �      �      �      �      b                      �	      �	      �	      �	                      `
      d
      h
      v
                      �      �      �      �      �            p      v      �      �                      �      �      �      �      �      0      �                    `       f       \"      f"      �#      �#      E$      E$      �$      �$      B)                      �            �      �      �      �      �                  0             *       f       s       �       �       #"      \"      f"      s"      f#      �#      �#      �#      Y%      �%      �%      �%      �%      �%      2&      �&      �&      �&      �'      �'      �(      �(      ,)      B)                      �      �      �      �      s"      T#      $      2$      J'      �'                      N      a      ~      )      %      "%      &      $&                      �      �      �      �      �      �      �       �       �       �!      �&      '      �'      �(                      �      �      �      �      �      #      �       �       �       �       �       �       !      !      !      �!      �'      �(                      (      1      ;      @      T      T      Y      �      �      �      �      �      �&      �&                      2$      E$      E$      E$      E$      e$      p$      �$      '      1'      �(      !)                      2$      E$      E$      e$      p$      �$      �(      �(                      _)      f)      �)      �)      �)      K*      `*      �*      �*      �*      �*      �*      �*      �*                      _)      f)      �)      �)      �)      8*      `*      �*      �*      �*      �*      �*                      &+      [+      ^+      e+      p+      �+                      0+      [+      ^+      e+      p+      �+                      �+      �+      P,      �,                      :-      �-      �.      �.      /      /                      �-      .      P.      �.      �.      	/      /      �/                      �-      .      P.      s.      �.      �.                      �.      �.      �.      	/      /      �/                      /      ,/      2/      �/                      �       >      �      �                                                    %      )      �      �      �                      P      �      �      �                      �      �      �                            �      �      �      �      �      �                      (      [      �      �      �      o	      �	      �	      �	      �	                      �      �      �	      �	                      �      �      o	      �	                      �	      l
      �
      �                      ;
      B
      B
      l
      �      �                      ;
      B
      �      �                      �
      �
      �
      �
                      �
      �
      �
      �
                      �
      �
            �      �      �                      �
      �
                                   @      b      o      �      �      �                      �                   �                      �      �      �      �             ^                      x      {      �      �      �      �                      `	      �	      
      
                      �	      �	      �	      �	                      @
      @
      N
      R
      U
      Z
                      ~
      �
      �
      �
      �
      C      `      v      �      �                      �
      �
      �
                  !                      �      �      �            0      X                            C      l      �                      �      �      �                            �                                        h      �      �      �      �      Z      p      �      �      �      �                            �      �      �      �      �      �      �      �      �                            7      �             (                      �      �      �      �                      �      �      Y      Y      �      �                      �            �      �      �      �                      �      �      �      �      �      �      �      �      �      �                      Y      _      c      q                      �      �      �      �                            )      �      �                      V      Z      ]      �                      0      :      <      >      C      C      G      [      �      �      �      �                      _      _      a      r                      �             p!      �!                      G       z       �       �       �       !      �!      �!                      `"      �"      �"      �"      #       #      0#      H#                      P#      P#      W#      [#      a#      f#                      �#      `$      �$      &      0&      �'      �'      0(      �(      �(                      �#      ($      �$      �%      �(      �(                      �#      $      	$      ($      3%      �%                      `&      �&      �&      �&      �'      0(      �(      �(                      �&      p'      �'      �'                      0(      j(      z(      �(      �(      �(                      @*      @*      [*      d*                      B*      E*      d*      g*      k*      #+      8+      �+                      �*      +      	+       +      H+      P+      `+      �+                      �+      �+      �+      �+                      �+      1,      5,      [,                      -      Y-      `-      `-                      u-      x-      �-      �-      �.      �.                      �-      �-      �-      �-      �.      �.                      
.      .      .      .      .      .                      6.      <.      =.      W.                      �6      7      7      ;7      ?7      A7                      �7      �7      �7      �7      t8      y8                      �7      �7      �7      �7                      �9      �9      �9      �9      �9      �9      �9      :                      :      :      :      ":                      ,:      0:      8:      h:      p:      x:                      �:      �:      ;       ;      ,;      �;                      V<      |<      �<      �<                      B=      K=      Q=      r=                      >      >      >      >      >      !>      5>      9>      =>      @>      C>      G>      G>      O>      S>      V>      ^>      b>                      $>      '>      (>      />      9>      =>      @>      C>      G>      G>      O>      S>      V>      ^>      b>      f>                      u>      y>      }>      �>      �>      �>      �>      �>      �>      �>                      y>      }>      �>      �>      �>      �>      �>      �>      �>      �>      �>      �>                      �>      �>      �>      �>      �>      �>      �>      �>      �>      �>                      �>      �>      �>      �>      �>      �>      �>      �>      �>      �>                      @      �@      E      �E      �E      F      3H      jH      jH      oH      oH      I                      0E      8E      =E      LE      QE      WE      hE      hE                      8E      =E      \E      hE      �E      �E                      `H      dH      jH      oH      �H      �H      �H      I                      �@      �@      F      �F                      �@      �@      F      AF                      �A      �A      �A      *C      *C      �C      8D      E      �F      �F      �G       H                      �A      �A      8D      DD      �F      �F                      �A      C      PD      E      �G       H                      �A      �B      �D      �D      �D       E      �G       H                      �B      �B      �G      �G                      3C      PC      TC      �C                      �C      �C      �C      �C                      �C      �C      �C      �C      D      D                      �F      �F      �F      PG                      G      G      G       G                      PG      TG      cG      mG                      �G      �G      �G      �G      �G      �G                      �J      �J      �J      /K                      |K      �L      �L      �L      M      M                      �K      �L      �L      �L      M      M                      �K      �K      �K      �L      �L      �L      �L      �L      M      M                       M       M      :M      FM      hM      kM                      pM      }M      �M      �M                      iN      �N      pP      �Q      R      R      US      `S                      �N      �N      �N      �N      �N      �N      �N      �N      �N      �N                      �N      �N      �N      �N      �N      �N      �N      �N      �N      �N                      pP      pP      �P      �P      �P      �P      �P      �P      �P      �P      �P      �P                      �P      �P      �P      �P      �P      �P      �P      �P      �P      �P                      �P      �P      �P      �P      �P      �P                      @T      @T      IT      PT      ST      UT      �T      �T                      �W      �W      �W      �W      �W      �W      �W      �W      �W      �W      �W      �W                      �Y      ?Z      �Z      �Z                      �[      �[      �[      �[      �[      �[                      \       \      (\      1\      5\      :\                      �\      �\      �\      ]      P]      U]      `]      �]      �]      �]                      �]      �]      �]      �]      ^      6^                      �]      �]      �]      �]      6^      C^      G^      y^      �^      �^                      >^      C^      G^      p^                      �]      �]      y^      �^      �^      �^                      �^      �^      �^      �^                      5_      5_      9_      >_      B_      G_                      �_      �_      �_      �_      �_      �_                      ;`      A`      C`      F`      O`      S`      Z`      i`      n`      r`                      `a      ca      ea      ia      la      a                      �b      �b      �b      �b      �b      �b      �b      c                      �b      �b      �b      c                      �d      �d      He      h      h      2h      8h      �j                      �d      �d      �e       f      hg      h      h      2h      8h      �h      �h      �j                      �d      �d      h      2h      8h      �h      �h      yi                      �d      �d      �d      �d      h      h                      Nh      �h      �h      Di                      �d      �d      hg      h      yi      sj      xj      �j                      lg      �g      �g      �g                      �g      �g      �i      sj      xj      �j                      �g      �g      �i      Cj      xj      �j                       f      �f      �h      �h                      (f      �f      �f      �f      �h      �h                      0f      �f      �f      �f      �h      �h                      �j      k      k      -k                      `k      k      �k      �k                      �k      �k      �k      �k                      l      &l      .l      7l      Tl      ]l      cl      hl                      l      &l      .l      3l                      m      m      Mm      Um      �m      �m      �n      Vo      ]o      �o      �o      [p      `p      ep      mp      op      tp      {p                      �n      �n      �n       o      o      o      @o      Go      �o      �o                      �n      �n      ko      �o                       o      o      o      $o      ]o      do      �o      �o                      o      o      $o      ,o      do      ko      �o      �o                      m       m      6m      =m      bm      bm      rq      tq      �q      �q      �q      �q                      jm      rm      �m      �m                      �m      �m      �m      On                      �m      �m      On      �n                      �m      �m      �n      �n                      [p      `p      ep      mp      {p      �p      �p      �p                      �p      &q      /q      3q      0�      9�      ?�      D�                      &q      /q      3q      Eq      x�      ��                      �r      �r      �z      �z                      �r      �r      �r      s      $s      0s                      s      $s      0s      Ys      is      us                      Ys      is      us      �s      �s      �s                      �s      �s      �s      �s                      pt      �t      ��      ȃ                      pt      �t      ��      ��                      �t      �t      ��      ȃ                      �t      �t       u      �u      �      �                       u      �u      �u      �u                      �t      �t      �~      �      a�      e�      �      �      �      0�                      �t      �t      a�      e�      �      �                      �~      J      W      �      �      0�                      �u      dv      pv      �v                      �v      �w      �      �      X�      _�                      Ey      �y      �y      (z                      Ey      Qy      Uy      ]y      my      wy      �y      �y      �y      �y      �y      �y                      ]y      my      �y      �y      �y      �y      �y      �y      �y      �y                      (z      �z      <�      :�      @�      J�      ^�      c�                      <�      1�      @�      J�                      A�      E�      K�      O�      V�      Z�      ^�      ^�                      E�      K�      ��      �      @�      J�                      ��      ƈ      Ɉ      ۈ                      �      �      @�      J�                      �z      �z      X~      �~      �      a�      X�      p�      �      a�      _�      ȇ      �      .�      �      D�      ��      �                      �z      �z      
�      �      ��      ��      ��      '�                      !�      !�      ِ      �                      5�      y�      ��      ��                      P�      W�      Z�      h�      k�      q�                      ��      ِ      �      ��      ��      ��      �      ��                      �      t�      �      ��                      �      #�      '�      9�                      E�      t�      �      ��                      #�      #�      2�      >�                      #�      2�      J�      T�      \�      d�                      X~      �~      ��      n�      ��      ȍ                      ��      ׌      ݌      �      �      �      ��      ȍ                      ��      �      �      �       �       �      ��      ��                      �      0�      X�      p�                      ��      �      (�      3�                      �      .�      �      �                      �      .�      �      �                      ��      ��      �      �      �      �                      "�      ��      ��      ��                      ĕ      �      �      C�      G�      ��                      ��      ��      ��      �                      }�      ��      ��      ǘ                      ƙ      ޙ      =�      G�                      ��      '�      G�      [�                      ��      ��      ��      ��      ��      ՛                      G{      G{      \{      h{                      G{      L{      P{      \{      t{      �{                      �{      �{      �{      |                      H|      �|      M}      U}                      L|      W|      Z|      \|                      p|      �|      �|      �|      �|      �|                      �      ��      ��      2�      7�      D�      ��      ��      e�      ��                      �      9�      <�      H�                      �      �      �      0�                      ��      ��      ��      ��      ��      ��      e�      ��                      �      �      Q�      X�      ��      <�                      �      $�      $�      '�                      ��      ��      a�      ��                      Ƃ      ؂      a�      ��                      �      �      �      0�                      Y�      ��      J�      ]�                      b�      z�      J�      ]�                      ��      Q�      ��      �      .�      ;�                      ��      ��      �      �                      ��      Æ      ȉ      �                      Æ      ܆      ��      ȉ                      ܆      �      ��      ��                      ;�      L�      L�      L�                      �      ��      D�      ^�                      D�      L�      Q�      t�                      ^�      b�      i�      m�      t�      
�      
�      &�      &�      h�      h�      ��      ��      ]�      ]�      ��      ��      `�      �      ��      ��      ��      ��      *�                      ��      ��      ��      ��      ̜      �      ��      ѡ                      n�      ��      (�      8�       �      *�                      ��      
�      
�      &�      &�      ��      �      h�      h�      ��      ��      ]�      ]�      ]�      ��      `�      �      ��      ��      (�      8�      ��      ��      ��      ��      ��      Щ       �                      ɝ      ӝ      ۝      �      �      
�      
�      &�      &�      ��      �      h�      h�      ��      ��      ��      ��      `�      �      ��      �      (�      8�      ��      ��      ��      Щ       �                      &�      &�      &�      =�      x�      (�                      x�      ��      ��      ��                      ؞      ��      �      h�      h�      ��      ��      ��      ��      @�      �      ��      �      x�      8�      ��      ��      ��      Щ       �                      �      
�      �      $�                      ��      ��      ��      ��                      П      �      ��      �                      -�      :�      :�      Y�      `�      ��      �      h�      h�      ��      ��      ��      ��      @�      �      x�      p�      ��      ��      ��                      G�      L�      ��      ��                      ��      ��      Ǡ      Ϡ                      ��      ��      ��      �      8�      @�                      �      �      #�      )�      /�      3�      9�      <�      M�      g�                      ��      ��      ��      ��                      |�      ��      ��      ��      N�      _�      b�      p�                      å      ǥ      ˥      �      ��      �                      W       e       p       }       �       �                       �       �       �       �             Q      R      _      h      t      y      �                      �      g      �      �      g      n                      w      �      �      �      !      $                      �      �      !      #                      �      �      �      �      �      !      $      0                      �            	                            @      j      n      p                                  (      &                             �      (      �                      H      i      (      H      K      O                      w      �      �      �      �      �                      �       �       �      �                      �       J            !                      �      �      �      C      �             p      �                      P      �             +                      `      �             +                      �      P      �      �                                   �      C      �      �                                   �      p      �      �                                   �      _      �      �                                   V      d      h      �                      `      d      h      h      n      �                      �      �      �      �            �                      u	      �	      �	      �	                      u	      y	      �	      �	      �	      �	                      �	      �	      �	      �	      �	      �	      �	      
      
      �
      �
      �
      	      :      I      P      T      V      Z      ]      b      �      �      �      �      �      �      ]                            '      7      t                      ;VF     YF     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     6ZF     YZF     ZZF     uZF     vZF     �ZF     �ZF     �ZF     �ZF     [F     [F     +[F     ,[F     T[F     T[F     �[F     �[F     �[F     �[F     �[F     �[F     �[F     �[F     \F     \F     T\F     T\F     z\F     z\F     �\F     �\F     �\F     �\F     �]F     �]F     [^F     [^F     �^F     �^F     O`F     O`F     w`F     x`F     +aF                     maF     �cF     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     6ZF     YZF     ZZF     uZF     vZF     �ZF     �ZF     �ZF     �ZF     [F     [F     +[F     ,[F     T[F     T[F     �[F     �cF     �cF     �cF     �cF     �cF     �cF     �cF     dF     dF     :dF     �[F     �[F     �[F     �[F     �[F     �[F     �[F     \F     \F     T\F     T\F     z\F     :dF     ndF     ndF     �dF     �dF     �dF     �dF     eF     z\F     �\F     �\F     �\F     eF     FeF     FeF     �eF     �\F     �]F     �]F     [^F     �eF     afF     afF     �fF     [^F     �^F     �fF     RgF     �^F     O`F     RgF     �hF     O`F     w`F     x`F     +aF     �hF     �iF                     y�F     ?�F     E�F     F�F                     ƄF     ��F     ��F     ��F                     �F     ��F     ��F     ��F                     {kF     �}F     �}F     �}F     �}F     k~F     l~F     ;�F     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     <�F     r�F     r�F     ÀF     ÀF     րF     րF     �F     �F     .�F     6ZF     YZF     ZZF     uZF     vZF     �ZF     .�F     {�F     {�F     ǅF     ǅF     �F     �cF     �cF     �cF     �cF     �cF     �cF     dF     :dF     �F     �F     �F     ��F     ��F     ��F     ��F     ��F     ��F     ܉F     ܉F     �F     �F     7�F     �[F     �[F     �[F     �[F     :dF     ndF     ndF     �dF     �dF     eF     7�F     |�F     |�F     �F     �F     ��F     ��F     ��F     eF     FeF     ��F     4�F     4�F     f�F     f�F     ��F     ��F     V�F     V�F     �F     �F     a�F     b�F     x�F     x�F     ��F     F     ��F     ��F     r�F     r�F     ʙF     ʙF     �F     �F     �F     �F     N�F     N�F     �F     �eF     afF     �F     ��F     ��F     ��F     ��F     ��F     ��F     םF     ؝F     9�F     9�F     W�F     X�F     �F     �F     ��F     ��F     `�F     `�F     ��F     ��F     ��F     ��F     ݤF     ݤF     ��F     ��F     3�F     4�F     ��F     ��F     ��F     ��F     ?�F     @�F     ��F     ��F     �F     �F     E�F     F�F     }�F     ~�F     ɮF     ɮF      �F      �F     6�F     6�F     T�F     T�F     ��F     ��F     I�F     I�F     f�F     f�F     ��F     ��F     ͵F     εF     �F     �F     D�F     D�F     Z�F     Z�F     ��F     ��F     ��F     ��F     �F     �F     ��F     ��F     ҿF     ҿF     (�F     (�F     ��F     ��F     �F     �F     ��F     ��F     B�F     B�F     Q�F     Q�F     `�F     `�F      �F      �F     ��F     ��F     ��F     O`F     w`F     �hF     �iF                     ��F     ��F     &YF     �YF     ZF     5ZF     ��F     ��F     ��F     �F     6ZF     YZF     ZZF     uZF     �F     l�F     l�F     ��F     �cF     �cF     �cF     �cF     �cF     �cF     dF     :dF     �[F     �[F     �[F     �[F     :dF     ndF     ndF     �dF     �dF     eF     eF     FeF     �eF     afF                     ��F     '�F     r�F     ÀF     ÀF     րF     րF     �F     �F     .�F     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     <�F     r�F     (�F     R�F     6ZF     YZF     ZZF     uZF     vZF     �ZF     �F     l�F     R�F     ��F     �cF     �cF     �cF     �cF     �cF     �cF     ��F     ��F     ��F     ��F     ��F      �F     dF     :dF      �F     r�F     l�F     ��F     r�F     ��F     ��F     �F     �F     �F     �F     L�F     L�F     ��F     ��F     I�F     J�F     k�F     l�F     ��F     ��F     ��F     ��F     ��F     ��F     �F     �F     M�F     �[F     �[F     �[F     �[F     :dF     ndF     ndF     �dF     M�F     ��F     �dF     eF     ��F     ��F     ��F     ��F     �F     ��F     ��F     ��F     ��F     ��F     ��F     ��F     eF     FeF     ��F     ��F     |�F     �F     ��F     ܉F     �eF     afF     �hF     �iF     ��F     #�F     4�F     f�F     f�F     ��F     ��F     V�F     V�F     �F     �F     a�F     b�F     x�F     x�F     ��F     F     ��F     �F     ��F     FeF     �eF     ��F     ��F     �F     N�F     ��F     ��F     ��F     םF     ؝F     9�F     9�F     W�F     X�F     �F     �F     ��F     ��F     `�F     `�F     ��F     ��F     ��F     ��F     ݤF     ݤF     ��F     ��F     3�F     ��F     r�F     r�F     ʙF     ʙF     �F     �F     �F     N�F     �F     afF     �fF      �F     6�F     6�F     T�F     T�F     ��F     ��F     I�F     I�F     f�F     f�F     ��F     ��F     ͵F     εF     �F     �F     D�F     D�F     Z�F     ��F     ��F     Z�F     ��F     ��F     ��F     4�F     ��F     ��F     ?�F     @�F     ��F     ��F     �F     �F     E�F     F�F     }�F     ~�F     ɮF     �fF     RgF     ��F     �F     �F     ��F     ��F     B�F     B�F     Q�F     Q�F     `�F     ��F     ҿF     ��F     �F     `�F      �F      �F     ��F     �F     ��F     ҿF     (�F     RgF     �hF     ��F     ��F     O`F     w`F                     $�F     �G     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     r�F     ÀF     ÀF     րF     րF     �F     �F     .�F     6ZF     YZF     ZZF     uZF     vZF     �ZF     �G     G     G     ,G     ,G     �G     �cF     �cF     �cF     �cF     �cF     �cF     dF     :dF     �F     ��F     ��F     ��F     ��F     ��F     �G     )G     *G     	G     �ZF     �ZF     �ZF     [F     [F     +[F     T[F     �[F     	G     4G     �F     7�F     4G     \G     ��F     ܉F     \G     �G     �G     �G     �G     �G     �G     G     G     G      G     JG     JG     �G     �G     �G     �[F     �[F     �[F     �[F     �G     �G     �G     �G     �G     �G     �G     
G     :dF     ndF     ndF     �dF     �dF     eF     |�F     �F     �[F     �[F     �[F     \F     T\F     z\F     
G     MG     �F     ��F     NG     pG     pG     �G     �G     �G     �G     G     G     3G     4G     NG     eF     FeF     4�F     f�F     f�F     ��F     ��F     V�F     V�F     �F     �F     a�F     b�F     x�F     x�F     ��F     F     ��F     z\F     �\F     NG     �G     ��F     r�F     r�F     ʙF     ʙF     �F     �F     �F     �F     N�F     N�F     �F     �G     �G     �G     �G     �eF     afF     ��F     ��F     ��F     ��F     ��F     םF     ؝F     9�F     9�F     W�F     X�F     �F     �F     ��F     ��F     `�F     `�F     ��F     ��F     ��F     ��F     ݤF     ݤF     ��F     ��F     3�F     �\F     �]F     �G     ~G     4�F     ��F     ��F     ��F     ��F     ?�F     @�F     ��F     ��F     �F     �F     E�F     F�F     }�F     ~�F     ɮF      �F     6�F     6�F     T�F     T�F     ��F     ��F     I�F     I�F     f�F     f�F     ��F     ��F     ͵F     εF     �F     �F     D�F     D�F     Z�F     Z�F     ��F     ��F     ��F     ~G     G     ��F     �F     �F     ��F     ��F     ҿF     ҿF     (�F     ��F     �F     �F     ��F     ��F     B�F     B�F     Q�F     Q�F     `�F     `�F      �F      �F     ��F     RgF     �hF     G     �G     ��F     ��F     O`F     w`F     �hF     �iF     �G     �G     �G     G                     �6G     17G     67G     77G                     r7G     8G     !8G     "8G                     �8G     l9G     q9G     r9G                     �9G     W:G     \:G     ]:G                     �;G     �;G     ^HG     aHG                     x?G     �AG     >HG     AHG                     �AG     ,BG     AHG     DHG                     ,BG     vCG     DHG     GHG                     vCG     /DG     GHG     JHG                     /DG     �DG     JHG     MHG                     �DG     �FG     MHG     NHG                     HG     >HG     aHG     bHG                     LIG     �IG     VG      VG                     7MG     YOG     �UG      VG                     YOG     �OG      VG     VG                     �OG     5QG     VG     VG                     5QG     �QG     VG     	VG                     �QG     |RG     	VG     VG                     |RG     �TG     VG     VG                     �UG     �UG      VG     !VG                     ߘG     u�G     z�G     ՙG                     ڙG     y�G     ~�G     ٚG                     ޚG     }�G     ��G     ��G                     �G     y�G     ~�G     ٭G                     ޭG     }�G     ��G     ݮG                     �G     ��G     ��G     ��G                     ��G     }�G     ��G     ��G                     ��G     ��G     ��G     ��G                     ��G     ��G     ��G     ��G                     ��G     ��G     ��G     ��G                     ��G     ��G     ��G     ��G                     ��G     ��G     ��G     ��G                     G     3VG     r�F     ÀF     ÀF     րF     րF     �F     �F     .�F     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     <�F     r�F     (�F     R�F     4VG     ZVG     ZVG     �VG     �VG     WG     WG     UWG     VWG     |WG     |WG     �WG     �WG     XG      XG     �XG     �XG     �XG     �XG     YG     YG     _YG     `YG     �YG     �YG     �YG     �YG     �ZG     �ZG     4[G     4[G     �[G     �[G     �[G     6ZF     YZF     ZZF     uZF     �[G     �[G     vZF     �ZF     �F     7�F     �[G     \G     \G     �bG     �bG     
cG     
cG     �iG     	G     4G     �iG      jG      jG     �pG     �F     ��F     ��F     ��F     ��F     ܉F     �cF     �cF     �cF     �cF     �cF     �cF     ��F      �F     dF     :dF     �pG     �pG     �pG     �wG     �[F     �[F     �[F     �[F     �wG     �wG     �wG     xG     xG     -xG     .xG     |xG     |xG     �xG     �xG     �xG     �xG     �|G     �|G     �|G     �|G     '}G     (}G     ��G      �G     1�G     2�G     [�G     \�G     3�G     �F     ��F     :dF     ndF     ndF     �dF     M�F     ��F     �dF     eF     4�G     e�G     f�G     ��G     ��G     g�G     g�G     c�G     �G     �G     d�G     ��G     ��G     y�G     z�G     S�G     T�G     *�G     *�G     �G     �G     ڔG     ڔG     ��G     ��G     ��G     ��G     ?�G     ?�G     ��G      G     JG     ��G     }�G     ~�G     W�G     X�G     .�G     .�G     �G     �G     ިG     ިG     ��G     ��G     ��G     ��G     C�G     C�G     ��G     ��G     ��G     ��G     [�G     \�G     2�G     2�G     �G     �G     �G     �G     ��G     ��G     ��G     ��G     G�G     G�G     ��G     4�F     f�F     f�F     ��F     x�F     ��F     ��F     r�F     r�F     ʙF     �F     a�F     ʙF     �F     �F     �F     �F     N�F     F     ��F     N�F     �F     eF     FeF     ��F     ��F     ��G     ��G     ��G     _�G     `�G     6�G     6�G     �G     �G     ��G     ��G     ��G     ��G     ��G     ��G     K�G     K�G     ��G     ��G     ��G     ��G     
�G     
�G     T�G     T�G     ��G     �F     l�F     ��F     ��F     ��G     �G     �G     �G     �G     ��G     ��G     �G     �G     c�G     �G     �G     c�G     ��G     ��G     Y�G     Y�G     ��G     ��G     �G     �G     \�G     \�G     ��G     ��G     P�G     P�G     ��G     ��F     ��F     ��F     ��F     ݤF     ��F     4�F     ��F     ��F     ��F     ��F     ?�F     �F     ��F     @�F     ��F     b�F     x�F     ��F     �F     `�F     ��F     ��F     ��F     �F     E�F     ��F     םF     F�F     }�F     ��F     `�F     ��F     ݤF     ��F     3�F     ~�F     ɮF     �eF     afF     �hF     �iF     ��F     #�F     ��G     ��G     ��G     ��G     ��G     ��G     ��G     I�G     I�G     ��G     ��G     ��G     ��G     8�G     8�G     ��G     NG     �G     ��G     ��G     ��G     0�G     0�G     ��G     ��G     w�G     w�G     �G     �G     ��G     ��G     f�G     f�G     �G     D�F     Z�F     ��F     ��F     ��F     �F     �F     ��F     ��F     ҿF     Z�F     ��F     εF     �F     ��F     ͵F     ҿF     (�F      �F     6�F     9�F     W�F     f�F     ��F     6�F     T�F     �F     D�F     FeF     �eF     �G     ��G     ��G     ^�G     ^�G     ��G     ��G     ��G     O`F     w`F     �G     ~G     ��F     ��F     `�F      �F      �F     ��F     Q�F     `�F     B�F     Q�F     I�F     f�F     T�F     ��F     �F     ��F     ��F     B�F     afF     �fF     ~G     G     �fF     RgF     RgF     �hF     G     �G                     �H     H     YF     %YF     H     -H     .H     ZH     ZH     hH     hH     vH     vH     �H     �H     �H     �H     �H     �H     2H     2H     @H     @H     RH     RH     wH     xH     �H     �H     
H     
H     $H     $H     HH     HH     H     H     �H     �H     �H     �H     �H     �H     �H                     1H     \H     �H     �H                     �H     �H     �H     �H     �H     H     H     $H     $H     5H     6H     �H     �H     <H     <H     sH     tH     �H     �H     �H     �H     H     H     aH     bH     vH     vH     �H     �H     �H     �H     H     H     -H     .H     MH     NH     mH                     nH     �'H     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     6ZF     YZF     ZZF     uZF     vZF     �ZF     �cF     �cF     �cF     �cF     �cF     �cF     dF     :dF     �cF     dF     �[F     �[F     �[F     �[F     :dF     ndF     ndF     �dF     �dF     eF     �dF     �dF     eF     FeF     FeF     �eF     �eF     afF     afF     �fF     �fF     RgF     RgF     �hF     O`F     w`F     �hF     �iF                     �'H     $)H     YF     %YF     &YF     �YF     �YF     ZF     ZF     5ZF     <�F     r�F     6ZF     YZF     ZZF     uZF     vZF     �ZF     �ZF     �ZF     �ZF     [F     [F     +[F     $)H     M)H     T[F     �[F     �[F     �[F     �[F     �[F     �[F     �[F     �[F     \F     M)H     �)H     T\F     z\F     z\F     �\F     �)H     *H     �\F     �]F     *H     �*H     �*H     +H     +H     �,H     O`F     w`F     x`F     +aF                                                    � @                    @                   �,H                    -H                   �J                    �K                    �K                   �K                  	 (�K                  
 8�K                   ��K                    �K                                                                                                                                                                                                                                             ��                     �K                 	 (�K             (     �J             ;     0@             =     `@             P     �@             f      �K            u     (�K            �     0@             �     @�K     0           ��                �      �K             �     `�K             �     �,H             �    ��                �    ��                     #@                ��                $    �@     >       T    �@            m   ��                v    �-H     �       �   ��                ��    `@     1       �
   �@     H       �    �@            �     @     k       �    p@     X       �    �@     z       �    P@     /       �    �@     �           0@                P@     #       ,    �@     �       I     0H     �       ^    `@     �       }    ` @     \       �    � @     7      �     "@     �       �    �"@           �    �#@     �       �    @$@     �           �$@     >       3    %@     u      V    �&@     <       m    �&@     �       �    p'@     (       �    �'@     -       �    �'@     m       �    �3@     #       �    07@     }       �     ;@               pQ@     \       +    �0H     �       B    Ђ@     y      f    P�@     &       �    ��@     &       �    P�@     �       �     �@     D       �    p�@     D       �    ��@     �       �    P�@     �           ��@     �       A    P�@     �       ^    �@     �       y    ��@     �       �    ��@           �    p�@     >      �    P�@     �      �     �@           �    ��@     F      �     �@     C	         ��                   ��                %   ��                0    ��@     3       ?     �@     �       ]    ��@     �       r    `�@     �       �    @�@     �      �    ��@            �    �@            �     �@            �    0�@            �    @�@            �    P�@     G       �    ��@     M       �    ��@            
     �@                �@     (       (    @�@     \      ;    ��@     8       6    ��@     8       C     �@            M    0�@            W    @�@     �      e     �@     +      q    `�@     �       �    �@     �       �     >H            �    ��@     �      �    ��@     �      �    `�@     !       �    ��@     
       �    ��@            �    ��@     �       �    ��@     )      �    ��@     S       
    0�@            !    P�@           4    P�@     �      O     �@           V    0�@     �       f    ��@     �       x    `�@     �       �    P�@            �    p�@     �       �    P�@     	      �    `�@     W       �    ��@     T      �     �@     �      �     �@     Y      	    `�@     R       	    ��@     	       0	    ��@     �      H	    ��@     X      `	     �@     �       n	    ��@     -       �	    ��@     0       �	    ��@     9       �	     �@     &       �	    P�@     �      �	    A            �	     A           �	    @A     �      �	    �	A     �       
    �
A           !
    �A     
      B
     A     4      Z
    @A     /       j
    pA     |       z
    �A     �       �
    �A           �
    �A     f       �
    PA     ]       �
    �A     �       �
    �A     7       �
    �A     <       �
     A     :           @A     7           �A     7       *    �A     R       6     A     U       E    �A     �       N    A     �       ]    �A     �      n    �A     �      �    P!A     �      �    �-A     �      �    pCA     �      �    `EA     �      �     GA                @JA     �           0KA     �      -     MA     ?      ;     7H     $       L     7H             a    @XA     �      q    �6H     $       �    �`A     c      �    `cA     �       �    `dA           �    peA           �    �fA     7       �    �fA     l      �    0jA               PkA     
           `kA            (    pkA     k      6    �lA     �
      C    @<H     �      T    `7H     �      a    pwA     b       r    @AH     p       ~    �wA     ~       �    `xA     R       �    �xA     �       �     ?H            �    ��A     �      �    P�A     �      �    @�A     �       �     BH     P           �AH     @       &    �AH            A    �AH            Z    PBH            p   ��                HA    @�A     )       x    p�A            �    ��A     1       �    ��A            �    ��A            �    ��A     �       �    ��A     n       �    �A                0�A                @�A     �            ��A            2    ��A     x       A    p�A            P    ��A     M       b    ��A           �    ��A     Q       �    @�A           �    `�A     T      �    ��A     �      �    p�A           �    ��A     �      �    @�A               P�A     P       %    ��A           �    ��A     �      3    ��A     �      A    p�A     Q      N    ��A     p       `    @�A     �      k    �FH     �      w    @�A     n       �    ��A     &      �    ��A     �      �    ��A     :      �    ��A     3      �     �A     �       �    ��A     
       �     PH     �       �    ��A     �       �    ��A     J	           ��A     %       S�     �A     �           ��A           #    ��A     �       3    � B     �       E    `B     �      S    `B           j    pB     �      {     B     c       �    �B     1       �    �B            �    �B     <       �     B     C       �    pB     H       �    �B     9       �     B     �           �B     Y          B     �       *    �B           7    �B     �      D    PQH            W    `QH            m    �PH     (       �    �PH            �    �PH            �     QH     P       �   ��                �    �B            �    �B     	       �    �B                  B     ;       /    @ B     F       E    @6B            [    � B            w    � B            �    � B     3       �    !B     
       �     !B     !       �    P!B     A       �    �!B     
       �    �!B     
           �!B     
           �!B     
       )    �!B     
       <    �!B     
       M     "B     	       a    "B     
       t     "B            �     TH            �    @"B     �       �     #B     
       �    0#B            �    P#B            �    `#B     x       �    �#B                �#B     (            $B     �       +    �$B     T       9    @%B     �      O    �&B     Q       ^    0'B     ~       p    �'B     o       �     (B     �      �     dH     P       �     ,B     
      �    0-B     �       �     .B     ;       �    `.B     �      �    01B               @5B     �           �5B     K       6    `6B     �       B    7B     &      W    @8B            m    `9B     D       �    �9B     �       �    �:B     �       �    @;B     D      �    �<B     >      �    �=B     Q       �    0>B     �          0@B     �           �@B     �      $    �BB     Z       7    �BB     W       K    PCB     �
      Y    0NB     V       h    �NB     �      y    @PB     �       �    �PB     �      �    pSB     �       �    �cH     P       �    TB     �       �    �TB     g       �    0UB     �      �     ZH     �	          �XB     �      $    @[B     G       6    �[B     7       I    �[B     b       [    @\B     q       u    �\B     r       �    @]B     ^      �    �`B     U      �     dB     Y       �     eH     �       �    `dB     �       �     eB     �      �     iB     E&          �QH                 XH     �      /     RH            C    �VH     L      V     VH     �       o    `fH     P       �     fH     @       �     gH     (       �    �fH            �    0gH            �    �fH                �fH                �fH            -    �eH     (       B   ��                M    p�B     K       d    ��B            r    ЏB     x       �    P�B            �    `�B            �    ��B     1       �    ��B            �    АB     .       �     �B            �    �B     
            �B     M           p�B     �      *    @�B     u      >    ��B     �      L    ��B     c      b     �B     �       q    �B     
       �    �iH     `       �     �B     <       �    `�B     4       �    ��B     Y       �     �B     9       �    @�B     �      �    �jH     �	      �    �jH                �jH     (       '    PjH            <    @jH            S   ��                Y     �B     V       g    ��B            u    ��B     h       �     �B     �       �    ��B     5       �    �B     #      �     �B     �       �     �B     �           ��B     �           0�B     H           ��B     �      >    P�B     u       Z    оB     �       l    ��B     
       |    �vH     0       �    пB     �       �    p�B     �       �     �B     t       �    ��B     q       �     �B     2      �    `�B               ��B     �          0�B     B          @uH     t       0    �tH     P       I    �vH            a   ��                j    ��B                ��B     1       �    ��B            �    ��B            �    ��B     �       �    ��B            �    ��B     _       �     �B     _       
    ��B                ��B     Q       0    ��B     6       >    0�B     �      L    �B     /       \    @�B     �       o    ��B     �          ��B           �    ��B     
       �     |H     P       �     �B     %       �    0�B            �    P�B     "      �    ��B     �      �    0�B                PC     6            �C     �      ,     �wH     �      9     �|H            P     �|H            i     `|H     (       }    ��                �     �C             �     �C            �     �C     /       �     �C     �       �     �C     L       �     �C     i      �     PC     l       �     �C     
       !    �}H     0       !    �C     �       .!    pC     �       <!    @~H     �       Q!    @C     k      _!    �}H     P       r!    �H            �!    �H            �!    `H     4       �!    @H             �!     H             �!     H            �!    �~H            "    �C     A       $"    �}H            7"   ��                ="      C            K"      C            Y"    @ C     y       m"    � C     �       �"    �!C            �"    �!C            �"    �!C            �"    �!C            �"    �!C            �"    �!C     N       �"    @"C     �       �"    @#C     =      #    �&C     �       #    0'C     
       1#    ��H     @       >#    @'C     �      S#    �(C            a#     )C     h       z#    p)C     U       �#    �)C     �       �#    ��H             �#    `�H             �#    @�H            �#    `*C     �      �#    ��H     4       $    ��H     4       $    0,C     �      %$    ��H            4$    ��H            E$     �H            Y$     �H            q$    BC     E      $     �H     P       �$    ��H            �$    ��H            �$   ��                �$    `DC     �       �$    `�H             �$    ��H     �       �$    @EC     �       �$     FC            �$     FC             �$    @FC            %    `FC     y       %    �FC     �       *%    �GC            =%    �GC     G       M%     HC     �      \%    �IC     �       m%    PJC     )       |%    �JC     �       �%    KC     
       �%    ��H     0       �%     KC     y       �%    �KC     g       �%    LC     �       �%    �LC     �      �%    `OC     �       &    @PC     '      &     �H            &    pSC     4       :&    �SC     �       O&    pTC     �      h&     �H     �      x&    `ZC     4      �&    �pC     �      �&    ��H     P       �&    �kC     �       �&    0lC     I       �&    �lC     d      �&    �yC     I      '    @�H             '    0�H            '    ЇH            +'   ��                2'     �C     �       A'    ��C     "       T'    ��H            `'    ��C            u'    ��C     �       �'    ��C            �'    ��C            �'    ��C            �'    ��C     3       �'     �C     $       �'    P�C     `       �'    ��C     �       (    P�C     R      (    ��C     $       ,(    ��C     (       :(    �C     '      M(    @�C     W      [(    ��C     �      t(    ��C     P      �(    ИC     :       �(    �C     $       �(    @�C     I       �(    ��C     �       �(    `�C     $       �(    ��C     e        )     �C     �       )     �C            %)     �C     3       :)    `�C     �       N)    �C            a)    0�C            p)    P�C     	      )    `�C     !      �)    ��C            �)    ��C            �)    ПC            �)    �C     �       �)    ��C     	      �)    ��C            *    ��C            !*    СC     !       0*     �C            E*    �C     	       Y*     �C            l*    @�C     �       �*    �C     �       �*    ��C     �       �*    @�C     �       �*    ФC     x       �*    P�C     &       +    pD     (       +    ��C            :+    ��C            T+    ��C            e+    ��C           y+    �C     �       �+    ��C     -      �+    ��C     �      �+    P�C     
       �+     �H     `       �+    `�C     E      ,    ��C     /       ,    �C     V       1,    @�C     �      G,    0�C     t       [,    ��C     u       m,    0�C     �      �,    �C     �       �,    ��C     �       �,    p�C     X       �,    йC     �       �,    ��C     �       �,    @�C     P      -    ��C           '-    ��C     �       :-    @�C     B      L-    ��C     �      ]-     �C           s-    0�C     
      �-    @�C     q      �-    ��C     )       �-    ��C     1       �-    0�C     (       �-    `�C     -      �-    ��C     J      �-    ��C     �       �-    ��C     )      .    ��C     
       /.    ��C     �      A.    ��C     J       S.    @�H     D       d.     �C     Z      v.     �H            �.    �H            �.    �H            �.    ��C     J       �.    ��H     ,       �.    ��C     �       �.    ��H            /    `�H     <       /    ��C     t       //     �H     L       J/    @�C     (      e/    p�C     K      �/    ��C           �/    @�H     P       �/    ��C     �      �/    `�H     �       �/    ��C     v      �/     �C     	      �/    �C     �       �/     �C     �      0    ��C     �       #0    p�C     j      60    ��C     2      I0      D           \0    @D     V       l0    �D     U       0     D     ?       �0    @D     ?       �0    �D     \       �0    �D     n      �0    PD     Q      �0    �D     &       �0    �D     �       1    �D     r        1     D     �      61     �H            O1     �H            k1    �D     B       �1    ��H     T       �1    @D            �1    PD            �1    `D     �       �1     �H     �       �1    ��H            �1    ��H            2    ��H            $2    `D     (      32     �H     <       K2    @�H            b2    �$D     �       t2    P%D     +      �2    �)D     
      �2    ��H            �2     �H     �       �2    ��H            �2    x�H            �2    ��H            �2    `�H            3    p�H            %3   ��                /3    �3D     �      K3    P5D            f3    p5D     �      �3    7D     �       �3    �7D     w       �3    �7D     w       �3    @8D     3       �3    �8D            �3    �8D            4    �8D             4    �8D     �      =4    p:D     �       Q4    @;D     H       d4    �;D            w4    �;D     �      �4    �H            �4    p=D     m      �4    �ED     �	      �4    �OD     8      �4    �QD     �      5    �TD     �      .5    �VD     C       C5    �VD            Z5    �VD     5      w5     \D     U      �5    �`D     <       �5    �`D     "      �5    �aD     }       �5    pbD     
       �5    ��H             �5    �bD     �      6    @dD     \      $6    �fD     Q       ?6     gD           b6    jD     I       }6    `jD     K       �6    �jD     �      �6    prD           �6    �sD     P      �6    �vD     �      
7    �yD     ?      7    �|D     �      77    ��D     f       T7    �D     �      d7    ��D     4      t7    0�D     �      �7    �D     �      �7    ��D            �7    ��D     =      �7    �D     Z      �7    P�D     �      8    @�D     �       )8    0�D     g       =8    ��D     l       S8    �D     Z      p8    p�D     �      �8    @�D     M      �8    ��H            �8   ��                �8    ��D     �       �8    p�D     �       �8    @�D     �      9    �D            #9     �D            99    0�D            O9    @�D     9       ]9    ��D     9       k9    ��D     �       z9    ��D     �      �9    @�D     Q       �9    0�D     u       �9     �D     V       �9    ��D           �9    P�D     �       �9    `�D     �       �9    @E     �       �9    �E     �       :    ��D     m       #:     �D     �       6:    ��D     C      Z:     �D     �      �:    ��D     #      �:    ��D     �       �:     �D     t       �:    ��D     Q       �:    ��D     �      �:    ��D     �       ;    ��D     �       ;    ��D     O      C;     �D     �      W;    p�D     "      f;    ��D     �      };    � E     �       �;    pE     4      �;    ��H            �;   ��                �;    �E     �       �;    �E     �       �;    pE     �       �;    PE     �       �;    �E     �       <    �E            <    �	E     a       <    @
E     �       <    0E           )<    PE     �       .<     E     B       B<    PE     !      V<    �E     �      j<    @E            ~<    PE            �<    `E     �       �<    �E           �<    E            �<     E            �<    0E            �<    @E     !       =    pE            =    �E            )=    �E     �      1=    `E     +      9=    �E     \      L=    �'E     2      \=    0+E     9       i=    p+E     /       }=    �+E     $      �=    �-E     S       �=   ��                �=    0.E            �=    @.E            �=    P.E     !       �=    �.E            �=    �.E            >    �.E           >    �/E     /       %>     0E     �       6>    �0E     h       O>    ��H     0       ^>     1E     {      q>    �3E     �      �>    6E            �>    �6E     �      �>    @;E     )       �>    p;E     G       �>    �;E     9       �>     <E     �      �>     BE            �>     BE            ?    0BE            #?    @BE     p      <?    �EE     *       J?    �EE           c?     HE     $       q?    0HE     S       �?   ��                �?    �HE     �      �?    `NE     �       �?    �NE     R       �?    @OE     ~       �?    �OE     2      �?     RE     �       �?    �RE            �?    �RE            �?    �RE            @    �RE            @    SE     .      "@    @TE     A      0@    �UE     �      J@    pWE     b      R@    ��H     D       _@    @�H     L       f@     I     x       m@    �I     x       t@     I     |       {@    �I     |       �@     �H            �@     �H            �@    �qE     �      �@    �sE     �      �@    @uE     	       �@   ��                �@    `yE     c       �@    �yE     �       A    `{E     �       A     �E     ,      (A    �~E     L       <A   ��                DA    P�E     )       [A    ��E     f      jA    �I     �       xA    ��E     p       �A    `�E     c       �A    ЇE     �       �A    ��E     c       �A    0�E     $      �A    `�E     /      �A    ��E     	       �A    ��E     �      �A    p�E     �       B    p�E             B    ��E     q      3B    �E     �       BB    ��E            QB    �E             dB    ��E     E      }B    ��E     )       �B    ШE     e      �B    @�E     O      �B    ��E     0       �B    ��E     �       �B    ��E     0        C    �E     H       C    @�E     �       0C    �E     0       @C     �E     P       KC    p�E            VC    ��E             gC    ��E     1       }C    �E     1       �C    0�E     %       �C    `�E            �C    ��E            �C    ��E     d       �C    �E            D     �E     )       D    P�E            1D    `�E            KD    p�E     �      dD    p�E           tD    ��E     �      �D    `�E     �      �D    0�E     f       �D    ��E     q       �D     �E            �D    @�E     (       �D    p�E     �       �D     �E     g       E    ��E     �       E    ��E     �      %E    ��E     �       AE    @�E     Y       SE    ��E     �       hE    0�E           xE    @�E     ]      �E     �E     �       �E    �E     �       �E    ��E     x      �E    @�E     �      �E    жE     �      �E    ��E            �E     �E     x       
F    ��E     $      F    ��E            2F    ��E     T       HF    @�E     J       _F    кE     8      pF    `�E            �F    ��E     d       �F    ��E     J       �F    �E     �       �F    ��E           �F    `!F            G    �E     �       G    �I     P      G    p�E     c       9G    �E     x       MG    `�E     h       dG    пE     {      yG    P�E     �       �G    0�E            �G    P�E     	      �G    `�E     �       �G    `�E     �	      �G    `�E            H    ��E            %H    ��E            ?H    ��E            [H    ��E     2       mH    ��E     5       �H     �E     h       �H    ��E     o       �H     �E     >       �H    @�E     Q       �H    p�E     �       �H    P�E     `      �H    ��E     j       I     �E     i       8I    ��E     �      MI    ��E     �       bI    0�E     �       yI    p�E     6      �I    ��E     �      �I    ��E     '       �I    ��E     '       �I    ��E     <        J     �E     �       J    ��E     F      2J    0�E     '       KJ    @�E     �      hJ     �E     }       �J    ��E            �J    ��E     U       �J     �E     b       �J    p�E     h      �J    ��E     �       �J    ��E     �       	K    @�E     x       K    ��E     X       -K     �E     ;/      DK    @I            WK    I            jK     I            }K    0I            �K    �I     X       �K   ��                �K    �/F     7       �K    �/F     �       �K    P0F     �       �K     1F            �K     1F     #       L    P1F     
       *L    �I             ;L    `1F     �      [L    �2F           lL    4F     �      }L     I     (       �L    @I     U       �L    �I     (       �L    �I     @       �L   ��                �L    �6F     &       �L    �6F     V       
M    @7F            M    P7F            M    `7F            &M   ��                1M   ��                8M   ��                GM   ��                OM   ��                [M   ��                lM     MRF             }M     qRF             �M     �RF             �M     �RF             �M     SF             �M     SF             �M     SF            �M   ��                �M   ��                �M   ��                N   ��                N    J            #N   
 8�K            LN    "J            ]N    �J            �N   ��                N    �J            #N   
 @�K            LN    �J            �N   ��                N    �J            #N   
 H�K            LN    �J            �N   ��                �N   ��                N    �J            #N   
 P�K            LN    J            �N    J            �N    J            O    J            .O    �,J            SO                   sO    H,J            �O    O,J            �O    V,J            �O    `,J            �O    p,J            �O    {,J            �O    �,J            P    �,J            (P    �,J            :P    �,J            MP    �,J            aP    �,J            tP    �,J            �P    �,J            �P    �,J            �P    �,J            �P    �,J     	       �P    �,J     	       �P    �,J            Q    �,J     	       )Q    0,J            RQ    8,J            {Q    @,J            $    Z}F     /       �Q    �}F            �Q   ��                N    �-J            #N   
 X�K            LN    �-J            �Q    �.J            R     /J     	       "R    /J     	       9R     /J     	       PR   ��                �N    0/J            �N    1/J            O    2/J            .O    �DJ            N    �/J            #N   
 `�K            LN    �/J            `R    @�K            �R    ��F     �      �R    `�K             �R    ��K            S    ��F     o       =S    �F     �       `S    ��F     ?      �S    �DJ            �S    �F     r      5T    �DJ            �T    �DJ            �T    �DJ            �T    �DJ            �T   ��                �T   ��                N     EJ            #N   
 h�K            LN    EJ            �N    EJ            �N    EJ            O    EJ            .O    *bJ            �T    mEJ            U    ��K            <U    /bJ            kU    4bJ            �U    :bJ            �U    @bJ            V    ObJ            :V    XbJ            lV    hbJ            �V    xbJ            �V    �bJ            W    �bJ            ;W    �bJ            ~W    ��K     x       �W    @�K     x       �W    ��K     x       �W    *G             X    *G            #X    6G     �       FX    6G     �       iX    8�K            �X    nG     *       �X    �G            �X    �G            $Y    �
G     �       �Y    G     *       �Y    DG            Z    dG            IZ    SG     �       �Z    �
G            /[    EG            $    �G     �       �[    �G            �[   ��                �N    �bJ            �N    �bJ            O    �bJ            .O    ؋J            N    %cJ            #N   
 p�K            LN    7cJ            �[    ��J            �[    O�J            �[    V�J            \    `�J     	       \    p�J            0\    x�J            E\    ��J            [\    ��J            p\    �G     �       �\    ��J            �\    ^!G            �\    r!G     0       �\    �:G     �      �\    �"G     b       ]    Z#G     [       9]    tHG     �      k]    ��J            �]    ЊJ            �]    ؊J     	       �]    �J            �]    ��J     
       �]     �J     	       �]    �J     	       	^     �J            ^    (�J     
       7^    8�J     	       N^    H�J            d^    P�J            y^    X�J     	       �^    h�J            �^    p�J            �^    v�J            �^    }�J            �^    ��J            �^    ��J            _    ��J            "_    ��J            6_    ��J     	       M_    ��J            a_    ��J     	       x_    ��J            �_    ȋJ            �_    ЋJ            �_    ��J     	       �_    �J            �_    ��J            L`    ��J            �`    ��J            a    ��J            da   ��                ua     �J            �a    �J     	       �a    @�K            �a    �J            �a    �J            �a     �J            �a    (�J            	b    0�J            b    8�J            5b    @�J     	       Lb    I�J            ab    P�J            wb    X�J            �b    `�J     	       �b    i�J            �b    p�J            �b    x�J            �b    ��J            �b    ��J            c    ��J            &c    ��J            <c    ��J            Qc    ��J            gc    ��J            }c    ��J            �c    ��J            �c    ǕJ            �c    ΕJ            �c    ՕJ            �c    ��J            8M   ��                �c   ��                �N    �J            �N    �J            O    �J            d    `�K            1d    h�K            Yd    ��K     �      rd    H�K            �d    P�K            �d    X�K            �d    w�J            �d    {�J            e   ��                N    ��J            #N   
 x�K            LN    ��J            )e     �J            pe    ȗJ            �e    `�K            �e    p�K            $f    x�K            `f    "�J            �f    �J            fg    ��J            �g    ��J            xh   ��                N    0�J            #N   
 ��K            LN    B�J            �h    y�K            �h   ��                N    ��J            #N   
 ��K            LN    J            �h    ĝJ            �h    �'H     J        i    ,(H            !i    ��H             ;i    
/G     #       Di    `:@     �       Vi  "  FeF     J       �i    ZkF             �i  "  ��G     �       Ej  "  Q�F            �j    6H     H       �j    -G            �j    p8F            �j    p�H            �j    �H            k    P�@     |       k  "  ��G     �      �k  "  �iG     *       �k    'H     �       �k     @             �k    ��G     S       �k    pNF     o      (l  "  &YF     \       Dl    �H            ]l  "  �G     �       �l    �F     n       �l    ��F     >       m  "  vZF     V       "m  "  C�G     d       �m    �H     �       �m    �I     @       �m  "  �G     2       Rn  "  ��G     �      �n  "  �\F     �        o  "  �[F     4       Co  "  �xG     N       bo  "  [^F     U       �o    ��H     (       �o    �@@     �      �o    *kF             �o    �H     p       	p    @gH     P       $p    `)@     P       .p    ��H            Hp     6@            Zp  "  �cF            �p    �G     #       �p    ��K            �p    PuE           �p    ~H     �       �p    P�H            �p  "  |xG     )       q    @I     h       q    D$G     /       q  "  VWG     &       5q    z@     +       Lq  ! 
 p�K     @       oq     �H             �q    ,H     *      �q    кH            �q    0�H            �q    ��H     h       �q    l	H     3       �q    �OF     (       r    ��K     (       �8   G     �       (r    �H            :r    �K            Ar    U%G     �       Jr  "  6ZF     #       br    ��H     H       xr    ��H            �r    H     /       �r  "  ��G     �       s  "  �F     R       3s    �H            Ls    Y(G     7       Vs    0x@            fs    ��H            s    /@     �       �s    @�F     �      �s  "  ��F            �s  "  �[F     4       �3   t,G     I       3t  "  �G     "       �t  "   �G     1       �t  "  H            u  "  ��F     (       Lu    ��H     (       au    <
G     B       hu  "  ��F     7      Xv    ��H     h       kv    0�@     �       �v  "  R�F     S       �v    �@     �       �v    `V@     �       �v    b
H     @      �v    =H     C       �v    w@     �       w    �?F     �       #w    ��H            5w  "  eF     *       �w    �<@            �w  "  �wG     1       �w  "  �F     �       Wx    p}@     �       lx    pGF     +       x  "  ڔG     �       �x  "  4VG     &       'y  "  .�G     �          EjF     �       �y    �F     T       �y    p�@     q      �y  "  ʙF     D      :z  "  �G     1       �z  "  ��G     �       �z    ��@     1       �z    �Z@     +       ��    �G     �       �z  "  @�F     d       *{    �UF     >       2{    ��@     �       H{  "  �H     =       m{    P�@            ~{  "  �G     �       �{   �H     W       |  "  ��F           �|    ��H     (       �|    0�H            �|    G     4       �|    p�H            �|    @�H     (       �|    ЧH            }  "  ��G     �      u}     a@     =      �}    @�H     )      �}  "  �G     G       �}  "  �F     +        ~    H     2       	~    p�@     �       ~  "  �G     -       2~    ��@     g       �$    �kF     $       ?~    �'H            \~  "  L�F     w       �~    �<@     �       �~    �H            �~    �@H     �       �~  "  ~�F     K       8    ��I           E    ��H            W  "  �cF     )       �   ,G            �  "  ��F            �    �H     (       �    `�H            �    �H            4�     �H     (       I�    ��H     �       c�  "  z�G     �       ��    ��H            ��  "  �[F             �    ��@     x       +�    �F     �       2�  "  ��F     )       u�    0�H            ��    
H     +       ��    ��F     H       ��    ��@            ��  "  |WG     <       Ɓ    �S@     a       ف    p�H            �    �FF     1       �    d�F     S       �    ��H     h       '�  "  �QF            -�     �H     P       G�    ��H            `�  "  ��F            K�     �H     (       `�    y@     }       q�    llF     9       y�     }E     $      ��    ��F     V       |$   ;uF     +       ��    ��H     (       ��    �H     2       ��    �F     S       ��    
�F     S            �H     �      ԃ    йH            �    sF     �       ��     MF     o      !�    @�H     (       6�    �R@     S       P�    �@     F       c�    ��@            ��  "  �F     V      m�    �H            ��    @�H            ��    �U@     6       ��  "  ҿF     V      ��     �H     h       ��  "  �YF     �       ��  "  P�G     W       ��  "  �F     )       B�  "  Y�G     U       ��    �%G     3       ��   �WF     c       ��    @�H            ��  "  [F     )       �  "  8�G     �      F�  "  .�F     M      d�    ��H     (       y�    �>@     �       ��     tF           ��  "  �H             Ɉ    �H     .       ш  "  ܉F     0       �    �H            5�  "  ��F     �      �  "  $)H     )       \   eG     �       `�    ��@     9      {�    Y*G     �       ��    @�H     (       ��    0|E     *       ��  "  z\F     *       �     �H     (       *�    �)G     /       3�    e@     �      F�    ��F     S       P�     �H     h       c�    Pv@     �       s�     4@     w       ��  "  �G     �       �  "  ��G     �       ��     �H     (       ��  "  ~�G     �       �  "  �xG     N       9�    �F     �       c�    0�H            |�  "  b�F            ��    ��H            ׍    �H            �    ��H     (       ��    �s@     �      �  "  �G     �      P�    �F@     �      _�    0�H            y�    �H            ��    �H            3�    *,G            ��    ��F     �       Ɏ    0J@     3       ێ  "  �H     +       �  "  �G     �       ��    ��H            ��    `�H            ŏ  "  ��G     U       �    ��H     x       �    ��@     o       .�    @�H     (       C�  "  �@     "       �    �iF     Z       `�    LaF     !       z�    0�H            ��     m@     �       ��  "  �@     I       ��  "  ��F     �        �    �G           �    �K             �  ! 
 0�K     @       T�    �I             e�    ��H     (       z�  "  �G     #       �    �l@     /        �    ЦH            2�    �I     ��      F�    �G     5       O�    �0G     �       V�    ��H            o�    ��H            ��  "  ÀF            ��    ��H            ��  "  �G            ��  "  �F     7      ��  	 0�K             �    nH            �    ��H     (       )�  "  ��G     W       f�  "  dF     ,       ��     �H     (       Ɣ    �{@     6       ڔ  "  �dF     &       �  "  NG     "       �1   -G     �       ��    0~E     �       ȕ  "  ��G     Y       �  "  HH     7       ,�    ��K            7�    ��H            Q�   EH     g       j�    ��F     V       r�    �=@     �       �    P6@            ��    �H            ��    �(@     \       ��    ~
G     5       ɖ    ��F     Q       і  "  ��F     �      ��    �H     +       �    H�H            ��  "  �G            ��  "  (}G     �      �    ��H     �      ��  "  xH     {       ;�    �F     S       D�  "  ��G     �       ��  "  �H     P       �    �rF     +       ��    P�H            �    �0G            �  "  G            ��     �H     h       ��    ".G     2       ƚ    пH            ߚ    �H     /       �    ��H     (       ��  "  {�F     L      �    p�H            3�    kH     2       :�    ��F     �       W�  "  ��G     �      ��  "  K�G     d       �    �zF     �       	�    G     +       �    ��@            .�    �R@     ;       J�    �P@     �       5�    �rF     *       Y�    ]�F     S       b�    �H            t�  "  �pG     �      ��    @�H     (       ֜  "  H            �    ��K            ��    ��H     �       �    @�H              �  "  ��G     �      b�    ��H     (       w�     �H     @       ��    s$G     �       ��    �mF     +       ��    t�F     u       ֝    P�H            �  "  \�G     �       l�  "  G     *       ��  "  �[G     O       Ϟ    ��H     (       �    �y@            �    0�F            
�    @[@     �       �    �H     3       '�    @(@            3�  "   G     *       z�    ��H            ��     j@     �       ��    nF     G      ��     �@            ��   ��K             ğ    �H            ݟ  "  �[G            ��    �H            �     �H            !�    �H            ;�    ��H             U�  "  tH     -       ��    =	H     /       (3   ?)G     x       ��    ��H     (       ��  "  �G     (       O�  "  NH            k�  "  VWG     &       ��  "  ��G     �      �    Px@     B       ��    �rF     +       �    f�F     ?       "�    �y@     h       4�    )�F     V       <�  "  �|G     1       f�  "  G     *       ��                  ��  "  �H     =       ݢ    JxF     .       �    ��@     6      �   WF     6       �  "  ZVG     H       (�    �yF     3       1�    ��H            C�  "  �@     "       `�    �@     �      z�  "  $H     $       �  "  vZF     V       4�     GF     '       G�     �H            Y�  "  �ZF            ��    ��H             ��  "  RgF     �      �  "  @     �       =�  "  *G     �      ݥ    �QF            ��    �5G            �    ��H            !�    0�H            :�    +�F     V       B�    �)G     /       J�    �2@     D       `�    �N@     c       r�    �F     /       ��    ��H            ��    �H            Ǧ  "  ɮF     W       ,�    �H     7       4�    �G            ;�    �uH     �       L�    Е@     �      ]�    ��@     |       s�  "  �G            ��    `dH     �       ̧    �X@            �  "  �F            ��    `OH     �       �  ! 
 ��K     P       $�  "  �G            ¨    ��H            Ԩ  "  
G     C       '�  "  YG     S       F�  "  
cG     �      ��    JH     �       ��  "  ��F     1       ��     �@     �      ��  "  �F     O       ߪ    ��H     (       �    �GF     ,       �    xxF     =      �    �H            2�  "  \�G     �       o�    I�F     �       v�  "  ��F     C       ī    ��H     8       ֫    0�H            �    �H     3       ��    p(@            �  "  \�G     �      V�  "   RF            ]�  "  WG     M       |�    P�H            ��    P|@     (       ��     �H     h       ��    ��H            Ь  "  *H     �       L�    �(G     7       U�  "  ؝F     a      ?�    �rF            E�  "  ,G     �      ޮ    �I             �  "  9�F            ϯ    ��F     m       �  "  �F     �      0�    �[@     �      E�    �Q@     g       a�    ��K            f�    ��H            �  "  �F            а    @�H             �    ��K            ��    �qF     #        �  "  �@     "       �  "  .xG     N       2�    �H            L�     �H     (       a�    ��K            d�    PF@     i       w�  "  �[F     E       ͱ    �H     /       ձ    ��H            �  "  x�F     I       .�  "  H     
       ��    ��@     ?       ��    �I@     Q       ��    05G     [       Ȳ    ��H     (       ݲ    }�F     V       �    �/@     �      ��    �I             =    � @             �    �P@     ^       �    ��H     h       /�  " WWF     ;       G�  "  ��F            "�    ��H            4�    �L@     �       F�     �H     (       [�  "  �H            9�    PI@     ~       K�    ��I           X�    �H     �       j�    �m@     �       |�  "  I�F            ]�    �lF     J      d�  "  �G     �       ��  "  �G     "       0�    �X@            @�    F0G     /       H�    ��H     (       ]�    `�K     �	      q�    нH            ��    o@            ��    �H     /       ��    `�H     0       ��    08F     7       η    P�H            �    vF           �    ��F     S       ��    ��H     (       �  "  ��F     1       �     �H           �  "  �eF     �       J�    ��F     �       l�    �D@     �       c    ��K            |�  "  T�G     �       ��    ��K            �    H�K            �  "  �iG     *       B�  "  ?�G     d       ��    �|@            ��    @�H            Һ    �|@            �    �H            ��    ��H            �  "  hH            ]�    /G     �       d�    Щ@     x      �    ��H     �       ��    ��H            ��    `K@     �       ��  "  :@     2       ɻ    0HF     k       �    ��@     f       �  "  ��F            �  "  0�G     �      \�    ]@           x�  "  <H     7       ��  "  r�F     P       	�    �U@     p       �    p�H            0�  "  ��G     �      r�    p7F     �       ��    �H     p       ��  "  2H            ؽ    �QF     (       ��    p�H            �    3H     /       �    мH            @    �qF     V       4�    dRF             J�    �8F            Y�    P�H            k�  "  εF            Z�  "  r�F     X       <�    ��K            F�    ��D     :       Y�    P�H            s�  "  $H     $       �    lF     3       �  "  RH     %       A�  "  l~F     �      U�     W@     �      f�    `�H            w�    ЯH            ��    `�H             ��    �2@     �       ��  "  
�G     J       ��  "  4�G     1       ��    ��H     (       
�  "  �}F             �    �H            7�    �	H     f       ?�    оH            X�    �x@     ^       g�    ��H            ��    {kF     -       ��    p�@     #       ��     �K            �8   �G     �       ��    �+G     P       ��    ��F     S       ��  "   XG     c       ��  "  ��F     *       ��    ��I            �    @)@             �  "  ��F            �    tH     Q       �    pIF     �       9�  "  �G            ��    @�H     @       ��    ��H            �    P�H            "�  "  �F     �      �    �G     ;       
�    ybF           :   -/G     .       �  "  �YG     .       /�    6$H     �       L�     �H     (       a�  "  x`F     �       ��    pJ@     i       ��    �pF     +       ��    @h@     �      ��    `�H     @       ��  "  �ZF     )       #�    pyA     :0      -�    $G     /       5�    `�H     0       O�    0�H            h�    ��@     F       s�    ps@            ��     �K     (       ��  "  .H            ��     �H     (       ��  "  ��F     7      ��  "  6�G     �       >�   EWF            Z�  "  ��G     �      ��  "  6H     �      ��     �H     (       ��    P�H            �    �H            �    �@     6       .�    �n@     F       Ms    i'G     x       D�    �{@     4       [�  "  �ZG     L       w�    �|H     �       ��    B�F     �       ��    �RF             ��     E     �      ��    �8F            ��  "  ��G     �      "�    ��H     (       7�  "  �bG     *       r�    ��H     (       ��    �G     r       ��  "  .xG     N       ��  "  �H     K      �  "  ��F     C       f�    ��H            �    0�@     �      ��  "  .H     ,       ��    ��H            ��    ��@            ��    P�H            
�  "  �G            ?�  "  �[F            f�  "  �H            :�    �2G     6       C�     �@     9      T�    8G     U       t�    �gH     P       ��    ��H            ��    �@     3       ��    |�F           ��  ! 
 ��K     P       ��    <H     /       �    p�H            �    �J     p      2�    �Z@     C       N�    0SF     R      8�    ��G     Y       i�    ��H     (       ~�  "  ��F     �       d�  "  �ZF            ��    �H            ��    @I     H       ��    �D            ��    @�@     !       ��    �|@            �    �K            �    �N@     �       !�  "  �WG     g       ?�  "  :@     2       S�    ��H            e�    P�H            ~�    ��H            ��     �@            ��    ,aF            ��    P�H            ��  "  �G     �      �    лH            ,�    X#H     �       I�    p6@     A       X�  "  b�F            ��    p�H            ��  "  �H            ��    ��A     �       ��    `s@            �&     @     &       ��    ��F            �  "  ZH            B�    �0G            I�     �H     (       ^�    yH     �       e�    ��H     8       w�    �`@     f       ��  "  +H     �      ��  "  @�F     d       :�    p�H            Q�    �pF            S�   F(H     f       f�     k@     F       s�  "  ��F     N       ��    аH            ��     I            ��    иH            �  "  ��F     �       t�  "  �[G     *       ��     ~@     $      ��  "  c�G     W       �  "  G     �      p�    �|@     .       ��  "  �H            c�    ��F     .       l�  "  (�F     �      ��     �G     %       ��     �H            ��    ��H            	�    ��F     h       >�    -�F     V       F�    @�H     (       [�  "  �H            ��  "  �pG     *       ��    E�G     �       ��    P�H            ��  "  �@     �       ��  "  �H     $       ��  "  ǅF           ��    @T@     6       ��    `5@     !       ��    ��H     (       ��    ��K            ��    0
H     2       �    ��H             �  "  RF            (�    �HF     �       C�    @?@     ^      U�    ��G     �       ]�    �O@     �       �l    ��F     �      p�  "  @H            ��    �n@            ��  "  �H     $       Q�    ��K            o�     �H     @       ��  "  �G     W       ��    �G     E       ��  "  F     �       ��    0@     &       ��  "  T�G     W       ��  "  ��G     Y       �  "  �H            ��    �4G     [       ��  "  4[G     S       �  "  �pG     *       ?�    ��F     J       G�  "  g�G     �       &�    �{F     �       i�    @z@     1      ~�  "  4�F     2       ��    (�K            ��    ��F     *       ��  "  �G     -       ��    �E@     �       ��    �(@     V       ��  "  ��G     U       7�    �!H     �       T�    YF            a�    ��H            {�  "  ��F            ��    pKF             ��  "  �F            �  "  ��G     �       ��    p�H            ��  "  �VG     e       ��    <@     �       ��    VH     ,       ��  "  HH     7       �    ��H            2�    DrF     +       �   <�G     r       @�  "  ZZF            X�    ��K            b�  "  ��G     �      ��    ��H     (       ��    �H            ��    uG     �       ��  "  �}F             ��    +@     �      ��    P�@     x       �    ��H            /�    p�H            H�    �WF           ��    �!G     �       j�    �w@            ��    �KF     I      ��    @�@     V       ��    �JF     �       ��    ��F     V       ��    P�H            ��    `�@     V       �  "  �H             /�    �H     /       7�  "  ��F             �    �H     2       (�    0�H            A�    ��G     �       I�  "  V�F     �       %�    �1@            ;�  "  �H            ��  "  pG     0       �    �vH     P       1�    ��H     H       C�    @@F     F       R�    ��H     (       g�    TH     .       n�    Pk@     �       ~�  "  \G     3       �  "  `�F     �      ��    �@            �  "  (�F     *       �    �UF     m       =�  "  l@     -       V�  "  	G     +       p�  "  ZZF            ��    �/G     2       ��  "  \G     �      ��  "  �xG     �      -�  "  Z�F     H       �    ��F     E       J�    ��H     h       ^�  "  ��F     j       @�     �H     (       Z�    @�D     �      '3   �&G     x       p�  "  w�G     �      ��    @:@            ��    ��H            ��    `�H     �      ��    ��@     c      	�    `�H            �     �H     (       0�    �I     P       K�  "  M)H     E       ��    apF     +       ��  "  �\F     J       �  "  �)H     }       ��    P�@     �       ��  "  ��G     �      �     I            �    p�H            0�  "  �XG     6       J�    @I     @       \�    0S@     S       v�    �G     Q      |�     �K             ��    *H     3       ��    �KF            ��  "  J�F     !       �    �)@     Q      �    [/G     *        �    �iF     F        �  "  ��G     W       ^�  "  ��F            C�    pD@     p       R�    
@     �
      W�    ��H     (       l�    ��F            ��    `|E     �       ��    	H     /       ��  "  �bG     *       ��    G     i       ��    @�H     (       ��    �$H     �       �    ��H            6�    0�H            P�    �pF     "       V�    p�H            o�    ��G     3       w�    @�H     (       ��    0�H            ��    ��H            ��     �H     �       ��    ��H            ��  "  �H            ��    'G     3       	�     �K            �    �JF             �  "  րF     B       e�    ��F     �      :�    �-@     !      T�    u0G            ]�    ��H     (       r�    �G     U       ��  "   RF            ��  "  YF            ��    @{H     �       ��    �l@            ��  "  @H            ��    G     �       ��    К@     �      �  "  
H            Y�    \,G            a�  "  �G     �       ��    @�H            ��  "  �G     0       �  "  �F     4       ��  "  �F            ��    ��H            ��     �H     H       ��    P�K            ��    p�@            �  "  
H            X�    �F     V       `�    bH     3       h�     �H            ��  "  .H     ,       ��  "  `�F     (       �    0G     /       �    ��F     V       �  "  6ZF     #       .�  "  ��F            �    !G     +        �    &G     x       �    ��F     V       �     �@     %      3�  "  t@     8       L�    @�H     (       a�  "  t@     8       3   �,G     "       z�    ��D            ��    #H     g       ��     �H            ��  "  �G            ��    �l@            ��  "  ZF            �    0�H            $�  "  ��F     j       �    @�@     .       �    6G     ;      .�  "  T\F     &       o�    ��G     r       v�  "   �F     r       ��  "  vH     P       ��  "  ��G     �       t�    ��@           ��    H     �       ��  "  �[F            ��  "  B�F            4�    �GF     +       I�  "  �H     |       ��  "  �XG     Q       ��    �RF             ��    ��H            ��    `I     P       ��  "  ��G     U       *�  "  ��F     #      k�    @�H     (       ��    �,H             ��  "  f�G     �      ��  "  H            ��  "  7�F     E       3�  "  ��G     �      ��    P@     c       ��  "  ~G     �       �     �H     x       2�    *G     D       8�  "  ��F     �      �3   � G     �       �3   +3G     �           �H            2    p�@     /       @    �H     ]       K    ��H     (       `    ��F     �      �    GlF     %       �    '}F     3       �  "  ��F            Z�    rF     )       w   ��@            �   �H            �   �H     h       �  �(H     .       �   � H     m       � "  �F     R        "  \F     C       U "  �G     a       �   ��H             "  �YG     	       "  �fF     U       �   �4@     Y       �   z4G     [       � "  4G               k�F     S       " "  �@            E   0�H            ^   @�H     (       s "  2�G     )       � "  D�F            ]   zG     x       z   @R@     E       �   �K            � "   jG     �      �   �H             "  X�G     �       �   ��@     O       �   0�H            �   ��H            �   Q�K            �    �H     (       �   P�H            �   �pF     Z        "  �dF     C       Y   ��H            s "  <H     7       �   �H     R       �   �H            �   �6@     d       �   `�@               �X@               �7@     �      6 "  :dF     4       x    �H     �       � "  �wG            �    �H     0       �   P�H            � "  I�G     �      1	 "  `YG     O       Q	 "  *�G     �       �	 "  �H            �	   0�@     �       
   �,G     $       �   �uF     /       
   �5@     [       /
 "  G�G     d       �
   `�@     Z      �
   �5@     #        3   �.G     +       �
 "  ��G     �       7    @H     `       Q "  r�F     Q       t "  �F     �          ��H            2 "  ݤF             "  �YG     .       2   y+G     "       8 "  �XG     6       R   �:F     �      d "  �H     P       � "  �QF            �   P�H            �   pY@     L      �   �5G               ��@     V        "  l�F     %       n   pJF     3       � "  `�G     �        "  f�F     H       �   D,G             "  vH     P       Z "  �|G     )       �   0�@            � "  X�F     �      n   `�H             �   0�H            �   �.G     .       �   V�F     S       �   maF           �   ��I            �   p�H            �    |@            �   ��@     ,       �   ��F     h          nG     I       +    HF     %       N    l@     �       g "  �YF     �       �   0Y@     :       �   �T@     �       �   0o@     *      � "  M�F     I       + "  ^�G     �      m   �.G     /       t "  &YF     \       �   P�@            �   0�H            �    �H     x       � "  �F     L       � "  H     G      {   H8G     ;      �   ��H            �   �H     @       �   ��H            �   !H     3       � "  xG     )       
 "   �F     �      �   �uF     /       � "  4�F     2       ) "  T�F     1          �H     3        "  �H            t   حH            �   @6@            � "  ��G     �          $�F     �       A   '�F     V       I   �@     3      U   ��H     0       o   �H@     �       �  �VF            �   �/G     2       �   �>@     &       �    |@     '       �    �K             � "  afF     �       L   YF            e   �J@     u       w   ��K             | "  vH     X      �  H     :          �8F     �         `xE     �       2 "  l@     -       K   ��K            c "  �G     <      �   �H            �    �D            �   ��H     (       �   ��H     (          �4@     y        "  ��G     �      [   �#G     `       c "  <�F     6       �   �	G     R       � "  r�F     P       � "  4�F     a      �   �H     8       	   ��H     8       # "  r�F     Q       F   LG     3       N "  �F     �      9   ��H     (       N "  ��G     W       �   �5G     D       � "  4G     (       � "  ZF            �   ��H               �H            ( "  ~�F     K       y   �/G     .       �   p�H            �    I     P       �   ��H     (       �   `�@     �       �   ��H            � "  �]F     �       n    `I     H       �    ��H            �  "  G            D!   ��H            V! "  ިG     �       ;�    orF            �! "  �}F     �       �!   p�@     >       �!   D G     �       0"   $�F     �       T"   �H            x" "  ��G     �      �" "  ��G     �      ##   ��F     *       ,#    �H     0       F# "   �F            $   ��H            7$   ЫH            I$   �%H     �       f$   Y@            {$   fuF     +       �$ "  ��F     1       ^% "  ndF     E       �%   @�H     (       �%   �3@            �%  ~H     f       �%   G     2       �% "  ��F           +&   �F     S       M�    �'G     x       4&   ]H     /       ;&   ШH            U& "  JG     G       �&    �H            �& "  tH     -       '   �kF     $       ' "  f�G     )       E'   ��F     K       M'    �H     0       g'    �H     (       |'   �@     �       �'   G@     �      �' "  f�F     '       �'   0L@     �       �'   �5G            �'   ��F     +       ( "  NG     J       x(   @�H     (       �( "  2�G     �       )   0�D            !)   �@F     M      4)   SG            ;)   �:G     2       J) "  T[F     ,       �)   ��H     0       �)   61G     �      �)   PF     �       �) "  $H            * "  �cF     )       N* "  ��G            *   �H     /       �* "  RH     %       �*   0V@     '       �*   H     m       �*   ��@     6      �* "  ��F            �+ "  �^F     �      2, "  6�F            - "  �hF     �       U-   �jF     <       \- "  :dF     4       �- "  �cF     (       �- "  �G     �       c.   ��K            {. "  (�F     *       �.    �H            �.   9�F     Q       �    �(G     x       �.   ��H     0       �. "  H            �.    x@     (       /   �1@     �       /   �kF     $       /   �H           </ "  d�G     ;       T/ "  �G     W       �/ "  �cF            �/   �H     3       �/    �H     x       �/   ��H     (       0    �H             0 "  �@     -      A0   �@     3       X0   `�H            j0   P�@     h       �   �uF     &       q0 "  ��F     �       }$   uF     *       �0 "  ��G     �      1   X H     i       #1  ;VF     6       81   `�@     2       F1   �S@     6       W1 "  xH     {       �1   �+G     %       �1   PGF            �1 "  ��F     O       �1    iH     �       �1  qVF     �       �1 "  O`F     (       2   ��H            '2    �K            02 "  ��F     }       �2   �I     P       �2   �M@     �       �2  �H     a       �2    �H     (       �2 "  �[F            3   �-G     +       &3   6'G     3       /3 "  ��G     J       C3   ��@            V3    y@            d3   @�H     @       ~3    �H     h       �3   �3G     �       �3   @�H     (       �3   ��K            �3   .+G     K       �3   �H     \       �3 "  f�F     '       �3 "  ��F     �       N4 "  �F     I       �4   �H            �4   `(@            �4 "  �*H     W       !5 "  �[G     *       [5 "  0RF            c5   �"H     �       �5   @RF             �5   d&H     �       �5   MqF     U       �5  �(H     J       �5   ^|F     �       �5 "  l�F            �5 "  N�F     �       H6 "  �G     +       ^6   �H            w6   ��@            �6   ��H            �6   0�K            �6   P�@            �6 "  4VG     &       �6 !  `-J             +7 "  F�F     7      8   ��F     E       ?8   wF     1      F8 "  ��F     6       �8 "  ��G     �      �8   z"G     }       �8   `�H     (       9   ��@     	       9   .H     n       9 "  ��F            �9   �PF     �       �9 "  |�F     h      �9 "  ��F     *       :   T.G     .       : "  bH           �:   ��F     �      �: "  ,[F     (       ��    �yF     �       ;   �I            ; "  ��F     0       7;   �H             crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.5415 dtor_idx.5417 frame_dummy object.5427 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux graphics.cpp /home/computerfido/.local/share/lemon/sysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_keymap_us ftinit.c ft_default_modules ftbase.c hash_num_compare hash_bucket destroy_size find_unicode_charmap memory_stream_close ft_recompute_scaled_metrics ft_raccess_sort_ref_by_id hash_str_compare ft_trig_pseudo_rotate.isra.2 ft_trig_arctan_table ft_trig_pseudo_polarize.isra.3 ft_trig_prenorm.isra.4 ft_property_do _ft_face_scale_advances.isra.6.part.7 FT_Match_Size.part.8 FT_Outline_Get_CBox.part.13 FT_Vector_Transform.part.14 FT_Outline_Transform.part.15 FT_Outline_Get_Orientation.part.16 FT_Vector_Unit.part.18 destroy_charmaps.part.22 FT_List_Add.part.24 FT_List_Remove.part.25 FT_List_Finalize.part.27 FT_GlyphLoader_Done.part.19 ft_glyphslot_done destroy_face find_variant_selector_charmap.isra.10 ft_raccess_guess_table raccess_guess_apple_generic.isra.17 raccess_guess_apple_single raccess_guess_apple_double raccess_make_file_name raccess_guess_linux_cap raccess_guess_vfat raccess_guess_darwin_hfsplus raccess_guess_darwin_newvfs raccess_guess_linux_double_from_file_name raccess_guess_linux_netatalk raccess_guess_linux_double raccess_guess_darwin_ufs_export open_face hash_insert IsMacResource open_face_PS_from_sfnt_stream.isra.28 open_face_from_buffer ft_open_face_internal ftfntfmt.c ftlcdfil.c truetype.c tt_get_kerning tt_get_metrics_incr_overrides TT_Load_Glyph_Header tt_loader_set_pp ft_var_get_value_pointer TT_MulFix14_long_long Current_Ppem Read_CVT Write_CVT Move_CVT Direct_Move_X Direct_Move_Y Direct_Move_Orig_X Direct_Move_Orig_Y Round_None SetSuperRound Dual_Project Project_x Project_y Compute_Funcs Direct_Move Direct_Move_Orig SkipCode opcode_length Ins_MIRP Ins_DELTAP tt_size_init tt_driver_init tt_driver_done tt_face_get_location tt_size_reset tt_size_select tt_size_reset_iterator ft_var_apply_tuple Compute_Point_Displacement Ins_IP TT_Done_Context tt_glyphzone_done tt_size_done_bytecode tt_size_done ft_var_done_item_variation_store tt_done_blend Update_Max TT_Load_Context tt_size_run_prep TT_Hint_Glyph TT_Access_Glyph_Frame TT_Forget_Glyph_Frame ft_var_readpackedpoints ft_var_readpackeddeltas Current_Ratio Move_CVT_Stretched Write_CVT_Stretched Read_CVT_Stretched Current_Ppem_Stretched TT_Load_Simple_Glyph tt_slot_init tt_face_done tt_face_vary_cvt tt_face_load_cvt ft_var_load_avar ft_var_load_item_variation_store TT_Load_Composite_Glyph tt_property_get TT_Get_VMetrics tt_get_metrics tt_get_advances tt_get_var_blend Ins_Goto_CodeRange.part.5 Ins_UNKNOWN Round_To_Grid Round_To_Half_Grid Round_Down_To_Grid Round_Up_To_Grid Round_To_Double_Grid Round_Super Round_Super_45 Ins_JMPR Move_Zp2_Point Ins_MDRP.isra.48 tt_delta_interpolate.part.51 TT_Vary_Apply_Glyph_Deltas load_truetype_glyph ft_var_get_item_delta.isra.53 _iup_worker_interpolate.part.54 Ins_IUP tt_size_request ft_var_to_normalized.isra.56 TT_Get_MM_Var fvar_fields.5991 fvaraxis_fields.5992 tt_set_mm_blend gvar_fields.5865 TT_Set_Var_Design TT_Set_Named_Instance TT_Get_Var_Design TT_Get_MM_Blend TT_Set_MM_Blend ft_var_load_hvvar tt_hvadvance_adjust tt_vadvance_adjust tt_hadvance_adjust tt_apply_mvar tt_face_init trick_names.7681 sfnt_id.7710 tt_get_interface tt_services tt_property_set Normalize.isra.65.part.66 Ins_SxVTL Pop_Push_Count tt_loader_init TT_Load_Glyph tt_glyph_load tt_service_gx_multi_masters tt_service_metrics_variations tt_service_truetype_engine tt_service_truetype_glyf tt_service_properties type1.c t1_get_ps_name t1_ps_get_font_info t1_ps_get_font_extra t1_ps_has_glyph_names t1_ps_get_font_private T1_Get_Multi_Master parse_buildchar parse_private read_binary_data T1_GlyphSlot_Done T1_Driver_Init T1_Driver_Done T1_GlyphSlot_Init T1_Parse_Glyph_And_Get_Char_String T1_Parse_Glyph T1_Compute_Max_Advance T1_Get_Advances t1_allocate_blend parse_weight_vector parse_blend_design_positions parse_blend_design_map T1_Done_Metrics T1_Done_Blend T1_Load_Glyph T1_Face_Done t1_get_name_index parse_dict t1_keywords read_pfb_tag parse_blend_axis_types parse_subrs t1_parse_font_matrix mm_axis_unmap t1_services T1_Get_Track_Kerning t1_ps_get_font_value t1_get_glyph_name mm_weights_unmap T1_Get_MM_Blend T1_Get_Var_Design T1_Get_MM_Var t1_set_mm_blend.isra.2 T1_Set_MM_Design T1_Set_Var_Design T1_Set_MM_Blend T1_Reset_MM_Blend T1_Size_Get_Globals_Funcs.isra.4 T1_Size_Request T1_Size_Init T1_Size_Done t1_get_index T1_Read_Metrics check_type1_format T1_Open_Face T1_Face_Init t1_service_ps_name t1_service_glyph_dict t1_service_ps_info t1_service_properties t1_service_kerning t1_service_multi_masters cff.c cff_cmap_encoding_init cff_cmap_encoding_done cff_cmap_encoding_char_index cff_cmap_encoding_char_next cff_cmap_unicode_init cff_sid_to_glyph_name cff_cmap_unicode_char_index cff_cmap_unicode_char_next cff_get_kerning cff_ps_has_glyph_names cff_get_is_cid cff_get_cid_from_glyph_index cff_set_mm_blend cff_get_mm_blend cff_get_mm_var cff_set_var_design cff_get_var_design cff_set_instance cff_hadvance_adjust cff_metrics_adjust cff_get_standard_encoding cff_standard_encoding cff_fd_select_get cff_get_var_blend cff_done_blend cff_slot_done cff_driver_init cff_driver_done cff_cmap_unicode_done cff_vstore_done cff_slot_init cff_make_private_dict cff_index_done cff_get_cmap_info cff_get_ps_name cff_parse_real power_tens cff_get_name_index cff_charset_compute_cids cff_blend_check_vector cff_blend_build_vector cff_index_get_pointers cff_parse_integer cff_index_get_sid_string cff_get_ros cff_ps_get_font_info cff_ps_get_font_extra cff_size_get_globals_funcs.isra.7 cff_size_select cff_size_done cff_size_request cff_size_init cff_index_read_offset.isra.8 cff_index_access_element cff_index_get_name cff_index_init cff_get_glyph_data cff_free_glyph_data cff_slot_load cff_glyph_load cff_get_advances cff_subfont_done.part.12 cff_face_done do_fixed.isra.13 power_ten_limits cff_parse_font_bbox cff_parse_num.isra.16 cff_parser_run cff_field_handlers cff_load_private_dict cff_parse_vsindex cff_parse_maxstack cff_parse_cid_ros cff_parse_multiple_master cff_parse_private_dict cff_parse_blend cff_parse_font_matrix cff_get_interface cff_services cff_get_glyph_name cff_subfont_load cff_face_init cff_header_fields.6955 cff_isoadobe_charset cff_expert_encoding cff_expert_charset cff_expertsubset_charset cff_service_multi_masters cff_service_metrics_variations cff_service_ps_info cff_service_ps_name cff_service_glyph_dict cff_service_get_cmap_info cff_service_cid_info cff_service_properties cff_service_cff_load type1cid.c parse_expansion_factor cid_slot_done cid_driver_init cid_driver_done cid_get_postscript_name cid_ps_get_font_info cid_ps_get_font_extra cid_get_ros cid_get_is_cid cid_get_cid_from_glyph_index cid_slot_init cid_load_glyph cid_slot_load_glyph cid_face_done cid_parse_font_matrix parse_fd_array cid_get_interface cid_services cid_size_get_globals_funcs.isra.0 cid_size_request cid_size_init cid_size_done cid_face_init cid_field_records cid_service_ps_name cid_service_ps_info cid_service_cid_info cid_service_properties pfr.c pfr_cmap_init pfr_cmap_done pfr_cmap_char_index pfr_cmap_char_next pfr_get_advance pfr_face_get_kerning pfr_extra_item_load_stem_snaps pfr_extra_item_load_bitmap_info pfr_slot_done pfr_slot_init pfr_extra_item_load_kerning_pairs pfr_extra_item_load_font_id pfr_aux_name_load pfr_get_service pfr_services pfr_get_metrics pfr_glyph_close_contour.isra.0 pfr_get_kerning pfr_glyph_line_to.isra.3 pfr_glyph_load_rec pfr_slot_load pfr_face_done pfr_face_init pfr_header_fields pfr_phy_font_extra_items pfr_metrics_service_rec type42.c t42_get_ps_font_name t42_ps_get_font_info t42_ps_get_font_extra t42_ps_has_glyph_names t42_ps_get_font_private T42_Driver_Done T42_Size_Select T42_Size_Request T42_GlyphSlot_Done T42_GlyphSlot_Init T42_Size_Init T42_Face_Done T42_Driver_Init t42_get_name_index t42_parse_sfnts t42_parse_font_matrix T42_Get_Interface t42_services t42_get_glyph_name t42_is_space t42_parse_charstrings t42_parse_encoding T42_GlyphSlot_Load T42_Size_Done T42_Face_Init t42_keywords t42_service_glyph_dict t42_service_ps_font_name t42_service_ps_info winfnt.c fnt_cmap_init fnt_cmap_char_index fnt_cmap_char_next winfnt_get_header FNT_Size_Select FNT_Load_Glyph fnt_font_done winfnt_get_service winfnt_services FNT_Size_Request fnt_font_load winfnt_header_fields FNT_Face_Init fnt_cmap_class_rec winmz_header_fields winne_header_fields winpe32_header_fields winpe32_section_fields winpe_rsrc_dir_fields winpe_rsrc_dir_entry_fields winpe_rsrc_data_entry_fields FNT_Face_Done winfnt_service_rec pcf.c pcf_cmap_init pcf_cmap_done pcf_cmap_char_index pcf_cmap_char_next pcf_get_charset_id pcf_property_set pcf_property_get pcf_driver_init pcf_driver_done PCF_Size_Select PCF_Size_Request PCF_Glyph_Load pcf_seek_to_table_type pcf_driver_requester pcf_services PCF_Face_Done.part.0 PCF_Face_Done pcf_find_property.isra.1 pcf_get_bdf_property pcf_get_metric pcf_metric_header pcf_metric_msb_header pcf_compressed_metric_header pcf_get_accel pcf_accel_header pcf_accel_msb_header pcf_load_font pcf_toc_header pcf_table_header pcf_property_header pcf_property_msb_header PCF_Face_Init pcf_cmap_class pcf_service_bdf pcf_service_properties bdf.c _bdf_atol ddigits a2i _bdf_atos by_encoding bdf_cmap_init bdf_cmap_done bdf_cmap_char_index bdf_cmap_char_next bdf_get_charset_id BDF_Size_Select BDF_Glyph_Load _bdf_list_ensure _bdf_list_done _bdf_add_comment bdf_driver_requester bdf_services _bdf_atoul.part.0 _bdf_atous.part.1 BDF_Size_Request bdf_free_font.part.3 BDF_Face_Done _bdf_list_split empty bdf_get_font_property.part.5 bdf_get_bdf_property _bdf_add_property.isra.7 _bdf_properties BDF_Face_Init _bdf_parse_start bdf_cmap_class _bdf_list_join.constprop.11 _bdf_list_shift.constprop.12 _bdf_parse_properties _bdf_parse_glyphs hdigits nibble_mask bdf_service_bdf sfnt.c get_sfnt_table sfnt_is_postscript sfnt_ps_map sfnt_is_alphanumeric sfnt_get_name_id compare_offsets tt_cmap_init tt_cmap0_char_index tt_cmap0_char_next tt_cmap0_get_info tt_cmap2_get_subheader tt_cmap2_char_index tt_cmap2_char_next tt_cmap2_get_info tt_cmap4_init tt_cmap4_set_range tt_cmap4_next tt_cmap4_char_map_linear tt_cmap4_char_map_binary tt_cmap4_char_index tt_cmap4_get_info tt_cmap6_char_index tt_cmap6_char_next tt_cmap6_get_info tt_cmap8_char_index tt_cmap8_char_next tt_cmap8_get_info tt_cmap10_char_index tt_cmap10_char_next tt_cmap10_get_info tt_cmap12_init tt_cmap12_next tt_cmap12_char_map_binary tt_cmap12_char_index tt_cmap12_get_info tt_cmap13_init tt_cmap13_next tt_cmap13_char_map_binary tt_cmap13_char_index tt_cmap13_get_info tt_cmap14_init tt_cmap14_char_index tt_cmap14_char_next tt_cmap14_get_info tt_cmap14_char_map_def_binary tt_cmap14_char_map_nondef_binary tt_cmap14_find_variant tt_cmap14_char_var_index tt_cmap14_char_var_isdefault tt_cmap_unicode_init tt_get_glyph_name tt_cmap_unicode_char_index tt_cmap_unicode_char_next tt_get_cmap_info tt_face_get_kerning tt_sbit_decoder_load_metrics tt_sbit_decoder_load_byte_aligned tt_sbit_decoder_load_bit_aligned sfnt_get_interface sfnt_services tt_face_load_kern tt_face_free_sbit tt_face_goto_table tt_face_find_bdf_prop sfnt_get_charset_id tt_face_load_hmtx tt_face_get_metrics tt_name_ascii_from_other tt_name_ascii_from_utf16 tt_cmap14_ensure tt_cmap14_get_def_chars tt_cmap14_get_nondef_chars tt_cmap14_variant_chars tt_cmap14_char_variants tt_cmap14_variants tt_face_load_gasp tt_face_get_name tt_face_free_ps_names tt_face_free_name sfnt_done_face sfnt_stream_close tt_cmap14_done tt_cmap_unicode_done get_win_string get_apple_string tt_face_load_any tt_face_load_strike_metrics tt_face_set_sbit_strike tt_face_load_sbit tt_face_load_pclt pclt_fields.6515 tt_face_load_name name_table_fields.6457 name_record_fields.6458 langTag_record_fields.6459 tt_face_load_post post_fields.6510 tt_face_load_maxp maxp_fields.6443 maxp_fields_extra.6444 tt_face_load_hhea metrics_header_fields.6550 tt_sbit_decoder_load_image tt_sbit_decoder_load_compound tt_face_build_cmaps tt_cmap_classes sfnt_load_face tt_encodings.5191 tt_cmap2_validate tt_cmap4_validate tt_cmap6_validate tt_cmap8_validate tt_cmap10_validate tt_cmap12_validate tt_cmap13_validate tt_cmap14_validate sfnt_table_info tt_cmap4_char_next tt_cmap12_char_next tt_cmap13_char_next tt_face_load_cmap load_post_names tt_face_get_ps_name.part.8 tt_face_get_ps_name sfnt_get_name_index sfnt_get_glyph_name tt_face_load_font_dir offset_table_fields.6396 table_dir_entry_fields.6379 tt_face_load_generic_header header_fields.6427 tt_face_load_bhed tt_face_load_head tt_face_load_os2 os2_fields.6499 os2_fields_extra1.6500 os2_fields_extra2.6501 os2_fields_extra5.6502 sfnt_init_face woff_header_fields.5225 ttc_header_fields.5258 tt_cmap0_validate tt_face_load_sbit_image sfnt_get_ps_name hexdigits sfnt_interface sfnt_service_sfnt_table sfnt_service_ps_name sfnt_service_glyph_dict sfnt_service_bdf tt_service_get_cmap_info autofit.c af_sort_and_quantize_widths af_cjk_get_standard_widths af_cjk_hints_compute_blue_edges af_cjk_hints_init af_cjk_snap_width af_latin_snap_width af_dummy_hints_init af_indic_hints_init af_indic_get_standard_widths af_latin_get_standard_widths af_latin_hints_link_segments af_latin_hints_init af_autofitter_init af_autofitter_done af_warper_compute_line_best af_warper_weights af_glyph_hints_reload af_latin_hints_compute_segments af_axis_hints_new_edge af_glyph_hints_align_strong_points af_cjk_metrics_scale_dim af_cjk_metrics_scale af_indic_metrics_scale af_latin_hints_compute_edges af_latin_metrics_scale_dim af_latin_metrics_scale af_glyph_hints_done af_face_globals_free af_get_interface af_services af_cjk_compute_stem_width.isra.0 af_hint_normal_stem af_glyph_hints_save.isra.5 af_latin_compute_stem_width.isra.7 af_latin_align_linked_edge af_dummy_hints_apply af_cjk_hints_detect_features af_iup_interp.part.11 af_glyph_hints_align_weak_points af_loader_compute_darkening.isra.15 af_face_globals_new af_autofitter_load_glyph af_property_get_face_globals af_property_get af_property_set af_warper_compute.constprop.22 af_cjk_hints_apply af_indic_hints_apply af_latin_hints_apply af_cjk_metrics_init_widths af_cjk_metrics_init_blues af_cjk_metrics_check_digits.isra.17 af_cjk_metrics_init af_indic_metrics_init af_latin_metrics_init_widths af_latin_metrics_init_blues af_latin_metrics_init af_service_properties pshinter.c psh_hint_table_record psh_globals_scale_widths psh_globals_set_scale pshinter_get_globals_funcs pshinter_get_t1_funcs pshinter_get_t2_funcs t1_hints_open t2_hints_open ps_hinter_init psh_globals_new psh_globals_destroy ps_hints_close t1_hints_stem ps_hints_t1stem3 ps_hints_t1reset t2_hints_stems ps_hints_t2mask ps_hints_t2counter psh_hint_table_done ps_mask_table_done psh_hint_table_activate_mask.isra.3 psh_hint_table_find_strong_points.isra.4 psh_hint_table_init.isra.12 ps_mask_table_alloc ps_mask_ensure.isra.16 ps_mask_set_bit ps_dimension_add_t1stem ps_hints_stem.part.17 ps_mask_table_merge_all psh_blues_set_zones_0.constprop.26 psh_blues_set_zones psh_hint_align ps_hints_apply.part.21 ps_hinter_done ps_dimension_set_mask_bits pshinter_interface raster.c New_Profile End_Profile Insert_Y_Turn Split_Conic Split_Cubic Bezier_Up Bezier_Down Conic_To Cubic_To Sort Vertical_Sweep_Init Vertical_Sweep_Span Vertical_Sweep_Drop Vertical_Sweep_Step Horizontal_Sweep_Init Horizontal_Sweep_Span Horizontal_Sweep_Drop Horizontal_Sweep_Step ft_black_reset ft_black_set_mode ft_raster1_init ft_raster1_set_mode ft_black_done Line_Up Line_To Render_Single_Pass ft_black_render ft_black_new ft_raster1_get_cbox ft_raster1_render ft_raster1_transform smooth.c gray_raster_reset gray_raster_set_mode ft_smooth_init ft_smooth_set_mode gray_raster_done gray_hline ft_smooth_get_cbox gray_record_cell gray_convert_glyph_inner func_interface gray_convert_glyph gray_raster_render gray_set_cell gray_render_line gray_line_to gray_move_to gray_raster_new ft_smooth_render_generic ft_smooth_render ft_smooth_render_lcd ft_smooth_render_lcd_v gray_render_cubic.isra.0 gray_cubic_to gray_render_conic.isra.1 gray_conic_to ft_smooth_transform ftgzip.c huft_build inflate_blocks_reset inflateReset inflateEnd adler32 ft_gzip_stream_close ft_gzip_free zcfree ft_gzip_alloc zcalloc ft_gzip_check_header inflate_flush inflateInit2_.constprop.4 inflate inflate_mask border cpdext cpdist cplext cplens fixed_tl fixed_td ft_gzip_file_fill_output ft_gzip_file_io ft_gzip_stream_io ftlzw.c ft_lzw_check_header ft_lzwstate_get_code ft_lzwstate_stack_grow ft_lzw_stream_io ft_lzw_stream_close psaux.c afm_compare_kern_pairs PS_Conv_Strtol ft_char_table PS_Conv_ToInt skip_literal_string skip_string skip_procedure ps_parser_skip_PS_token ps_parser_skip_spaces ps_parser_to_token ps_parser_to_token_array ps_parser_to_int ps_parser_to_bytes ps_parser_init ps_parser_done ps_parser_to_fixed ps_parser_to_coord_array ps_parser_to_fixed_array ps_parser_load_field ps_parser_load_field_table t1_builder_done t1_builder_close_contour cff_builder_done cff_builder_add_point cff_builder_close_contour ps_builder_done t1_decrypt cff_random t1_cmap_std_done t1_cmap_standard_init t1_cmap_expert_init t1_cmap_custom_init t1_cmap_custom_done t1_cmap_custom_char_index t1_cmap_custom_char_next psaux_get_glyph_name t1_cmap_unicode_init t1_cmap_unicode_char_index t1_cmap_unicode_char_next t1_decoder_parse_metrics cf2_hintmap_map cf2_hintmap_insertHint cf2_glyphpath_computeOffset ps_table_release t1_decoder_done afm_parser_done t1_cmap_unicode_done ps_table_done afm_parser_init ps_table_new ps_table_add cf2_arrstack_setNumElements cf2_arrstack_push t1_builder_add_point PS_Conv_ToFixed ps_tofixedarray ps_builder_init cf2_getSeacComponent cf2_hint_init t1_make_subfont ps_decoder_init t1_builder_add_contour cff_builder_add_contour t1_builder_init t1_builder_check_points t1_builder_add_point1 t1_builder_start_point cff_builder_init cff_check_points cff_builder_add_point1 cff_builder_start_point t1_lookup_glyph_by_stdcharcode_ps t1_decoder_init cf2_decoder_parse_charstrings afm_tokenize afm_key_table afm_stream_skip_spaces.part.0 afm_stream_read_one afm_stream_read_string afm_parser_read_vals ps_builder_close_contour.isra.1 cf2_builder_moveTo cff_decoder_prepare cf2_glyphpath_hintPoint.isra.35 cf2_hintmap_build cf2_buf_readByte.part.39 cf2_stack_pushInt.part.43 cf2_stack_setReal.part.48 cf2_stack_pushFixed.part.44 cf2_stack_pushInt cf2_stack_pushFixed cf2_stack_popFixed cf2_stack_getReal cf2_stack_pop cf2_free_instance cf2_doStems.isra.54 cf2_glyphpath_pushPrevElem cf2_getT1SeacComponent.isra.58 cf2_glyphpath_closeOpenPath.part.60 cf2_glyphpath_lineTo cf2_glyphpath_moveTo cf2_glyphpath_pushMove cf2_glyphpath_curveTo cf2_doFlex t1_builder_check_points.part.61 ps_builder_check_points.isra.63.part.64 ps_builder_add_point1.part.65 ps_builder_start_point.part.66 cf2_builder_cubeTo cff_check_points.part.67 cf2_computeDarkening.part.71 t1_cmap_std_char_index.part.72 t1_cmap_std_char_index t1_cmap_std_char_next afm_parser_next_key.constprop.76 afm_parser_parse cff_decoder_init cf2_hintmask_read cf2_builder_lineTo cf2_stack_popInt cf2_interpT2CharString readFromStack.8234 readFromStack.8241 readFromStack.8239 readFromStack.8236 psaux_interface psnames.c compare_uni_maps ps_unicodes_char_index ps_unicodes_char_next ps_get_macintosh_name ps_get_standard_strings psnames_get_service pscmaps_services ft_get_adobe_glyph_index.part.0 ps_unicode_value ps_unicodes_init ft_extra_glyph_name_offsets ft_extra_glyph_names ft_extra_glyph_unicodes pscmaps_interface ftsystem.c ft_ansi_stream_close ft_ansi_stream_io ft_alloc ft_free ft_realloc ftbitmap.c fb.cpp filesystem.cpp ipc.cpp runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp syscall.c lemon.cpp _ZN3frgL8null_optE _ZN3frg15_to_string_implL12small_digitsE _ZN3frgL6endlogE _ZZN5mlibc17sys_anon_allocateEmPPvE8__func__ debug.cpp ensure.cpp essential.cpp stdlib-stubs.cpp _ZN3frgL9dont_lockE _ZN3frg9_redblack12_GLOBAL__N_1L15enable_checkingE _ZN3frg12_GLOBAL__N_1L15enable_checkingE _ZZN13AllocatorLock4lockEvE8__func__ _ZN12_GLOBAL__N_111mblen_stateE _ZZ6strtolE8__func__ _ZZ6rand_rE8__func__ _ZZ5abortE8__func__ _ZZ13at_quick_exitE8__func__ _ZZ10quick_exitE8__func__ _ZZ6systemE8__func__ _ZZ6mktempE8__func__ _ZZ7bsearchE8__func__ _ZZ3absE8__func__ _ZZ4labsE8__func__ _ZZ5llabsE8__func__ _ZZ4ldivE8__func__ _ZZ5lldivE8__func__ _ZZ5mblenE8__func__ _ZZ6mbtowcE8__func__ _ZZ6wctombE8__func__ _ZZ8mbstowcsE8__func__ _ZZ8wcstombsE8__func__ _ZZ14posix_memalignE8__func__ _ZZ8strtod_lE8__func__ _ZZN5mlibc7strtofpIdEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIfEET_PKcPPcE8__func__ _ZZN5mlibc7strtofpIeEET_PKcPPcE8__func__ _GLOBAL__sub_I_stdlib_stubs.cpp ctype-stubs.cpp _ZZN5mlibc20polymorphic_charcode7promoteEcRjE8__func__ _ZZ8iswctypeE8__func__ _ZZ8towlowerE8__func__ _ZZ8towupperE8__func__ environment.cpp _ZN12_GLOBAL__N_117empty_environmentE _ZN12_GLOBAL__N_118find_environ_indexEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_110get_vectorEvE6vector _ZGVZN12_GLOBAL__N_110get_vectorEvE6vector _ZN12_GLOBAL__N_110get_vectorEv _ZN12_GLOBAL__N_113update_vectorEv _ZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcb _ZZN12_GLOBAL__N_115assign_variableEN3frg17basic_string_viewIcEEPKcbE8__func__ _ZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEE _ZZN12_GLOBAL__N_117unassign_variableEN3frg17basic_string_viewIcEEE8__func__ _ZZ6getenvE8__func__ _ZZ6putenvE8__func__ _ZZ6setenvE8__func__ errno-stubs.cpp file-io.cpp _ZN5mlibc12_GLOBAL__N_1L24globallyDisableBufferingE _ZN5mlibc12_GLOBAL__N_116global_file_listE _ZZN5mlibc13abstract_file4readEPcmPmE8__func__ _ZZN5mlibc13abstract_file5writeEPKcmPmE8__func__ _ZZN5mlibc13abstract_file5ungetEcE8__func__ _ZZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeEE8__func__ _ZZN5mlibc13abstract_file4seekEliE8__func__ _ZZN5mlibc13abstract_file10_init_typeEvE8__func__ _ZZN5mlibc13abstract_file13_init_bufmodeEvE8__func__ _ZZN5mlibc13abstract_file11_write_backEvE8__func__ _ZZN5mlibc13abstract_file6_resetEvE8__func__ _ZZN5mlibc13abstract_file18_ensure_allocationEvE8__func__ _ZZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeEE8__func__ _ZN12_GLOBAL__N_110stdin_fileE _ZN12_GLOBAL__N_111stdout_fileE _ZN12_GLOBAL__N_111stderr_fileE _ZN12_GLOBAL__N_111stdio_guardC2Ev _ZN12_GLOBAL__N_111stdio_guardC1Ev _ZN12_GLOBAL__N_111stdio_guardD2Ev _ZN12_GLOBAL__N_111stdio_guardD1Ev _ZN12_GLOBAL__N_118global_stdio_guardE _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ5fopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ5fopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ5fopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_clES1_ _ZZ6fdopenENUlPN5mlibc13abstract_fileEE_4_FUNES1_ _ZZ6fdopenENKUlPN5mlibc13abstract_fileEE_cvPFvS1_EEv _ZN3frg9constructIN5mlibc7fd_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEJRiZ6fdopenEUlPNS1_13abstract_fileEE_EEEPT_RT0_DpOT1_ _ZSt7forwardIZ5fopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _ZSt7forwardIZ6fdopenEUlPN5mlibc13abstract_fileEE_EOT_RNSt16remove_referenceIS4_E4typeE _GLOBAL__sub_I_file_io.cpp stdio-stubs.cpp _ZZN13ResizePrinter6expandEvE8__func__ _ZZ6removeE8__func__ _ZZ6renameE8__func__ _ZZ8renameatE8__func__ _ZZ7tmpfileE8__func__ _ZZ6tmpnamE8__func__ _ZZ7freopenE8__func__ _ZZ6setbufE8__func__ _ZL9store_intPvjy _ZZ5scanfE8__func__ _ZZ6sscanfENUt_10look_aheadEv _ZZ6sscanfENUt_7consumeEv _Z8do_scanfIZ6sscanfEUt_EiRT_PKcP13__va_list_tag _ZZ7vfscanfENUt_10look_aheadEv _ZZ7vfscanfENUt_7consumeEv _Z8do_scanfIZ7vfscanfEUt_EiRT_PKcP13__va_list_tag _ZZ6vscanfE8__func__ _ZZ7vsscanfE8__func__ _ZZ8fwprintfE8__func__ _ZZ7fwscanfE8__func__ _ZZ9vfwprintfE8__func__ _ZZ8vfwscanfE8__func__ _ZZ8swprintfE8__func__ _ZZ7swscanfE8__func__ _ZZ9vswprintfE8__func__ _ZZ8vswscanfE8__func__ _ZZ7wprintfE8__func__ _ZZ6wscanfE8__func__ _ZZ8vwprintfE8__func__ _ZZ7vwscanfE8__func__ _ZZ5fgetsE8__func__ _ZZ6fgetwcE8__func__ _ZZ6fgetwsE8__func__ _ZZ6fputwcE8__func__ _ZZ6fputwsE8__func__ _ZZ5fwideE8__func__ _ZZ5getwcE8__func__ _ZZ8getwcharE8__func__ _ZZ5putwcE8__func__ _ZZ8putwcharE8__func__ _ZZ7ungetwcE8__func__ _ZZ7fgetposE8__func__ _ZZ7fsetposE8__func__ _ZZ8getdelimE8__func__ _ZZ14fgets_unlockedE8__func__ _ZZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ _ZZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modEE8__func__ string-stubs.cpp _ZZ7strxfrmE8__func__ _ZZ8strtok_rE8__func__ _ZZ6strtokE5saved _ZZ6wcstodE8__func__ _ZZ6wcstofE8__func__ _ZZ7wcstoldE8__func__ _ZZ6wcstolE8__func__ _ZZ7wcstollE8__func__ _ZZ7wcstoulE8__func__ _ZZ8wcstoullE8__func__ _ZZ6wcscpyE8__func__ _ZZ7wcsncpyE8__func__ _ZZ7wmemcpyE8__func__ _ZZ8wmemmoveE8__func__ _ZZ6wcscatE8__func__ _ZZ7wcsncatE8__func__ _ZZ6wcscmpE8__func__ _ZZ7wcscollE8__func__ _ZZ7wcsncmpE8__func__ _ZZ7wcsxfrmE8__func__ _ZZ7wmemcmpE8__func__ _ZZ6wcschrE8__func__ _ZZ7wcscspnE8__func__ _ZZ7wcspbrkE8__func__ _ZZ7wcsrchrE8__func__ _ZZ6wcsspnE8__func__ _ZZ6wcsstrE8__func__ _ZZ6wcstokE8__func__ _ZZ6wcslenE8__func__ _ZZ7wmemsetE8__func__ allocator.cpp _ZZ12getAllocatorvE16virtualAllocator _ZGVZ12getAllocatorvE16virtualAllocator _ZZ12getAllocatorvE4heap _ZGVZ12getAllocatorvE4heap _ZZ12getAllocatorvE9singleton _ZGVZ12getAllocatorvE9singleton _ZZN16VirtualAllocator3mapEmE8__func__ _ZZN16VirtualAllocator5unmapEmmE8__func__ charcode.cpp _ZZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEEE8__func__ _ZZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEEE8__func__ _ZZN5mlibc16current_charcodeEvE15global_charcode _ZGVZN5mlibc16current_charcodeEvE15global_charcode _ZZN5mlibc22platform_wide_charcodeEvE20global_wide_charcode _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstateE8__func__ _ZZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstateE8__func__ charset.cpp _ZZN5mlibc15current_charsetEvE14global_charset guard-abi.cpp _ZN12_GLOBAL__N_15Guard6lockedE _ZN12_GLOBAL__N_15Guard4lockEv _ZN12_GLOBAL__N_15Guard6unlockEv af_mlym_nonbase_uniranges getwchar FT_Done_GlyphSlot _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvjNS_14format_optionsERT_ longjmp _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEEEbPT_ stpcpy putchar FT_Done_Memory af_khms_nonbase_uniranges af_cyrl_titl_style_class FT_Stream_ReadULong _ZN3frg15do_printf_charsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN11PrintfAgentI13BufferPrinterEC1EPS0_PN3frg9va_structE _ZN5mlibc7charset8to_upperEj _Z12GetVideoModev strcpy _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN3frg14format_optionsC2Ev af_osma_dflt_style_class _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN5mlibc13abstract_file4tellEPl unsetenv _ZN3frg8optionalIiEC2ERKS1_ _ZN3frg16do_printf_floatsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN5mlibc7charset8is_alnumEj t1_builder_funcs _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorppEv _ZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEPKc _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC2EPS3_ _ZN3frg8optionalIiEC2IRivEEOT_ _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_iiic af_knda_script_class FT_Request_Metrics setjmp af_latp_uniranges cff_cmap_unicode_class_rec FT_DivFix af_lisu_nonbase_uniranges ft_validator_init _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD2Ev tmpfile mousePos FT_Stream_OpenGzip _ZN5mlibc7charset8is_alphaEj af_tibt_uniranges _ZN3frg8optionalIiEaSES1_ ps_parser_funcs vscanf _ZN13BufferPrinterC1EPc FT_Stream_ReleaseFrame _ZTVN5mlibc20polymorphic_charcodeE af_limb_nonbase_uniranges strtok_r af_mymr_dflt_style_class af_copt_dflt_style_class tt_cmap_unicode_class_rec wcstok _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer af_adlm_uniranges stdout vsprintf _ZN3frg8optionalIiEC2Ev pshinter_module_class af_bamu_uniranges wcstof _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg17basic_string_viewIcEC2EPKc af_grek_sups_style_class vswprintf FT_Stream_Close af_gujr_dflt_style_class FT_Vector_Transform_Scaled _ZN5mlibc13abstract_file4readEPcmPm _ZSt4moveIRPcENSt16remove_referenceIT_E4typeEOS3_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemC1EPS3_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC2Ev _ZN11PrintfAgentI13BufferPrinterEclEPKcm _ZN5mlibc8code_seqIwEcvbEv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE8allocateEm af_sund_script_class ungetc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12insert_rightEPS7_SC_ tt_cmap6_class_rec FT_Stream_ReadUShortLE _ZN3frg17basic_string_viewIcE10find_firstEcm FT_Init_FreeType ft_module_get_service strerror _ZN5mlibc10sys_accessEPKci FT_Raccess_Guess FT_GlyphSlot_Own_Bitmap af_glag_uniranges _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ FT_Reference_Face _ZN11PrintfAgentI13StreamPrinterEclEPKcm _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ FT_Stream_ReadUShort _Z10lemon_readiPvm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN13StreamPrinterC1EP17__mlibc_file_base _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN5mlibc13abstract_file14update_bufmodeENS_11buffer_modeE FT_Get_Sfnt_Name _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE15_construct_slabEi _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10deallocateEPvm _ZN3frg11_fmt_basics9print_intI14LimitedPrinterlEEvRT_T0_iiic ft_mem_qalloc FT_Set_Debug_Hook _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC2Emmi syscall FT_Stream_ReadUOffset _ZN5mlibc20polymorphic_charcodeC1Ebb FT_List_Finalize _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ _ZN5mlibc8sys_openEPKciPi _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvNS_10escape_fmtENS_14format_optionsERT_ af_kali_script_class af_cyrl_subs_style_class fileno_unlocked af_orkh_nonbase_uniranges af_olck_script_class af_nkoo_uniranges _ZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE FT_Load_Glyph af_blue_strings _ZN3frg6formatIcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg3maxImEERKT_S3_S3_ wcstoull FT_Vector_Polarize _ZN5mlibc7fd_fileD1Ev ft_mem_alloc _ZN5mlibc15current_charsetEv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushERKS1_ FT_Done_Face af_cyrl_sups_style_class tt_driver_class _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC1ENS3_10frame_typeEmm ft_mac_names af_cher_uniranges _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EEclEv _ZNK3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4sizeEv af_cyrl_nonbase_uniranges af_osge_uniranges _ZN5mlibc13wide_charcode7promoteEwRj af_tavt_script_class af_latn_nonbase_uniranges _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ af_deva_dflt_style_class _ZN3frg8optionalIiE13storage_unionC2Ev ft_mem_dup getenv _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE4freeEPv af_kali_dflt_style_class wcslen iswcntrl ft_mem_free _ZN13BufferPrinter6appendEc FT_Lookup_Renderer af_taml_dflt_style_class _Z12lemon_map_fbP6FBInfo iswpunct tt_cmap2_class_rec _Znwm af_tibt_nonbase_uniranges af_cakm_dflt_style_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10get_parentEPS7_ af_copt_script_class FT_Stream_ReadAt strtold FT_Stream_OpenLZW isblank af_cyrl_script_class wcstoll iswalpha iswblank af_script_classes af_shaw_dflt_style_class bsearch _Z12DrawGradientiiii10RGBAColourS_P7Surface af_armn_script_class FT_Face_GetVariantsOfChar FT_New_Memory_Face FT_Library_SetLcdFilterWeights _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_insertEPS7_ af_latn_sinf_style_class af_buhd_uniranges FT_Render_Glyph _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_insertEPS7_ tt_cmap12_class_rec _ZN3frg14format_optionsC1ERKS0_ _ZN3frg11_fmt_basics9print_intI13BufferPrinteryEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPvEERS4_T_ _ZN3frg11_fmt_basics9print_intI14LimitedPrinterjEEvRT_T0_iiic vsscanf _ZN5mlibc13sys_clock_getEiPlS0_ af_kali_uniranges _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPKcEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI13StreamPrinteryEEvRT_T0_biiic _ZN5mlibc7strtofpIdEET_PKcPPc af_goth_script_class ft_synthesize_vertical_metrics qsort _ZN5mlibc13utf8_charcode12decode_stateC2Ev wcsrchr _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockE10reallocateEPvm af_mlym_dflt_style_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11rotateRightEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIPvEERS4_T_ FT_GlyphLoader_CheckPoints fgets af_sylo_script_class ft_lzwstate_reset _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKcNS_14format_optionsERT_ af_orkh_script_class vwprintf _Z13AddNewWindowsv iswxdigit tt_cmap4_class_rec ps_property_get FT_GlyphLoader_Prepare _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ af_avst_script_class _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ _ZN3frg8optionalIiEC1IRivEEOT_ _ZN5mlibc13abstract_file13_init_bufmodeEv af_osge_dflt_style_class _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC2Ev af_grek_c2sc_style_class af_armn_uniranges af_lisu_script_class ps_property_set _ZN3frg11_fmt_basics12print_digitsI13ResizePrintermEEvRT_T0_biiic FT_Get_Kerning af_osma_nonbase_uniranges af_hani_nonbase_uniranges af_glag_dflt_style_class _ZN5mlibc13abstract_fileD2Ev FT_Get_Char_Index _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED0Ev _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ af_latn_sups_style_class af_taml_uniranges _ZN3frg11_fmt_basics9print_intI13ResizePrinterjEEvRT_T0_iiic ft_smooth_lcd_renderer_class ft_mem_realloc af_latn_script_class _ZN8ListNodeIP8Window_sEC2Ev _ZN5mlibc9PanicSinkclEPKc af_grek_smcp_style_class FT_Outline_Reverse _ZplRK8Vector2iS1_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14size_to_bucketEm setvbuf __TMC_END__ _ZTVN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEE t1_decoder_funcs af_orya_script_class _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE3endEv FT_Outline_Translate af_sinh_uniranges ft_adobe_glyph_list renameat perror af_sund_dflt_style_class af_none_dflt_style_class _ZN3frg10bitop_implImE3clzEm af_khms_uniranges _ZN3frg16intrusive_traitsIN5mlibc13abstract_fileEPS2_S3_E5decayES3_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_leftEPS7_SC_ __DTOR_END__ _ZN5mlibc7charset17is_ascii_supersetEv af_hebr_script_class _ZN3frg11_fmt_basics9print_intI13ResizePrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsENS_8endlog_tE af_cakm_script_class FT_Stream_ExitFrame _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE5_emitEPKc _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratoreqERKSA_ ft_lzwstate_done _ZN3frg17basic_string_viewIwEC2EPKw _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC2Ev dragOffset af_nkoo_nonbase_uniranges _ZN5mlibc8sys_seekEiliPl islower FT_Done_Size ft_validator_error _ZN5mlibc20polymorphic_charcodeD1Ev FT_MulDiv __fpurge tolower _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E12replace_nodeEPS7_SC_ _ZN5mlibc20polymorphic_charcodeD0Ev af_dsrt_nonbase_uniranges _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC2ES6_ _ZN11PrintfAgentI14LimitedPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE af_blue_stringsets _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC2ERS1_ iswlower _ZN3frg11_fmt_basics9print_intI13ResizePrinterlEEvRT_T0_iiic _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ system af_latn_ordn_style_class feof _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratordeEv tt_cmap14_class_rec fgetws af_cyrl_dflt_style_class wcspbrk af_osma_script_class _ZN5mlibc7strtofpIfEET_PKcPPc af_cyrl_sinf_style_class wcstol _ZN5mlibc13abstract_fileD1Ev _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterjEEvRT_T0_biiic _ZN3frg16do_printf_floatsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE malloc remove FT_GlyphLoader_CheckSubGlyphs FT_Face_GetVariantSelectors FT_Set_Charmap iswspace af_geok_uniranges _ZN3frg13printf_formatI11PrintfAgentI13ResizePrinterEEEvT_PKcPNS_9va_structE af_geok_script_class _ZN13AllocatorLockC2Ev mainFont pcf_driver_class af_lao_nonbase_uniranges _ZN3frg11_fmt_basics12print_digitsI13ResizePrinteryEEvRT_T0_biiic af_cari_script_class af_indic_writing_system_class vsnprintf strtoll _ZN5mlibc13abstract_file18_ensure_allocationEv af_geor_dflt_style_class _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC2Ev _ZN13ResizePrinter6appendEPKcm af_telu_script_class FT_Stream_Read _ZN5mlibc7fd_file2fdEv FT_Get_SubGlyph_Info wcsncmp FT_RoundFix _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIcEERS4_T_ af_sinh_nonbase_uniranges FT_Get_Advance strtoul FT_List_Add __dso_handle af_latn_smcp_style_class _ZN3frg8optionalIiEcvbEv af_cprt_dflt_style_class af_saur_uniranges af_shaw_nonbase_uniranges af_thai_nonbase_uniranges _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED1Ev wcsstr af_beng_script_class _ZNK3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorneERKSA_ _ZN5mlibc8code_seqIKwEcvbEv _ZN13BufferPrinterC2EPc _ZN3frg15do_printf_charsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE FT_Stream_Seek mktemp _ZN5mlibc13abstract_file5purgeEv FT_Stream_TryRead ispunct _ZN11PrintfAgentI14LimitedPrinterEclEPKcm _ZN3frg5_list19intrusive_list_hookIPN5mlibc13abstract_fileES4_EC1Ev __mlibc_errno _ZN5mlibc20polymorphic_charcodeC2Ebb wctomb FT_New_Size _ZN5mlibc12sys_libc_logEPKc _ZN13StreamPrinter6appendEc wcstombs af_sund_uniranges _ZN8ListNodeIP8Window_sEC1Ev FT_Set_Default_Properties _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ _ZN3frg8optionalIiEC1ERKS1_ _Z10lemon_openPKci af_limb_uniranges _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD1Ev af_autofitter_interface _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_biiic _ZN4ListIP8Window_sE8add_backES1_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5eraseENS9_8iteratorE _Z11SendMessagem13ipc_message_t clearerr_unlocked af_hebr_uniranges af_avst_dflt_style_class isspace vwscanf FT_GlyphLoader_Rewind FT_Get_Sfnt_Table _ZN5mlibc13abstract_file7disposeEv af_latn_titl_style_class af_tfng_dflt_style_class _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_iiic mempcpy fflush pfr_driver_class FT_New_GlyphSlot FT_Stream_ReadULongLE _ZSt4moveIRPN5mlibc13abstract_fileEENSt16remove_referenceIT_E4typeEOS5_ cff_driver_class ft_property_string_set _ZN13AllocatorLock6unlockEv t1_driver_class _ZTVN5mlibc7fd_fileE _ZN3frg11compositionINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEE3getEPSA_ af_orkh_uniranges _ZN3frg6formatIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN14LimitedPrinter6appendEPKc _ZN3frg13printf_formatI11PrintfAgentI14LimitedPrinterEEEvT_PKcPNS_9va_structE _ZN5mlibc7charset8is_digitEj _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5isRedEPS7_ FT_GlyphLoader_CopyPoints _ZN3frg11unique_lockI13AllocatorLockE6unlockEv af_lao_script_class _Z10lemon_seekili mbstowcs _ZN5mlibc22platform_wide_charcodeEv _ZN3frg11_fmt_basics9print_intI13BufferPrinterlEEvRT_T0_iiic putenv _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED1Ev af_deva_uniranges af_kali_nonbase_uniranges wmemcpy FT_FloorFix _ZN11PrintfAgentI13BufferPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZdlPv _ZN13StreamPrinter6appendEPKcm af_latb_dflt_style_class FT_Stream_GetUShortLE tt_cmap8_class_rec af_none_uniranges _ZN3frg11_fmt_basics14format_integerImNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ vswscanf _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E16remove_half_leafEPS7_SC_ _Exit _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE9push_backES6_ ps_table_funcs _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11predecessorEPS7_ _ZN5mlibc13abstract_file5ungetEc _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8allocateEm FT_Outline_Decompose FT_Face_GetCharVariantIndex drag af_sinh_dflt_style_class _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4dataEv af_taml_nonbase_uniranges backgroundColor abort _ZN4ListIP8Window_sEixEj _ZN3frg8optionalIiEC2EOi af_ethi_nonbase_uniranges af_guru_script_class fb FT_Set_Pixel_Sizes _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ wcscoll af_beng_uniranges _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frame8containsEPv _ZSt4moveIRN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessEENSt16remove_referenceIT_E4typeEOS8_ FT_Atan2 FT_Get_Charmap_Index ftrylockfile af_none_script_class isxdigit FT_Vector_NormLen t1_cmap_classes FT_Get_CMap_Format tt_cmap10_class_rec _ZN5mlibc10sys_getpidEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_rootEv af_mlym_uniranges FT_Get_Glyph_Name af_glag_script_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC1Ev FT_Select_Charmap ft_sid_names _Z12getAllocatorv FT_Outline_Render _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10get_parentEPS7_ strtol _ZN3frg11_fmt_basics9print_intI13StreamPrinterlEEvRT_T0_iiic _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEEC1Ev FT_Property_Set fsetpos af_cprt_script_class __mlibc_rand_engine af_grek_titl_style_class FT_Outline_Transform wcstod af_hebr_nonbase_uniranges FT_New_Memory af_cyrl_smcp_style_class mblen iswprint af_hani_script_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E7isBlackEPS7_ af_latn_uniranges _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEPKc _ZN5mlibc13abstract_file6_resetEv FT_Request_Size _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ lastKey active _ZN11PrintfAgentI13BufferPrinterEC2EPS0_PN3frg9va_structE _ZN3frg16do_printf_floatsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE FT_Stream_GetULongLE af_osma_uniranges FT_Stream_GetULong af_goth_dflt_style_class af_cyrl_ordn_style_class _ZSt7forwardIR16VirtualAllocatorEOT_RNSt16remove_referenceIS2_E4typeE rename FT_Raccess_Get_DataOffsets bdf_driver_class af_copt_uniranges FT_Face_Properties _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm FT_New_Library _ZNK3frg17basic_string_viewIcE4dataEv _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterjEEvRT_T0_biiic _Z22RemoveDestroyedWindowsv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC2Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC1ES5_ FT_Get_Module af_latn_c2sc_style_class _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterjEEvRT_T0_biiic FT_Stream_Open strrchr _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3getEv _Z14ReceiveMessageP13ipc_message_t af_cari_dflt_style_class wcscpy af_knda_dflt_style_class memcpy_sse2_unaligned FT_Bitmap_Init af_dsrt_uniranges _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_nodeEPS7_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E5firstEv mouseData af_shaper_get_elem af_tfng_nonbase_uniranges _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ strtod _ZN3frg15aligned_storageILm456ELm8EEC1Ev _ZN3frg7mt19937clEv FT_Remove_Module af_lao_uniranges af_cans_nonbase_uniranges af_latb_uniranges FT_GlyphLoader_Reset _ZSt4swapIbEvRT_S1_ _ZN11PrintfAgentI13ResizePrinterEclEPKcm af_tfng_script_class _ZN3frg7mt19937C2Ev af_khms_dflt_style_class wmemchr af_grek_c2cp_style_class FT_Stream_Skip af_adlm_dflt_style_class atof FT_Get_Font_Format environ fputs_unlocked iswgraph _ZN13BufferPrinter6appendEPKcm _ZN3frg17basic_string_viewIcEC1EPKcm t1_standard_encoding FT_MulFix _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_leftEPS7_ _ZN16VirtualAllocator3mapEm _Z16memcpy_optimizedPvS_m _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iteratorC1ES6_ af_cjk_writing_system_class af_nkoo_dflt_style_class af_cprt_nonbase_uniranges _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10rotateLeftEPS7_ strcat __ensure_warn _ZN13ResizePrinterC1Ev _ZN5mlibc7charset8is_printEj af_mymr_script_class _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4item6appendEc FT_Get_Next_Char rand_r FT_Get_Advances af_deva_nonbase_uniranges _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EEclEv TT_RunIns vprintf af_beng_nonbase_uniranges af_latn_pcap_style_class FT_List_Up FT_Outline_Get_Orientation closeButtonSurface _ZN5mlibc8code_seqIcEcvbEv af_shaw_script_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_leftEPS7_SC_ _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN5mlibc14sys_libc_panicEv _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterlEEvRT_T0_biiic _ZN5mlibc13utf8_charcode12decode_stateclERNS_8code_seqIKcEE af_dsrt_script_class af_orkh_dflt_style_class af_bamu_dflt_style_class FT_Attach_File FT_Outline_Get_Bitmap FT_Stream_ExtractFrame _ZN13ResizePrinter6appendEc winfnt_driver_class _ZN5mlibc7fd_file5closeEv memset32_sse2 ft_lzwstate_io FT_Bitmap_New _ZN11PrintfAgentI13ResizePrinterEclEcN3frg14format_optionsENS2_15printf_size_modE af_geor_script_class _ZN11PrintfAgentI14LimitedPrinterEC2EPS0_PN3frg9va_structE af_bamu_script_class fseek _ZN3frg8optionalIiEC1EOi _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE6decodeERNS_8code_seqIKcEERNS3_IjEER15__mlibc_mbstate _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEED2Ev af_cans_dflt_style_class FT_Stream_ReadFields _ZN3frg7eternalI16VirtualAllocatorEC1IJEEEDpOT_ af_avst_nonbase_uniranges ft_hash_str_insert af_armn_dflt_style_class _ZSt7forwardIRiEOT_RNSt16remove_referenceIS1_E4typeE _ZN3frg8optionalIiE13storage_unionD2Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC2Ev getdelim FT_Vector_Rotate _ZN5mlibc7fd_file7io_readEPcmPm cff_cmap_encoding_class_rec af_cyrl_c2sc_style_class FT_GlyphLoader_New _ZN5mlibc13abstract_file4seekEli _ZTVN5mlibc13abstract_fileE wcstold af_arab_dflt_style_class ft_standard_glyph_names FT_Get_TrueType_Engine_Type _Z8DrawCharciihhhP7Surface af_osge_script_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E6removeEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemD2Ev af_telu_uniranges psnames_module_class af_shaper_buf_create FT_Vector_From_Polar FT_Stream_ReadChar stdin FT_Load_Sfnt_Table _ZN13BufferPrinter6appendEPKc _ZN10win_info_tC1Ev af_sylo_uniranges af_grek_sinf_style_class af_grek_uniranges FT_Vector_Unit _ZN5mlibc8InfoSinkclEPKc af_tavt_dflt_style_class _ZN3frg11_fmt_basics12print_digitsI13BufferPrinterlEEvRT_T0_biiic af_latn_subs_style_class _ZN5mlibc7charset8is_spaceEj FT_Stream_Free _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE8freelistC1Ev af_olck_dflt_style_class _ZN5mlibc8code_seqIjEcvbEv TT_New_Context FT_Outline_Embolden _ZN5mlibc13abstract_file10_init_typeEv _ZN3frg7eternalI16VirtualAllocatorE3getEv ferror af_latb_script_class strstr af_arab_uniranges FT_Outline_Check _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_biiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameC1Emmi af_latn_dflt_style_class __cxa_pure_virtual FT_Load_Char _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_NS_14format_optionsERT0_ af_avst_uniranges ps_builder_funcs af_vaii_dflt_style_class _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE16_ensure_capacityEm _ZN11PrintfAgentI13StreamPrinterEC1EPS0_PN3frg9va_structE FT_Raccess_Get_HeaderInfo _ZN3frg11_fmt_basics9print_intI14LimitedPrintermEEvRT_T0_iiic _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_biiic FT_Stream_GetUOffset _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_EC2Ev iswctype _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEmEEvRT_T0_biiic strcoll af_geor_uniranges af_dsrt_dflt_style_class _ZN5mlibc7fd_file14determine_typeEPNS_11stream_typeE isupper af_gujr_script_class _ZN3frg15aligned_storageILm8ELm8EEC1Ev _ZN11PrintfAgentI13ResizePrinterEC2EPS0_PN3frg9va_structE strncmp af_hebr_dflt_style_class _ZN4ListIP8Window_sE6get_atEj _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC2ES7_ _ZN5mlibc7strtofpIeEET_PKcPPc FT_Get_Renderer ft_hash_str_lookup af_nkoo_script_class library wmemset af_grek_dflt_style_class _ZdlPvm _Z18memset64_optimizedPvmm FT_Select_Metrics strncpy FT_Sfnt_Table_Info _ZN3frg15aligned_storageILm1ELm1EEC2Ev FT_Vector_Transform _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEEC1ES7_ program_invocation_short_name af_dummy_writing_system_class _ZN3frg11_fmt_basics9print_intI13StreamPrinteryEEvRT_T0_iiic _ZN5mlibc7fd_file7io_seekEliPl _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS6_12partial_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ FT_Done_FreeType _ZN3frg11_fmt_basics9print_intI13StreamPrintermEEvRT_T0_iiic _ZN3frg17basic_string_viewIwEC1EPKw _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_EC1Ev funlockfile _ZN13ResizePrinter6appendEPKc _ZN11PrintfAgentI13ResizePrinterEC1EPS0_PN3frg9va_structE isascii _ZN3frg4swapERNS_8optionalIiEES2_ FT_Stream_EnterFrame _ZN3frg11unique_lockI13AllocatorLockEC2ERS1_ windowCount towupper _ZN5mlibc7fd_fileD2Ev FT_Set_Char_Size FT_MulDiv_No_Round _ZN3frg11_fmt_basics9print_intI13StreamPrinterjEEvRT_T0_iiic _ZN5mlibc7charset8is_graphEj __cxa_atexit af_cari_nonbase_uniranges _ZNK3frg17basic_string_viewIcE4sizeEv _Z8DrawRectiiii10RGBAColourP7Surface _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE14bucket_to_sizeEj _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clImEEDaS2_ af_sylo_dflt_style_class _ZN13StreamPrinter6appendEPKc FT_Set_Transform strtok _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE6bucketC1Ev af_latn_c2cp_style_class at_quick_exit _ZN3frg8optionalIiED2Ev mouseDown _ZN3frg11_fmt_basics12print_digitsI13StreamPrinterlEEvRT_T0_biiic af_khmr_nonbase_uniranges af_orya_uniranges fdopen _ZN3frg7mt19937C1Ev FT_Matrix_Invert ft_glyphslot_alloc_bitmap af_cyrl_c2cp_style_class af_guru_dflt_style_class _Z19__frigg_assert_failPKcS0_jS0_ FT_Get_Sfnt_Name_Count _Z15DrawBitmapImageiiiiPhP7Surface ft_hash_num_init _Z8DrawRectiiiihhhP7Surface isalpha af_osge_nonbase_uniranges ft_hash_str_init _ZN5mlibc13utf8_charcode12decode_stateC1Ev wcscspn _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9successorEPS7_ wcstoul af_telu_dflt_style_class strncat _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E6removeEPS7_ ft_corner_orientation _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEE3getEv _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE8iterator1hES6_ pfr_cmap_class_rec sfnt_module_class FT_Bitmap_Done af_latp_script_class wcschr FT_Outline_Copy _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE5beginEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10rotateLeftEPS7_ FT_Cos _ZN3frg10escape_fmtC1EPKvm _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev _ZN3frg3minImEERKT_S3_S3_ _ZN3frg8optionalIiED1Ev fread _ZN3frg13printf_formatI11PrintfAgentI13StreamPrinterEEEvT_PKcPNS_9va_structE _ZN11PrintfAgentI13StreamPrinterEclEcN3frg14format_optionsENS2_15printf_size_modE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E14aggregate_pathEPS7_ _ZN5mlibc7fd_fileC1EiPFvPNS_13abstract_fileEE tt_cmap13_class_rec _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E11insert_rootEPS7_ af_writing_system_classes af_shaper_get_cluster _ZN3frg11_fmt_basics12print_digitsI13BufferPrintermEEvRT_T0_biiic ft_glyphslot_set_bitmap af_goth_nonbase_uniranges af_style_classes FT_Get_Sfnt_LangTag af_tfng_uniranges af_tibt_script_class t1_cmap_standard_class_rec _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ strtoull _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvjNS_14format_optionsERT_ _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ FT_GlyphLoader_CreateExtra _ZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE cff_decoder_funcs af_sund_nonbase_uniranges _ZN14LimitedPrinterC2EPcm cff_builder_funcs FT_Face_GetCharsOfVariant fopen __bss_start wcsncat _Z8DrawRect4Rect10RGBAColourP7Surface _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEixEm FT_Matrix_Multiply putwchar _ZN3frg11_fmt_basics9print_intI14LimitedPrinteryEEvRT_T0_iiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_nodeEPS7_ FT_Select_Size main af_ethi_script_class _ZN5mlibc13abstract_file9_save_posEv ft_lzwstate_init wcsspn _ZN11PrintfAgentI14LimitedPrinterEC1EPS0_PN3frg9va_structE ftell af_saur_script_class _ZN5mlibc7charset8is_lowerEj af_bamu_nonbase_uniranges af_buhd_nonbase_uniranges srand af_ethi_dflt_style_class strxfrm af_cher_script_class af_vaii_nonbase_uniranges af_beng_dflt_style_class af_hani_uniranges af_goth_uniranges _ZN5mlibc8code_seqIKcEcvbEv vfwprintf font_default _Z5floord _ZN13AllocatorLock4lockEv FT_Matrix_Multiply_Scaled clearerr af_arab_script_class _ZN5mlibc7fd_file8io_writeEPKcmPm _ZdaPv _ZnwmPv t42_driver_class FT_Outline_Get_CBox _ZN3frg15aligned_storageILm1ELm1EEC1Ev fclose FT_Add_Module _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC2EPNS_9slab_poolIS1_S2_EE getchar _ZN3frg11_fmt_basics14format_integerIiNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ af_vaii_uniranges _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE1hES6_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE5clearEv _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E8get_rootEv af_cari_uniranges autofit_module_class _ZN5mlibc10infoLoggerE FT_List_Remove _ZN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEC1EPNS_9slab_poolIS1_S2_EE isgraph wcsncpy af_cakm_nonbase_uniranges _ZN3frg7eternalI16VirtualAllocatorEC2IJEEEDpOT_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10frame_lessclERKNS3_5frameES7_ fgetpos isalnum _ZN3frg8optionalIiEC1Ev _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E8get_leftEPS7_ tmpnam isprint FT_Outline_New_Internal _ZN4ListIP8Window_sED2Ev af_buhd_script_class _ZN4ListIP8Window_sED1Ev ps_hints_apply _ZN5mlibc16current_charcodeEv af_knda_uniranges _ZNK3frg17basic_string_viewIwE4sizeEv FT_Outline_Done _ZN3frg14format_optionsD2Ev af_latp_dflt_style_class _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11insert_rootEPS7_ FT_List_Insert fread_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE5_emitEPKc strcmp _ZN3frg17basic_string_viewIcE10sub_stringEmm _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC1IJRS2_EEEDpOT_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ FT_Set_Renderer _ZN5mlibc7charset9is_xdigitEj _ZN3frg8optionalIiE13storage_unionC1Ev _ZN3frg9_redblack15null_aggregator9aggregateINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEEEbPT_ _Z11lemon_writeiPKvm _ZN5mlibc13utf8_charcode12encode_stateclERNS_8code_seqIcEERNS2_IKjEE _ZN14LimitedPrinter6appendEc memset64_sse2 af_glag_nonbase_uniranges t1_cmap_unicode_class_rec _ZN3frg11_fmt_basics9print_intI13BufferPrinterjEEvRT_T0_iiic _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE7reallocEPvm af_mlym_script_class _fini _ZN3frg11_fmt_basics12print_digitsI13BufferPrinteryEEvRT_T0_biiic _ZN13AllocatorLockC1Ev _ZN3frg6formatIPvNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg15do_printf_charsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE FT_Get_CMap_Language_ID _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEiEEvRT_T0_iiic ft_raster1_renderer_class fgetc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E10fix_removeEPS7_ af_thai_dflt_style_class FT_Angle_Diff strerror_r af_adlm_script_class _ZN5mlibc13abstract_file11_write_backEv strtof strtod_l _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9get_rightEPS7_ FT_Get_X11_Font_Format af_khmr_dflt_style_class af_mymr_nonbase_uniranges __cxa_guard_release strcspn _ZN3frg17basic_string_viewIcEC1EPKc _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg5_list14intrusive_listIN5mlibc13abstract_fileENS_13locate_memberIS3_NS0_19intrusive_list_hookIPS3_S6_EEXadL_ZNS3_10_list_hookEEEEEE11iterator_toES6_ af_thai_uniranges _ZN13ResizePrinter6expandEv _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEjEEvRT_T0_iiic FT_GlyphLoader_Add flockfile _ZN3frg13locate_memberIN5mlibc13abstract_fileENS_5_list19intrusive_list_hookIPS2_S5_EEXadL_ZNS2_10_list_hookEEEEclERS2_ iswdigit _ZN4ListIP8Window_sE10get_lengthEv af_geok_dflt_style_class af_deva_script_class _ZN11PrintfAgentI13BufferPrinterEclEc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E1hEPS7_ FT_Face_GetCharVariantIsDefault stderr _ZN3frg13printf_formatI11PrintfAgentI13BufferPrinterEEEvT_PKcPNS_9va_structE af_lisu_dflt_style_class _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ ft_mem_strcpyn af_gujr_uniranges af_olck_uniranges _ZN5mlibc11panicLoggerE af_vaii_script_class af_tibt_dflt_style_class srandom _ZN3frg6formatIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ af_none_nonbase_uniranges _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEEC1Ev _ZN16VirtualAllocator5unmapEmm af_guru_uniranges ft_glyphslot_free_bitmap FT_Open_Face FT_Property_Get ft_glyphslot_preset_bitmap _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC2EPS3_ af_arab_nonbase_uniranges _ZSt4moveIRiENSt16remove_referenceIT_E4typeEOS2_ af_cyrl_uniranges af_latb_nonbase_uniranges _ZN3frg11_fmt_basics12print_digitsI13StreamPrintermEEvRT_T0_biiic _ZN14LimitedPrinter6appendEPKcm _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ _ZN3frg15aligned_storageILm8ELm8EEC2Ev FT_Attach_Stream putchar_unlocked ft_service_list_lookup _ZN3frg16do_printf_floatsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE FT_Stream_New ft_hash_num_lookup _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ tt_default_graphics_state _ZN3frg9_redblack11hook_structC2Ev _ZN3frg9_redblack11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS6_10frame_hookEEENS5_10frame_lessENS0_15null_aggregatorEE6insertEPS6_ af_cher_nonbase_uniranges _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E9get_rightEPS7_ _ZN13ResizePrinterC2Ev fputc _ZN14LimitedPrinterC1EPcm FT_Bitmap_Convert _ZN3frg7eternalINS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2IJPNS_9slab_poolIS2_S3_EEEEEDpOT_ _Znam af_cher_dflt_style_class FT_Done_Library feof_unlocked FT_List_Iterate _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4backEv _Z24CreateFramebufferSurface6FBInfoPv _ZZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E_clIjEEDaS2_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E14aggregate_pathEPS7_ getchar_unlocked _ZN3frg7eternalINS_9slab_poolI16VirtualAllocator13AllocatorLockEEEC2IJRS2_EEEDpOT_ _ZN11PrintfAgentI14LimitedPrinterEclEc FT_Sin _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12replace_nodeEPS7_SC_ af_mymr_uniranges af_tavt_uniranges fwide iswupper __ensure_fail t1_expert_encoding af_grek_pcap_style_class FT_Stream_GetChar FT_List_Find _ZN5mlibc13abstract_file5flushEv fflush_unlocked _Z13lemon_readdirimP12lemon_dirent FT_Outline_Done_Internal _ZN3frg14format_optionsC2ERKS0_ FT_Library_Version FT_Render_Glyph_Internal FT_Outline_EmboldenXY _ZN3frg6formatINS_10escape_fmtENS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ _ZN3frg11_fmt_basics12print_digitsI13ResizePrinterjEEvRT_T0_biiic fputws _ZN3frg14format_optionsC1Ev FT_Hypot af_hani_dflt_style_class ft_smooth_lcdv_renderer_class _ZN3frg11unique_lockI13AllocatorLockE4lockEv _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17decode_wtranscodeERNS_8code_seqIKcEERNS3_IwEER15__mlibc_mbstate fwrite_unlocked af_olck_nonbase_uniranges af_latin_writing_system_class af_buhd_dflt_style_class wmemcmp _ZN11PrintfAgentI13StreamPrinterEclEc _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11rotateRightEPS7_ lldiv _ZN3frg11unique_lockI13AllocatorLockEC1ERS1_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E5isRedEPS7_ wmemmove _ZSt7forwardIPN3frg9slab_poolI16VirtualAllocator13AllocatorLockEEEOT_RNSt16remove_referenceIS6_E4typeE af_geok_nonbase_uniranges ft_validator_run _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clIjEEDaS2_ _ZN5mlibc13abstract_fileC2EPFvPS0_E isdigit FT_CMap_New af_guru_nonbase_uniranges FT_Get_Track_Kerning _ZN5mlibc13sys_anon_freeEPvm fwrite FT_Match_Size FT_Stream_GetUShort _edata _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ _Z19__mlibc_do_finalizev FT_Get_First_Char _end _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE17encode_wtranscodeERNS_8code_seqIcEERNS3_IKwEER15__mlibc_mbstate _ZN5mlibc9sys_closeEi FT_Bitmap_Copy FT_Gzip_Uncompress _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10deallocateEPvm af_saur_dflt_style_class af_shaper_get_coverage af_sinh_script_class af_telu_nonbase_uniranges ft_hash_str_free _ZN3frg11_fmt_basics12print_digitsI14LimitedPrintermEEvRT_T0_biiic vfscanf _ZN3frg14format_options15with_conversionENS_17format_conversionE rewind _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEC2ES5_ _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E16remove_half_leafEPS7_SC_ af_knda_nonbase_uniranges af_orya_nonbase_uniranges _ZN3frg9_redblack11hook_structC1Ev freopen _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E10fix_removeEPS7_ af_grek_script_class _ZN3frg11_fmt_basics9print_intI13ResizePrinteryEEvRT_T0_iiic fgetc_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIiEERS4_T_ _ZN3frg14format_optionsD1Ev af_grek_ordn_style_class af_cans_uniranges _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE5frameC2ENS3_10frame_typeEmm ungetwc af_copt_nonbase_uniranges t1_cmap_expert_class_rec af_limb_script_class FT_Vector_Length af_lao_dflt_style_class _ZN3frg11_fmt_basics14format_integerIjNS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEEEvT_NS_14format_optionsERT0_ psaux_module_class af_orya_dflt_style_class _ZN3frg3getINS_5_list10locate_tagENS_13locate_memberIN5mlibc13abstract_fileENS1_19intrusive_list_hookIPS5_S7_EEXadL_ZNS5_10_list_hookEEEEEEERT0_PNS_11compositionIT_SA_EE af_lisu_uniranges _ZZN3frg14do_printf_intsI14LimitedPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E1_clImEEDaS2_ _ZN3frg7mt199374seedEj FT_New_Face _ZN5mlibc7fd_file17determine_bufmodeEPNS_11buffer_modeE _ZN5mlibc13abstract_fileC1EPFvPS0_E _ZN5mlibc20polymorphic_charcodeD2Ev _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinterlEEvRT_T0_biiic _ZN3frg15do_printf_charsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE towlower af_tavt_nonbase_uniranges _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E1hEPS7_ af_geor_nonbase_uniranges af_khmr_uniranges _ZN5mlibc7charset8is_upperEj FT_Reference_Library llabs _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E7isBlackEPS7_ _ZN3frg6formatIPKcNS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvRKT_RT0_ af_thai_script_class FT_GlyphLoader_Done _ZN5mlibc9sys_writeEiPKvmPl setbuf _ZN5mlibc20polymorphic_charcode7promoteEcRj iswalnum wcscmp af_latp_nonbase_uniranges _ZN3frg8destructIN5mlibc13abstract_fileENS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEEEvRT0_PT_ af_adlm_nonbase_uniranges _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEED2Ev atoi _ZN11PrintfAgentI13ResizePrinterEclEc iscntrl af_gujr_nonbase_uniranges af_khms_script_class ft_mem_qrealloc _Z10DrawWindowP8Window_s _ZN3frg11unique_lockI13AllocatorLockED2Ev FT_Get_Name_Index ferror_unlocked _ZN5mlibc13abstract_fileD0Ev _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEviNS_14format_optionsERT_ af_taml_script_class _ZZN3frg14do_printf_intsI13BufferPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clImEEDaS2_ af_shaper_buf_destroy FT_Bitmap_Embolden fileno fgets_unlocked _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsENS_8endlog_tE ft_standard_raster getline _Z10surfacecpyP7SurfaceS0_8Vector2i _ZN5mlibc13utf8_charcode12decode_state6cpointEv _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIPKcEERS4_T_ _ZSt4moveIRbENSt16remove_referenceIT_E4typeEOS2_ wcscat _ZN3frg15aligned_storageILm456ELm8EEC2Ev FT_Get_Module_Interface strspn FT_CMap_Done _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE10slab_frameEXadL_ZNS7_12partial_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_12partial_hookEEES9_E11predecessorEPS7_ _ZN3frg11_fmt_basics12print_digitsINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEjEEvRT_T0_biiic _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E9successorEPS7_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4item6appendEc strlen _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemC1EPS3_ _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsIjEERS4_T_ _ZZN3frg14do_printf_intsI13StreamPrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structEENKUlS2_E0_clIjEEDaS2_ program_invocation_name _ZN3frg10escape_fmtC2EPKvm af_cakm_uniranges toupper ft_grays_raster _ZN5mlibc13utf8_charcode12decode_state8progressEv FT_Stream_OpenMemory ft_corner_is_flat atoll _ZN5mlibc7charset8is_punctEj _ZN3frg8optionalIiEdeEv _ZN3frg11_fmt_basics9print_intI13BufferPrintermEEvRT_T0_iiic _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemD1Ev wcsxfrm ft_smooth_renderer_class af_cans_script_class af_saur_nonbase_uniranges _ZN4ListIP8Window_sE9remove_atEj FT_Add_Default_Modules af_cprt_uniranges FT_Tan _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE11_find_frameEm _ZN3frg14do_printf_intsI13ResizePrinterEEvRT_cNS_14format_optionsENS_15printf_size_modEPNS_9va_structE strchr _ZN5mlibc8sys_exitEi ft_mem_strdup FT_Activate_Size _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockEC1ERS1_ fputs _Z11lemon_closei _ZSt4swapIPcEvRT_S2_ t1cid_driver_class _ZN5mlibc17sys_anon_allocateEmPPv _ZN3frg3maxIiEERKT_S3_S3_ af_limb_dflt_style_class font_old _ZN3frg13format_objectINS_19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemEEEvPKvNS_14format_optionsERT_ t1_cmap_custom_class_rec FT_Get_Postscript_Name _ZN5mlibc8sys_readEiPvmPl af_ethi_uniranges _ZN3frg8optionalIiE13storage_unionD1Ev fgetwc vfwscanf _ZSt4swapIiEvRT_S1_ ft_hash_num_insert FT_Stream_Pos af_grek_nonbase_uniranges tt_cmap0_class_rec vasprintf af_khmr_script_class fbInfo fputc_unlocked strchrnul _ZN3frg11unique_lockI13AllocatorLockED1Ev _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE4pushEOS1_ _ZN3frg6vectorIPcNS_14slab_allocatorI16VirtualAllocator13AllocatorLockEEE3popEv af_shaw_uniranges FT_CeilFix _ZN3frg11_fmt_basics9print_intINS_19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemEmEEvRT_T0_iiic _ZN11PrintfAgentI13StreamPrinterEC2EPS0_PN3frg9va_structE _ZdaPvm _ZN5mlibc7charset8is_blankEj memcpy_sse2 _ZN5mlibc7charset8to_lowerEj aligned_alloc __cxa_guard_acquire posix_memalign _ZNK3frg17basic_string_viewIcEeqES1_ _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE16_construct_largeEm _ZN5mlibc7fd_fileD0Ev af_grek_subs_style_class FT_Library_SetLcdFilter af_cyrl_pcap_style_class windows FT_Outline_New _ZN13StreamPrinterC2EP17__mlibc_file_base _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE10tiny_sizesE _ZN3frg9_redblack16tree_crtp_structINS0_11tree_structINS_9slab_poolI16VirtualAllocator13AllocatorLockE5frameEXadL_ZNS7_10frame_hookEEENS6_10frame_lessENS0_15null_aggregatorEEES7_XadL_ZNS7_10frame_hookEEES9_E12insert_rightEPS7_SC_ _ZN5mlibc7fd_fileC2EiPFvPNS_13abstract_fileEE mbtowc _ZN3frg19stack_buffer_loggerIN5mlibc8InfoSinkELm128EE4itemlsINS_10escape_fmtEEERS4_T_ _ZN3frg11_fmt_basics12print_digitsI14LimitedPrinteryEEvRT_T0_biiic vfprintf af_sylo_nonbase_uniranges ft_lcd_padding strpbrk _ZSt4moveIRN3frg14slab_allocatorI16VirtualAllocator13AllocatorLockEEENSt16remove_referenceIT_E4typeEOS7_ _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN3frg9slab_poolI16VirtualAllocator13AllocatorLockE4freeEPv _ZN3frg17basic_string_viewIcEC2EPKcm fputwc _ZN5mlibc28polymorphic_charcode_adapterINS_13utf8_charcodeEE24decode_wtranscode_lengthERNS_8code_seqIKcEEPmR15__mlibc_mbstate _ZN5mlibc13abstract_file5writeEPKcmPm _ZN3frg19stack_buffer_loggerIN5mlibc9PanicSinkELm128EE4itemlsIjEERS4_T_ afm_parser_funcs _ZN5mlibc18generic_is_controlEj af_armn_nonbase_uniranges  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .tbss .init_array .ctors .dtors .data.rel.ro .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                               � @     �                                     !              @            �+                            '             �,H     �,                                   -              -H      -     
s                             5             �J     �
     T%                            ?             �K      �                                   E              �K      �                                  Q             �K     �                                   X             (�K     (�                                   _             8�K     8�     x                             l             ��K     ��     `                              r              �K      �     `                              w      0                �     +                             �                      P�      8                             �                      p                                   �                      �     ��                            �                      |�     ��                             �                      �     ��                            �                      �f$                                   �      0               �f$     �y                           �                      ��'     �                            �                      ��9     ��                                                  ��;     ��         &                	                      ��<     Q;                                                  ��=     �                              