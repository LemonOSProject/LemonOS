ELF          >    � @     @       ��          @ 8  @                   @       @     �4      �4                    @       @@      @@     h      �             �+  �+  �     H��    UUH��������I  ����    �hL@ H=hL@ t�    H��t	�hL@ ��f��ff.�     @ �hL@ H��hL@ H��H��H��?H�H��t�    H��t�hL@ ���ff.�     @ �=)K   uwUH�'K  H��ATA�@@ S�@@ H��@@ H��H��H9�s%f.�     H��H��J  A��H��J  H9�r��0����    H��t
� ,@ �<���[A\��J  ]��ff.�     @ �    H��tU��L@ � ,@ H������]����D  ����UH��AWAVAUATSH��hH�}�H�E��@����t:H�E�H�   H��H�E�H� H�¸ M@ A�    A�    H�ƿ   ��(  �  �    � �    ��%�� �    H�u�H���   H�u��v������I��H�    ����L!�H	�H��H�Ή�H�       H	�H��H��H��H��H�ι M@ ����  �    � �    ��%�� �    H�U�L���   L��H�    ����H!�H��I��H�U��R�҃���H�� L���H	�I��L��L��L��L��H��H�ι M@ ���Y  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H���/  H��p���H�E��@������H��x���H�    ����H!�H	�H��x���H��x�����H�       H	�H��x���H��p���H��x���H��H��H�й M@ ��H��H���  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�    H�E�H���   H�E�H��H���f
  H�E�H�U�H�    ����H!�H��H�E�H�E��@������H�� H�U���H	�H�E�H�E�H�U�H��H��H�й M@ ��H��H����  �    �@�@   �ǉ�%�� �  @ ���E�   �E�   H�E�H���   H�E�H��H����	  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H�й M@ ��H��H���A  H�E����   ����H�E����   ����H�E�H��H��h M@ A��   A��   ��   H���  H���E�   �E�   H�E�H���   H�E�H��H����  H�E�H�E�H�U�H�� M@ A�    A�    H���   �0%  H�e�[A\A]A^A_]�UH��SH��  ��L@ �{  H��F  H��F  H��H��H��F  H���F  �H��F  f�HH���0  H��H�E�H�E�H�H�HH�vF  H�wF  H�PH�HH�pF  H�qF  H�@ H�nF  �XF  �NF  ��H�H���  H�FF  H�E��PH�E��@�u�h�   A�    A��   �щ¾    �    ��  H��A�    A�    �    �    �    �   �$  H��p���H���  H������H����  fǅ����d fǅ����d fǅ����
 fǅ����
 H������H��H�Test WinH�0�@dow ǅ����    H������A�    A�    �    �    H�ƿ   �{#  �	,@ A�    A�    �    �    H�ƿ   �S#  �    �,@ ��  �E��E��   �(M@ ���-  ��D  ��D  h M@ h�   A��   A�@   �щ¾    �    �  H��H������A�    A�    �    �    H�ƿ   ��"  ������9E���  �������E��E�    �E�;E���  �E� H��p���H���j  �E�Hc�H��p���A�    A�    �    H�ƿ   �a"  H������H�E��E�    H��p���H���~  9E�����t.�U�H��p�����H���r  H� H9E�����t�E���E���Eۃ����  ��   �  H�E�H�E�H��p���H��x���H�PH�HH������H������H�PH�H H������H������H�P(H�H0H������H������H�P8H�H@H������H������H�PHH�HPH������H������H�PXH�H`H������H������H�PhH�HpH������H�Px���������   H�E�H�U�H�H�E��@��H�E��@
��H�E����   H�E����   H�U�H��p���H��H���  �E��7����E�    �E�;E�}*�U�H��p�����H���  H�E�H�E�H���|����E��΋E��   �(M@ ���  ��7  �qB  ��Љ}7  �{7  �ZB  ��)Љg7  �DB  �������u  �2B  �����c  � B  H��p���H���d  ���Ẽ}� �=  �U�H��p�����H���R  H�E���6  H�E����   9��  ��6  H�E����   H�E��@���9���   ��6  H�E����   9���   ��6  H�E����   H�E��@���9���   �U�H��p�����H����  H��H��p���H��H���#  �U�H��p�����H���  H�E�H�E����   �P�46  9�|RH�E��@����uD�6  H�E����   )
6  H�E����   )��ȉ�@  ��@  ��@  �	�m��������@  ��th��5  ��@  )�H�E����   ��5  ��@  )�H�E����   H�E����   ��yH�E�ǀ�       H�E����   ��yH�E�ǀ�       �J@  ����t�=@  ��t�2@   �*@  ��t�@  ������u�@   �@   � @  ��t0h M@ j A�    A��   �2   �2   �,  �    �  H����?  ������t0h M@ j A��   A�    �2   �2   �,  �2   �d  H���E�    H��p���H����  9E�������   �E� �E�    �E�;E�}sH��p���H���8  �E�Hc�H��p���A�    A�    �    H�ƿ   �/  H������H�E��U�H��p�����H���`  H� H9E�����t�E���E���Eǃ���t�U�H��p�����H���U  �E��5����5�3  ��3  h M@ j A�    A��   �   �   ���^  H��H�    ����H!�H�É�H��H�E�H�ھ M@ H���A
  �?���UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]ÐUH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H�}�u�H�E�@9E�r
�    H� �3H�E�H� H�E��E�    �E�;E�sH�E�H� H�E��E���H�E�H�@]�UH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �]
  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��H�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]ÐUH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H���;  H�E���D  L�J�H��taI��vH�t$�fnL$�I��1�I��fp� f�     H��H��H��I9�u�H��H���H�<�I)�H9�t�7M��t�wI��t�w�D  ATUH��SH��H����t]H��tGH��t>H�l$�~D$H��1�H��fl� H��H��H��H9�u�H��H���H��H9�tH�+H��[]A\��     I��H��H��A���  M��t�H�+I��t�H�kI��t�H�kI��t�H�kI��t�H�k I��t�H�k(I��t�H�k0H��[]A\�H��H	�t��  �AUI��ATA��I��UH��SH��L)�H��H��H���  M��uH��[]A\A]��    H��I�4H�| L��[]A\A]�  D  SH���(   ��  H�T$H�     H�P�T$H�X�P�T$�P[�ff.�     f��,�f��1��*�f/���)���     SD�\$L�T$��y�1���y�1�A��E��E��M�J��A��D	�A	���~LA;r}F�\�D�\�D  ��~'A�B9�}���A�B��9�~���H�E��D9�u�9�t	��A9r�[�fD  D��SE������AQ��A��P�T���XZ[�H��I��H��A��H�� ��H�� ������� AWf��AVA��AUA�ՍRAT��A��USL��H��A�@
�L$J�, �B>��I����*�������L$D��    D�y�E������   D;s��   A�D�D��G�t,��D$@ E����   D�CE9���   D��D��D�\$�UD  D�S L�[G��D��E��G�M��L�KD�A�HE�	D�A�HH�{D�D9�t?D�C����A9�~0���xD�L �HH�H�A��u��9u��?u�D9�u��    D�\$E)�9t$t��9s�>���H��[]A\A]A^A_�ff.�     @ AWD��AVAUA��D��AT��A��U����SH��8H�\$p��y�1�E��yE�E1���  ;{�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$� A��D9s~nf���L$D��D���A*Ǻ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P�w���XZD9�u�H��8[]A\A]A^A_ÐAWD��AVAUA����ATA��U��D��S��H��8H�\$p��yA�E1��y�1����  ;s�  D��f��������f��f��E�����*�f��A���*�D��E��E1��*����*��t$�\�f���A*��|$ �^��t$(�$f���*��\��^��D$f���A*��\��^��D$�@ A��D9s~nf���L$D��D���A*ǹ   D��A���Y��XL$ �D,��L$�Y��XL$(S�YD$E���XD$ �D,��,�E����P����XZD9�u�H��8[]A\A]A^A_Ð�NH��H�� ����   AVAUATUS�O��)���~qI��I���,�    E1��f�     A�E)�D9�~KA�FA�M��    A��Hcҍ4�    A�E Hc�Iv�<�B�#A�����Hc�I}����E9f�[]A\A]A^�ËNA��AUH�� ATL�VUSH�_����   �G)Ѕ���   D�f��E1�f.�     E��~d�G��D)�~X1�E�)��    �G��D)�9�~:D��A���Hc�A��A��A��A���   uA���D�H���D�f��D9�|��NA��A9�}
�G)�D9��[]A\A]�f.�      H���   HD���  ff.�     @ ��  ff.�     �k
  ff.�     �����ff.�     �K
  ff.�     �;
  f.�     �UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��L��H��~7fHn�fo%�@ f��fs�f��fs�f��fs�f��f H����H��]�UH��H��H��L��H��~%fHn�fo%�@ f��fs�f��f H����H��]Ð�����������                AW�B��A��AVAUE��ATU��SH��H��`F@ �D$A��L�t$P�L$H��D$�Z A��@��   A�� ��   A����   A���  A���0  A���Z  A����  H�뀃�9l$��  D�#E��y�A��AVD���   RD�L$�   ��D�D$�Z���_AXA��@�w���A��AV�   ��RD�L$A��   D�D$�&���Y^A�� �N���A��AVA��   RD�L$�   ��D�D$�����XZA���%���A��AVA��   RD�L$�   ��D�D$�����A[XA�������A��AVA��   RD�L$�   ��D�D$����AYAZA�������A��AVA��   RD�L$�   ��D�D$�W���_AXA�������A��AV�   ��RD�L$A��   D�D$�#���A��Y^�}���A��AV�   ��PD�L$A��   D�D$H�뀃������XZ9l$�T���H��[]A\A]A^A_�ff.�      AWI��AVAUATUSH���?@��tEA��A��E��A����fD  H��D��D��E���t$HA���I��A���M���A�?XZ@��u�H��[]A\A]A^A_� H��H��E1�E1�H�t$1ɿ   H�D$    �i  H�D$H���f.�     D  H��H��E1�E1�H�T$1ɿ   �2  �D$H���f�     Hc�E1�E1�1�1ҿ   �	  f�     H��H��H��Hc�L�D$H��E1ɿ   ��  �D$H���D  H��H��H��Hc�L�D$H��E1ɿ   �  �D$H���D  H��Hc�E1ɉ�L�D$Hc��   �  �D$H���f�     H����E1�Hc�L�D$1��X  �D$H���ff.�     @ H���7���H��H��H���W���H��H���{���ff.�     ����ff.�     H�������1�H���H��1������   ��u��H���D  ������1�H����ÍGP1�S�5�+  �����9�+  C�+  ��H����
  f��H��HM@ @�X��+  H�     H�@    H�@     �X�@(   H[��     H��HM@ H�n,      H�[,      H�     H��@M@ �?+     H�     H��8M@ �#+      H�     H�,      H��+      H��+      �f.�     AWAVAUI��ATUSH���D  1�H��+  A�   ��	  M�e 1��	  M��t�H��+  H����  H��+  I�mHH����  �S�KA�   A��A)�I9���  ��)�L9�v
H�l+  I��H9�s$H�CH����   �P�HH�É�)�L9�w�H9�r�H�S H���@  H��H)�H��(H9���  H�J�rH��t%H��H)�H��(H)�H9���   H��H�J�rH��uۋCH�D�H)�H)�H9��8  H�CH���t���A��t#D�������H�CH����  H��Q���A��uH��*  H����  E1��3���f�D������H�CH���r  H�H���(���H�T$�~D$H�H�L$H�F(H��`�F����D�f�D$D�n�F�H�JH�^�H�H�BA�D$(H��CH��@M@ L ��u<H���   �F�1��  H��H��[]A\A]A^A_ËP�HH��E1��[����    �   H)�Hƃ�H���D  �P�HH��E1�E1��(���@ H�2H�H(H�JH�P(A�T$(D�`DH�@0    �@@���H�X8D�hHSH��@M@ L"L�"H��8M@ L9"LC"H��`H��L�"��uH�ź   �P�1��9  �2����   H)�HЃ�H����D���)���H�)  H���V���1�1��   �����H�C(�C@���f��H�C C(A�D$(CH��@M@ D�cDL D�kHH�[8L� H��8M@ L9 LC H��`H��L� ��u7H�ݸ   �C�1��  ����H�C(H�H�S0H�C �C@���H�C(    닸   H)�HÃ�H���ff.�     �H����   SH�G�H��H)�H�� HC�1��  �C�H�s�=���u~�K�H�{�H��@M@ H��H)
�OH�S�)���H�K؃�(�G�C�ޭ�H��tH�
H�H����   H�QH�W H��'  H��tnH��t�w�Q+Q)�9�}H�=�'  1�[�   ��H�~'  ����� ���� t
f=��t<�u�H�V'  1�[�n  fD  H�P'  ��    H9=Q'  H�GtKH9�tVH�H��tH�BH�GH��tH�H��HM@ �W�wH)�Y  1�[�  �H�W �5����    H��&  ��    H��&      � ��SHc�H�������H��t1�1��     � �QH��H9�w�[�ff.�     @ AUATUSH��H��H����  I��H����  H�G�H��H)�H�� HC�1��T  �E�H�U�=����2  D�e�M9��e  1��>  L���6���H��I����  H�CI�L$�H9�H�E��H9������  H���v  H��1�H��H��H��H��H��fD  �oD H��H9�u�H��H���H��H��    H��L�H�I�<�H9�t'A��H�W�H��vA�PH���PH��vA�P�PH��H��H��   H��H�4L�$�H�M��t��I��t�V�PI��t�V�PH�������H��H��[]A\A]�f.�     ��H��$  ����� ���� tHf=��tB<�t>1�1���  H��H��[]A\A]��    D�j 1�H����  H��H��[]A\A]�@ H��$  �fD  �[���1��l���@ H��H��[]A\A]����fD  H��H��H�4�   1��    ��T H��H9�u������ H�������H��L�B�H����   I����   �t$�I��H��I���I�fnD$�f`�fa�fp� f�H��L9�u�H��H���H�8I)�H9���   @�1M����   @�qI��t|@�qI��tr@�qI��th@�qI��t^@�qI��tT@�qI��tJ@�qI��t@@�qI��t6@�q	I��	t,@�q
I��
t"@�qI��t@�qI��t@�qI��t@�q�H���e���ÐH��H���  H�NL�B�H9�H�H@��H9���@���   I����   M��1�I��I��L��H��H���oH��H9�u�M��I���J�<�    H�>H�M9�tH�	H�I����J��   H�H�H��v�>H��H��H���y�H��t)�<@�<H��H��tD�D�D�D�H��t�V�Q�f�L��H��L��   1��    H�<H�<H��L9�u��u���f�H���f.�     �I��SH��H��H��L��L��L���i[�fD  1��ff.�     f�H��xM@ �  1�� H��Hc�E1�E1�H�T$1ɿ   ����H�D$H����     1��f.�      H�9  H���t3UH��S� @@ H��D  ��H��H�H���u�H��[]�f.�     ��J����  /snake.lef /dev/mouse0        zR x�        ����I    A�CD  (   <   ����   A�CM�����      h   ����2    A�Cm      �   s����   A�CH�   �   ����-    A�Ch      �   ����    A�CL      �   ����V    A�CQ       ����"    A�C]       $  �����    A�CE��       H  R���-   A�C(        l  `���k       <   �  �����    B�A�D �G0U
 AABI[ AABL   �  L���k    R�E�H �D(�M0R
(A ABBHD(M� A�B�B�        l���3    A�q      ,  ����          @  �����    A��  $   \  ���     D�LG FAA      �  ���       H   �  ���Q   B�F�E �H(�G0�A8�GP"8A0A(B BBB   T   �  (���o   B�E�B �H(�G0�F8�Dpxa�FxApI8A0A(B BBB  T   <  @���o   B�E�B �H(�D0�F8�Gpxa�FxApI8A0A(B BBB  <   �  X����    T�B�B �A(�A0�}(A BBBA�����4   �  �����    H�F�E �A(�� ABB           P���             \���          4  X���          H  T���          \  P���          p  L���       �   �  8���R   B�K�B �E(�A0�C8�DP�XI`XXBPPXH`ZXAPPXJ`XXAPPXJ`YXAPPXJ`YXBPPXJ`XXBPPXH`^XAPLXH`aXAPN8A0A(B BBBT   ,  ����m    B�E�B �B(�A0�A8�D@cHMPWHA@I8A0A(B BBB        �  ���1    D l    �  0���'    D b    �  H���          �  T���+    D f    �  l���+    D f    �  ����'    D b      ����!    D \    (  ����    DI    @  ����    DI    X  ����          l  ����          �  ����    DK     �  ����0    DV
FM          �  ����h    F�a     �  ����v       H   �  `����   B�B�B �E(�A0�A8�DP�
8D0A(B BBBA,   8  ����m   J��
�Hm�[�B
�F    h  ���1    D�l   t   �  (���P   B�B�A �A(�G0_
(D ABBKo
(D ABBHR
(D ABBEd
(D ABBK         �   ����            ����         $  ����    D�U          D  ����          X  ����          l  ����(    D c    �  ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ��������        ��������                                               1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d                                                                                                                                                                                                                                                                                                  <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             @     �      �@     I       @     2       P@     -       ~@            �@     V       �@     "       @     �       �@     -                      ,    a       �@     �                                       ]       �  �  	  0               �  
5   �  �  int �   �  ]   �  W  p   =  �  �     ;   �        �   �  
�   7  w    ;  w   bpp d     w   
 �   �   �   �  �  �  (|  x C    y 	C   7  C   ;  C     C   P  
Q   H  	|  `  

Q     	Q   �  
  �   �  x 	C    y C    �  	�  
�  �  s   �  	�  |�  c  x d    y d   7  d   ;  d     w   �  c  Z  �   l  �  t�  l  \  �
    �  s  �   _ �  �  �  	�  �  �  	�  	  �  	�  $  	�  C   �  �    �  �  	@@@     .  �;"    <�   �  =s  pos >�  ��   ?"  � �  fb B
|  	�L@     �  D�   	�L@     �  F�  	 M@     )   z  �    G  Hj  	(M@     ,  I�  	@B@        J"  	+M@     �  K"  	,M@     ]   L�  	0M@     G  �  6  D   
    �   5    %  0  �  C    �  !u  E  K  �   �  -   `  k  �  �   �  >%  �  �  �  �   �  N<  �  �  �  �  �    �  X�  �  �  �  �  �    �  bO  �  �  �  �   �     l�   C       �   �   p�  �  0  ;  �  �      �  �  T  Z  �   Q  �V  �  s  y  �   �  �   �  �  num ��   T �   	�  
�  	�  �    |   	       
  obj �  �   *         T �   	�  
    =  �@     -      ��  �  �  �Hpos p�   �D U  v  �h!obj z�  �X"�@     	       �   �  r�  �P #�@     8       !i x�   �d  K  �  @     �       �  �  �  �Hobj -�  �@ �  .  �X $�       %�     &  ]  C  �@     "       �L  '  �h (�  k  �@     V       ��  �  �  �Xpos N�   �T U  Q  �h#�@             !i S�   �d  (�  �  ~@            ��  �  �  �h )�  �  �  %�  �   &�  v    P@     -       �%  '�  �h *B  cC   @     �      ��
   �  e�  �� �  mC   �\ �  o�  ��~ �   p�  �P h   rs  ��} �   ~C   ��#@     �       �  �C   ��}"�@     �      o	  !j �C   �L#�@     �       �  �
"  �K �   �s  ��| �   ��  ��"�@     N       K	  !i �C   �D #G	@           !win ��  ��   "^
@     9       �	  !i �C   �@#m
@     $       !win ��  ��  "@     \      �	  !i �C   ��+    !win ��  ��  #�@     �       !i �C   ��#�@     �        �  �	"  ��#�@     �       !j �C   ��#�@     m        �   �s  ��| �   ��  ��~      	s  
�
  $O  �
  �
  %�  �
   &�
  z  �
  @     2       ��
  '�
  �h ,�  N  @           �  win N�  �� �  ^�  �� -�    �  �@     I       �Z  l 0Z  �hr EZ  �` .�   N    �  �@     �@     +  src/gfx/sse2.asm NASM 2.14.02 ��@              %U   :;9I  $ >  $ >  :;9   :;9I8   :;9I8  ;   	 I  
& I     :;9n  .?n4<d   I4  I  ! I/   <  4 :;9I?<  4 :;9I?  4 :;9I?  :;9  .?:;9n2<d   I  .?:;9nI2<d   :;9I82   :;9I82  / I  .?n42<d  .Gd@�B   I4   :;9I   4 :;9I  !4 :;9I  "  #  $.G:;9d   % I4  &.1nd@�B  ' 1  (.Gd@�B  ).Gd   *.?:;9I@�B  +U  ,.?:;9n@�B  -.?:;9nI@�B  . I   %  . @   '   s  �      /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/gfx/window /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include /home/computerfido/Desktop/Lemon/FakeSysroot/usr/include/lemon  graphics.h   main.cpp    window.h   list.h   stdint.h   fb.h   surface.h   types.h   stdio.h    G 	�@     
�ff!.  tt!.�  	@     � Lt<ZK
�H<
t&!#'�
<E$:D�
</#�1tQ�#<<T�bXh�
<f.�4�#<�:�
.J�j�
<6#��'�5 
�7N9�<'.)�<.�0&�N�	0GJ	t����1u<6:Kf<f(<�
v	9%�������	�*(!?
9*f�� t
�K�+�* t ��<<tKK +mt'����)��= lX� t � u �k>f��f��tf � ��"u%�* f�uf�, �9 fG �; �  .Y �f fM �t �� f� �� �h .�)v�<f5 J; t& <K+f �7.Df9�J�v v.
�%�,ff.�,ff.��( J��( J�� J	�w  �" t fK	uw�0tfK0( t �	�K t��+�<<tKxfft& J q<�4)  	@     �*  	P@     ����  	~@     � 
�u  	�@     � �t* X�� t* � �h�  	�@     �  	@     ,�#��tY�����  	�@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K �    '   �       src/gfx/sse2.asm      	�@     !>==?LLKK0=!$!>==?LLKK0=!#!>==>K0Y�KYKYKYMKL1="#!>==>K0Y�KYMKL1=""��            prev mouseDown uintptr_t _ZN4ListIP8Window_sE8add_backES1_ uint64_t _ZN4ListIP8Window_sEC4Ev dragOffset testWindow handle_t next long long int windowHandle windowInfo fb_info_t _ZN4ListIP8Window_sE10get_lengthEv ListNode mouseDevice Vector2i active remove_at _ZN4ListIP8Window_sE9get_frontEv stdin _ZN8ListNodeIP8Window_sEC4Ev List<Window_s*> uint16_t linePadding _ZN10win_info_tC4Ev this _windowCount keymap_us GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions _ZN4ListIP8Window_sE9remove_atEj temp get_front long unsigned int _Z10DrawWindowP8Window_s width short unsigned int depth _ZN4ListIP8Window_sE8get_backEv _ZN4ListIP8Window_sEC2Ev ListNode<Window_s*> bool stdout decltype(nullptr) FBInfo operator[] windowFound vector2i_t fbInfo long double title pitch /home/computerfido/Desktop/Lemon/Applications/Init _ZN4ListIP8Window_sEixEj current _ZN8ListNodeIP8Window_sEC2Ev _ZN10win_info_tC2Ev operator+ _ZN4ListIP8Window_sE6get_atEj surface_t unsigned char node short int info main.cpp 10win_info_t clear uint32_t _ZplRK8Vector2iS1_ get_length _ZN4ListIP8Window_sE9add_frontES1_ buffer _ZN4ListIP8Window_sE10replace_atEjS1_ _ZN4ListIP8Window_sE5clearEv add_back drag IOFILE replace_at get_at stderr add_front renderPos fbSurface uint8_t DrawWindow windows renderBuffer flags handle _ZN4ListIP8Window_sED4Ev mousePos ~List height main mouseData get_back ownerPID                 *@     ]@     f@     g@                     @     �@     �@     @     @     P@     P@     }@     ~@     �@     �@     �@     �@     @     @     �@     �@     �@                                                    � @                   � @                   ,@                   	,@                    ,@                    @@                   @@                    @@                  	 �L@                  
                                                                                                                                                                                                                           ��                      @@                  @@             (      ,@             ;     � @             =     @             P     P@             f    	 �L@            u    	 �L@            �     �@             �    	 �L@     0           ��                �     @@             �     �4@             �     �+@             �    ��                �    ��                     � @                ��                #   ��                /   ��                @     �@             Q     !@             l     x@                  �@             �     �@             �     �@             �    �@            �   ��                �   ��                �   ��                �   ��                b   ��                �    � @     h       �    dL@            �    `L@               	 pM@               	 hM@               	 `M@            .   	 XM@            ;   	 PM@            N   ��                W   ��                a   ��                m   	 HM@            y    � @             �    �@     o      �    @B@            �   	  M@     (       �   	 8M@            �    @+@            �    � @     v       �    p+@            F   	 xM@              "  �@                @@     +           0@     o      D  "  �@     "       a     *@           h  "  �@     I       {   	 @M@            �   hL@             �   @@             �   	 0M@            �    �@     '       �    p!@     �      �    @@             �  "  �@     "       �  "  @     �           �@     1             @              "  �@               	 ,M@            $  "  �@     V          	 �L@            �    � @             =    `+@            K    @@@            U  "  @     2       i    �@     k       �    �&@     1       �    @             �   	 (M@            �     @            �    0@     k       �    8@             �    p@     +       �    �@     R      �  "  @     2       �    � @                  @                �+@     (         "  �@            %    `@     �       @    �&@     P      H    �@             m   	 +M@            w    �@     Q      �     @     �       �    @@     m       �  "  P@     -       �   	 hL@             �    �@                  )@     �       '    @     �      ,    `F@            9    �@            C  "  �@            J    �@             X    ,@             ^  "  ~@            �    �+@            �  "  �@            �    �@     3       �    P @     0       �    hL@             �   	 �M@             �  "  P@     -       �    �@     '       �    @               @     �       �    0 @            /     @            ;  "  �@     -      \    `B@            e   	 �L@            l  "  �@            t    �@     !       �    �@             5    @ @            �    �@     �       �     %@     m       crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4699 dtor_idx.4701 frame_dummy object.4711 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux graphics.cpp /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp runtime.cpp src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret bigzero text.cpp font.cpp fb.c filesystem.c allocate_new_page l_pageSize l_pageCount l_memRoot l_bestBet l_warningCount l_errorCount l_possibleOverruns memory.c syscall.c _liballoc.c l_allocated _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface mousePos renderBuffer l_max_inuse syscall liballoc_init liballoc_unlock _Znwm lemon_read _Z12DrawGradientiiii10RGBAColourS_P7Surface _ZN8ListNodeIP8Window_sEC2Ev memcpy _ZplRK8Vector2iS1_ l_inuse __TMC_END__ __DTOR_END__ dragOffset lemon_open malloc __dso_handle _ZN8ListNodeIP8Window_sEC1Ev _ZN4ListIP8Window_sE8add_backES1_ lemon_map_fb lseek _ZdlPv drag _ZN4ListIP8Window_sEixEj liballoc_lock keymap_us _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm calloc memcpy_sse2_unaligned mouseData _Z16memcpy_optimizedPvS_m memset32_sse2 lemon_write _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev liballoc_alloc _ZdlPvm _Z18memset64_optimizedPvmm realloc _Z8DrawRectiiii10RGBAColourP7Surface mouseDown _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main font_default _Z5floord _ZdaPv memset64_sse2 _fini _ZN4ListIP8Window_sE10get_lengthEv liballoc_free _Znam _Z24CreateFramebufferSurface6FBInfoPv access _edata _end _ZN4ListIP8Window_sEC2Ev lemon_seek _Z10DrawWindowP8Window_s _Z10surfacecpyP7SurfaceS0_8Vector2i lemon_close _ZN4ListIP8Window_sE9remove_atEj font_old fbInfo _ZdaPvm lemon_readdir memcpy_sse2 _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                  � @     �                                     !             � @     �       A+                             '             ,@     ,                                    -             	,@     	,                                    5              ,@      ,      �                             ?              @@      @                                    F             @@     @                                    M              @@      @      H                              S             �L@     hL                                     X      0               hL      +                             a                      �L      �                              p                      sM                                    �                      �M      �                             �                      8Y      �                             �                      \      �                             �                      �c                                    �      0               �c      c                            �                      7i                                    �                      Gi      �                                                    j      @         @                 	                      Xx      �                                                   �      �                              