ELF              ��4   �7      4    (           � ��(  �(           �(  �����   �        �W  ��  �                 �    UU���}  VW�����_^�Y  �    �i���f�f�f�f�f��,�=,�t$�    ��tU���h,��Ѓ��Í�&    f�Í�&    ��&    ��,�-,����������t(�    ��tU���Ph,��҃��Í�&    �t& �Í�&    ��&    ��=@� ugU�D���V���S����딸����9�s�v ���D����D�9�r��'����    ��t��hО�Q~�����@��e�[^]�Í�&    ��&    ��    ��t'U���hH�hО�~������	�����&    f�������L$����q�U��Q��  f�`�/ �E� �ĸ��P�  ����h`��  ���ȸ��P�  ���E�<
tơ(�Pjj�E�P�  ��������tك�hĞ�a  ����U��S���v  �5  ��h   ����  ���E�}� u�    �%�E�U�P�E�   �E�P�E��@   �E�]���U��S���  �â5  �E�    ���u��u�  ���E��}� y�    �$���u�u��[������E�}� t�E���    �]���U��S���  ?5  �U�R�U���u����  ���    �]���U��S���  5  �U�R�U�U�U��R�u�u����  ���E��E��]���U��S���B  �4  �} t,�U�R�U�U�U��R�u�u����  ���E��E�����]���U��S����   �4  �M�U�R���uQR����  ���]���U��S����   P4  �U�R��jj R���  ���]���U���   &4  �    ]�U���   4  �    ]�U��S���q   �3  �URjj�UR���������]���U��S���I   ���3  ���u�-  ���E�E��ujP�u��������E�9�u�    �������]��Ë$Ë$�U�������y3  ǀ\      ǀ`      ǀ0      ǀ4       ����    �B    ����    �B    ����    �B    ǀd      ǀh      ǀl      ǀp      ǀt      ǀx      �]�U����@����2  �E�    ��U�E�ЋU��E��E�;Er�E��U����	����2  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS��������2  �E���E�E���0   �E�    ��Ѕ�u��0   �E�    ���E����0   �E�    �����E䋃4   9E�s	��4   �E���u��T  ���E���jj �u���������}� u%��d  ��h  ���� ��d  ��h  �    �l�E��     �E��@    �E��U�P��0   �E�E��P�E��@   �E��@    �E��@�ƿ    ����P� �������Q�E��e�[^_]�U��WVS��L�`������0  �E�    �E�    �E�    �E�    �E�E��E� �-  �}� u5��d  ��h  ���� ��d  ��h  �  ��j�������  ��\  ��u-���u��9�������\  ��\  ��u��  �    �{  ��\  �E��E�    ��`  ���C  ��`  �P��`  �@)ЉE��E�    �E����    ;E؉�E��
  ��`  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ�`  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u��\  �E��E�    �|  ���u��'������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ����P� �������Q����0�x����P� 9Ɖ��s�Ɖ�����0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    ����P� �������Q����0�x����P� 9Ɖ��s�Ɖ�����0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���X  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    ����P� �������Q����0�x����P� 9Ɖ��s�Ɖ�����0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    ����P� �������Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u��\  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������Y  �    �e�[^_]�U��WVS��,�,����ñ)  �} u#��d  ��h  ���� ��d  ��h  �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx��l  ��p  ���� ��l  ��p  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u��t  ��x  ���� ��t  ��x  �c  �  �E��@�E�����P� �M��I�ο    )�������Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ��\  9E�u�E܋@��\  ��`  9E�u
ǃ`      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋�����P� �M܋I�ο    )�������Q�E܋@��P�u��z  ���G��`  ��t=��`  �P��`  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉�`  ��  �e�[^_]�U��S������5'  �U�U�U�U��R���%������E��E��Pj �u��-������E��]���U��S���e������&  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E���
  �E���E�E�@=���tz��l  ��p  ���� ��l  ��p  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u��t  ��x  ���� ��t  ��x  �
  �    �_�E�@�E�E�;Er�E�U�P�b
  �E�;�X
  ���u��������E���u��u�u����������u��������E�]���U���������%  �E�    ��E��U��E�� ��u�E���U��S���������S%  �E�    �E�    ��U�EЋM�U�� ��E����u������9E�|ԋU�E��  �E�]���U����j����$  �E�    ��U��EЋM��U�� ��E��E�9EwߋU��E��  ���U��S���%����ê$  ���u�	������EЃ��uP�$������E�]���U�������p$  ��E�P�U� ��u�    ��E� �U8�u܋E]�U�������5$  �E�    �(�E� �U8�u�E�E��E�P�U� ��u�E���E� ��u΋E��U��S���_������#  �E�    ��E��E� ��t"�E�P�U� ����P�u�4�������uЋE�]���U��S�������Ñ#  �E�    �)�E� ����P�u���������t�E���E�E��E� ��u͋E�]���U��VS������=#  �} t�E��|  ���|  ��u
�    �   ��|  ��|  ���uP�
�������E���u�u�G������EЉ�|  ��|  9Euǃ|      ��|  �/��|  � ��t��|  �  ��|  ����    ��|  �E�e�[^]�U�������y"  ��E�E�E��E� 8�u
�E� ��uދE� �ЋE� ��)�]�U�������-"  �E�    ��E��E�E�E��E� 8�u�E� ��t�E�9EwҋE� �ЋE� ��)���U��VS�J������!  ��E�E�E� ����P�  ���ƋE� ����P��  ��9�u
�E� ��u��E� �ЋE� ��)Ѝe�[^]�U��VS���������[!  �E�    ��E��E�E�E� ����P�  ���ƋE� ����P�{  ��9�u�E� ��t�E�9Ew��E� �ЋE� ��)Ѝe�[^]�U��S���P������   ���u�4���������P��������E���u����������Pj �u��  �����u�u�� �������]���U��S�������j   �M�U��j j j QRj���C  �� �E�]���U��S������4   �U��j j j j Rj���  �� ��]���U��S���y���   �]�M�U��j S�uQRj����  �� �E�]���U��S���@����  �]�M�U��j S�uQRj���  �� �E�]���U��S�������  �]�M�U��j SQ�uRj���f  �� �E�]���U��S�������W  �]�M�U��j S�uQRj���-  �� �E�]���U��S������  ���u�u�u����������]���U��S���i����  ���u�u�u���������]���U��S���=����  ���u�u�u���������]���U��S�������  ���u�u���������]���U��S�������q  ���u���������    �]���U��S���������F  ��j �u�������E�}� t���u���������    ��   �]���U��WVS�t����  �E�]�M�U�u�}�i�[^_]�U��S���I����  ��$����R�u���������]���U��S�������  ��$����R�u���������]���U�������x  �}/~�}9~�}`~�}z~�}@~�}Z�   ��    ]�U������9  �}`~�}f~�}@~�}F�   ��    ]�U���}���  �}z����]�U���d����  �}@����]�U���K����  �}/~�}9�   ��    ]�U���$����  �}/~�}9~�}`~�}f~�}@~�}F�   ��    ]�U��������k  �E�E����U�������U  �E��!��]����]�U������7  �} t�}	u�   ��    ]�U������  �]�U���w���   �]�U��S���g������  ���u�~�������t���u�I�������u�   ��    �]���U��� ����  �E��_]�U�������  �E�� ]�U�������  �    ]�U�������k  ��@��  �    ]�U��S�������J  �M�U��j j j QRj���#����� �E�]���U������  �    ]�U����x���  �E�E���E��P�U��U��E�P��U��u�E��U��� �@����  �E�E��E�E��E�E��"�E��P� �M���Q�E��E��m�E�E�}�w؋E�E���E���E���E��E��m�E�E��}�wދE�E���U��E�ЋM��U��� ��m�E�E�}� uۋE�á�����t6U��S�������&    �v �Ѓ�����u��[]Í�&    ��&    ������  
Lemon:  > test1234

         zR |�         ����    D Gu Cu|       @   }���]    A�BD�U��     d   ����c    A�BD�[��     �   ����4    A�BD�l��      �   ���@    A�BD�x��      �   !���J    A�BD�B��     �   G���1    A�BD�i��        T���.    A�BD�f��     <  ^���    A�BP�     \  R���    A�BP�      |  F���,    A�BD�d��      �  N���Q    A�BD�I��    �  {���          �  k���          �  [����    A�B��      ����7    A�Bs�     ,  ����r    A�Bn� ,   L  Q���8   A�BF���+�A�A�A�   ,   |  Y���4   A�BF���'�A�A�A�   ,   �  ]���~   A�BF���q�A�A�A�       �  ����K    A�BD�C��        ����f   A�BD�^��   $  ���1    A�Bm�      D  %���a    A�BD�Y��    h  b���H    A�BD�     �  ����>    A�BD�v��     �  ����8    A�Bt�     �  ����P    A�BL�     �  ����S    A�BD�K��       ���V    A�BD�N�� $   4  M����    A�BB����A�A�   \  ����I    A�BE�    |  ���_    A�B[� $   �  S���q    A�BB��i�A�A�$   �  �����    A�BE��|�A�A�    �  ����k    A�BD�c��       B���6    A�BD�n��      4  T���2    A�BD�j��      X  b���9    A�BD�q��      |  w���9    A�BD�q��      �  ����9    A�BD�q��      �  ����9    A�BD�q��      �  ����,    A�BD�d��        ����,    A�BD�d��      0  ����,    A�BD�d��      T  ����)    A�BD�a��      x  ����+    A�BD�c��      �  ����J    A�BD�B�� (   �   ���*    A�BC���`�A�A�A�     �  ����/    A�BD�g��        	���/    A�BD�g��     4  ���?    A�B{�     T  3���3    A�Bo�     t  F���    A�BU�     �  ?���    A�BU�     �  8���'    A�Bc�     �  ?���?    A�B{�     �  ^���    A�BU�       W���    A�BZ�     4  U���'    A�Bc�     T  \���    A�BL�     t  L���    A�BL�      �  <���G    A�BD���     �  _���    A�BQ�     �  T���    A�BQ�     �  I���    A�BP�     	  =���    A�BY�      8	  :���6    A�BD�n��     \	  L���    A�BP�     |	  @���8    A�Bt�     �	  X����    A�B��     ����    ����                                            ��                                                                                � � �GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o                      t�          ��          ��          ��          О          ��          ��          ��          ��     	     @�     
                           ��   ��         ��      (   О      ;   ��      =    �      P   P�      f   @�    
 u   D�    
 �   Ё      �   H�    
             ���   ��      �   ��      �   p�      �            ��  ��                  ��           ��           ��  ��    
 )  ��    
 3  ̸    	 >  и    	 J   �    
 Y  �    
 f  �    
 y  ȅ7     �  ��r     �  q�8    �  ��4    �           ���  �    
 �           ���           ���           ���           ���           ��           ��           ��             ��  ��      /  ��/     7  �    
 C  =�a     %  $�    	 J  �    
 V  ��*     ^  ��     l  )�     U  @�    
 |  ��9     �  ��     �  `��    
 �  �     	 �  ȝ�     �  �    
 �  ,�    	 �  ��     �  �/     �  &�6     �  ��     �   �     �  ��     �  ��4    �  �       ��    	   ��G       ]�'     #   �     
 *  n�     1  ʙ,     7  4��     C  �?     f  t�      L  �     Z  \�P     b  [�K     |  ��,     i  �>     p  �1     v  ǘ9     $  (�    	   ��&     �  ĸ    	 �  r�,     �  ��     �  d�_     �  F�6     �  ��H     �  Öq     �  ��f    �  U��     �  �     �  ��]     �  [�3     �  ��@        ��k       �c       ,�     
 �  ��8       ��       @�.     $   �     	 ,  Q�4     3  ?�     ;  �?     C  ��     K  ȸ    	 X  �I     _  ��      e  ��V     �   �    	 m  |�     {  ��,     �  ��'     �  ŃJ     �  J�J     �  ,�     	 �  D�     
 �   �9     �  &�     �  ��S     �  �1     �  ��)     �  �     �  \�2     �  $�8     �  Q     �  9�9     �  �+     v  ݎ~     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp fileio.c l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 string.c p.1056 filesystem.c syscall.c stdstreams.c stdout.c ctype.c _liballoc.c memory.c _GLOBAL_OFFSET_TABLE_ putchar l_allocated strcpy l_max_inuse syscall liballoc_init liballoc_unlock lemon_read isblank currentDirectory _stderr l_inuse __TMC_END__ __DTOR_END__ lemon_open islower tolower feof malloc __x86.get_pc_thunk.ax __dso_handle ispunct isspace _stdin fflush lseek strncasecmp isxdigit liballoc_lock strrchr calloc strcat fseek lemon_write promptStringStart isupper strncmp liballoc_alloc strncpy strcasecmp realloc strtok __x86.get_pc_thunk.bx fdopen isalpha fread strdup fopen __bss_start main ftell _stdout fclose isgraph isalnum isprint promptString strcmp _fini strcspn liballoc_free fputc isdigit fwrite access _edata _end lemon_seek iscntrl strspn strlen toupper lemon_close strchr fputs lemon_readdir  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment                                                     t�t                     !         ���   !                 '         ���                    -         ���                    5         О�  �	                 ?         ���(                    F         ���(                    M         ���(                   V         ���(  l                   \         @�,)                    a      0       ,)  +                               X)   	     6         	              X2  �                               K7  j                  