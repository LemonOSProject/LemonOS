ELF          >    �@     @       x�5         @ 8  @          @       @ @     @ @                              X      X@     X@                                          @       @     �\	     �\	                    `	      `i      `i     �      �                    (`	     (`i     (`i     P      P             /lib/ld64.so.1     "                                         !                                                                  	         
                                                                                       	                                                                                        '                      .                      4                      ;                      B                      P                      W                      _                      f                      l                      �     �@            s                      z                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                      �                       libc.so longjmp strcpy setjmp memmove getenv qsort memcpy malloc __mlibc_entry strtol strrchr strcat fseek memchr strstr strncmp strncpy realloc __cxa_atexit memcmp isalpha fread fopen memset ftell fclose isprint strcmp sprintf strlen toupper free _start �ai                   �ai                   �ai                   �ai                   �ai                   �ai                   �ai                   �ai                   �ai        	           �ai        
           �ai                   �ai                   �ai                   �ai                    bi                   bi                   bi                   bi                    bi                   (bi                   0bi                   8bi                   @bi                   Hbi                   Pbi                   Xbi                   `bi                   hbi                   pbi                   xbi                   �bi                    �bi        !           �+  �F� �     �5�W) �%�W) @ �%�W) h    ������%�W) h   ������%�W) h   ������%�W) h   �����%�W) h   �����%�W) h   �����%�W) h   �����%�W) h   �p����%�W) h   �`����%�W) h	   �P����%�W) h
   �@����%�W) h   �0����%�W) h   � ����%�W) h   �����%�W) h   � ����%�W) h   ������%zW) h   ������%rW) h   ������%jW) h   ������%bW) h   �����%ZW) h   �����%RW) h   �����%JW) h   �����%BW) h   �p����%:W) h   �`����%2W) h   �P����%*W) h   �@����%"W) h   �0����%W) h   � ����%W) h   �����%
W) h   � ����%W) h   �����H��@ �t���@ ��ti H=�ti t�    H��t	��ti ��f��ff.�     @ ��ti H���ti H��H��H��?H�H��t�    H��t��ti ���ff.�     @ �=�h)  uwUH��h) H��ATA�`i S� `i H��`i H��H��H9�s%f.�     H��H�mh) A��H�bh) H9�r��0����    H��t
�0�H �|��[A\�2h) ]��ff.�     @ �    H��tU��ti �0�H H���C��]����D  ����UH��SH��   L�EԸ   �    �    �    �    L���i�Eԉ�h) �E�    ��ui �Q  9E�������   �E� �E�    �th) 9E�}cH��P���H���  L��P����   �M�    �    �    L���iH�E�H�E؋E�ƿ�ui ��  H� H9E�����t�E���E���E����t�E�ƿ�ui ��  ��\) �E��E����H�Ĩ   []�UH��SH��   L�E̸   �    �    �    �    L���i�Ẻ�g) �E�    ��g) 9E��2  �E� H��P���H����  L��P����   �M�    �    �    L���iH�E�H�E��E�    ��ui ��  9E�������   �E�ƿ�ui ��  H� H9E�������   �E�ƿ�ui ��  H��P���H��X���H�PH�HH��`���H��h���H�PH�H H��p���H��x���H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�Uȉ��   �E��	�E������E������   ��   ����H�E�H�E�H��P���H��X���H�PH�HH��`���H��h���H�PH�H H��p���H��x���H�P(H�H0H�U�H�M�H�P8H�H@H�U�H�M�H�PHH�HPH�U�H�M�H�PXH�H`H�U�H�M�H�PhH�HpH�U�H�Px�Uȉ��   H�E�H�U�H�H�E��@��H�E��@
��H�EЉ��   H�EЉ��   H�E�H�ƿ�ui �  �E������QZ) �H�Ĩ   []�UH��H�� H�}�H�u�H�M�I����tH�M��I���H�M��I�Ƀ��M�H�M�H���   H�M��I�ɉ�H��H�    ����H!�H	�H�ʋM�H�� H�։�H	�H��H�M�H��H��H��H��H��H���W  ��UH��AUATH�� H�}�H�u�H�E؋@����t�    ��   �E��E�    �E�E�H�E�H���   H�E�H��H���i  I��H�E��@����L��H�    ����H!�H	�I��H�E��@����H�� L���H	�I��H�E�L��L��L��L��H��H��H���  �H�� A\A]]�UH��AWAVAUATSH��   H�}�H�E��@�����  H�E��@����t6A�@ui H�E�H� H��H�E�H�   H�¸   �    �    L���i��  �    � �    �ǉ�%�� �    ���E�   �E�    H�E�H���   H�E�H��H���L  H��@���H�E��@����H��H���H�    ����H!�H	�H��H���H��H�����H�       H	�H��H���H��@���H��H���H��H��H�й@ui ��H��H����  �    � �    �ǉ�%�� �    ���E�    �E�   H�E�H���   H�E�H��H���  H��P���H��X���H�    ����H!�H��H��X���H�E��@������H�� H��X�����H	�H��X���H��P���H��X���H��H��H�й@ui ��H��H���7  �    � �    �ǉ�%�� �    ���E�    H�E��@�����E�H�E�H���   H�E�H��H����  H��`���H�E��@������H��h���H�    ����H!�H	�H��h���H��h�����H�       H	�H��h���H��`���H��h���H��H��H�й@ui ��H��H���n  �    � �    �ǉ�%�� �    ��H�E��@�����E��E�   H�E�H���   H�E�H��H���  H��p���H��x���H�    ����H!�H��H��x���H�E��@������H�� H��x�����H	�H��x���H��p���H��x���H��H��H�й@ui ��H��H���  A�    A�*�2   D���A��D��%�� �  @ A�Ļ    �`�`   �ǉ�%�� �  ` ���E�   �E�   H�E�H���   H�E�H��H���#  I��H�E��@����L��H�    ����H!�H	�I��L����H�       H	�I��L��L��L��L��H��A�@ui D���H��H���F  H�E����   H�E��@��Ѓ���H�    ����L!�H	�I��H�E����   ����H�� D��H	�I��L����ui �@ui ��  H�E����   ����H�E����   ����H�E�H��H��h@ui A��   A��   ��   H���'  H���E�   �E�   H�E�H���   H�E�H��H����  H�E�A�@ui H�E�H� H��H�U��   �    �    L���i��H�e�[A\A]A^A_]�UH��ATSH���   �(ui �M  H��]) H��]) H��H��H��]) H���]) �H��]) f�HH���  H��H�E�H�E�H�H�HH��]) H��]) H�PH�HH��]) H��]) H�@ H��]) ��]) ��]) ��H�H���J���H��]) H�E��PH�E��@�u�h�   A�    A��   �щ¾    �    �0  H���   A�    �    �    �    �    D���i� �F �"�F �����H�E�H�}� u
�   �"
  H�E��   �    H�������H�E�H������H�E�H�E��    �    H�������H�E�H�H���w���H�E�H�u�H�U�H�E�H�Ѻ   H���7���H�E�H��H�E�H�E��@��\) H�E��@��\) ��  �'���H��\) ��\) ��\) H�M�A��ui I�ȉщ¾    �    �  A�4�F �   �    �    �    �    L���i�    �F�F �g  �E��E��   �hui ���  ��[) ��[) A�@ui D�:Q) �щ¾    �    �  �Q) ��t,��[) ��[) A�@ui D�Q) �щ¾    �    �  �E�    ��[) 9E�}%�E�ƿ�ui �	  H�E�H�E�H��������E�����P)  �E��   �hui ����  ��P) �Q[) ���Љ{P) �yP) �8[) ���)ЉeP) �[P) ��y
�MP)     �KP) ��y
�=P)     �3P) ��Z) 9�|��Z) �P) �P) ��Z) 9�|��Z) �P) ��Z) ����   ��O) ��O) ��Z) H� [) )щʉ��   ��O) ��Z) H��Z) )щʉ��   H��Z) ���   ��yH��Z) ǀ�       H��Z) ���   ��yH��Z) ǀ�       �.Z) �������}  �Z) �����k  �
Z) ��ui ��  ���E�}� �J  �E�ƿ�ui ��  H�E�H�E�H�5O) H����������  �E�ƿ�ui ��  H�ƿ�ui �%	  H�E�H��Y) ��N) H�E����   �P��N) 9���   H�E��@������   H�E����   H�E��@��ЍP�|N) 9��vN) H�E����   ��9�~h�[N) H�E����   H�E��@��ȃ�9�}DHǅp���   H�E�H�@tH���u���x�����p�����h�����`���H���o  H��0��  ��M) H�E����   )�M) H�E����   )��ȉ�X) ��X) ��X) ��   Hǅp���   H�E��@����t0��M) H�E����   )ЉE��M) H�E����   )ЉE��4�lM) H�E����   )Ѓ��E�VM) H�E����   )Ѓ��E��E�H�� H�E�H	�H��x���H�E�H�@|H�E�H�E�H�@tH���u���x�����p�����h�����`���H���X
  H��0��	�m�������W) ����t��W) ��t��W)  �W) ���\  �mW) �������G  �[W)  �UW)  H��W) H��t!H��W) H�5oL) H���������t�   ��    ����   �PL) H�iW) H����   Hǅp���   H�NW) �@����t6�L) H�7W) ���   )ЉE܋ L) H�W) ���   )ЉE��:��K) H�W) ���   )Ѓ��E܋�K) H��V) ���   )Ѓ��E؋E�H�� H�E�H	�H��x���H��V) H�@|H�E�H��V) H�@tH���u���x�����p�����h�����`���H����  H��0H�qV) H��t!H�eV) H�56K) H��������t�   ��    ����   Hǅp���   H�,V) �@����t6��J) H�V) ���   )ЉEԋ�J) H��U) ���   )ЉE��:��J) H��U) ���   )Ѓ��Eԋ�J) H��U) ���   )Ѓ��EЋE�H�� H�E�H	�H��x���H��U) H�@|H�E�H��U) H�@tH���u���x�����p�����h�����`���H���  H��0H��0���H���Z  H�������0  H��@���H=�  ��   H=� u�H�U) H����   H��H��������hi �E�H��P���H��t�Ẻ��������t�Ẻ��~����E�H��H���H��H��t(H��H�����H��tHǅp���   �E�H�H��x����Hǅp���   �E�H�H��x���H�}T) H�@|H�E�H�nT) H�@tH���u���x�����p�����h�����`���H���  H��0�(H��H���H��u�0����H��H���H��u� ����������������H) ��H�    ����L!�H	�I�ċ�H) ��H�� D��H	�I��L��`hi �@ui �:  �!S) �S) ������H�<S) H�E�H�@H��H����  �7F) �-F) �5cH) �YH) A�@ui D�UH) ����
  �"���H�e�[A\]�UH��H���}��u��}�u'�}���  u��ui �   ��bi ��ui �@&@ �������UH����  �   ����]�UH��H�}�H�u�H�U��
H�U��ʉ�H�    ����H!�H	�H�U��JH�U��Rʉ�H�� ��H	�]ÐUH��H�}�H�E�f�   H�E�f�@  H�E�f�@  H�E�f�@  �]�UH��H�}�H�E�H�     H�E�H�@    H�E��@    �]ÐUH��H�}�H�E��@]ÐUH��H��H�}��u�U�H�E���H���   ��UH��H��0H�}؉u�H�E؋@��tH�E؋@9E�r	H�E���   H�E�H� H�E��E�    �E�;E�s)H�E؋@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@H�E�H�E�H� H��t H�E�H�@H��tH�E�H� H�U�H�RH�PH�E�H�@H��tH�E�H� H��tH�E�H�@H�U�H�H��}� uH�E�H�H�E�H�H�E؋@�P�H�E؉PH�E؋@9E�����tH�E�H�PH�E�H�PH�E�H������H�E��ÐUH��H�}�H�E�H�     H�E�H�@    �]�UH��SH��(H�}�H�uп   �K  H��H�    H�C    H�C    H������H�]�H�E�H�     H�E�H�@    H�E�H�U�H�PH�E�H� H��uH�E�H�U�H��,H�E�H�@H��tH�E�H�@H�U�H�H�E�H�PH�E�H�PH�E�H�U�H�PH�E؋@�PH�E؉P�H��([]�UH��H�}�u�H�E�@��tH�E�@9E�sH�E�H� H��uH�E�H� H�@�KH�E�H� H�E��E�    �E�;E�s)H�E�@9E�sH�E�H� H��tH�E�H� H�E��E���H�E�H�@]�UH��H��H�}�H�E��@��tH�E��    H���2�������UH��SH�}�H�E�    L�E�H�M�   �    �    �    L���iH�E�[]�UH��SH�}��u�L�E�H�M��   �    �    �    L���i�E�[]�UH��S�}��   D�E��    �    �    �    D���i�[]�UH��S�}�H�u�H�U�H�M�H�u��   D�E�H�Uп    D���i�E�[]�UH��S�}�H�u�H�U�H�M�H�u��   D�E�H�Uп    D���i�E�[]�UH��S�}�H�u؉U�H�u�   D�E�H�M؋U�    D���iH�E�[]�UH��S�}�H�u�H�U�H�M�H�u�!   D�E�H�Uؿ    D���iH�E�[]�UH��SH�}�L�E�H�M�   �    �    �    L���iH�E�[]�UH��SH�}�H�E H�E�H�E(H�E�H�E0H�E�   L�E�H�M�H�U�H�u�    L���i�[]�UH��H��H�}�H�}� uH�E�   H�E�H��������UH��H��H�}�H�}� uH�E�   H�E�H���`�����UH��H��H�}�H�E�H����������UH��H��H�}�H�u�H�E�H����������UH��H��H�}�H�E�H���������UH��H��H�}�H�u�H�E�H���m������UH��H�}��u�H�U�H�E�H�P�H�U�H������tH�E��U�H�E��ڐ]�UH��H��0H�}�H�u�H�U�H�E��H��t(H�E�H�P�H�U�H������toH�E�H�U�H�H�E���H�E؃�H�E�H�E�H+E�H�E�H�E�H��H��H�M�H�E�H��H���  H�E�H�P�H�U�H������tH�E�H�U�H�H�E��ؐ��UH��H��0H�}�H�u�H�U�H�E��H��uH�E���H��tH�U�H�M�H�E�H��H�������   H�E؃�H�E�H�E�H+E�H�E�H�E��H��uH�E���H��t H�E�H��H��H�M�H�E�H��H���  �H�E�H��H��H�M�H�E�H��H���E  H�}� t'H�U�H�E�H�4H�U�H�E�H�H�E�H��H��������UH��H�� H�}�(   ����H�E�H�E��@    H�E��PH�E���E��H�E��P�E��H�E��P�E��H�E��P�E��H�E��PH�E�H�U�H�PH�E���UH��SH��H��H��H�M�H�]�H�U؋U؋E�9�|/�E؋M��U��9�} �U܋E�9�|�E܋M�U��9�}�   ��    []�UH���E��E��,��E��*E�f/E�v�E�����E�]�UH��H�� I��H��L��L��H��H�u�H�}��U�H�M��M��U��u�E�L�E��}�M��A�����  ���UH��H��@�}܉u؉UԉM�D��D�ɋE�ỦʈUȈEă}� y�E�E��E�    �}� y�E�E��E�    �E������E���	��E�	�   ��E�H�EH�@H�E��E�    �E�;E���   �U��E��H�E�@9�}u�U��E��H�E�@�E�U܋E��H�E�@9�|H�E�@+E���EԉE�}� ~,�E�HcЋM܋E�ȉ�H��    H�E�H��E���H��������E��l������UH��H�� �}��u��U�M�D�E�L�M��E����E�D���E�D���M��U�u��E��u�W������H�����UH��H��P�}̉uȉUĉM�L�E�L�M�H�E�H�H�UҋP�U��@f�EދE܉�HE��E��E��Eă��P��H����*��������E�E����E��E��E�    �E�   �E�    �E�;E���  �U�E��H�E��@9���  �E�    �E�;E��k  �U��E��H�E��@9��T  �E������E��E�Љ�H�E�H�� <uT�E������E��E�Ѓ���H�E�H�� <u,�E������E��E�Ѓ���H�E�H�� <��   �UȋE�Љ�H�E��@�E��ЋM̋E���E�ЉE��E������E��E�Љ�H�E�H�H�E�H�P�E�H����E������E��E�Ѓ���H�E�H�H�E�H�@�U�����H����E������E��E�Ѓ���H�E�H�H�E�H�@�U�����H������E������E�)E��E��E�E��E��F������UH��H��0�}�u�U�M�D�E�D�M؃}� y�E�E��E�    �}� y�E�E��E�    �E�    �E�;E��  �U�E��H�E�@9���   �*M��E����*��E����*��\��*U��^��Y��E����*��X��,����*M��E����*��E����*��\��*U��^��Y��E����*��X��,�D���*M��E����*��E����*��\��*U��^��Y��E����*��X��,����U�E��<�U��E��uQE��A���Ѻ   �������H���E���������UH��H�� I��H��L��L��H��H�u�H�}��U�M�L�E��M��U��u�E�D�E�}�H���u�E��A�����   H�����UH��H��0�}�u�U�M�D�E�D�M؃}� y�E�E��E�    �}� y�E�E��E�    �U�E��H�E�@9�~H�E�@+E���E�E��E�    �E�;E��  �U�E��H�E�@9���   �*M��E����*��E����*��\��*U��^��Y��E����*��X��,����*M��E����*��E����*��\��*U��^��Y��E����*��X��,�D���*M��E����*��E����*��\��*U��^��Y��E����*��X��,����U�E��4�U�E��uQE��A���   ������H���E���������UH��H��0H�}�H�u�H�U��E�    H�E��@9E���   H�E�P�E�)�9E���   �U�H�E��@�H�E�@9�~H�E�P�E�)��H�E��@�E��E���H�H�U�H�JH�U��R�U���Hc�H�4H�U�H�JH�U�RD�E܋}�D����U����Hc�H�H��H�������E��E������UH��H��@H�}�H�u�H�U�H��L��H��H�E�H�UȋU��E��H�E��@9�~H�E��P�E�)���EȉE��UċE��H�E��@9�~H�E��P�E�)���ẺE�U؋E��H�E�@9�~H�E�P�E�)���E��E��E�    �E�;E���   H�E�P�E�)�9E�}v�E���H�H�U�H�J�uċU��H�U��R����Hc�U���Hc�H�H�4H�U�H�JH�U�RD�E܋}�D����U����Hc�H�H��H��������E��k������UH��H�}�H�u�H�U�H�E�H�@H�E�H�E�H�@H�E��E�    H�EЋ@9E���   H�E؋P�E�)�9E���   �E�    H�EЋ@9E���   H�E؋P�E�)�9E���   H�EЋ@�E��E��H�H��    H�E�HЋ ��=�   vWH�EЋ@�E��E��H�H��    H�E�H��ŰE��H�E؋@�ЋE�E��H�H��    H�E�H����E��I����E������]�UH��H�r?) H����  �X?)     �]�UH��SH��(�B?) ����H�=C?) �  ������t*L��i �    �    �    �    �    L���i�^  H�5�i H�=�i ����H�E�H�}� u*L��i �    �    �    �    �    L���i�  H�E�   �    H���%���H�E�H�������H�E�H�E�    �    H�������H�E�H������H�E�H�U�H�u�H�E�H�Ѻ   H���c���H�E�H������H�U�H�D>) H�u�L�A>) �    H���D�  �Eԃ}� t%L�i �    �MԺ    �    �    L���i�QH��=) �   �    H����?  �EЃ}� t%L��h �    �Mк    �    �    L���i�
��=)    H��([]�UH��SH��8H�}���=) ����H�=�=) �K  ������t*L��g �    �    �    �    �    L���i�^  H�E�H�5�g H���U���H�E�H�}� u*L�ah �    �    �    �    �    L���i�  H�E�   �    H���j���H�E�H������H�E�H�E�    �    H���D���H�E�H�������H�E�H�U�H�u�H�E�H�Ѻ   H������H�E�H�������H�U�H��<) H�u�L��<) �    H��艾  �Eԃ}� t%L��g �    �MԺ    �    �    L���i�QH�D<) �   �    H���2>  �EЃ}� t%L�8g �    �Mк    �    �    L���i�
��;)    H��8[]�UH��SH��x���u��U���D��D�ɈE��ЈE����E��ȈE��E���������u
�    �!  ��;) ��u�;�����;) �����   �e��E�    �}���   �E������E��H���ni H���E��E�    �}�L�E��y;�E��M��U��}�u��D�E�}�D��uPA��A�й   �   �T���H���e�E�뮃E��v����   �d  �E������E���	��E�	�   ��E�H�EH�@H�E�H�M�H��:) �   H��H���j�  �Ẽ}� t7L�f �    �M̺    �    �    L���i�d:)     �    ��  �E�    H�\:) H���   ���   �E�9���  �U��E�Ѕ���  �U��E��H�%:) H���   ���   �   )����H�E�@�E��E�    H��9) H���   ���   �E�9��*  �U��E�Ѕ��  H��9) H���   H���   H��9) H���   ���   �E��ȋE�ȉ�H�� <�u*�U܋E�ЉE�Љ�H��    H�E�HE؉�  H�Y9) H���   H���   H�D9) H���   ���   �E��ȋE�ȉ�H�� ���b  H�9) H���   H���   H� 9) H���   ���   �E��ȋE�ȉ�H�� ���*��Qd �^��E��U܋E�ЉE�Љ�H��    H�E�HЋ �E��E�%�   �E��E���%�   �E��E���%�   �E��E��*�f(��YM��*U���c �\E��Y��X��,��U��*�f(��YM��*U���c �\E��Y��X��,���	��E��*�f(��YM��*U���c �\E��Y��X��,���	ЉE��U܋E�ЉE�Љ�H��    H�E�HE�����E�������E��D���H��7) H���   H���   H��H�]���UH��SH��xH�}��u��U���D��D�ʈE��ȈE��ЈE��J7) ��tH�O7) H��tH�;7) H��u������#7) ���ub�E�    H�E�� ���  �}��u��M��U�D�E�E�D�A��H�E�� ��H���uA��A��D�։������H���E�H�E���E������E���	��E�	�   ��E�H�EH�@H�E��E�    H�E�� ����  H�E�� <
��  H�E�� ����������u
H�E��[  H�E�� H��H�J6) �   H��H�����  �Ẽ}� t2L��a �    �M̺    �    �    L���i��5)     �  �E�    H��5) H���   ���   �E�9���  �U�E��H��5) H���   ���   )ЍPH�E�@9��~  �U�E��H��5) H���   ���   )ЍPH�E�@�E��E�    H�i5) H���   ���   �E�9��  H�J5) H���   H���   H�55) H���   ���   �E��ȋE�ȉ�H�� <�u-�U��E�E�E�Љ�H��    H�E�HE܉�  H��4) H���   H���   H��4) H���   ���   �E��ȋE�ȉ�H�� ���e  H��4) H���   H���   H��4) H���   ���   �E��ȋE�ȉ�H�� ���*���_ �^��E��U��E�E�E�Љ�H��    H�E�HЋ �E��E�%�   �E��E���%�   �E��E���%�   �E��E��*�f(��YM��*U��g_ �\E��Y��X��,��U��*�f(��YM��*U��8_ �\E��Y��X��,���	��E��*�f(��YM��*U��_ �\E��Y��X��,���	ЉE��U��E�E�E�Љ�H��    H�E�HE���E�������E��1���H�"3) H���   H���   H���E�ЉE�H�E��c������H�]���f�UH��H��H��H��fof H��H����H��]�UH��H��H��H���o� H��H����H��]�UH��H��H��~2fHn�f��f��fs�f��fs�f��fs�f��fH����H��]�UH��H��H��L��H��~ fHn�f��f��fs�f��f H����H��]�f.�     f�U�`�F H��S���F H��D  H��H���\�  H�3H��u�H��[]�ff.�     f�USH���p�F H��  ����H���I  ����>  fD  �� �?  ��	�6  H��1��%�    ��:t#�LH��H��H���   �  �Hc���u��D< �>:��   H9���   H��1�H���&fD  ��=t%���   H��H��H=�   ��   �Hc���u�Ƅ<�    �9=��   H9���   H��1�H���!���	t'��  H��H��H=�   ��   �U Hc����u�Ƅ4   �E ��t<	u8H9�t3H��$  H��$�   H��H�t$�D  �}  t�UH�E�������H�Ę  []�fD  H���� ��   �������   �6�����   �D  AUATI��USH���C H��tiL��H��H���r  A�Ņ�uDI�,$���F �`�F fD  H��H���T�  H�3H��u�I�<$����H��D��[]A\A]�D  H���hC ��fD  H��A�   [D��]A\A]�ff.�     �H��tSH��C  H���*C 1�[�fD  �!   �f.�     H�71�H���t# H��H��H��H)�H�
H���u��D  �ff.�     @ Hc��H��H��H)���H�H��H��H)�H��H��H��H����H�H��H��H)�H����H���     �9����     ATUH��SH��L�f H�|$H�|$�V�M1�H��I���     H�;H��t'H�t$�U��uH��I9�v�E��I��H�;H��u�H��H��[]A\�D  ATI��UH��SH�FH��H��tH����I�D$H�@xH��tH����H�sPH�EH��t	H����H�EH�CP    H��H��[]A\���     H�wPH��t\HcGHH��H��@ H��H9�w;H��zcinuu�D�BA�� 
 t	A��   u�H���   1�� H��xcinutH��H9�v�&   �D  H���   1��fD  SH�7H��H��t
H�G8H���PH�    H�C    H�C0    [ÐH���   HcNH��H��H��?H�� �  H���   H��H��H��?H���H�FH��H��?H�� �  H�����H�H�F H���   H��H�H�� �  HcVH��H�� H���H�F(H���   H��H�H�� �  H��H�� H���H�F0��     ������f9|�����ff.�     �H�6H�?�8t1��H�����������H���ff.�     f�H�H�USH��  ��|�   f.�     L��H��H��  Z I��H��H��  ��|�H��1���� A�   � f�H��L)�M�H)�M�H��t4H�,� �F �HO�M�I��I��H��y�H��L�M)�H�M�H��u�H�[L�]�H��  - �&f�H��H��H��  Z H��H��H��  - �I���k���H��I���`����L�H�USL��H��I9���   H9���   I�ӻ  Z H��1���� A�   �$fD  H��M�L)�H�M�H��t4H�,� �F �HN�O�I��I��H���H��M)�L�H)�M�H��u�H��xQH��L�H���H�[]�1�H9�}�H��H��  ��L��H��I���l����H�һ  � H��  L�I��HN�H���M���f��   L�H)�H��H���H��H�[]�D  L�L��   D��D����M��AI���M��AI�	��҃�)эB�����I��I��L�L��@ �   )�I��I��L�L��@ H���  H��A��H����A���   H����   AWE��AVL�wAUI��ATI��USH��H���GD�L$I�,�I9�r�&�    I��L9�vI�H��H� H�x�������u�L9���   I�>H�H�@@H��tq�8�F ��H��teE��t8H� H��tXI�>�L$H��L��[L��]A\A]A^A_��f��   �f.�     H�@H��tI�>H��L��L��[]A\A]A^A_��fD  �   H��[]A\A]A^A_�@ �!   �f.�     �   ��f�     H�H����   H�x(��HDx ��t`�B��    H�T��#D  H��H��xGH�� H��H��H�F�H9�t.H�H��y�H��H��x�I��I)�L��H��H��H��H�F�H9�u�1�ÐI��I)�L��H���ݐ�$   �f.�     SL�^A�ҋFM�م�t&H�9��8��8I��L�@$L��I��?H��H��I��M)�H�^�FI�؅�t&H�9��8��8H��H�p$H��H��?H��H��I��I)�M��uwH��ME�I�� I�� I���I���tTM��tO�G8��~HH�w@�P�1�H��� H��H�FH�� H���I9�uH�H�� H���L9�t,E��u'H�GH�� H9�uʸ   [� H��MD���    1�H��t�H�9[�ff.�     �L�WfE��teH�GI��H�8H�HI�H��I��I��I9�v0@ H�H9�HO�I9�LL�H�PH9�HO�I9�LL�H��I9�w�H�>L�NH�NL�F�@ E1�E1�1�1�H�>L�NH�NL�F�fD  ATI��I��UL��H��SH�� H���T���H�$�   H��   ���   H�t$H��   ���   H�|$H��   ��   L�D$I��   ��   �EI��$(  I��$  L�]����u(H��H��?I��?H��H��I��H�U@H�uHH�}PL�EXH��t\H�yhH���Qp��tE<uAI��$  H��tH�SH��u�)f�H�RH��tH�J�y ltuou�H��H�yhH���Qp��u�H�� []A\ø   ��f�     HcHcWSHcLcNLcFH��L��L��HcNH��H��?H��M��H�� �  I��?M��[H��I��?Hc�K�� �  H��H��H��?H�H�H�K�� �  H��Hc�H��1 �  H��H�H�H�G�@ ATUSH�oH�_H��H�H9�s I��@ H��tL��H���@���H��H9�w�[]A\�f�SH��H�wH�[�� H�G    �4���[H�H��H��H�H�GH��H��H�G�@ AWAVI��AUATI��USH���GHH�wP��~T1��    H�,�L�,�    H�E L���   H�EH�@H��tH����H��L��H��A�WI�t$PJ�.    A9\$H�H��tL��A�VI�D$P    A�D$H    H��[]A\A]A^A_�H�GH�F    H�H��tH�pH�w� H�7H�w��     H�H�VH��tH�PH��tH���    H�H��u�H�G� AWI��AVAUATUSH��H�H��t6I��H��I��fD  L�cM��tH�sL��H��A��H��H��L���UM��u�I�    I�G    H��[]A\A]A^A_� H��H��H��?H��8�  f1��f.�     H����  f1��D  H��f1��f�     I��I�й   H��yH�߹����H��yH����I��H��yH����I�и���M��tI��L��1�H��H�I��H��H�ڃ��HD��@ I��I�й   H��yH�߹����H��yH����I��H��yH����I�и���M��tH��1�I��I��H��H�ڃ��HD��f.�     Hc�Hc�H��H��H��?H�� �  H��H��H��A�   H��y	H��A�����H��y	H��A��H�ٸ���H��tH��H��1�H��H�H��H��H��A���HD��H���G  H���>  LcHcNAWAVAUATLcfUHcnSLcLcOHcWL��M��M��L��I��L��M��L��L��I��?I��H��?I��O��* �  H�D$�I��?M��I��I��?L��J��; �  Mc�H��?O��3 �  H��I��H�D$�I��HcGHc�Mc�I��?H��L�J��" �  H��H�H�\$�H��Hc�H��M�� �  H�\$�H��?H��I��H��?M�� �  H��9 �  [H��( �  I��H��Mc�H��Mc�Hc�M�H�L�]L�NH�A\A]H�NA^A_H�F��    �ff.�     @ H����  L�GH�7L�OH�WIc�Hc�H��Lc�Ic�I��I��I��I��?I��?J�� �  N�� �  H���   I��Hc�Mc�L)���   I��H����   H��H����  I��I��J�1�H��H��H�GM����   I��1�K�I��I��H����   H��H�GM���a  I��1�K�I��H�H���0  H��1�J�I��H�G1��@ ��    H��H��H����   I��I��J�1�H��H�GM���r���I��L��1�L)�I��I��H��y?L��H��H�GM��y=I��L��1�L)�I���2  f.�     I��L��1�L)�H��I��L�OM����   I��1�K�I��H���/���H��H�H����   H��1�J�I��H��yH��H�G1��I��M��I��J�1�I��H��H�GM�������I��L��1�L)�I��I���:����    H��L��1�H)�I����    I��L��1�L)�I���i���@ H��L��1�H)�I��H���n���H�G1�ÐI��I��M��I��J�1�I������fD  I��L��1�L)�I��H������H�H������H��L��1�H)�I�������     �   �f.�     H���  H���  AWI��H��AVI��AUATUSH��H��(L�H�/L��H��L�L$�]���L�sM�cL��H�$L��L���C���H��M�{L��H�D$L���,���L��M�kL��H��L������L�sL�L$L��H�D$L��L�������H�[L��L��H�D$H�������L��L��L��H�D$ �����L��H��L��I�������Hl$L�$$H�T$Ld$I�I�kHT$ M�#I�SM�sH��([]A\A]A^A_��    �ff.�     @ H����  SL�1�L�OL�WL��L�_H��������H��?H��L1�H)�L��H��?H�T$�H��L1�H�L$�H)D$�L��H��?H��L1�H�L$�H)D$�L��H��?H��L1�H�L$�H�L$�H)D$�H��H9�H��uH��H9�tH�H9�~�H��H9�HO�H��H9�u�H�����bH���Z  aL��M��L��I��I��M��H��M��H)�M��H��H��?M�H1�M�H)�K�H9�tH�H��H��2�   [��    1�[�@ H��H��A-  H���N�yA-H��H��H��H��H��H��H��xzH��1�H�7H��H��t�M����   I��1�I�0H��I��M����   I��1�I�1H��I��M��xyI��1�I�2H��I��M��xDI��1�I�L��H��I�������D  H��H��1�H)�H��H���|���f�     1��D  I��H��1�L)�H��H��I������fD  I��H��1�L)�H��H���@ I��H��1�L)�H��H���P���f�     I��H��1�L)�H��H������f�     H��t{H��tvAVI��H��AUI��ATUSH�/H��H�6H�������L�kI�sL��I��L������H��I�sL��I��M�����L��I�sL��H������L�#H�H�k[]A\A]A^� �ff.�     @ H�H�WA�   A�ɉЅ�y	A��A�����A�   ��y
��A�������E���T  ���<  AUATUSA9��U  ����D��ھ����A��1����A��H��I9�@�Ń�A)�E���@  D��A����A9��  D����¹   )�f�     A�ȉ�E����A����E��D��A��A��D��A�A���  AI�D��   A����	��A�Յ�D����  DI�A��D����  �D��H��H��A���HD�H���H��H��A���HD�E����H�WD�D����  AH���   E���~   A�L$��   []��D��A\A]����@ A��D��Mc�L��f���tA��Mc�L�_���    D���������@ ����D������@ ��)�A������������     ��)�[]��A\A]� H��1�H��H)�H����H��?)��fD  I��H�L�I��?L1�L)�I��I��?L1�L)�H9���   H�4vH��H�H��H��?H1�H)�H��H��?H1�H)�H9�~kH�IH��H�H�H1�I��L��H��?I)�I1�I)�M9�~#K�@H��L�H�H)�H��H9������@ K�IH��L��� H�<H��H��v���H�RH��H�� H��t{H����   �Gt<H��  H�H��   H�FH��(  H�FH��0  H�FH��8  H�F 1�� 1�1�H�F    f�1�H�F    f�VH�F     �f.�     �#   �f.�     �   �f.�     H��tk�GtEH��p  ATA����UH��SH����   ��ufD��@  H��t'H��H  H�U []A\��    H��t+H�    1�Ð[1�]A\�f�     �#   �f.�     1��ff.�     f�H��t1��Gt��Q  ƇP  �D  �#   �f.�     1��ff.�     f�H��tH���   H�H�@@H��t�C�F ���1��ff.�     f���ff.�      �G    H�G�GP    H�G`H�G H�GhH�G(H�GpH�G0H�GxH�G8H���   H�G@H���   H�GHH���   H�GPH���   H�GXH���   �f.�     USH��H��H�w H�/H��tH���UH�s(H�C     H��tH���UH�s0H�C(    H��tH���UH�s@H�C0    H��tH���UH�sXH�C@    H��tH���U�C    H�C�CP    H�C`H�C H�CX    H�ChH�C(H�CH    H�CpH�C0H�C    H�CxH�C8�C    H���   H�C@Hǃ�       H���   H�CPHǃ�       H���   H��[]�ff.�      USH��H��H�/�����H��H�EH��H��[]��ff.�     f�H��t��f�     �ff.�     @ H�GH�O �G`    Ǉ�       H��HG(H��H�GpH�G0Hр H�OhH�OH�HH�GxtH�G@H�HWHH���   H���   �GPH�@H��HGXH���   �f�     H��tS�O�Wb�G`fG�f�W���   WPf��~&H�Wx�p�H�BH�4p�
fD  H��f
H��H9�u��,���@ ��    H��tsAUI��ATUH��SH���GH�_ ��t2��L�d��     H�3H��tH���UH�    H��L9�u�I�] H��t	H��H���UI�E     H��[]A\A]�D  ��    H������H�H��H�B�    HD�H���ff.�     @ H�����U���H�H��H�B�    HD�H���ff.�     f�H�����   ��t�fD  H��p  H���  H��`  H9�I��LM�I9�LL�L)H9�HO�H9�HO�H��h  H)WH��x  H��X  H��H9�HN�H9�HO�HwH9�HL�H9�HL�HW�H��h  H��x  H��X  H9�I��LM�I9�LL�L)H9�HO�H9�HO�H��p  H)WH���  H��`  H��H9�HM�H9�HL�H)wH9�HO�H9�HO�H)W��     �   �f.�     �   �f.�     H��t[�   H��tVH��   H��X  H�VH��`  H�VH��h  H�VH��p  H�V H��x  H�V(H���  �f.�     �!   �f.�     H��tSUH��SH��H��t5H��H�?H��u�(H��H�;H��tH��茤����u�H�CH��[]�D  H��1�[]��    1��D  H�w@H�WH�OP�GT    �ff.�     f�������f.�     H���wT�   �o���ff.�     @ H��t;ATU��SH�G0H��L�g8H��t�Ѕ�uI�D$H��L��[]A\��fD  []A\� �ff.�     @ H��(  H��tL�P��tDSH���   H��H��tH�GH���   H���PH��(  �PHǃ�       ����P[�fD  HǇ�       �ff.�     �ATUSH�GH��H���   H�EL�eH���   H��t��H���`���H��(  H��tH�E H� ��tL��A�T$Hǃ(      []A\�H�>H��t�s���H��(  H�    �� ���   ltuo��  AWAVAUATUSH��(H����  H�H�RH��I�Ճ�?��?H��I��H��I��I��A��H���   H�t$�����H�L$H�|$H�T$ I��I����?��?I��I��H�L�I�M�H�L$H�$H�D$H�|$H�ƃ�?H��H�H�H�փ�?H�D$H��L�N�.H�T$ A���)  A����  A�   A���G  H��?H��?L�$H��H��H��H��H�4L�I�H��J�'I��L)�I)�A����   H��A��u
O�IA�   H���  A���   ��I�� ���E���   A�   @��A���   	�H�� ���E���   ��fE���   	�H���  E���   A���   ��H��([	�]A\A]A^A_�fD  �   �f.�     E1�1�E1�1��i����H�@A�   H�xH����M���f�     �   H�|$L���^���H�L$H�|$A�   H�D$H�T$ ������    H�� H��H��I��H��I��L$H�I9�t~H��L�R H��H��L��L)�H��H��L�L�H9�twI��I)�H�xA�   H��H����� �   H�|$L������H�L$H�|$A�   H�D$H�T$ � ����    ��?��?H�D�H��/I���h���fD  ��?A��?J�|�H��H���n���D  I�p�9����    H�QA�   �P���f�     UH��SH��H������H���   H��[]ÐH���   USH��H�WH���   H���   H�hH��t"H�AH9�u�T H�PH9�tH��H��H��u�H��[]�D  H�QH�G(H��H��t��H������H�EH��H��H��[]��@ �H���   ��ff.�      AVAUI��ATUH��SH���   H��L�bH��tH���   ���	@ �+���H���   H��u�H��tH���   L��H�꾀G@ ����Hǃ�       H�C`H��tH����H��H������I�D$hH��tH����L���   M��t!I�D$0L�kM�t$8H��tL����A��   tCH���   H�EHǃ�       H��tH����H�EHǃ�       H��H��[]A\A]A^��@ L��L��A�V�@ H��tcH���   �@0    H��tXH�H�H�NH�HH�NH�HH�NH�HH�NHNtR�@0   H��tdH�2H�zH�p H�x(H�JH
t�H0��    H�    H��H�@    H�@    H�@   H�>   u�H�~   u��f�     H�@     H�@(    �ff.�     @ H��tH���   �@x1��D  �#   �f�H����   ATUSH���   H��twH���   �Px�J��Hx1���~	[]A\�@ H�M H��u�MD  H�IH��t?H;yu�L�eH��H��H�} �v���L��A�T$H��H��L������[1�]A\�f�     [�#   ]A\�fD  �#   �f.�     H����   AUATUSH��H�/H����   L���   M����   H���   H��u�[ H�IH��tOH;yu�M�l$H��H��H���   �����L��A�UH9��   t:L��H��L�������1�H��[]A\A]��    H���$   []A\A]��     H���   Hǅ�       H��t�H�@H���   �@ �$   �f��#   �f�     �"   �f�     �Gt���u���|���@ �#   �f��   �f.�     H�WH�GI��I)�H��y
H9�HM�I��H��u&H�gfffffffK�@H��H��H��?H��H��H��H)�H�W H�OH�w8H��H��?H�H��H��L)�H)�H��H��?H�O(H�H��H�G0�H��Hw@H���   H�VL�NL�B I��fD�AM�A I��fD�A�G��   ���   H��xIH����   H��H��H��H�1�H��H�A M����   H��I��1�H��L�H��H�qH�A(�2���f�H��  �H��tH��H��H��H)�1�H��H��H�A M��xv����H��t^�f.�     �H�A    H�A(   ��L�I0H�H�A8    H�A@H�QH� L��H�A ���H�   ����H��?H!�H���H�A(H�q�����H��  �H��t�H��I��1�H��L)�H��H�qH��H�A(�b���f�AUATUSH���   H�GL�c��t&D�.H��H��H�~L�FA����  D���$�@�F �H�{ H�C    H���H�CH    I)�A�L$8���H�H�C    H�C(   []A\A]� D���   ���   H���   A)�Mc�H��H��?H1�H)�L��H��?I1�I)��AI����t&H�9��8��8H��L�P$L��I��?H��H��L)�I�ӋAM��t&H�9��8��8I��H�H$H��H��?H��H��H)�I��H���P  M����  ����H��tH��L��1�H��H��H�H��H��H�K M���X  M����  ����M���	  H�{(A���   E��tfH�{ L�C(�!�H�{ L�C(H����  L�C L���     ���   Hc�Mc�H��L��H��L��H��?H��?L�� �  M��  �  I��I��I�� I�� L��H��I��I��fD�[fD�S[]A\A]�J���f.�     ���   ���   )�Hc�I���b���D  ���   I���h����H�uxL���   H+uhL+Mp�5����     M��x[����M��tL��L��H��H��H�1�I��H�C(H�C L��L���Y���I��������H�K(H��L��L���>���I������fD  H��  �M��t�L��L��H��H��H)�1�I��H���f.�     H��  �H���;���L��H��H��H��H)�1�H��H��H������H��  �M���/���L��L��H��H��H)�1�I��H��H������M���G���H�{(I���;��� L��L��1�H��H��H�I��H������� H9�}H�K(H��I������@ H�{ I�������1�E1������f.�     H��tK�GtE��x19w8~,H���   Hc�H�@H���   H��t2H���   ��f�     �   �f.�     �#   �f.�     H���g���1�H���H��t[H��tfH�~ x_H�~ xX��   ��wASH��H��H���   H�GPH�@    H���   H�@H���   H��t*��H��[�f��#   �f.�     �   �f.�     H�CH����H��u@�t,�   ��u�H�L$H��������u��t$H��������@ �#   �f�     H�������1��y����H��(H��toH��HDָ@   H��@HL�H��@HLЅ�t7E��DD�H�t$H���$    H�T$�L$D�D$�����H��(�f�     E��uA�H   �H   �fD  H���D���ff.�      H��(��t(��Dց���  ���  G�������  G����@ ��u1�@   �@   H�t$H���$    H�T$H�D$    �0���H��(É���    H���g  M���n  H���   I�     I�@    H�@H���   H���,  ATA��L��UL��SH���Љƅ���   A����   L���   HcE IcQ H��H�H�� �  HcUIcA(H��H��Hc�H�M H�H�� �  H��Hc�I��H�}A����   A�Af��w6H��H����   H��G�z�GL�PL��H��L��H)�H��H�H��H�M A�Af��w2H��H���   H��G�z�GH�xH��H��H��H)�H��L�I��H�� I�� H���I���H�M L�E[��]A\� 1�[]��A\��    1���� �#   ����     �   ��f�     H��G�z�GA�   I)�L��H��I)�I��I�I��I���x���f�H��G�z�G�   H)�H��H��H)�H��H�H��H������ H��tkH��tvL���   I� H�@@H��tsAUI���O�F ATI��U��SH��L��H����H��tH� H��L���L��H��[]A\A]��D  H���   []A\A]ø#   �f.�     �   �f.�     �   �f.�     H��tk��tG��cinutoH�GPH��tnHcWHH��H9�s"H�;ru�/�    H�9rt H��H9�w�   Ð�WH�   ��u�� H���   1��fD  �#   �f.�     �{��� �&   �f�H��tFH�H��t>�PH��~4H�pPH;>t+�J��   H���D  H��H9|��t��H9�u��D  1�ø�����ff.�     @ H��t+H���   H��tSH�PH��H���R;C r1�[��     1��ff.�     f�ATI��USH��H��t@H���   H��H��t1H�  t*�t$fD  H�CH�t$H���P ;E s�1҅�t
�T$�1�1�M��tA�$H��H��[]A\��    UH��SH���D$    H��tJH��H���   H��t;H�{  t4H�G1��P;C r�D$    H�T$1�H���?����D  �D$��t�1�H��t�T$�U H��[]�ff.�     ��t	H����   ��tz�N�E1�H��H��H��<@ H=fdcl��   H=deesutH�BH���   H��tD� ��AH��FtH��H9�t+H�H=kradu�H�BH���   H��t%�8�FpH��H9�u�1��f��Ft������    �Fp��f.�     �   �f.�     �   �f.�     H��tK�GtEH��t@H���   H�BPH���t/UH��SH��H��H��t&H�@H��t8H��H��H��[]���    1��D  H���   H�H�@@H��uH�BP����H��1�[]�@ �W�F ��H��tH���   H�BP��    H���   H�@P������ff.�     @ H����   H��tj��tf� ��H;G }c�GtUL���   I�@PH���tDU��SH��H��H��t\H� H��tH����H��[]���    I�@P����H���   []�@ �   �f��   �f.�     �#   �f.�     H���   H�H�@@H��t��L$�W�F H�$��H�$�L$H��tH���   H�FP�e����H���   H�@P�����t���ff.�     �H��tkH���   H�B8H���tZSH��H��tH� H��t$H��[�� H���   H�H�@@H��uH�B8����1�[Ð�b�F ��H��tH���   H�B8��    1��D  H���   H�@8�������    H��t[�GtUH���   H�H�@@H��tBU���w�F SH��H��H����H��tH�@H����H��[]���    H��1�[]��    1��ff.�     f�H��t[�GtUL���   I�H�@@H��tbAVM��AUI��ATI��UH���w�F SH��L����H��t,M��L��L��H��H��H� []A\A]A^��#   �f.�     [�   ]A\A]A^�f��   �f.�     �#   H��tv�Gt}L���   I�H�@@H��teAUI��ATI��U���w�F SH��L��H����H��t!M��H�L$L���H���PH��[]A\A]� H���   []A\A]��     ��    �   �f�H��t[H�H��tSH���   H�H�@@H��t@S���F H��H��H����H��tH��H�����uH�$H��[� H��1�[��     1��ff.�     f�H��tTSH��H��H�H��t;H���   H�H�R@H��t(���F ��H��tH��H�����uH�D$H��[�D  H��������H����f�H����   AUATUSH��H�_PH��tdH��t_HcGHH��I��L�$�L9�r�:f.�     H��I9�v'H9+u�H���J���H��t�H�I���   1��fD  �   H��[]A\A]�H���&   []A\A]ø#   �f.�     H��tTUHc�SH�,�H��H��H9�w�4@ H��H9�v'H�;�   u������H��u�H�H��[]�fD  H��1�[]�1��@ H��tH���   H��t	�xcinut1�� ATI��UH��SH��H�wP�H�g���H��t"H�PH���   D��H��[L�B(��]A\A��@ [1�]A\�f�     H��t@UH��SH��H��H�wP�H����H��tH�P��H��H�J0H����[]��H�������[]Ã����    H��t3SH��H�wP�H�����H��tH�PH���   H��[H�R8��1�[�@ 1��D  H��tKUH��SH��H��H�wP�H����H��tH�PH���   H��H�J@H����[]��f�H��1�[]��    1��ff.�     f�H��tKUH��SH��H��H�wP�H�#���H��tH�PH���   H��H�JHH����[]��f�H��1�[]��    1��ff.�     f�H��t+H�H��tH���    tH���   1���    �#   �f��$   �f.�     H��tEH��  H��tH�H��tH�HH�    H��t!H�A;p u�@ H�A9p tH�IH��u�1�� H��tH�
��    �ff.�     @ H��t-H��  H��t!H�B;p u�@ H�B;p tH�RH��u�1���f.�     AUATUSH��H��tQH��tL�GH�_I��L�,�L9�r�7�    H��I9�v'H�+L��H�E H�x�Ą����u�H��H��[]A\A]�f�H��1�[H��]A\A]�H������H��tH� H�@(H���fD  1�H���f�     H����   AUATI��UH��S��H��H�H�@@H��ta��H����tF��tBH�EH�X�@L�,�L9�s,D  H�;H9�tH�H�@@H��t
L����H��uH��I9�w�1�H��[]A\A]�@ �   1���    1��D  H����  H��t0�WH�GH��H��H9�sH;wu��    H90tH��H9�w�"   �@ AW��AVAUATUSH���OH�z�H9�v H�HH��H�H�H9�w�L�6L�fH��H�B�    L�nI�M��tI;�$0  ��   �uW�u3I�F8H��tH����H��L��A�UH��1�[]A\A]A^A_�f.�     H�SH��t�H�{ H�پpl@ �����@ I��$  H��u뚐H�mH��t�H;]u�H�CM�<$�xHltuot~I��$  H������L��A�WI��$  H��u�qf.�     H�@H��t^H�P�z ltuou�H�I��$(  H� � ����    IǄ$0      �����    �!   �H�{hH���u���H�@p�P(�i���1��D  E1�A�   ����f�E1�E1��u���D  A�   A�   �_���ff.�     @ H��t���  1�Ð�!   �f.�     H��t+D�OD�G�GH��tD�H��tD�H��t���     1�E1�E1���fD  H���=  ���  �P�1����  ���  AWAVAUATI��USH��(H�D�H�D$��F H�T$H�D$    H�$H�D$D��E����   H�$1�L�(��    H��D��A9�vOI�\�L�3M��tI�~L���À����u�A�t�H�C H��t�H�x�����H�C H��u�E�|$H��D��A9�w�H�$H�$H�T$ H9��s���E��t���L��I�t�����A�D$��u�H�D$L��H���PH��(1�[]A\A]A^A_��     �H�$H�$H�L$ H9�u��ø!   �@ H����������tH��u�f.�     ��H���8  �D  H��t;H�����F ����H��t 1Ҿ��F H���I���H��t� H���D  1�H��Ð1��ff.�     f�H��t{L���   �   M��t���   pmoct�D  9��   v��H�vH��LЋ0�2�P��PH�L$A��PA�H�PH�H�PH�QH�P H�QH�@(H�A1��fD  �   �f.�     H��t3H��t.H��t)M��t$;w s�GtH��p  H��  H��t��@ 1��D  H����  H����  AWAVAUATUSH��   f�? �^ L�v(��  H�G� f�D$f���7  H�T$E1�M��H�4$H�|$H�D$(    L�d$L�D$L��H��M�t$L��H��L�I�I�I�NH��H�L$HH�D$H��H��H��L)�L)�H�T$@L�L$@H�D$HL�T$HH�} H�uL�L$0L�T$8M�T$M�A�������  ����   H�$L�\$ H�|$@H�t$���ufI9���   L�\$ L��M��M��A�FL�����  <��   H�G��H�t$H��L)�H�D$pH�GH�|$pH��L)�H�D$xH�$�P��toH�Ĉ   []A\A]A^A_�D  ��H��H��C�L)�L)�������  H�H�H��H��H��?H��?H�H�H��H��H�|$@H�t$HI��I������f�I��L��H9��2���M��H�$H�t$H�|$@�P�  �    H�G H9��c  A�F��<�S  H�G��L�0H��L)�H�D$PH�GH��L)�H�D$XH�G H��L)�H�D$`H�G(H��L)�H�D$hH�$H�@L9��{  H�W0H�t$`H��L)�H�T$pH�W8H�|$PH��H�L$L)�H�T$xH�T$p�Ѕ������I��L�������     H�G��H�WH��H��H��L)�L)�H�T$0H�t$8L9���  H�G L� H�(��E�VM�fH��H��H��L)�A��L)�H�D$`H�L$hA���n  E���=  L�t$0�pfD  H�D$`H�T$hH�D$0H�T$8L9���   I��I���I��A�$H��L)��H�D$`I�wH��H��L)�H�L$h���   ����   H�T$0H�t$8H�H�H�|$0H��H�t$pH��?H�H��H��?H��H�H�T$pH�T$H��H�D$xH�$�P���N����j���f�     M��H�$H�T$H�t$@L���P���B���H�D$D�\$��D$(A����9���   H�|$H�D$(H�WH��H�D$(�<Bf�|$f��������    �   �����fD  H�|$@H��H�t$H�.���D  H�$H�T$H�t$`H�|$0�P�������M��L�������    �   �1����� �   �M��L�t$0����M��H�L$H�T$@H�t$`H�|$P�������    H��t[�wD�1���fD	�tN��~EE��~@H�1������D  �G9�~(9�~$H����A9����    9ֺ   E��fD  �   �f.�     H��tSH��tN�   �9uSH9�tFUH��SH��H��H�Wf��uXH�f��u7�C �U �����	ЉE H��1�[]�D  �   �f�1��D  ��    H�}H�sH��`w���fD  H�~H�sH���Gw��H�}H�SH�s�5w��� H����   H����   USH��H�/H����   H���F t=H�vH��tH���UH�sH�C    H��tH���UH�sH�C    H��tH���U�    1�H�C    H�C    H�C    �C     H��[]��     �!   �f.�     �   �f.�     �   ��f�     H��tH��t�!�����ff.�     @ H��t)D�GH�GE��~1� ��H0��HPH��D9�|�ÐH����   f�? ��   AW1�E1�AVUSf�H�WA��Hc�L�BH�GH��H��L��H�L��H��H�H9�s,H�L�ZH��H��L�pL�xL�r�L�z�H�XL�XH9�r�H�WH�
H�H9�s@ ��2H��H��@�p��JH9�r�A���A�JA��9��_���[�w ]A^A_�Ãw �ff.�      H��tH��t&H��t	�|���@ �   �f��!   �f.�     �   �f.�     H��tCH��h�BH�$�P��D$    ��v<u�D$   H��tH��t)H������H��h�@ �   �f��!   ��f�     �   ��f�     H��tH��t������ff.�     @ H��tH��t�a�����ff.�     @ AWAVAUATUSH�� H�$    H�D$    H�D$    H�D$    H���F  f� �;  H��I�������H�$H�D$H9��/  H�t$H�T$H9��  ��A�   I�k��H��E��Hǉ���H��H�	�1�����A)�DH�)���A���A)�DH�f����   I�C��L�m1�L�XM�$S1�fD  H�D��H��H��H�H�0L�pH��D��I��9�|UA��Hc�A)�H��I�H��I��H�M�fD  H�D��L�xH��H��D��I��H�L��M)�I��I��H�H��I9�u΍SL��M9�tI���r���f��   H��t@ 1�H�� []A\A]A^A_�H�� �   []A\A]A^A_�ff.�     H���   H��H��AWH��?AVH��?AUH�H�ATH��H��UH��SH��pH	�H�L$0H�D$Hu1�H��p[]A\A]A^A_�@ H�|$P������D$\����  H�D$Pf�8 L�p~�H�D$(    E1�M��E��H�D$PH�|$(E1�D��L�$$E1�E��M��H�@�D$X����H�D$    H�D$     D�x1�H�D$    I��D���tD  Hc�Hc�H�|$`D�L$H��H��L�L�H�
H�RH+H+PH�L$`H�T$h�=���D�L$A��M��tH�D$`H�|$hM��uR��H�<$I��M�ՍED9�AMĉ�9��  ;\$X�  ;l$X�u���H�D$ H�|$L�T$H�D$`H�|$hM��t��L$X��yH�$L�|$ �\$XH�L$L�l$Ic�Lc�H��H�L$@Hc$I��H��H��?H�T$Hc�I��H�T$8L��L��H��?M�� �  H�T$I��H�� �  Mc�H��Hc�I�I������  I��L�H�T$8H<$H�D$H�T$@I��   H��H��?H�� �  H��Hc�H��H��?H�� �  �T$\H��H����<  H)�H��H�$M9�Lc<$HcD$0Ic�MO�D�L$@I��Ic�H��H��H��?H��H�� �  H��?H��L��2 �  I��A9��   H�t$0L��L�D$8����L�D$8D�L$@H�|$HH�t$0Hc�H��I��L�<0H��H��?H�� �  H��A9���   I��H��H�|$L��D�$虸��D�$L�f�Hc�H��L�L:HB�SA9ى�AN�9�u�H�D$`H�|$h�����H�D$PH�D$(M��E�qH�L$(� 9����������f�     H�D$HL�|$0�@ H)�H�\$H�$�����    H�$H�|$L��D�L$8����D�L$8HD$H�S��� H�$L��L�D$8�Ϸ��D�L$@L�D$8�����H�|$P�   f�? ���������   ÐH��������     AVI�։ʹ   AUH��ATI�����F USH��0��À� �ۅ��4  ��txH�l$L�m�
   H�t$L���-n���E H�D$�8,��   L9���   H��L�pI9�u�L���
   H�t$��m���ǉD$,H�D$� ���   L9���   L�t$�A�~A�A�F����   ����   A�NA�v��xy��xu9�q9�mE�F9�eA���  w\E�NE�VA���  @��A���  A��D�u9���  w1A�T$@E�D$DA�D$HE�T$LA�L$PE�L$TA�t$XA�|$\��    �   H��0��[]A\A]A^�@ ���F �   H����À� �ۅ�uL����   �ϢF �   L���   ��� ��u�A�D$8   �   H��0��[]A\A]A^�f.�     �բF �   H����À� �ۅ�tD��F �   H����À� �ۅ�uX����   A����    H�A�D$`�.���f�     ��uLA�A�D$<����fD  A�>t"�   ������     �   �����fD  A�D$8   �����f�1��
   L����k��H��A�D$<���� �
   1�L����k���_���ff.�     �I���   ���F I����� ����tR���F �   L����� ����t'�բF �   L����� ����u\A�H<�
�@ A�H8�
�f�     A�H@�
A�HD�JA�HH�JA�HL�JA�HP�JA�HT�JA�HX�JA�H\�J��     �   �f.�     AWI��AVI��AUM��ATM��UH��S1�H��H�T$�ef.�     I�F(H��t1�1�1�L����H��u_I�F    A��    H��M�D� H��H�T$H��L��L��H�����F A��H��H��	t3H�E     M��u�A��    �fD  A��U   H��H��H��	u�H��[]A\A]A^A_� 1�H��t�Gt��0  �ff.�     H�7H�WH�G    H�G@    H�G(    H�G0    ��     H��tH�G0H��t���ff.�     @ UH��SH��H��H�G(H��t1�1���H��uH�kH��1�[]� H9ws�H���U   []�ff.�      H��xSUH��SH��H�_H�G(H�H��t"1�1�H����H��uH�]H��1�[]��    H;_v�H���U   []�fD  �U   �f�H�G�ff.�     AUATUSH��L�gI9�v=L�G(I��H��H��H��M��t8A��I��I�41�H�uM9�rH��[]A\A]��     H���U   []A\A]�I)�H�7H��L9�LF�H�L���Uh��� H��H��H�w�q����U1�SH��H�GL�OL9�s"L�W(H��I��H��M��t!H��H��A��H��HkH��H��[]��    I)�L9�LF�HL��H��L��L����g�����     SH��H��tH�( tH�6H��t
H�G8H���PH�    [�D  L�G(H�WM����   �U   H9���   AUATUH��SH��H��H��~lL�g8L��A�T$H����   H�sH�H��H��H���S(H�3I��H9�vXH��tL��A�T$1�Lk�U   H�s@H�H�    H�sHH��[]A\A]�@ H�    �   u�H�w1�1�A��H�3I��H�s@H�1�H�sHLkH��[]A\A]�D  H�O�U   H9�s*H)�H9�r"H�H�H�G@H�H�H�GH1�H�w��    ��    H�    �@   �`���ff.�     @ UH��SH��H��������uH�S@H�U H�C@    H�CH    H��[]�ff.�     �SH�( H��tH�7H��t
H�G8H���PH�    H�C@    H�CH    [�f.�     H�W@1�H;WHsH�BH�G@���     H�W@1�H�JH9OHv�H�������B�	�H�W@�f�     H�W@1�H�JH9OHv�BH�������B�	�H�W@��     H�W@1�H�JH9OHv��JH������	��J�	�H�W@�f�H�W@1�H�JH9OHv
�H��ȉ�H�W@ÐH�W@1�H�JH9OHv�H��H�W@�D  UH��SH��H��H�G(�    �D$ H�wH��tL�   H�T$��H��t�E U   H��1�[]�f.�     H�s�D$H��H�sH��[]��     H9wv�H��0�ڐUH��SH���    H�wH�FH;GsKH�G(H��H��tW�   H�T$��H��u-H�sH�T$������B	�H��H�sH��[]��    �E U   H��1�[]��     1�H��Ht��@ AVI��AUM��ATI��USH��H��0H�F(H����  1�1�L��H����H����  L�c�   L��H��H�T$�D$    �����ŉD$���4  �|$ �k  �D$���^  �T$���Q  D�L$E���B  �L$�����t$D�D$A�����Hc�	��D$I�u 	��D$��	��D$Hc���	��T$	��T$��	��T$H���D	�E��D	�D�L$A��D	�Hc҅���  H9���  H��H)�H9���  H��������L�I��M)�M9���  L�L)�L9��{  L�H�KH�H9��h  I�L�H9��Y  H�C(I�u H���  1�1�L��H����D�D$H���  L�cA���   L��H�T$ H��D�D$/�D$    �4����ŉD$����   1��   �   1��     �T ��E�:TE�H��H��u�	���   H�CH�hH�C(H����   1�1�H��H����H����   H�k1�H�t$H�߉D$�����l$��u1H��H��xjI�H�C(H����   1�1�L��H����H��u$L�cM�&H��0��[]A\A]A^�@ L;c�����H��0�U   [��]A\A]A^�f�H��H)�H9��X���H��0�   [��]A\A]A^�D  H;V�8����H;k�?����U   �;���L;c�t����ff.�     �UH��SH���    H�wH�FH;GsKH�G(H��H��tW�   H�T$��H��u-H�sH�T$�B�����	�H��H�sH��[]��    �E U   H��1�[]��     1�H��Ht��@ UH��SH���    H�wH�FH;GsSH�G(H��H��tW�   H�T$��H��u5H�sH�T$��J�R����	�	�H��H�sH��[]��     �E U   H��1�[]�1�H��Ht��@ UH��SH���    H�wH�FH;GsCH�G(H��H��tG�   H�T$��H��u%H�sH�T$�ȉ�H��H�sH��[]��    �E U   H��1�[]�1�H��Ht���@ AVAUATI��U��SH��H��H�t$�b����T$��u	9�t�   H����[]A\A]A^�f�H�t$H���3����T$��u�H�CH�hH�C(H����   1�1�H��H����H����   H�kH�t$H���D$    �����T$��u�f��t�D��E1��,f�1�1�H��H����H��uNH�k�D$    A��E9��P���H�t$H�������T$���<�����t@H�CH�hH�C(H��u�H;kv�H���U   [��]A\A]A^�D  H;k�M�����@ H�t$H���;���H�ŋD$���y���H�t$H�������T$���`���Hc�I�,$�����    H��H�    H��tL�¾  �d���@ �Q   �f.�     H��H�    H��tL�¾ �4���@ �Q   �f.�     UH��SH���    H�wH�FH;Gs;H�G(H��H��tG�   H�T$��H��uH�sH�T$�H��H�sH��[]� �E U   H��1�[]��     1�H��Ht���@ H���G  H���N  AUE1�ATI��UH��SH�^H���s�H�W@�F�<��   ���$�h�F f.�     �C�L�L;EH��  �U   E��t:H�}( t#H�u H��tH�U8�D$H���R�D$H�E     H�E@    H�EH    H��[]A\A]��    �B�JH������	��J�	ȹ   f�     ��tH����H��K��s�L�@���/  @���  @����   H�H���s��F�<����H�U@1��1���f.�     ��JH������	��J�	ȹ   뀋1�H���s��� �1�H��ȉ��_����    �BH�������B�	ȹ   ���8����     �H�������B�	ȹ   ���������   H��������    �s�H���������k���H�U@A�   ����D  �����f�     ������f�     f�������     @��t L�������f��   �f.�     �(   ��K�L��s&�uT��t��2@�1�t��T�f�T��fD  H�2H�1��H�|2�H�|1�H�yH���H)��H)���H�։��H��|����2���1�T��T��i��� H��H��H������H�$H����     H��H��H������H�D$H����    H��H��H�t$H��H�$   H�D$    ����H�$H�T$�   H��H��yH�ھ����H��yH����H������H��tH��H��H��H�1�H��H��H�ڃ��HD�H���f�H��H	�u1��D  H��L�T$H�<$H��H�t$L���c���H���[���H�D$H��ÐH��t����fD  �ff.�     @ H���G  H���>  USH��H�H�OH��H�$H	�H�L$��   L�\$I��H��H��L������H��L�҉������H�$H���|   �[��H��H��   @H�T$H�� H����   �[��H��H��   @H�� ����   �M��   ��H�H�0H��?H�H��?H)�H)�H�Ή�H��H��H�3H�CH��[]�@ H��&$����H��H��   @H�T$H�� H��H���|���H��&$����H��H��   @H�� H�څ��t�������H��H��H�3H�SH��[]�f.�     �ff.�     @ H����   SH��H�H�OH��H�$H�L$H��tjH�|$ uH�H��H1�[H)��@ L�T$H��L��耘��H����v���H�$H��xM�[��H��H��   @H�� ��U�ۉ�H����[����    H��H��H��?[H��H1�H)��f.�     H��&$����H��H��   @H�� H�څ�~��K��   H��H����[H�H��H���@ 1��ff.�     f�H��H�<$H��H�t$�����H���fD  H����H�������   H����   ATUSH��H�H�H��H�$H	�H�|$tUL�T$H��H��H��L���]���H��A���R���H�<$H��xA�[��H��H��   @H�� E��xID��H��H�D$H�;H�E H��[]A\�D  ��    H��&$����H��H��   @H�� H��E��y�D�������ff.�      H��tH�7H��H�G    �����     �ff.�     @ H��H)�H= L�}f�H  hH= L�|�ÐH-  hH=  � �ÐUH��SH��H��H��~/�WH��H��tDH��1�H����U��H��1��E H��H��[]�D  1�H����Ѓ��E H��H��[]�fD  �@   ��f�     UH����   SH��H��H�T$�u����T$��uH�H�E H����[]�ff.�     f�AVAUATI��UH��SH��H��H���D$    �U��L��I���U��H�T$H��I�t�����T$��un�/   H��H���&T��I��H��tNI��H��H��I)�I�mI�V�eT��B�D3 L��H���T��H��H����S��H��H��[]A\A]A^�f�     � �� H��1�H��[]A\A]A^�fD  UH�ֺ�F H��SL��H��H�?����H��tH�E 1�H�    H��[]� H���@   []�ff.�     �UH�ֺ��F H��SL��H��H�?�����H��tH�E 1�H�    H��[]� H���@   []�ff.�     �AWI��H��AVI��AUM��ATI��U�
   SH���T��H=���wI�?H�pH�T$H�������l$��tH����[]A\A]A^A_�@ H��L��H���bR��H�H���c   �/rsrf�CI�I�E     �AWI��H��AVI��AUM��ATI��U�
   SH���S��H=���wI�?H�pH�T$H�������l$��tH����[]A\A]A^A_�@ H��L��H����Q��H�H��H�/..namedH�H�fork/rsrH�C�c   f�CI�I�E     �ff.�     H��t[H��tVUH����  SH��H��H�T$�{���H�D$��u&H�   
   H�H�J�B   ǂ�     H�U H��[]� �   �f.�     AVAUATUSH��H�    H���  H����   L�7I��H��H�T$�P   L�������D�l$H��E��uBL�p8��tIH�CH�SH�E    H�E@    H�U H�EH�E(    H�E0    L�u8I�,$H��D��[]A\A]A^Ð�u<I�V���   H�{  ��   H��L���ҋD$H�k ��t�H��u(A����    H�sH����� H�S�D$H�U ��t�I�VH��L��1���D�l$�w���@ H��A�   [D��]A\A]A^�f�H��A�!   [D��]A\A]A^�f.�     �D$   �fD  ATUH��SH��PH�t$(H�T$H�t$�D$   �y����Å�u@H�|$H��tIH�� �l���H�l$��H��tH�E0L�e8H��tH����H��L��A�T$H��P��[]A\��     H��P�Q   ��[]A\�AVH�ֺ�F M��AUI��ATUH��SH��L�'L�������H��tSL��H��H��H���2�����t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      AVH�ֺ�F M��AUI��ATUH��SH��L�'L���(���H��tSL��H��H��H��������t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      AVH�ֺ�F M��AUI��ATUH��SH��L�'L������H��tSL��H��H��H���������t&�D$H��L��A�T$�D$H��[]A\A]A^�fD  I�] H��[]A\A]A^��    H���@   []A\A]A^�ff.�      H����   ATUSH�� L���   M����   H��I�|$H�T$H���������unI�D$L�d$H���   �   H��tL��H����L�d$1�H�{  t�+���M��t1I�T$0I�\$8H��t�D$L���ҋD$��u�D$L��H���S�D$H�� []A\��    H�� �"   []A\�f.�     �#   �f.�     H��t+H��HH�t$H��H�D$     �$   �����H��H�D  �   �f.�     ATI��USH��H��H�GH��(  H���   �B�tIH���   H��tH���UHǃ�       H�T$L��H�������H���   �D$H��[]A\��     ���B���     H���'  H���   H���  AWAVAUATUH��SH��H��(L�hH�@H�T$H�pXL���z���I�ċD$��tH��tH�E     H��([]A\A]A^A_� I�\$H�T$�P   L���   �D$    I�GM�wH�$I�GL��I�$�����T$I������   I��$(  I�H� ��ttH�$H���   H����   L���ЉD$��uvH���   I�T$L���   H���U���L�e H��([]A\A]A^A_�@ �   �f.�     �#   �f.�     H�T$��   L��L�D$�i����T$��t!�T$L���E���L��L��A�U�D$�����f�L�D$L�0I� �D$    �4����     �D$�D����    AWAVAUATUSH��8���   =stibteA��H��(  H��H���BJud=ltuo�*  H��t6L��  M��t*M�EA;@ u�$  @ M�EA9@ �  M�mM��u�A�   ��E1�H��8D��[]A\A]A^A_�L�nD�vL�D$ H�L$H�D$(    H�T$D��L���������$  1�L���~�������   I��p  H�D$�EH�D$H�ڋt$L��I���   ��  A�ǅ�uEL�D$ H�L$D��L��H�T$�+�������   H��(  �t$L��PH���������  ��t�I���   脪��ǃ�   ltuoL��(  L��  M������� 1�D��H��L��A�PxA�ǅ������<��������   H�������H��  M��tI�EH��u����D  H�@H�������L�@A;P u�I��딋��   =ltuo�?����d���ǃ�   stibI���   �ȩ���f��� H��H��t(H�OH��tH���   H�z��H������f.�     �   �f.�     H���  AWAVAUATI��USH��(H���    �P  H���   H���@  H�߉�L���   A������H�{8��H�C0    H���H�Ch    )��Hp1����H�Hǃ�       I�E    I�E    I�E    I�E     ƃ�    I��$�   Hǃ�       H�Bǃ�       Hǃ�       L��0  ��ǃ�         ��   Hǃ�       E�Hǃ       Hǃ      Hǃ       ǃ�       H�Cp    H�Cx    Hǃ      Hǃ      @��t�����
������  @ E�M��t���  uI�D$%   H���  H�B��I��$�   D��H�����   ������  ���   ltuo��  A��A��A��   A��E����  Hǃ�       H�CPH���   ��    ujA�D$tbI��$�   H�CpH�z H���J  H��H��H���J  H�F H��H�CpH�CxH�r(H���E  H��H��H���E  H�B H��H�CxE����   M��$�   A�t$0��tvH�C���   H���   H�@H��(  H��t;W t'H��  H��u�   H�@H����  H�x;W u�H�GI�L$ L��H���PX��H���   L��$�4����$H��(  D�s�hH��u_@��uY���   =pmoctL=stibtE������u1���   @�����tH��(H��[]A\A]A^A_�r���f�1�H�߉$�â���$H��(��[]A\A]A^A_��    �#   ��Hǃ�       H�ChH���   �R���D  A��A��   u$I��$�   H�x H��V  H�������D  @�� ��  H�H�    ��  ��H�@@�����L$H����  H��D�\$�C�F H�$��H�$D�\$H�Ǿ/�F D�\$H�$��C��H�$D�\$H��t�z8t�|$�<  I�D$��(���I��$�   ����fA��$�   �	���I��$X   �����I��$h   �  �����D  L���������������A��A��A��   A��@�������L�CXH�C0L�S8H�{`L��H�SHH�D$H���I��L�T$H�4$H�s@H�B?I���H���I��I���E���  H�CHH�D$H�4$L�S@I�D ?L�T$L�{`H���H�sXH)�H�C0I�D:?H���L)�H�C8H�CPH�� H���H�CPH�ChH�� H���H�Ch�J���@ �#   ���H�H� ��������I�D$A��I��$�   A���tK@��uEH�B��D�\$D���@D�$H�����   D�$D�\$����u���   stib�����I��$�   D�\$D��H��A��M��$�   D�L$H��L��A�B0L�T$A�B0    �$I�H�@(�PL�T$D�L$���$D�\$A�B0�o����H��H��H��������    H)�H��H������@ H��H��H��������    H)�H��H������@ ��ltuo����@����   ���������   M�D$(M�L$ H���   �������1��    ��L��L@H��9�|������fD  H���h�������f.�     H�<$H+T$H�CHH���L�{`H�{XH�|$H)�L�S@H�t>?H�C8H���L)�H�s0�����L��L��$�4���A�t$0�$�=���1�����H���g  AWAVAUATUL��SH��M���]  H�G A��A��1�A�A��I������9���D9������   ����   E����   H���   H�@H���   H��t*A����   I��D��D����L���Ѕ���   <��   �   A��    uuA��   �   E��A��DD�Mc��"@ H���   I��H�ȃ�H�E H��A9�tPD���L���u�����u&I��$�   A��u�H���   I��H���� �   H��[]A\A]A^A_�@ A��tRH��1�[]A\A]A^A_ÐD���������@�������f�     �#   �f.�     �   �f�     H��D��D��H��[I��$�   ]A\A]A^A_�|���ff.�     �H����   H����   ;w ��   AUA��ATI��U��SH��H��H���   H�@H���   H��t<��t,M����   D��H���Ѕ�tN<tH��[]A\A]��    ������t�H��M����D��H�ߺ   []A\A]����fD  �   �f�@��u�H��H���   ��L��[�   ]A\A]隀��f.�     �#   �f.�     �   �f.�     H��t;U��SH��H��H���   H��tH�G�P;C �Ƹ    C�H����H��[]�p����#   �f.�     AWI��AVAUE��ATI��USH��8H�oH�_H�D$,�T$H�uHH��H��H�L$L�L$������T$,I�ƅ��0  L���   �|$ H���   I�$I���   tI�N   H�T$,��   H������I�ǋD$,����   M���   I�Gh    E��~<H�L$A�U�H��H��H��fD  H��I�h uH�8rcniuH�HI�OhH9�u�H�E`A�Gt����H����   �T$L�D$D��L��I�<$��I���   �D$,I�$����   H��L���[���H�EhH��tL����M��t	L��H���SM��t	L��H���SH�D$pH�     �D$,H��8[]A\A]A^A_�f�H��tsH��H��E1������H�EhH��u��f�I���   I�$L���=y����t<&t�D$,�f���@ H�D$pL�0�D$,��t�H��L��譂��H�EhH���N����S��� H�EhH���Z���1����Q���f�H���  H���  H���   H����   AWAVAUATI��USH��H��L�pH�    H���   H�T$I�vPH�������t$I�Ņ�t$M��t	L��H���U�D$H��[]A\A]A^A_� H�T$�   H���f����L$I�ǅ�tM��t�L��H���U� I�] H�T$�H   H���2����T$��u�I�EPI�FpH��tL���ЉD$��u�M�,$H���   L��M�o�����D$���c���� �"   �f��#   �f.�     �   �f.�     H���O  H���N  H�~ 
  �   �+  AWAVAUATUH��SH��(�GH�4$�D$���f  ��L�fH�_L�l� �D  H��I9�t?L�;L��M�7I�~�:����u�H�$�   I�VH9Q��   L��H��菶���E�D$�|$L�m �0   �D$    wxL�4$H�T$L��I�v�����H�ËD$��uXI�H�kL��L�kL�3�uq�tH��0  �tH�SH�$H�@0H����  H���ЉD$���?  �U�J�MH�\�H��([]A\A]A^A_�f�     ��    �!   �f��   �L�e H�T$�   L���D���I�ǋD$����   H�M��A�ƋBHH�S�C =ltuou@H�BpH�T$H�@H��t.H�shL���ЉD$����   H�T$H�BpH�@ H�CpH�BPH�CxI�_H��  L������H��  H��u�   fD  H�@H����   H�P�z ltuou�|$H��(  ��t	E����   H�3�|$H��H����������    M��ua�D$H�3�t"H�CH��t�xHltuouH�{hH��tH�@p�P(H��L��A�U�D$�����D$�{���L�/�D$    ����1��d���L��L��A�T$�|$�h���fD  SH��H��~�W1�H�������[�D  1�H����у��[�ff.�     @ SI��H��H��H��?H��H��?��H���uH��y�   A�H��L��[� H��tKH��tF�����
   H�H��H9�|�H��H��H��uNL�$H��L��1�A�RL�$H��I�������@ 1�M��t�L�$L��L��A�RL�$E1�L��A�H��[�H��L�L$L��L��L�$A�RL�$L�L$H��LE�H��ۃ�@�D���ff.�     AVI��AUATM��UH��SH��H��L�L$�D$    �����I�ŋD$��u
M��tI9�|A�$H��L��[]A\A]A^�D  L)�1�H��H��I��I�|- �>6���D$���     SH��E1�1Ҿ   H���GH�?L�L$� �[���H��H�C@�D$��uVH�sL�C �C�SH��Hs(H��H��H�spH�s0I�H�H�L�ChL�CH�SHH�J�4FH���   H�sxH���   H��[�AWAVAUATA��USH��H��(�G�WbD�L�/�D$    ��D9�w,�G�O`�W�A�1�D9���   H��([]A\A]A^A_�f��n������  �N  D��L�G A��   L�L$L��H��L��H�D$�W����t$H�C ����   L�C(H�T$L��L��L�L$�   �)����L$H�C(����   �{ �  H�s�C`�k�S�H��A�D9���   �    A��A���A���  ��   L�C0L��D��L�L$�   ����H��H�C0�D$��uWD�cH�KH�SL�C H��HS(H��H�SpH�OI��{ H�SxL�ChtH�S@H�HsHH���   H���   �������H��輊���D$H��([]A\A]A^A_�f�     H��(�
   []A\A]A^A_�@ �D$H�{0�i��� L�C@C�?�L- L��L�L$�   ������T$H�C@��u�H�T$I��J�<0H��H�4�42��Ls@L�sH�����    USH�����   �WGPL��D$    �1�9�wH��[]�@ �^L�GXH��L�L$����0   L�׉��_���H��H�EX�D$��uŋMP�]H�IH��H�H���   H��[]ÐSH��E1�H����   1Ҿ   H�P   �   H��H��C    L�L$H�C�F@ H�C G@ �����H�C �D$H��[�f.�     H���  AUATUSH��L�'IcT$H��~3M�D$PI;8t4�J��   ��H����    H��I9|��t��H9�u�H��[]A\A]�1ۍJ�fD  H��Hc�L�L$�   I��$�   M�l���F����T$I�D$P��u�A�|$H�SD�G�9�~8Hc�H���H���H��H�9�tI�D$PH�t�D9�u߃�L�.H��9�u�E�D$HI9�$�   t:H�E H���   H�EH�@H��tH����H��H���SH��[]A\A]Ð��    IǄ$�       �f.�     AWAVAUATUSH��(�D$    H����   H����   L�*M����   M���   H��H��I��H�t$H�7H�T$L�������I�ƋD$��ulH�E H�UI�^I�H�CI�VH��tH�t$L���ЉD$��uvIcUHM�EPL�L$L���   �JHc������H��I�EP�D$��uGIcUH�rA�uHL�4�M��tM�4$H��([]A\A]A^A_��     H��(�   []A\A]A^A_�@ I�H���   I�FH�@H��tL����L��H��E1��S�D$M��u��D  H���7  AWAVAUATUSH��L�/H����   M����   �    H�A    H�A    H�A    �A     ����   9���   �
   ���  wkA��H��A��H��1�L�L$E1�L���   L�������T$H�C��u&L�L$E1�L��1Ҿ   L������H�C�D$��tB�K H��H�������D$H��[]A\A]A^A_��     H���   []A\A]A^A_�@ Ic�L�L$E1�1Ҿ   L���.���H�C�D$��u�fD�{fD�#�K � �!   �f.�     AWAVI��AUI��H��ATI��USH��H���j���D$    I��H� H��tL�h1�H����[]A\A]A^A_�@ H�T$�   L���N����l$��u�I�L� L�h�C;s���C�D  D�c�����E1�L��L�L$�   L�{ �D$    C�$�ȉK����1��=���H�C �D$��uaE��tcA�D$�M��M�l��    I�$H��tH�8H����i��I�$H�I��M9�u�M��t
L��L��A�V�D$��u�C�P���D  ������M��u���f�����ff.�     ������f�     AWI��AVM��AUATUSH��H��8H�H�L$H�D$H�F(D�L$H����   1�1�L��H����H����   L�{H�t$,H���D$,    �l����T$,��ux�D�`A���  ��   1�E��G�   fD  H�t$,H���3����T$,f�D$��u:H�t$,H�������T$,��u%M9�tl��A9�tTH�t$,H��������T$,I�Ņ�t�H��8��[]A\A]A^A_� H;V�I����U   ���    �   ��f�     �   �f�     �T$H�L$xH��Iǃ�Hc�H�H��H���
  w�H�C(H���l  1�1�L��H����H��u�H�D$xL�{1�L�L$,H�|$E1��   �D$,    H�������T$,I�Ņ��3���H�D$xH�0H���  L��E1��    1�1�L��H����H����   L�sH�t$,H���D$,    �����L$,I�ǅ���   H�CL�pH�C(H����   1�1�L��H����H��umL�s�D$,    M���  H�D$xA����� I��H��L�}�H�0L9�~wH�t$,H���[����t$,f�E ��u'H�CL�pH�C(H���:���L;s�E����D$,U   M��tH�D$L��H���P�T$,� ���L;s�e�����L;{������#����|$ u{H�D$xH�|$1�E1�L�L$,�   H������T$,��u�H�L$x1�H�9 ~#H��H�|$H��I|H�L$xH�<�H��H9�H�T$p�D$,    H��T����D$,   �G����@I@ �   L���(���n����     AWAVAUATI��UH��SH��H��   H�L�D$H�L$`L�D$hH�$����A��tH�Ĉ   D��[]A\A]A^A_��    L�t$xA�   H��H��AVA�TSOPL�l$xAUH�L$xH�T$p�����AYAZ���  AVE1�A�tnfsH��AUH�L$xH��H�T$p�����A��XZE���y���L��H�L$xH�t$pH�H��I��I��?I1�L9��`  H�E N�,�H�D$H�C(H����  D�T$1�1�L��H����D�T$H���?  L�kH�t$\H��D�T$�D$\    �����D�t$\D�T$I��E���  H���M  H=��� �1  H�L$L��H��H��D�T$�.  D�T$��A�ƉD$\�:  H�C(I��H����  1�1�L��H����D�T$H����  L�kH�|$H�T$\L��D�T$�D$\    �����D�t$\D�T$I��E���v  H�sL��H��H��D�T$�߽��D�T$��A�ƉD$\�F  A���F I��~A�<$OTTO��F LD�L�L$1�L��L��H��D�T$�  D�T$A��H�t$pH��tf�H�$D�T$H���PD�T$E���L  H�D$H�T$xH� H�����fD  I��L�|$xL�t$p�D$\   I���h  M����  H�E E1�E1�H�l$H�D$�xf�     1�1�H��H����H��uqH�kH�t$\H���D$\    ����D�T$\E����  H=��� ��   ���� I�L$H)�H9���   N�d I�EI9���   I��H�C(K�,�H��u�H;kv�L�t$pA�U   M��tH�$D�T$L��H���PD�T$E�������H�D$H� H�    ����f.�     L;k�W���A�U   H�������E���[����    L�t$pA�	   � I�D$H�l$H�D$0H���o  H�t$0H�|$H�T$\����D�T$\I��E����  E1�� �  1ɾ   fD�@�   1�L�d$@I��L�t$(I��L�l$8I��H�l$HH���D$$   �e  �1�1�L��L�D$H����L�D$H���e  L�CH��H�t$\�D$\    �x����|$\���@  H=���H�D$�/  H�t$\H���n����t$\�����  ���D$\
   ��   H�T$H�J�H���    HF�;D$$�n  H�|$0I�uH9���   L��G�4/H��C�T/L��H��C�T/L��H��C�T/���1  H�UH9��I  A�/�L�mI��A�D/A�D/ A�D/ A�D/ A�D/ �D$$H�D$@H9��  H�,H9��  H�sL�H���'����D$\��u3I�D$L;d$8�  I��H�D$(N��H�C(H�������L;C������D$\   H�D$L��H���PD�T$\L�t$p�T����    A�   M���C��������@ A�   �}���L;k�d��� H�t$pA�U   �`���H�t$p�V���fD  L�t$pA�
   �����I�H������H�t$pA�	   �%���H�t$pA�   �����L$\���E����8���@ H�t$pH�����������H��H�|$0L��L��H�PH�l$H�D$\
   H9������I�uA��A�DH9�r�H��A�L�L$H��H��A�#�F A�DH��H��A�DH��1�H��A�7L���
  L�t$pA������M�������H�D$D�T$L��H���PD�t$\D�T$�����H��H��L��L��H�l$H�D$\
   H�PH;T$0�F���A�?�A�D?�Q���f�AWH��AVH��AUATUSH��  H��H�D$X    A��H��?H�D$`    A����  H����  E��E1��tE1�H�~  A��H�T$H�T$XH��H��D�D$(H�L$H�|$�O����D$T����  H�H�D$ �E ��p  L�](M���c  I���A  ��l  D�E0L�M8H��L��D��H�D$hPH�L$H�t$hL�\$ �������D$dA[[L�\$�  M��H�|$ H�T$T�   ������|$T���%  L�D$`I���   L�@H�� tH����g��L�D$`H�|$ xH1�L��������D$T���{  H�|$`H��$   �����D$T���]  L�D$`H��$   I���   I�@�t+A���   f��y
��fA���   � uA���   fA���   ��  A�P8���  I�@@�z�H��H�H H��$fD  H�x xIH�x xBH��H9���  H�� �f��y��f�H�pH��yH��H�pH�pH��yH��H�pf��y�1�1�H�@    f�Pf�0H�@    H�@    � H�D$     ��E1�H�\$X��Qtg��tb��Ut]H��t4H�C0H�k8H��tL�\$H����L�\$E��uL�\$H��H���UL�\$H�t$`H��tH�|$ L��荀���D$T�	  @ �|$( ��  �T$T��u��D$T   널H�D$�D$T   H�X�@L�$�L9���  E1��   �    D�E0L�M8H��D��L��H�D$hPH�L$H�t$h�����D$dAYAZ���������E��t1H����F �	   H�H�r��� ��u=�   tjf.�     M���������H��I9��'  L�;I�� t��E �b���E1�E1��_����    �   H�Ĩ  []A\A]A^A_�f�     L�D$XI�@(H��tZ1�1�1�L��L�D$0��H��uJH�t$XL�D$0I�@    H�L$H�T$H�|$�D$T    �  �D$T����  ���;��� L�����D$TU   H�\$XM��H���  H�C(H��tL�\$(1�1�1�H����L�\$(H���X  1���   H��L�\$(H�C    H��$   H��H�D$0�7���L�\$(����   ��$   
�$j  
�$r  ��  ��$!  �P��� ��  ��$_   �  ��"   �q  ��$s   �c  ��$s  L�D$H��L�\$(H�L$H�|$�Hc�H��H��H������L�\$(�Ѓ��  ����  ��U��  �D$TH�\$X���H���H���"���H�C0H�k8H��tH����E������H��H���U�����fD  �D$T�����D$T    H�\$XH������������E u�D$TU   H�\$X�f���E1�E1�����H��$   H�D$0H�D$H�UH��E1�L�D$0L�L$tL�\$@H��$�   L�0H��H��A�   H�D$h    蘯��1�1�D�l$(��L�t$8D��L�l$0M��I��I�����   F�D�tE����   J����   Ǆ$�      H����  H�T$hH��$�   L��H��$�   �������t<Q��  ��utH�t$hK�T� L��L�D$H�L$����H�t$hH��t<H�N0H�V8H��t!�D$LH��H�T$0H�t$�ыD$LH�T$0H�t$�D$H���R�D$���  �۹   E�I��I��	��   L��H�����F ��1ۃ�����@��uһ   �����L�D$H�L$1�H��H�|$L�\$(�_���L�\$(������f�H�|$`�}�������I���   H�|$ H�    H�@    H�@    H�@   H�@     H�@(    �@x   �@p���   H�D$L� ����H��u�M���v���f.�     I�G�q����E �4��������L�\$@H��$�   D�l$(A��L�t$8H�]HM���    H�u H��tL��A�VH�E     H��H9�u�M��H�\$XE���3����D$T    H�\$X������   ����L���z|�������H�\$XE1�����H�\$XH�������H�C0H�k8H��tH����E�������H��H���U�D$T����ff.�     f�H��t3H��HA�   H�t$H���$   H�D$     ����H��H��    �   �f�H���7  AWAVI��AUI��ATM��UH���P   SH��XL�?H�T$L�D$L��H�$�/���H�ËD$����   L�D$H�+L�sH�C    H�C@    H�C(    H�C0`H@ �D$   H�\$0M��tL��L���D$
   �����H�D$8H�$E1�L��H�t$L��������uI�$H�b����H��X[]A\A]A^A_�@ H�S0H��t�$H���ҋ$�$H��L��A�W�$H��X[]A\A]A^A_�D  �$H��L��A�W�$H��X[]A\A]A^A_�f�     �   �f.�     AWI��AVAUI��ATUSH��H��HH�H��L��H�L$H�D$��HO�H�FH�t$<H�$�=����T$<��uUH=1pytt]�D$<   I�G(H����  1�1�H�4$L����H����  H�$�T$<I�GH��H��[]A\A]A^A_�D  �T$<��u��f�H�t$<L�������T$<A�ą�u�I�GH�hI�G(H���c  1�1�H��L����H���>  A��I�o�D$<    �D$ ����  H��H������L�l$(1�H���D$' I��H��?H�D$�- I��1PYT�#  �|$ t	L9��K  ��;l$ �.  H�t$<L�������T$<I�ą��"���I�GL�pI�G(H����   1�1�L��L����H����   M�wH�t$<L���D$<    迴���T$<I�ƅ������H�t$<L��裴���T$<�������I�� DIC�B���I��I��H��H����  �D$'�0��� H�$I;G�X���f.�     �U   �P���fD  I;o�������@ M;w�N����U   �&���@ I��I��H��H���t  �D$' ����f�     ��   �����fD  L�l$(I��I�G�D$<    �   L9������H�ƺ   L)�L9������M�G(L4$M����   L�\$1�1�L��L��A��L�\$H���)���M�wH�|$H�T$<L���D$<    L�\$������T$<H�����k���L�\$I�wH��L��L������L�\$���D$<u^�|$' �#�F L��H��A�'�F �    L�L$L��LD�H��HN������D$<��������D  L9��V����z���f.�     H��t�H�D$H��H���P�T$<�������I��L�l$(�D$'����I��L�l$(�D$' ����ff.�     f�H��t;H��HH��L��A�   H�t$H��H�T$H���$   H�D$     �����H��HÐ�   �f.�     A�   ����D  AW�   AVAUATUSH���D$   H��thH��tc�Gt]��0  9�vR��H��H  H��1�H��H��CL�sf��tM��tC���f�E �Cf�E�Cf�E�CL�u�Uf�E1�H��[]A\A]A^A_�f�     L���   1���E1�L���   L�L$�   L���8����T$H�C��udM�E(L�{M��tI1�1�L��L��A��H��upH�CM�}�KH��L��L���D$    軧���D$��u@L�s�S�6���M;}v��D$U   H��tH��L��A�T$1�H�C    1�f�C����H�C���D$U   H�C��ff.�     @ AW�   AVAUATUSH���D$   H��tfH��ta�Gt[f��8  �   uL�   �� �  v?�� �  ;�P  s1H��X  H��H�vH�,�1��E L�uf��tM��t��L�31��SH��[]A\A]A^A_�L���   1���E1�L���   L�L$�   L��������T$H�E��uJM�E(L�}M��to1�1�L��L��A��H��umM�}�M L��L��H�U�D$    �I����D$��t)H�EH��tH��L��A�T$1�H�E    1�f�E �F���L�u�U �9���M;}v��D$U   ��D$U   H�E�ff.�     f�SH��E1�H����   1Ҿ   H�P   �   H��H��C    L�L$H�CpF@ H�C`I@ �����H�C �D$H��[�f.�     H��t�g�     �ff.�     @ AUATI��UH��SH��H��~CI��H���WI��H��tJ1�M��uA�$H��L��[]A\A]ÐH��L��H������I����D  E1�H����Ӄ����     �@   �f�     ATI��1�UH��SH��H��tH�����H�PL��H��H��[]A\�N���ff.�      H��v:���t3H�T��@ ���t!H��H���G�H9�u�� 1��> ���D  H��1�� �> ��ÐH��t#H�H��tH;pu� H9ptH�@H��u��1���@ H��tH��t�U����ff.�     @ H��tH��tH�H�    H�FH��tH�0H�7�@ H�w��f�H��tH��t��T����ff.�     @ H��t1H��t,H�H��t$H�VH�PH��t!H�H�H�    H�FH�0H�7�f�     H�G��f.�     H����   AUATUH��SH��H����   I��A��H�˅�t
�   H��ttI��  I��  H��u�}D  H�vH��toH;nu��L����} ltuotsH�EL�hhE��t>E�a�I��I��I��D  H��L9�tH�SH�3H��A�Յ�t�H��[]A\A]� H��1�[]A\A]� H���   []A\A]��     H�EI��(  L�hhE��u���f.�     �!   �f.�     H��tKH��tFATI��UH��SH�?H��u�"f�H��H��tH�_L���Յ�t�[]A\�fD  [1�]A\�f�     �   �f.�     H��tH��t�AS����f.�     D  H��p  H�    H�A    H��tSH�����   H�H�1�[�f�1��ff.�     f�H�H���   H�@hH��t}H�L�BM��tqSH��H�� HcW`H�D$    H��H�$HcWdH�D$    H�xH�T$1�A�Ѕ�u'�$�{l Hǃ0      �C`�D$�Cdu�Cl�ChH�� [�f�     �ff.�     @ H��X  �   H�J
H9�`  rw������B	�f�G<�B�����B	�H��H�G@�B�����B	�H��H�GH�B�����B	�H��H�GP�B�����B	H��X  	�H��H�GX1��ff.�     @ HcG`H�w@H�HcOdH)�H���   H��H��H��zx(tXH�Gp1�H�Gx    H���   HǇ�       H��8  Hc�0  H��H  Hc�4  HGXH��@  H)�H��P  �fD  H��  H��t���)   A����.   H�Gp��H�Gx    H���   HǇ�       A��t�������Hc��s���1��l���@ H��pglh�s  vqH��srts�T  �.  H��oxps�1  ��   H��r  H��sxbs�  ��   H��x  H��oybs��  H��t  �    H��sybsHD��D  H��7psg��  �e  H��dlch��  �
  H��9psg��  ��  H���  H��csah��  H���  �    H��alchHD�� H��v  �    H��oxbsHD��H���  H��oyps�C  ��  H��|  H��syps�)  H�Ǆ  �    H��ortsHD��f.�     H��nrcv��   ��  H��  H��sdnu��   �S  H��   H��csav��   H��  �    H��focvHD���    H���  H��nrch��   ��   H���  H��srcht}H���  �    H��csdhHD��fD  H��2psg�S  vY1�H��4psg��  ��  H��5psg��  H��6psg�  f���  vH���  H���@ H��  ��     H��0psg��  �  H���  �    H��thpcHD��D  H�Ǫ  �    H��fochHD���     H��z  �    H��sxpsHD���     H��   �    H��odnuHD���     H��  H��csdv�S���v2H��  H��pglv�=���H���  �    H��tghxHD��fD  H��  �    H��srcvHD����    1�f���  �����H���  H���@ 1�f���  	�����H���  H�� �@ 1�f���  
�����H���  H��$�@ f���  �����H���  H���fD  f���  �q���H���  H���fD  f���  �Q���H���  H���fD  1�f���  �/���H���  �H���  ��     1�f���  ����H���  H���@ H��~  ��     H���  ��     H���  ��     1�f���  �����H���  H���@ H�Gǀ  ����1��ff.�     @ Hc�Hc�H��H��H��?H��    H���f����  ��     H���  H���@ H���  H���@ H���  H��@ H���H���   �@x��(t��#tHV(�
�fD  ��+   u�H��HV(H��HFH�
�f�     H���H���   �xx(tH��H��HFHHHV(�
�fD  ��+   tڀ�,   tр�-   u��� ��H��HVH
Ð��H��HVHJ�H��H��xHк    HH�� H)к    H��HO���     �Љ�%�   ��@t��   =�   �)  =�   �  H��H��H  �Ѓ�0����   ~k�� ��   ��0ucH�vH��H�HHI�H��
����   ��Hc�H��H��H�BHH�H��H��H��H��P  H��H  H��X  �f.�     1Ʌ�t�H��P  H����u��@�     ��udf����H����0H��H  ���S���H��H�NHI�H��
���g���H�V��w����    H��H��?H�H��	���@������    H��H  �����@ ���Hc�H��H  �����@ H��"  H��$  Hc�Hc�H��H��H�H��H��?H��    H��H���     H��  H��   Hc�Hc�H��H��H�H��H��?H��    H��H���     H���ff.�     �H���ff.�     �H��&  ��"  f�� @�N  ��(  L��$  f�� @��   H��H��H��I��H�H��H���  f�� @��   f��$   @�$  HǇ�  0	A f��   @��   f��    @��   HǇ�  p	A H���  HǇ�  �A HǇ   �A H= @  tkH�  H=�  wHǇ�   @  HǇ�      �fD  L���  f�� @�[���f��   @HǇ�  �	A �j���HǇ�  �	A �t���@ f��&   @tef��(   @u�HǇ�  0A HǇ   �A �}����    H��H���  ������     HǇ�  �	A ����HǇ�  �	A �����HǇ�  �A HǇ   �A HǇ�      �ff.�      H���  Hc��  H��  H���  H9�}-H���  ����  �� �F ���  ��xHc�H�H9�};�G�   �   �D  L�@L9�~��t��   )򉗜  Hc�H�H9�|�1��@ AWAVAUATUSH��H��L�6��  fD9��   �/  H�vH���  H�NH��H9��  f9WT�	  H��H  H��8  H�D$H���  ��  ��  I��H��X  H��H)�H)�HH�H9�P  ~H��H��M��HH�I��A��L���   H��HSXH��L�
L�RI�f��n   I��uM��&  D���k�����(  D��H�I�M��T���H�I�0I�H���   M�PI�xH�4L�
H�|L�RI�PI�0H��L)�L)����  H���   H��I����  L�H��HC`H�QH�1H+PH+0���  ��D   H��tL��L��H��L1�LH����  H����H����  @����   ��n  f9�l  uL��L��L)�L)�HH�H;D$MO�H�L$L��H�����  ���  H�L$��tM����   H9�HL�H)�A��H��H��H���   ���  ��  f��  ���  tfD��  fD��  H��[]A\A]A^A_�fD  ���   t��C�   f��  ���  t��fD  1�E1������fD  L��M��x(Hк    HH��D����    H��H9�HO��C����H)к    H��HO�����ff.�     �AVAUATUH��SH����  L�m M����  I��H�s8A�   �   �E H�����  H��H����<q��   L�F <rID���`  H�H��I9�tWI��M9�r=H����   H�C0H�~�H�{8H�T��f9STw����   H��t�I���C�   M9�s�H�s@[]A\A]A^�@ ��H�A�H��H�Ή�HI�H�*�b  H���   H��H��xx(tXH�sH��H�����  H�s8�`����    H���>����    ���   t�C�   1�H�C8    H�s@[]A\A]A^Ð��+   t���,   u6���   tf��(   ����L�Cp��H��A� ������e���D  ��-   H��������H�s8����ff.�     f������Ƈ�    H���   1�HǇ  �����ff.�     @ �Gx(   1��fD  �ff.�     @ H���  A��I9���   f���   L���  t<��M��LƋL�^ȉ�I��M9���   H���  H9�sb�    1���    �L��L�^��A���FD	�M�H��I��M9�wD�FE��D�FA��E	�E��H���  H�M�H9�r�L9�sH��I9�u�)Ɖ2� 1�1��2ÐL9�w�D����fD  �v�A���W��� USH��H�/���   �  H�G H�WƇ�    L�G(H�GhH�G0H�W`H�GxH�G8L�GpH���   H�G@H���   H�GHH���   ��   f����   �Obf����   H����P  ��   H���   Mc�I��H��H��?H�� �  H���� ���H�H�GxH���   I��H��H��?H�� �  H���� ���H�H���   H���   Ƈ�   L��L��H��?I��  �  H���� ���H�H���   @����   1�H��[]�@ Ƈ�   @��u�����f9�sIH�Spf���   H��H���   �@��Hǃ�      H���   ǃ  ����H�C`H�CX1���    H�Khf���   H��H��Hǃ�      H���   �H@��H���   ��    H�����   H������? �@���{b���   H�Ch��Hc��@��HcSh�KbH�CpH���   H��H�H�� �  �S`H���� ���H�H���   �����    SH��H�?H���   �Gu,H��p  H�S���   ��t�����H���   [�f�     �;\��H��1��q���1�[�ff.�     f�H��H��   �N���1�H����    �����   AWf�� @I�׸   AVI��AUM��ATI��U��S1�H���9@ 1�H��H��HN�H9���   H��HI�H9���   H����=����A9vP��I��H��t�I�vH�4�H��tcH9�t�f��t�I�<�H9�~PI�L� H9�}FH9�~)H)�H)�H�ǃ��=��A9w�H��[]A\A]A^A_�@ H��H)�H)�H��H���y���@ H��1�[]A\A]A^A_ø   ÐAWAVAUI��ATI��UH��S��H��H��&  H��u!H��(  H��uMH��[]A\A]A^A_�D  I�D$D��H���  H��I��N�48��<��I�T$H��(  I�N�4:H��t�I�D$H��H���  L��L�t��<��I�T$L�H�DH��[]A\A]A^A_�fD  AWAVAUATI��UH��S��H��H��&  H��t.H�D��H���   �@x��(��   ��#��   I�D$(L�H��(  H��tSH�E H���   �xx(u��+   ��   I�D$I��H���  H��I��N�l0�<��I�T$L�J�D2I\$(�H��[]A\A]A^A_��    ��+   �r���I�D$M��H���  H��I��N�48H�L$�;��I�T$H�L$I�N�4:�8������,   �`�����-   u��R���D  AWAVAUATUH��SH��(��  ��  ���  �  �_VD�_TH�WHD�PD�wRL�OXf�\$H�_hL�W`L�gxD���   H�\$H�_pH�\$fD9��%  H��T$H��fD�yf�QH�T$fD�q
H�Q H�T$L�QH�Q(L�a0fD�i8fD�YL�IfA� H��I�L�H�t$I�RI�2H+PH+0���  H���  H��&  H��I���v:��H�t$L��H�H��(  H���  �W:��H�E H��(1�[]A\A]A^A_�f����   D���   H���   D���   f�D$H���   D���   L���   H�D$H���   L���   L���   H�D$��D���   fD9���������   t�G�   1�fA� H��(�   []A\A]A^A_�f�     AWAVAUATUSH��H��(H��0  H9W ��   f��l   ��  �GT��   f9���   L�cXH����  I�Hk`f;��   �a  H��H��   H��A�   H�PH�0I+T$I+4$���  H�D$��  H��H��H��   H�PH�0H+UH+u ���  H��0  H�D$�   �    ���   H�C8��   Hǃ0     H�C@H��([]A\A]A^A_�f�     f��n   ����f��p   ����f9�s�L�ghH����  I�Ho`f;��   �  H�D$    E1�H�D$    H�C8H���s���H�S0H��H�C8L�<����   D9�wV���   ��   �C�   H��([]A\A]A^A_� �C�   �%���@ H�D$    A�   H�D$    �fD  D��I�$M�T$H��L���  E����   H��H��   H�L$H�VH�6L)�H)�H��A��H�L$I��H��   H��H�QH�1H+UH+u ���  1�I��M��tH�|$ L����   L)�A��H���   H�����  H�C8H��0  H�W�H��0  H��������D��� H���   L���  H�L$H���  H�H�2H�RI9�t_)�D)�Mc�Hc�Hc�Hc�I��H��H��H��H��?H��?H��0 �  H��: �  H��H��H��Hc�Hc�A��H�L$I���	����    L)�������     H�T$H�t$L��H�D$�I6��L�T$H������@ H���  H���  H��H��   M�$H�0H�PM�D$H���  H9�t[D)�D)�Hc�Hc�Hc�Hc�E1�H��H��H��H��H��?H��?H��> �  H��H��
 �  H��H��Hc�Hc���H�D$���� L)�L)�H��E1���H�D$����USH��H��H�oH�w0Ǉ       H�������H�C0    H���  H��H�C(    ����H���  H��Hǃ�      Hǃ�      ����H�C    H��H��Hǃ�      ǃ�      H�    H��[]�d���@ USH��H�/H��tvH�w0H��H���C���H�C0    H�s(H���/���H�C(    H�sH������H�C    H�sH������H�C    H�s H�������H�C     H�    H�C    H��[]�D  USH��H��H�H��  H���   H��t����Hǃ      H���  H������H���  H��Hǃ�      Hǃ�      �m���1�H���  Hǃ�      f���  �����H��   H���>���H��  H��Hǃ       �$���Hǃ�       Hǃ      Hǃ      Hǃ      Hǃ  ����H��[]�fD  SH������ƃ�    [�ff.�      AUATUSH��H��H�vL���   H��tl���tVE1�f.�     D��L��A��H�,@H��H�t.�t���H�CL��H�H�@    H�p�Y���H�sH�D.    D9#w�L���?���H�C    H�sH��tA�C��t*1�D  A��L���J�4�����H�sJ��    9kw�L�������H�C    H��[]A\A]�f�AVAUATUSH���  H����  L���   H�CI��H�sL��(����H�C    H�sL������H�C    H�s(L������H�C(    H�sL���p���H�s8H�C    H��tJ��t6D�m�1�I��I��D  H�t.L���;���H�s8H�D.    H��L9�u�L������H�C8    H�sHH��tLL���D���H�CHL��H�p0�����H�CHL��H�@0    H�p(�����H�sHL��H�F(    �����H�CH    H�sXH��tLL�������H�CXL��H�p0����H�CXL��H�@0    H�p(����H�sXL��H�F(    �s���H�CX    H�s`H��t8H��L������H�C`L��H�p(�F���H�s`L��H�F(    �2���H�C`    H�spL������H�Cp    H���   L������H��L��Hǃ�       []A\A]A^�����f�     []A\A]A^��    L�1�M9�r�D  ATI��L��UH��L��SI��H��   H��M�$L�L$�A���I�$�D$��uH�+H��[]A\�f�     UH��SH��H��H�7H�WH����  ���   ���  ���   ���  ��  ���  ��  ���  H��   H���  H��  H���  H���   H���  H���   H���  H���   H���  H���   H���  H���   H���  H���   H���  H���   H���  H���   H���  H���   H��   H���   H��  H���   H��   H��  H�BXH�H���  H�HH���  H�HH���  H�HH���  H�H H���  H�H(H���  H�@0H���  ��  ���  ��  ���  H��(  H��  H��0  H��  H��8  H��  H��@  H��   H��H  H��(  H��0  H��P  H�{PH���H��  H��X  H��   H��`  H��(  H��h  H��0  H��p  H��8  H��x  H��@  H���  H��H  H���  H��P  H���  H��X  H���  H��`  H���  H��h  H���  H��p  H���  H���  H���  H���  ���  f��8  H���  H��@  H���  H��H  H���  H��P  H���  H��X  H���  H��`  H���  H��h  H���  H��p  H��   H��x  H��  H�CH    H���  ��Hǃ�       )����   1����H�L�SHL�KPL�CXH�{`H�shH�KpL���   H�SxL���   L���   H���   H���   H���   H���   H���   L���   H���   L���   L���   H���   H���   H���   H���   H��   H�C(H�{�   H�K0H�t$H�D$���  L�@ ����H�T$H�S(���   H��[]��    ���  H�{�   H���  D���  H�t$H�D$�[����T$���  ��u�L��  L��  ǃ      L��  L��   H��(  H��0  L���   H��8  H��@  L���   L���   L���   H���   H���   H���   H���   L���   L���   L���   L���   H���   H���   H���   H��   L�[HL�SPL�KXL�C`H�{hH�spH�KxH���   ƃ`   H��[]�f�     AUATUH��S��H��L�/H���   H��H���   tIM���  Hc�1�1�L���  @ Ic�H��H��H��?H��0 �  H��H�I�ЍQH��H;��  r�L��  H��L��L���;�������  AƄ$`   A��$�  I��h  I�D$     I��p  AǄ$�      I��$  I��$   IǄ$(      IǄ$0      H����  1ɾ   ��  H�       @H�   @   @fA��$(  I��$   I��$  AǄ$l    fA��$p  IǄ$0     H��P  I��$   H��X  I��$(  H��`  I��$0  H��h  I��$8  H��p  I��$@  H��x  I��$H  H���  I��$P  H���  I��$X  H���  I��$`  H���  I��$h  H���  I��$p  H���  A��$�  ���   A��$�  I��$  I��$  ��  A��$�  ��  A��$�  H��   I��$  H��(  I��$   H��0  I��$(  H��8  I��$0  ��  H��@  H��H  H��[]A\A]�f.�     I��$�  L��I��$�  IǄ$�      AǄ$x     A���  ����f�     AWAVAUA��ATUSH��H��H�H���   H���   H�GL��  M��~���   H���   H���T���H���   H�SH��  H��P  H��  H��X  H��   H��`  H��(  H��h  H��0  H��p  H��8  H��x  H��@  H���  H��H  H���  H��P  H���  H��X  H���  H��`  H���  H��h  H���  H��p  E���!  H�RXH�JH�RH���  H���  ���   H��H�L�H�9H�W H���H�H�L�H�9H�W H���H�H�L�H�yH�W H���H�QH�T�H�BH�� H���H�BM����   �}x(�r  ���   H���   H��H�t�H�|�H�spH�{xH�t�H�|�H���   H���   H�t�H�|�H�T�H��8  H��@  H�H�RH��H  1�H��P  H��[]A\A]A^A_�f.�     H��  H�CL�ppD���  L���   L���  L��0  L��  L���   L��(  L��  L���   L��  L���   L��   H���   H��(  H���   H��0  H��   H��8  H��  L���  H��@  L���  HǇ�      Ǉx     L�_HL�WPL�OXL�G`H�whH�OpH���   H���   H��   �   f��p  H�H�WxH���   H���   L���   L���   L���   L���   H���   H���   L���   L���   L���   L���   H���   H���   Ǉl    Ǉ"   @  Ǉ&   @  Ǉ   @  Ǉ@     HǇ0     H�G     Ǉ�      ���  H��  ��t���   ������h  ��A
��A��}x(�����H��  1���+   �x���H��[]A\A]A^A_�f����   H���   Hǀ�     Hǀ�     H���C���H���   ������    ATH��A��UH��SH�_0H���p����t[]A\�fD  D��H���]r����u�H�S@H��X  H�SH[H��`  ]A\�ff.�      H�0�s���    AWAVAUATI��UH��SH��H��(L�o8�    �D$    �s��H�$��������   D���\  D��H9���   A�NL�L$E1�1Ҿ   L��豣��H�$�D$����   D�31�1�E��tD  L���Hs��H�$A�ǉ؃�L�,BE����   A��L��D$�s�����fA�m E��thH�4$D�l$��L�<FA��@ I��D9�t?L�����r�����fA�/A9�w�H�$H��([]A\A]A^A_� H�$    ��fD  D���X���A9��O�����D  A��L��A�ǉD$�r���fA�m E��t�H�$D�l$��L�<BA��@ I��D9�t�L����lr���fA�/A9�w��f���A��L���1r��A����A��A	�D��H9�������R���f�AW��AVAUATUSH��(H�G8�D$    H�D$H9��F  ��I��L�L$E1�1Ҿ   H���
���I�ŋD$���  1ۅ�tkD  L���q��A��A��?����   �@ue9���   E1�f.�     L��A���tq���KH��H��I�D� ��E9�r9�wى�E9���   9�r�H��(L��[]A\A]A^A_��     9�vtE1�f�     L��A���4q���KH��H��I�D� ��E9�r�9�w���    9�v4E1�f�     I�D�     �CA����E9�r9�w���g���fD  H�|$L��E1��8����Y��� E1��N����     H���  H��u��$  f��uH���  H���  H���fD  ��"  H���  f��uH���  H���f�SH�����  �������A������Hc�Ic����H���  [�AUI��ATUH��SH��H��H���  L�$��]���L��H������H���  L�H��H��[]A\A]�f�     ATI��UH��SH������H���  H��H��J�����H�[]A\�UH��SH��H�������H���  H�Hc�H��[]H��H�H�� �  H��H���    SH���������  [H�H��H�H�� �  H���f.�     AWAVAUATUH��SH��(D�<H��X  L��`  L�gE��E���  A�D$A�T$`�D�A;D$�0  A���  ��  M�D$xI��I�<@C�D?H�H�I9���  ������A	�E��~fA� f����  I�PH�YH9�vP�qH�Y��A���qD	�fA�pf9�|(�x  f�H���C������C�	�f�f9��W  ��H��H9�w�E����  D�z�A���4  D��A�L$A�D$b�D�A;D$�~  H�EL�SHǀ      Hǀ       M9���  ��[��	�D���E ��   L��L)�L9���  H��  �   M��H�t$L�T$���  H���  L�$H�|$H�x�&���H��  �L$���  ���w  H�EL�$f��H���  L�T$L��  H��   t%L��L��L�L$L�$�����L�L$L�$�     M�D$pM�Mc�O�M9���  I�qI9��  A�I�@A����o  L��L��L)�L)�L�I��' H�~I9���   �W�H���P����?  H��H9�u�I�|$hI��I�I9���   L9���  M�L$pH��E1�L���8f�     L�YM9�wm���	�;  I�L��L� H��H��I9��6  �2@��uȃ�u�H�qL9�w0D��IA��D	�H��I�H����    H�AM�D$xI9�s�   H��([]A\A]A^A_�fD  �L�������A	�����f.�     1�D��L��H�$�ߜ��H�$�������묐1�E1��k���fD  1�A�wL��貜�����l����H��L��f�L�NM9��i����7H��H�I9��W�������   ����L�DfD  H���P�L9�u������    I)�L��������   ����1��9�    H�qL9�������	� uJH)�H��H�W��H��I��A�A�I9�v4A��uƨ u�H�qL9������D��IA��D	�H��H�H���fE�|$b1�fE�t$`H��X  ����L�������I���_���H��(  H�8�����H���  AUATUSH��H��H���  L���   H���   L��p  H��t	H���  ��M��tH��A�T$H���   H���  ��g��L���   Hǃ�      H��   I�|$8�M���H��   L��Hǃ       �g��H���  L���$���H��`  H��Hǃ�      Hǃx      �g��H��p  H���pg��H��HǃX      Hǃh      �����Hǃ�      H��[]A\A]�@ ��    AW�ravaAVAUATUSH��(H���   L���  �D$    H�L$L�k8H��A�D$0��@  �D$��tH��([]A\A]A^A_��     H�t$H����f���D$��u�H���Si��H��H���Hi��H��H�D$H��   tH���?h��H��([]A\A]A^A_�I�D$� H9�u�H��L�L$E1�I�־   1�L��臘���T$I��I�D$8��u�M��t�H�$    f.�     H��Hc,$�4h����fA�H��    H;D$��   L�L$E1�1Ҿ   L���#���I�G�D$��up1�fA�? tJfD  H��I��H����g��I�OI��H��H��H��J�1�g��I�OH��H��J�D1A�9��H�$I��H�$H9D$�L���������E�I�t$8���t>Lc�H�$I����H)�H��H�� �J�t>L���þ��I�t$8J�D>    I��L9�u�L��褾��I�D$8    ����fD  AWAVAUATUSH��H��   L���  H�n8�D$t    M��t,H���   t"H��I��H�L$x�ravc��@  �D$l����   �D$l    H�D$    E1�E1�H�D$    H�D$    H�t$H������L��H�������H�t$H������H�t$H���ݽ��L��H���ҽ��H���   1Ҿ`A ������D$lH�Ĉ   []A\A]A^A_�f�     H�t$xL���Cd���D$l���O���I�G@L��M�/H�D$�f��H=   tL���D$l    �e���&���fD  A�$L�L$lE1�1Ҿ   H������D�T$lI��E��t0L��E1��Me��H�D$    H�D$    H�D$    �����D  A�$L�L$lE1�1Ҿ   H��荕��D�L$lH�D$E��t&L��E1���d��H�D$    H�D$    ����@ A�$E1�H��L�L$l1Ҿ   �=���D�D$lL��H�D$E���,  �e��L���T$ ��d���T$ H�t$x��A��fA���A�ÉD$L��H�H9���  H�D$L)�H�H�L$(f���/  H��x  E1�1�H��L�L$l�   D�\$ 謔��I�ŋD$l����  H�D$    D�\$ H�D$8    �D$     fE����  H�l$PH�\$Xf.�     L���8d��L��f�D$0�+d����f���  ��%�  A;D$h�:  I�L$pH���,  A�$L��H��H����H�4�������@�  H�L$L�D$��L��L���e���H���D$0HD$(H�D$0H���,  I�I�W@H�|$(H)�H�T$@I�WHH��H)�H�H9�H�t$xHG�I�W@�� �*  �T$tH�\$�T$p��uH�D$X��x  L��H�L$(����H��H���;  H���2  H�|$8��t$pH�L$(�9  �~�1�Hc�L�D$X��u�Gf.�     H���4SI;�x  s$HcL� H��I��I��?J��	 �  H��Hc�IL� H�JH9�u�H�t$8H�|$P�$���H�D$8    H�|$PH������I�GHI�H�\$@H��H)�H�H9�HG�I�G@H�T$0�D$ �D$ H�T$(9D$L�!���H�l$PH�\$XH��x  H��t(H���  1�1�I�D� H   H��
��QH��H9�r�L���a��H�|$��}����k���f.�     H�|$8��1���H�D$8�����;����D$l   L���va��E1�H�D$    �&���A�$�������1�f�\$@��H�l$ L���a���ك�H��H��H�D� A�$9�w��\$@�������1��H�l$L���ha���ك�H��H��H�D� A9$w��\$@�i���H�T$pL��H�L$(�4����T$pH�t$xH�D$8H��H�L$(����A�$1���%��� L��� a�����H��H��I��A9,$w������H�D$XH;�x  �����H�������L�D$XHc�1�1�D  HcT� H��H��H��?H��
 �  H��Hc�IT� �wH��I;�x  r�����I�WHI�D�\$0M�o@H��H)�I)�H�H9�L��HG�I�W@H�T$t�L���M�L�L$lH��H�D$I�G@K�*H��x  L�T$(H�D$ I�GHH��L)�L9�   HG�E1�1�I�G@�����t$lL�T$(I��D�\$0�������H�D$ L)�H�D$(�e���H�l$PH�\$X�D$l   ����L���U_��H�D$    �����    AUH��ATUH��SH��H��L�f8� tvcH�L$��@  �D$��t)Hǃx      1�Hǃ�      H��[]A\A]�fD  H�L$L�L$E1�1Ҿ   L��H��H��x  �B���H���  �D$��u�H��x  H��H�4 � ]���D$��u�L���  H��x  M�d� M9�sH��I����^�����A�E�M9�w�H���_^�����   �D$�U���H��H�������E���ff.�      AWAVAUI��ATI��USH��8H���   L���  H��H�k8�Z���D$,��t*E1�L��H��輵���D$,H��8[]A\A]A^A_�f�     H�t$,H���s_���T$,��u�f��t�D$,   � H�t$,H���+d��H�D$�D$,��u�H�t$,H���1_��D�|$,��A�U E���r�����t���L�L$,E1�1Ҿ   H���΍��D�\$,I��E���F���E�U E��tA1�f���H�t$,H�߉T$I��H�$�c��H�$D�L$,H�E���	����T$��A9U w�H�t$H��L��sY���D$,�������H�t$,H���z^��D�D$,fA�EE�������H��H�t$,�Z^���|$,��A�U�������I�VA�M;
t�D$,   ����E1�1��Ⱦ   L�L$,H�������|$, I�E�]����D$    �D$A9E��   D�t$I�EE1�1�A�ML�L$,�   H��N��L�$葌��L�$�|$, I�����I�EfA�} N�4���   �$    H�t$,H���]���t$,f�D$�������H�t$,H���i]���L$,f�D$�������H�t$,H���K]���T$,�������H�T$H���$I��H���$H��I�F�A�EI�V�H�T$H��I�V�9��k����D$�����A�M E1�1�L�L$,�   H��誋���|$, I�E�$����$    �$A9E �����$H��I�4�Lk�MuL��}W���D$,�������H�t$,H���\���|$, ��A������H�t$,H���f\���|$, ���D$�����H�t$,H���G\���|$, ��A�V�����;T$�����A;U�����E1�1��Ⱦ   L�L$,H���׊���|$, I�F�Q���1��:H�t$,H�߉T$��[���L$I�v�����|$, H��� ���A;E�������A�F9�w���A�E1�1�L�L$,�   H���e����|$, I�F�����1�A�A�F9�vPE1��>H�t$,H��D�D$�L$�T$�Y[���|$, ������T$I�vD�D$�L$f�VA��B�D;D$r��A�$�[���H�t$,H�߉L$�T$�Z���|$, �X����|$I�vf��L$f�~H������)�A9Fw����R���fD  AWAVAUE1�ATUSH��H�L��X  H��`  H�_H�<$L�` �   D  ��H�H9��9  A�N����  f����  A�v��	�I�v�ɉHA�N��A�N��	��ɉHfE���  �L�vE1ɉ��N��	�1�H��H��H�΃� H�HE��L�HH�x H�p(�/  E�}H��D������A������   I�~H9���   D��H�IH��H��   H�@    A�A�N��	�f�PA�v����A�v	������L9�}>��A�у�f��Ƀ����fA���������@��   ��H�H9�������    A�   H��D��[]A\A]A^A_��     ��@��   �L�vE1ɉ��N��	��~�vH����H��	�1�H��H�������fD  ��f����   A�v��	�I�v�ɉHA�N��A�N��	��ɉH�e���@ D�Q�IE������     �HA�NI�v�H�5���@ ���   �L�v���N��	��~H����H��A���~D	�D�NH��E��D�NH��A��E	�D�V�vM��A��I��D	�H��H������� �HA�NI�v�H����@ I��1��   E1ɹ   �����D���   H�$D�D$H�{0�GS��L��X  D�D$L�H)�H��   �O���f�     I���   �p�F ��� ����t�   ��    A�Hx�
Ð���   tH��p  ��   H��  ��f��h  �t6���  )�f����  ���  ����)�)�9�H�fA� �f�     ���  )�f����  ���  ��@ AWAVAUATI��US��H��H�G%  ���toH����   �   A��$�  t?��t9L��D�<L�t$L�l$���M��L��1�L���H�������D$H�E�D9�u�1�H��[]A\A]A^A_��     H��t{�   A��$�  tԅ�t�L��D�<L�t$L�l$fD  I��$p  ��M��L��1�L���H����  �D$H�E�A9�u��fD  �G��(����3���f�     �G��{����@ H���  H��t4H��t�8�>H��tH�pH�2H��tH�PH�M��tH�@I� 1��@ H��t�    H��tH�    M��t�I�     1��f.�     Hc�H��H�H���  H��t:H��   H9�|H���  1�H���  H���  ��x  ��G�   �   � �G�   �   � ���  H���  H��H��H9���   ���  �f�     H��(H9�vw:Hu�x t�Hc��  ;��  }e�JH���  H��I�����  ��x  H��  �
H�N�0H�JH�B   H�B�V���w)H�P� ���Aƀ�   ��    �G�   ��G�   ��G�   ���    H�B H��xH�    H���HH��fD  H)�    H���H��H��HO��f�     H��xH�2�    H���H�� HH��D  H)�H������H���H��H)�H��HO��@ H��xH��    H���HH��f�     H�к    H)�H���H��H��HO��fD  H�B?H��xH�    H���HH��fD  H)�    H���H��H��HO��f�     H�BH��xH�    H���HH��fD  H)�    H���H��H��HO��f�     L��P  H��X  H��H  L)�H�H��H��xH�H!�H��L�IH��@ H)�H!�J�I��H��H��IO��L��P  H��X  L)�H�H��H  H��xH�H�H��H��L�IH�� H)�H�H��H��L�I��H��H��IO��ff.�     H�H��uH�8 tAH��  H���  x1Hc��  ��~H��H��  H�R�H;BƇ�   H�> x� �G�   ��     H��@  H��H��@  H;�H  v��G�   �ff.�     f�f��&   t3H�H���   �xx(tf��H��H��   HE��t��H��   �f��(   t4H�H���   �xx(t9��H��H��   HHE��t��H��   ��@ ��+   u��D  ��+   t���,   t���-   u�� AWAVAUI��ATUSH��H����  f;��   �h  f9GT�^  ��H��L��8  H���  H��f��l   tf��n   �}  H���   HCXH��H�H�VH�6H+PH+0��I��H��P  H��~-H��X  H�L9�~H��H)�I9�~H��H��M��HH�I��f����  H��H����  ���   L��H�����  I�����  tM����   I��M9�MO���  H��   H��H�UH�u H��HC`H+PH+0���  L��A��H��H)�H���   ���  ��  f��  fD��  ���  tfD��  H��[]A\A]A^A_�f.�     ���   t��C�   �fD  ��M����   M��Iֺ    LH���=���M9�ML��1���f�     H���   HGhL���  H���  H�L�L�HH�2H�RI9��}   D)�D)�Mc�Hc�Hc�Hc�I��H��H��H��H��?H��?H�� �  H��: �  H��H��H��Hc�Hc���I���!���f.�     I)׺    M��M��LO���~����o����L)�L)�H����Hc��  H�H��H�L�� �  I��Mc������f�AWHc�A��AVH��I��M��AUA�Չ�H��AT)�E��UH�D1�SH��8�t$H�|$H�D$D�\$Ic�Ic�I�I�H��H��I�I�<I�M�$I��I��I)�M)�L9���   H��H)�L�L$(L)�D�T$$D�D$ H�$�!���H�$L��t$D�D$ D�T$$M��I��H��H��L��L�L$(I��D��E��A��9t$|^H�t$H�H�$I�6I�1H�t$H��L��D  L�H��H�H��H9�t%H�H9�~�L9�|`L�H��H��H�A�H9�u�@ H��H�������H��8[]A\A]A^A_� uH9�u�L9�uB1��t$9t$�f�����f.�     )�H�H�$I��I��?J�� �  H��H�H��]���L��M��I��H��H��H��L��I��H��D��E��A�������AWAVAUATUSH���   L���   ���   L���  Ǆ$�       M�e8�  M���  E��t:E�X�L�R1�I��I��D  M�I��L�M�LI��L�LH��I9�u�1�A9wx��   M���   ��nI�4�I94���   E��H�L$(�   L��$�   D��$�   L��E1�H�T$1�H�|$ L���Pz��D��$�   H�D$E��t^H�$    H�D$    H�t$L���p���H�t$L���c���H�4$L���W�����$�   H���   []A\A]A^A_�fD  �   ��L��L��$�   E1�1�L��   ��y����$�   H�$    H�D$���z����   E1�L��1�L��$�   L���y����$�   H�$���J���I���   L��H��H�,�H���mE����$�   ���!���H)�L��H���@G����$�   ������I�E A�E1�1�L��$�   �   L��I�]@H�D$8�y����$�   H�D$`���K  A�1�L��$�   E1��   L����x����$�   H�D$h���v  A�L��$�   E1�1Ҿ   L���x��H�D$0    H�D$H��$�   ����  L���`H��L����L$0�RH����H9��.  �L$0��f���f�T$X�҉�$�   ��H9��  H+\$8H�H�\$Pf����  E1�1�L��$�   L��   L���x����$�    H�D$@��  E1�1�L��$�   L��   L����w����$�    H�D$8��  H�D$0    ��$�    tEH�D$H�|$H�p��$�   �P�1�H��H��H�H��H�H�LH��H�LH��H9�u�f�|$X ��  ��$�   H�l$L�d$xH�D$X    �C�L��$�   ��$�   H��Ǆ$�       H��H��$�   �C���$�   �C���$�   �C���$�   L����F��L��D����F����f���k  ��%�  A;Gh�E  A�H�|$`H��H����I�OpH�4��R�����@��  L�D$HH�L$h��L��H�T$`����Lt$PI��L��$�   H����  I�U I�E@H�t$PH)�H��$�   I�EHH��H)�H9�vH��H�I�E@�� �Z  ��$�   H�\$0��$�   ��$�   D��$�   L��I���   ��AD�������$�   I���   L��H�D$p��AD�����H����H�|$p H��H��$�   �����  H����  H�����  1Ƀ�$�    H�4$H�|$t(� H�H��H�TH�D H�TH��H9�$�   u�1Ƀ�$�    Mc�t}���sH��;�$�   s_H�$�H�T$pH��H�Hc�I��H��H��?H��: �  H��Hc�HH��$�   Hc�I��H��H��?H��2 �  H��Hc�HP��9�$�   w�H�D$f�8 ��   f�D$P  E1�L��$�   H�\$H�D$PH�SD�BE9�|:H�$Mc�B�< ��  A�T$Hc��H�$H���|� ��  A��A9�}�A��H�\$f�D$P�D$Pf9�L��$�   1�1���$�    �!  H�|$8L�T$L�D$@L�L$ �"H�L�I� H���H��9�$�   ��   H�\E H�TEI� L�I+BI+TB9�$�   w���  9�$�   ��  9�$�   �z  9�$�   u�A���  u�L�H�� H�D$0    H�D$H    H�D$h    H�t$0L���К��H�t$`L���Ú��H�t$hL��趚��H�t$HL��詚��L����B������H�D$0    H�D$H    �Ǆ$�      H�D$0    �H�|$X�tH�t$XH�|$x�[���H�D$X    H�\$xH�t$pH���@���H��$�   H���0���I�EHI�U H��$�   H��H)�H9�vH��H�I�E@H��$�   ��$�   ��$�   H�\$P9�$�   �����L�d$xL��$�   J�4�    1�L�D$8L�L$@H�|$(�eI�H� H��   H��
HGI� H��   H�\$H��
HTGHKI�H�� �  H��H��HI� H��H�� �  H��H��HQH9�u�H�t$@L���C���H�t$8L���6���H�|$0��Z����H���A�? �"���E1�L���A��H�t$hD��A��H��H��H��A�D9�w؅������E1�L���mA��H�t$HD��A��H��H��H��E9'w������I�EHI�U I�m@H��H)�H)�H9�vH�H��I�E@I���   H��$�   L������I�] H�D$0I�E@H�D$PI�EHH��H)�H9�vH�+I�E@E1�1�L��L��$�   �   L����p����$�    H�D$8    H�D$@�����H�D$PE1�1�L��L��$�   �   L��H)�H�D$P�p����$�    H�D$8���������Ǆ$�      L�d$x�w���E1�A�? �����L���B@��H�t$`D��A��H��H��H��E9'w�����H�t$@L��胗��H�t$8L���v���H�D$0    ����H�t$@L���[���1�L���Q���H�D$0    �f���E��E�uE9�|QD��$�   Mc�D��L��E��� L�D$I��D�������D��I��E9���  H�$B�<0 t�A�v��z9�~�D����D��E��Hc�H�T$H��H�H�t H�H+
H�vH+rH��H	������L��H���HL I��HtH��D9���
HL Ht��H��A9�}�����1�Mc�H�|$8L�D$@L�L$ �L�H�I��H��H��A��9�$�   �����H�\$pM��H�4�Hc�H��$�   I��H��H��?H��
 �  Hc�H��I��Hc�H��H��?H�� �  H��Hc�9�$�   w�D9�$�   tqD9�$�   tQD9�$�   t;D9�$�   �f���A���  �X���H�H���L���A���   �x�������A���   u���A���  u�L�I������A���  u���A���  �*���H�I� �����A���  ������I���   H��$�   L������H�D$XH������E��I��D��$�   ��E�rD9�tF�zA9�|L�D$I��D��D������E��~.A�u�A9�%L�D$D��I��D���E���d��������E�������E�������ff.�     @ AWAVA��AUA��ATA��USH��H��  H�GH�/Ǆ$�       H�D$���  9�sf���  D�c(�C u`H�CH�@XH�pH�@H�D$H���   H�4$H�@hH��tXH�xH� H��$�   D�����$�   ����  H�Ĩ  []A\A]A^A_�f�H���   H�$   H�D$   H�@hH��u�H�S8D��H���0����K8�D$3 H�D$����  ���  H�C@    H�CP    H�CH    H�CX    L�S0L�;1�E1�E1�E1�f��$�   L��L�T$(fD��$�   fD��$�   fD��$  �8��1�D��L��M��p  H�D$ L��$�   H��$�   A��  H�SXD��L��L��$  H��$�   �g���H�D$ L�T$(H��L���7�����
  ��$�   ��$�   �{l �C`��$�   ��0  ��$  �Cd��4  u�Cl�ChǄ$�       E���  �s8H�߅�tf�{< ��  荗��D��H���B���H�E  �u
�E���  �   A�   D��H�     H��$�   1�H��$  H��$�   �H�H�CpH�;H��$  Ǆ$�   H��$�   H�CxǄ$�     H��$�   H���   H��$�   H���   H��$�   H��8  H��$�   H��@  H��$�   H��H  H��$   H��P  H��$  H��$�   H��$�   H��$�   H��$�   H��$�   H��$�   �������$�   ����  H��$�   H�CpH��$�   H�CxH��$�   H���   H��$�   H���   H��$�   H��8  H��$�   H��@  H��$   H��H  H��$  H��P  H����  ��uH��$   H+�$  H�� H���Ch��uH��$@  H+�$0  H�� H����4  �C ��   Hc$HcCpHct$H��H��H��?H�� �  H��H�H�CpHc��   H��H��H��?H�� �  H��H�H���   Hc�8  H��H��H��?H�� �  Hc�@  H��H��H�H��8  H��H��?H�� �  Hc�H  H��H��H�H��@  H��H��?H�� �  H��H�H��H  Hc�P  H��H�H�� �  H��H�H��P  Ǆ$�       �    �|$3 tH���   H��$�   H�@hH�xH� �P��$�   �L���L��$P  1��
   Hc�$�   L��H��$�   �H��S8L���3���K8L�{0�D$3H�D$    ���X���H���  H��tgHT$D��H����H  ��$�   ���W���H����X  H�߉�$�   ��P  D��$�   E���-����K8�������f�{< ���������f�H���   H�xh u�Ǆ$�      �����H��$�   L���28��D�苄$�   ����  H�fD;��  �.  A�ո   ;S8�Z  H��  �   M�苰�  H�xH���  H��$  H��$  ����H��  ��$  ��$�   ���  ���  H���  L��L���3����$�   ����   H��  H�KH�C�|$H���  D�L$~L��  H�q@H��   �A)�f���   �AD)�f���   �$H��HA(H��H�H���   H�q H�HQHH���   A��H�HA0H���   1�H���   H��   f��  �H���   H�H��� ����   ��9�w���   H��f���   �x����     ��$�   �D���@ �ۑ��D��蓐���C8H�t$H�ߍH�H���  H�T
D����H  ��$�   ������f�{< �  H����`  ��$�   ���n  H����P  L�cH�Ǆ$      H�spH�{xM�t$bI�T$hL���   M��I��J�4*J�|*H���   H���   J�t*J�|*H��8  H��@  J�t* J�|*(H��P  H��H  J�|*8J�t*0I�T$pB�2 I�T$pB�D2 I�T$pB�D2 I�T$pB�D2 H�;A��H�G  ���  �G���  E1�H�C I�t$hI��A����  M�E@���   H�CI�H�@XH�HH�PH�G  ��q  �G��g  I9�vUHc�Hc�H��LcH��L��M��I��?O�� �  I��Mc�L�P�LcP�L��M��I��?O�� �  I��Mc�L�P�I9�w����  ����  M����  ���
  f���   1�H��L�$�F���L�$��$  L��L��耊����$  ��$�   �������H�|$�`��������tyH��h  �����E��L���   H��h  f�C<H��t'E����  D���D  ����  H�R��H��u�H��L��H�L$�,���H�L$H����  Ǆ$�       H����P  �b���Ic�L��$  E1�1Ҿ   L���eb����$  I��������H�;�s(I�T$`E��H��H�$�	���H�;L�$��$  ���  ��uK�L)K+)H�� H���Kh��uK�T)0K+T) H�� H����4  �����������J�.J�T.��H�CpH�SxJ�D.J�T.H���   H���   �0	  J�D. J�T.(H��8  H��@  J�D.0J�T.8H��H  H��P  M���<�������f�I9������Lc�Lc�H��L�� HcH��H��I��I��I��?J�� �  H���� ��Hc�H�P�HcQ�I��I��I��?J�� �  H���� ��Hc�H�P�I9�w��z���H��H������D  H�pH�@H��u�L��H��H�T$�K���H�T$H������L�zH�D$H���p�@f�t$f�D$~��h  ��$�   �������H��   H��H�D$(��P  H�E  �u
�E��  H�D$E1�1Ҿ   L��$�   L�����   HǄ$      HǄ$       �D$ ��H��f��$  f��$  HǄ$(      ��_����$�    �h  E1�1�L��$�   L��H��$  �   H�D$@��_����$�    I���/  E1�1�L��$�   L��H��$  �   �_����$�    H�D$8��  L��$�   E1�1�L��H��$  �   �]_����$�    I���y  �D$ L�T$@L�\$8f�D$4H�D$L��H���   1��&HcOH��H��0H�J�HcO�H�J�A�fA�CH��H�4 ��M�L�f9D$4Ƌ|$ �    L�T$@f��IǍxf�D$ H�CpH�H�CxH�B�D$ H��A� f�H��H���   H��L�H�0H���   H�p�qA�fA�<SH��H��8  H��H��L�H�8H��@  H�x�AH��H��A�fA�4SH��H��H  H��L�H�2H��P  H�rH��$  D��A�fA�KL��D��$  L��$  L��$(  L��$   L�L$8����L�L$8����$�   �  H�D$1�L�T$@H���   �&�@tH��H��A�4
A�L
�p�HH��0H��f9T$4�H�D$ H��I�H�
H�RH�SxI�TH�KpH�
H�RH���   H���   I�T I�D0H�
H�RH��8  ���  H��@  H�H�@H��H  H��P  ��u"H��$  H��I�D�I+D�H�� H���Ch��u%H��$  H��I�D�I+D�H�� H����4  H��$  L��L�L$ ����H��$   L��HǄ$      ����H��$(  L��HǄ$       �փ��L�L$ L��HǄ$(      L��躃����$�    �<���H�S ����   Hc4$HcCpH��H��H��?H�� �  H��H�H�CpHc��   H��H��H��?H�� �  H��H�H���   Hc�8  H��H��H��?H�� �  HcL$H��H�H��8  Hc�@  H��H��H��?H��8 �  H��H�H��@  Hc�H  H��H��H��?H�� �  H��H�H��H  Hc�P  H��H��H��?H�� �  H��H�H��P  ���}  L�|$H�C0E���   L��E�gPH�D$ �C8�D$4����E���Y  �D$Mk�0H�l$�$A�E�D$xA�F�M��I��I�DM��Hk�0H�D$p�h�ED�D<$9��   E9��  H�u D��H��H��H��H�H�L�8H�XL+:H+ZL��H	��%  Ǆ$�       I��0L9l$p��  I���   I��H  E��4  I��8  I��@  E�^hH�D$HI�D$XH�T$`M��P  �T$xD�T$@B�4(E�T$H�L$P1�I�npI�^xH�|$XL��M���   L�L$hD�\$8D�T$�������$�   ����  I�L$XD�T$L��A��u_H�t$HH�|$XI�npH�T$`L�L$hI�^xI���   H�t$PD�\$8M���   I��8  �t$@I��@  I��H  M��P  E�^hA��4  A�t$�t$A9������I�nD��H��Hu H��$  �uD)�f��$  ��f��� f�t$8��  LcyHcY��7���D��	��z���f�|$8 t	����  I�V ���P���I�FH�pXHcFL��L��H��?M�� �  HcFI��H��Mc�H��H��?H�� �  H��Hc��A�����������I�H���   �xx#uI�� I���H�� H��������@ M������J�D. J�T.(H��8  H��@  J�D.0J�T.8H��H  H��P  ����A�T$`A�D$bL�$I��$�   f���   I��$�   f���   H���   I�T$pH���   H���   I�T$xH���   H��   1�f��  H�PH���q���H�C I�t$hH�;L�$I��A������H�qH��$  D�T$HH�L$@����H�L$@D�T$H�A�N���E1�����H��L��H�L$8H��$  ����H�L$8Ǆ$�       ����J�D. J�T.(H��8  H��@  J�D.0J�T.8H��H  H��P  �����H��$�   �   L��H�L$�7����$�    �e���H�L$L�xH��H������#���H�|$�"���H�Cǀ�   pmoc����Ǆ$�      H�l$����H�D$ H�l$L��I�F0�D$4A�F8H�D$(I��   A�F �Z����A�P����t$94$�C���M�fA�D$f���tA�T$b�TBA;T$�N  Ǆ$�       I�|$I�t$ H�CpH�SxH��H��H�H�TH���   H���   H�DH�TH��8  H��@  H�D H�T(H��H  H��P  H�D0I�D$(H�T8�8 I�D$I�T$(�D I�D$I�T$(�D I�D$I�T$(�D L�c0H��   L���!����$�   ���[����������H�l$�:���H�qH�yH�L$8�4��H�L$8H��H�q H�y(Hc�L���|4��H�L$8H�H��L��H��?M�� �  H��I��H��?Mc�H�� �  H��Hc�������p1�L����U����$�   ���d�������H�D$ H�C0�D$4�C8H�D$(H��   ����fE���4���H��  �'����     AW��E��AVH��I��I��AUATA��US��H��8H�L�N�M9�~H��L��I��L��M��I��I�vI�N�L�<L�,J� L��M��L�$L)�I)�M9�tvM9�tqH�D$    E1�A9�rML��L�T$I��E1�H���D  Hȃ�H�.A9�r&I���H��H�(I9�}�I9�jL���H�.A9�s�H��8[]A\A]A^A_�@ A9�r��H��L�8M9�|"@ IɃ�L�>D9�wƉ�H��L�8M9�}�O�L9�MO�M����f�E��t;�/Mc�D)�H�I��I��I��?J�� �  A�   H��H�H��<���f�     H�t$H�<$L�D$(H�L$ L)�H)�L�L$H�T$����I�~I�vI��L�D$(H�L$ L�L$H�T$�y���@ AWAVAUATUSH��HH�H���   �xx(��   f��   �  ���  �  H��  A�   H��H�D$ H��   H��H�D$(H��(  H��H�D$0��  I��E1�E1҉T$8f�     I��8  I���,AA��@  )ōB�9�F�A9�w0I��0  E��D��F�,t�   f���D�,��   ��9�v�A��A��fE9�  ~IA��  뒀�+   ������,   t	��-   u ��  ���  ��  Ƈ,  f��uH��H[]A\A]A^A_�H��  A�   H�D$ H��   H�D$(H��(  H�D$0�����D  �CA��A��9�vb�   fD  �L$8D9�vdD9�v_D��E��H�|$ �D$L�\$E��D�L$D�T$�t���D�T$D�L$L�\$�D$A��A9�w)I��0  D��D�,
t�A�T$�A�w9�v�E��A��A9�v�A9�t|A�w��9�w3�D$89�v+A9�s&A��D����D�L$H�|$ D�T$�����D�L$D�T$��tX�S�D9�rP�D$89�vHA9�sCD��A��D��D�L$H�|$ ����E��D�L$�T���H�t$(��H�|$ H��H�H+u@ E���.���A9�s@A��L��A�<H��I�H�I��J�|fD  H
H��H9�u�9�r���H��H9�s�E�������Ƈ-  f���$�������f�ATI��USH��H��H�?�GtIH��p  H�T$���   �Ņ���   �����H�;H���   L���F���H��@uH����[]A\�f�1���@ 1�H��������Ņ�u�H�CXA�T$�Hf9AGT$A�<$t��u�H   ���   �Ҿ   �����H���   H����[]A\�D  H�t$H���ێ��H����[��]A\�ff.�      AWAVI��AUATUSH��H�oH�|$�M H�]9�F�t$��t|I��D�f�E1��$fD  �"  K��    H��0I�GM9�tLI��H�sK�D� H��H9�H9CHMCH��H�CH9�~�H�sH)�H��0H)������H��K��I�GM9�u��M H�D$�\$L�`89��  ����)�I��H�I�T�fD  H�     H��H9�u�M��teE1�E�$A��vIM�T$D��A�   1�M�<�I�?I�RI�B I�JH9�~�e H��H�@H�P�H9�HA��A�pA9�u�A��I��D;m r�H��[]A\A]A^A_��    H)�H)�����K�������@ D��H��I�I�H�qA��I��I+rH)�H)������I�T$�HDI�D;m �1����M��t���t������AWAVAUI��ATUSH���   H���   L���  H�t$H���   H�D$Ǆ$�       M����  �D$@ E�'E1�D��A�MH�DH����L$8H�D$ H�[H��H�D$(��H��H�D$��A��H��H��    H�D$0M���}  H�|$ �*  I���  H�|$H��$�   H�p ��,��H����$�   ���  I���  H��H�P H�p蛁��H�T$(H�|$H��H�D$ D�AH�D H�H�AH�QH�E��t,A��H��H��I��N�Df�     H�>H��H�L9�u�H�t$Ht$0H�E��tpA�t$�H�|�H��=H��htdw��  H��zspo��  H��tnlsuH� ��F fD  H��H��0H9�t$H�p H�H��thgwu�H��H� ��F H��0H9�u�H�D$H���$�   H���   []A\A]A^A_�fD  H��$�   H��ravg��@  ��$�   ��t%H��$�   H��2FFCL��A��@  ��$�   ��u�H��$�   H��ravfL��A��@  ��$�   ���y���H���A��H��$�   � �F H��I���Y#����$�   ���J���H�|$H��$�   ��   ��$�   D��$�   ��*��H��I���  ��$�   ���	���B��   D��$�   9��D$@D�"�[���f�     H� �F ����@ H� ��F ����@ H�|$C��H�L$HH��$�   H�t Ht$(Ht$ I���  Ht$0H�|$H�p �A*��H��H�D$P��$�   ���j���H�T$ L� H�L$(I���  D�T$8L�L�
H�xE��H�L$HD�'�G����D�WH�WL�_H�|$I�4;t3�|$8L��    L�؃�H��H��L��    H�0H��L�H9�u���$�   H�D$HD$0I�L�E���  E�D$�K�D�L� L�I��H��0L9�u�H��H�L$XL�D$H���L�D$HH�L$X����$�   �}���H�D$PH�L$XH��$�   D�d$HM��L�pJ�D@"H�\$`I��L��I��@ L�� �F H���8!����$�   ���)���H��$�   H�C H��$�   H��H�SH��$�   H�SH��$�   H�S��$�   �S(H��H�C H�H���BH�C H�H���BH�H�S �PH��@ ��$�   fA�$H�CH9CH;C~H�CH�CI��H��0M9��:���D�d$HH�L$XH�\$`H�|$E1�1Ҿ   M���  L��$�   �`G��I�F(��$�   ���=���f��$�    �.  1�9D$8�  I��p  L��$�   �   L��L�t$8L��H��$�   ��(  ����  L��H��$�   �   L����(  ��tpA�   H�L$8H��$�   �   L����(  ��tK��$�   H�|$PH��HGH�WD�p�@   H� E��tA�L$�H�t�H�JH��H��0H�H�H9�u�I���   M���  �RAVML��H�L$8L�u8H��A��@  ��$�   �������H������H��$�   H��H�D$8�K����$�   �T$@��������   H���Y���T$@��$�   f��������������H��$�   �0   L���w&����$�    I�G`�h����   H�������$�   ���L���I�W`H��$�   H��H�T$@���H�T$@��$�    f�����H��$�   H�������$�    f�D$@�����H������I�O`�t$@L��Ht$8H�D$HH�Q�p�����$�   �������M�W`E1�1Ҿ   L��$�   L��A�
L�T$8��D��L�T$8��$�    I�B(�����H�t$HH��������$�   ���j���I�G`H���0��Hc������$�   ���F���I�O`H�\$8�L�q(H��H��L�H�D$@�OH������H��I��?��H��fA�F�2��A�vfA�F
��;s�"  ����Hk�HC;0�  I��L9t$@w�H�\$8�  f�I���  �x0 �f  H�|$PH�@(H�H��H�ǀ|$@L�l$`I��H�H�\$xE1�H���D�d$HH�D�H�D$XH��    H�D$hA�D$�I��H��   H�D$p�    H�t$XH�������$�   ���l���H���T��H����A�F�E��M�.H�D$p�T$HI�\ ��tH��I�����I�E�L9�u�|$@ udA�F��  H�D$`I�L��A���t$HI��H���  �I���H��Ld$h�|����$�   D9��S���D�d$HL�l$`H�\$x�����    H�������A�F�H��H�L$H����H�L$H����$�   ���������H���Q��L��I���&���L��H�������$�   ���\���f��$�    H�D$PH�@H��I���  H�@(H���W���� ���fD  A�   �S���H��$�   H�D$8����Ǆ$�      H�\$8H�������$�    �����I�G`�H�P(H��H��H�2L���6o��H��t� f�BH��H9�w�A���     �d����AWAVI��AUATI��U��S��H��   H���   L���  Ƈ�   �D$H    H�D$M���Z  M�}A�79�Fޅ�tJI�H   H=   ��  I�F�S�H���#�     H�8H��H��   H��   ��  H9�u�A��$�   uI���    ��  I�} �D$ �(  I�}H���S  ���e  I�H9�e  D�S�L�G�   I��� L�HI��M�<�L99��  L�ȉ�L��L9�u��D$    E1�M�D$A��  ��  A��A��D��L�M�E(I��9���  D�F�A�   A)�N��   E1�f.�     N�< N9<EE�I��M9�u�E����  H�9 ��  �BH��H���@ H��H�x� ��  ��9�r�A�u ��L��H���pu��@����  �|$ M�uI�MtA�] I��$�  ��9F(H�D$���$  �u�1���H��H��I��H�PH9�u��9�v&����)�I��H�I�T� H�     H��H9�u�H�D$L�h8M���>  ���N  �]��l$ M��L��H��H��L�fD  E�A��vLM�WH�} �   E1�I�RI�B M�JH9�~#��   �     I��H�@H�P�H9���   �΍ND9�u�I��H��I9�u�H�D$�l$ H�@H�H1��>�2  �q)�Hc�Hc�H��H��H��?H��2 �  H��Hc�H�I��H��H��09�vzI��H�yH��y���+q�fD  �   H�Ĉ   []A\A]A^A_ÐA��I��M�I�BI�1I+2H)�H)�����I�WJ*H�E �>���H�D$H�@H�H���G��� I��$�  AƄ$�  H��t<�D$����   ��u*H�|$�e��I��$�   L��IǄ$�      �ڭ���D$HI��$�  H�|$��d���D$HIǄ$�      �,����    I�<�������    9���  �F�A�   )�L�T�H��D  H�8 EE�H��I9�u�����f��D$   �1��� 1������D$H�������M��$�  ����A�   �D$   �Z���D  I��$�   L��舥���D$H�)���H�|$��L�L$HE1�1Ҿ   �<��I�E�D$H���Q���A�7�D$����H�|$��L�L$HE1�1Ҿ   �l<��H��I�E�D$H������A�7�D$   �g���I��$�   H�L$P�ravgH�x8H�D$H��H�|$L��A��$@  �D$L�������H�|$����H�|$H�T$X���F H�D$ �����D$L�������H�|$X   �   �����I�M�T$`f;�w����L$bH�|$PH��H��H��H��H9��W����L$rD�D$p��f��H�H���H��I��H9��-���A�uhH�t$xA�H1�I���   H�|$L�L$LE�ExE1�H�t$(�   �:;��I���   �D$L�������H�t$(H�L$ A�ExH�HL$PH�t$(�pH�L$0�D$r��   H�|$H�������D$L�������1҉l$<�݉����A;]x�   H�|$�,��I���   HD$(��H��H;D$0vЉ��D$L   �l$<�R E�������AƄ$�  ������1���1������H��1�1������H��1�1�A�   �D$   �������l$<H�|$�	���D$L�������A�Eh��un�D$H    A�7����H�|$H�����D$L�������1҉l$<�݉��	��A;]xw�H�|$�	��I���   ��H�%�� HD$(H��H;D$0v������L$`H�|$E1�1�L�L$L�   ���9��I�Ep�D$L���A���H�|$H�t$ Ht$h����D$L���!����t$`A�uhH�|$H��M���D$L�������1�L�t$M��A�܉l$ ��A;mhs@1�f�|$` t.H�|$�����T$`H����H���͍<I�Mp��H��9�w҃�� H�|$D��l$ M��L�t$�O���D$L�D$H���|���A�7������    AWI��AVAUI��ATUS��H��L���  L���   �D$    M����  I�nI�F�M 9�F�H����  ����  D�C�1�1�M�H�@ H��I�4�H94�t	H�4п   H�rL9�u�J�ȉ�I�UA����  ���   ��H��HUH�R�N��9�v5�Q�)�L��   1�f.�     I�4H94t	H�4�   H��I9�u�I�~ t	@���]  L�L$E1�1Ҿ   L���7��I�ǋD$��uNI���  �0 ��   I�VL���������u 1�L��L�������D$��uI�EH�̀����HD�I�EL��L���^���D$H��[]A\A]A^A_�fD  K�@H��HU9��H���D�A�E��A)�N�D�D  H�rH90tH�0�   H��H��0L9�u�����D  L���h���I���  �;���@ 1�������D$��uAM���  �"���D  1�L�L$E1��   L���6���T$I�F��u�M ����D  E1�����1�1��4������������ff.�     f�AV�   AUATU��SH��H��H���  H����   �K9�ro��t~L�j��L���   H��H��I�UL�t�H��p  H�T$A�v��   ��u3H�s0L���]��H�D$I�H��A�u H�C0������t*����    D�H��[]A\A]A^�fD  1�1�H��������S��H�c���H	�H�kH��[]A\A]A^Ð1��i�����u�H���  �/���f�     AUI��ATI��US��H��H���  H����   H�} ��   9] ��FM A���   t`��t H�}�q�1���H��H��I��H�PH9�u�9�v(����)�I��H�I�T�D  H�     H��H9�u�1�H��[]A\A]� ��t��Q�L��I�T��H�     H��H9�u��fD  1�������u�I���  H�} �H��� 1�1��   L���������,����ff.�     f�AUI��ATI��US��H��H���  H����   H�} ��   9] ��FM A���   t`��t H�}�q�1���H��H��I��H�PH9�u�9�v(����)�I��H�I�T�D  H�     H��H9�u�1�H��[]A\A]� ��t��Q�L��I�T��H�     H��H9�u��fD  1��q�����u�I���  H�} �H��� 1�1��   L���������,����ff.�     f�AW��AVH�@AUATUSH��8H�FH��H�XH�D$�@H�\$ ����H�\$(���l  H�D$    E1�I��I���    H�D$D��fA� H�t$H�@��I�GH���$  1�   E1��2@ H��H)�H��H)��_����    A�WA��H��H��A9�szH�H�SH9��H�sH9��H��H��A��H��?A��tH��u�H��t�I�} H�H�</H9�t�H9���   H9���   H9��t���H��H)�H��H)�H���а���s��� H�H�L$ H�l$A��Hl$(H�iH��H��H�H�� �  H��H�HD$H�D$D;`�����H�D$H��8[] �  A\A]��A^A_�fD  1�떸   �H��81�[]A\A]A^A_�@ ���  ��  AWAVAUATI��USH��H���  L�M`A�M�q(H��L�I9��g  1�1�L���  1�f�D$
f�T$f�L$�-�H��csdh�#  H��pglhfED$
f�D$
I��L9�vSL�M`I�6L���)^��A�N
A�VL��I��I�q����M��t�A�V�fA�U I�H��csahu�I��f�D$L9�w�D�t$D�|$D�l$
A��$�   ��A A��$�   I��$�   A��$�   A��$   A��A��$  fE��$�   )�A�fA��$�   Aŉ�fE��$�   f��E��E)�1�fE��$�   f��)�fA��$�   H��[]A\A]A^A_�WZ���    f�D$�����fD  ��    E1�E1�E1��7���f.�     AWAVI��AUM��ATA��USH��H���   H���   ���F �T$H�x����H���  1�L��I���d����Ņ���   M��D��T$H��L��A�W�Ņ�urH��  �dbk�H9���H=eurt��!ʹtsl�H9�����tH-   H�������  H���   �t$H�K   H�D$ ��x��M��D��H��H��A�W�Ņ�tH���   ��[]A\A]A^A_�f.�     L�c(M��tWA��F A��F �f�     I��M9�t7L��L���d��H��t�H�D$HL��@  H�D$(�  ��   �f�     H�|$H1��   f��    H��H�|$(L��@  �H��    ��  1�H�Ft�D$: �D$; �D$9 f�|$H�D$�l$<D�d$H��(  I��J� H��mgpf�Y  H��perp��   H�� tvc�'  f�D$�D$f;�   r��l$<�T$HH�L$(�h�F �ذF �|$9D�D$;D�L$:��H��0H��H9���   �@��uH�8 u���E��uH�x u���E��uH�x  u�����u��|@ �D$:��  A�   I��L�|$(1�L�d$M���$ I��I��0L9|$�6���H��(  I��h�F HD$H9Pu�H���c  A�I9�`�F u��A���u��l$<H�K    L�|$ H�L$(�xmdhH��M�g8L��A�҉D$D��uH�t$HH���  H�C���   H���   H�xh �_  H�t$ H��肜���Ņ�t<��v���H�L$(H�T$ �mgpfH����@  ���:  Hǃ`      HǃX      H�L$(H�T$ �perpH����@  ���k  Hǃp      1�Hǃh      H���   H�xh ��  H�C�t$����t����  HǃH  �/A HǃX  0 A Hǃ`  �4A Hǃh  �JA HǃP   0A ����M�������1�H���   H�0H��A�҅���   H��(  H�L$L���   L�dL��L��L�d$0������uyI���  1�D  L��I���d����I��w�H�d$0H�D$0H��t<A�   �   H�\$0��A)ĉ�L���}�����    �������D9�u��H�\$0L������L��@  �����@ ��  E1��D$9�f���fD  �ć  A�   �D$;�K��� L��   L��L�������D$D���  L��   A�GE�w��AΉ�A�G	�A��A������DG�f=� ��   D��E��f���L  I�V�H����  ��   H�L$H1�E1�L�L$D�   L��D�T$H�L$���)���T$DD�T$H��   ����   H�|$O�D7L�L9��  E�J�1�1��L�H��I�H9�rH��   A�t@�4�rI9�u�H�D$H��  L��  H��  �D$D����������m��� �   �`���fD  �D$D   H�|$ L�������Hǃ      �fD  H���  H�T$ �fylgH����@  ��<���  ������H���   H�xh ��  Hǃ�      H�L$(H�T$ �acolH����@  ��   �������f���   H�D$H�a  H=�� �  H��H���  �   H�S H�rH9�t	H9��  H�t$HH�|$ H���  �g���H���   ��t<��U�����������H���fD  1�����H�������Ņ��)���H�������>���H�t$HH�|$ H��`  H��X  ������Ņ������<����������L�L$DE1�1�1Ҿ   L���'��H��   �D$D���j���1�����H�t$HH�|$ H��p  H��h  �����Ņ������<�������y���Hǃ�      Hǃ�      �}���1��D$: �D$; �D$9 �{���H=�� ��   H��H���  �   �����s8���/���H���   �!���H���   ����E1�E1�E1�fD  H�T$DD��H���xc���L$D��tA�������M��A�   I��L;��  r�A�������M����   H�CH���H�C����H�D$H�� ���  �����H�D$H�� ���  �7���D��   H��(  H��H�|$ I��I��I������L9�sk1������   �    H�UH)�H��~
H9�HL�L�H�� I9�w�@��t4I9�wEH�C L�l$HH��H���  �y���H�|$ �l���H���  �����H�t$ H�vH��H�t$H)��H���  1�H��tH�B�H�C �2���H�T$(�   D��H��������������|$H.�����H�|$(���F �(\����������w���ff.�     U�   ��SH��H���[�����uH�SH�р΀����HD�H�SH��[]�f�     AWAVI��AUATA��USH��8H���   H���  H��@  L�k8@��t6�EPH�L$(H�ھRAVV��A�D$ E��t6H��8D��[]A\A]A^A_�D  �E@H�L$(H�ھRAVH��A�D$ E��u�H������H�t$ H��H�$�p���D�T$ A��E��u��   H������A�D$ ��u�A�   fA���{���H�t$ H������D�T$ I��E���]���H��H�t$ �����D�T$ H��E���?���H�T$ �8   L��E��tw�g��D�T$ I��H�EXE������H�$L��L��J�48�ߔ��A�D$ �������H��uQA���  E��t���EQA���  �����@ ���EAA���  ��������D�T$ I��H�EHE��t�����M���   H�4$�D$I�G8H�L��H�D$�����ƉD$$��tA���f���H�t$$L�������t$$�؅�u�H�t$$L��� ����t$$��A�U ��u�f����D�T$t�   �H�|$�   ��E1�L�L$$1�D�T$�"���t$$I�E0��u�A�M H�|$�   1�L�L$$E1��d"���t$$I�E(���W����ٸ   ��D�T$����E1��������$E;E ��   E1�1�H�t$$L��D�T$D�D$D�L$�T$�L$�����t$$��������T$D�L$���L$D�D$��A��D�T$	�A9�r�����A;E ����I�}(D��#$��Hk�IE;�����I�E0A�����^����    �D$$������A�������@ 1����   ��   AUATUSH��H��L���  M����   ��I�Մ�t;A�|$P ��   A�|$Q ��   I�t$XH�F0H��uFH�V�   9*vc1��K@ A�|$@ u1�����A�D$DL���  A�|$A tUI�t$HH�F0H��t��V �J�9�H�V(HF���,�H���  ������AE 1�H��[]A\A]�f.�     ��    A�D$D�ܐA�D$T��f�     �   ����A�D$TL���  �&���D  �   �����fD  1������f�     ATI��� �F UH��S�L���H��H��tH��[]A\�@ M��t�I�|$H��t徝�F �����H��t�H� H�@(H��t�[H��L��]H�@ A\��ff.�      U��H���   S�p�F H����À� �ۅ�t�   H����[]�fD  H�ׄ�u1���#t��(t�   H����[]��    �ExH����[]�@ �
   1��U����f�UH��SH��H��H�<$H��H�t$蓧��H�4$H�T$H��H�FHI�H��H��f�E H�BHI�H��f�H��[]�ff.�      f9��   v_f9��   vVD����I��L��   H��H��   M�M�@L+H�@L��L��H)�H	�t5���  tIL)�H��L��H	�uC1�� ���   �   t&�G�   �f�� @  H��H��H�I����1�H����H��L����L����fD  AW1�I��AVAUATUSH���   L�I���   �zx(�  M���  1�A��  A��+  fA��,  �   A��T  H��L�H�H��HC�H9�vH��   ���  HC�fA��T  IǇ0      IǇ@      f���  ���2   �2   Ƀ�2L�Hc�I���  �  H�I��8  I�P H��H��H��H9�s
I��8  H��I��H  A���  IǇ�      fA9��  ��  IǇ  �4A IǇ  �4A IǇ  P4A IǇ    4A L���aR��A��@  <w���$��F @ IǇ�  `QA D  I���  I���  E1�A�   I���  �Lc���A���  A�� �F A���  ���  H�H�H9��T  A�� �F I� ����H)�I�8�~  I�(����)  Hc�I�W8�� �F ��H�I�G@H9��.  M�G0AƇ�  A�G    I�,Ѐ���(%  D��B�$� �F H�E H9�|	H���R*  A���   ��%  H�E      I�G@A���  I�G ���|   I��I��@B �X%  I���  I���  H9��^  A��`   �����1��    L�JI9��J  D�LD�ȸ   D)�A���  �����H�U I��H  f�I�G Ic��  I��  �q���f�     I�H���  H���5  �IG8I�G@H9��   A�G�   ��   H���   []A\A]A^A_� A���   ��%  ��t1I�01�H��    A���  H��Hc����� �F ����f9�w�I�G8    �2����     J��,  I��8  � ���@ H���������L��H��H��������    IǇ  �A IǇ  �A IǇ  �A IǇ   �A �����    ��)  �������1�A�@ �������d  ������������    I�G@������    IǇ�  �RA ������     IǇ�  �QA �����IǇ�  `RA �����IǇ�  �QA ����IǇ�   RA ����IǇ�  �A ����IǇ�  �RA ����L���x���A�G@ ���h���=�   �@���A���  I���  H��H��H9�r� ���D  H��(H9������z t��rA8��  u�Ic��  A;��  ��   A��x  I���  H��I��  �H�N�2H�HH�@   H�P�F�����   H�RL���[���<�����A�G����f.�     H��L���S��A�G�����} �z#  A���   �t���A�G�   ��   �E���A���  1����4���A�G�   ��   �"����    A�G�   ��   �	���H�} �����H��L���Ж��A�G����L��A��  H�E A�G����H�U A�OTL�Ef9��   fD9��   H�}A���   H�uf9���  f9���  H�M fA9��   ��  I�G`��E��H�L$hI��H������H�T$ H��H�L�H�L�JH��H�|$XL�`L�D$`H��H�\$(H�I���   L�L$HH)�H�:H�H�\$H��H�8H�rH�@L��@   H�t$0H)�L��L)�L�T$PL)�H�|$H�t$8H�D$萕��H�t$H�|$�@   H���y���H�t$H�|$�@   H��b���L�L$HH�|$�@   H�D$@L��L)��C���H��H�L$hL�T$PH��?H��L�\$XL�D$`H����H1�I��H)�I��H��H�4PH�D$@H�H�H1�H)�H9���(  I���   I�W`M��   H�I�J�4HT$ I�HHHH�xHH�H��I�I�CHCHFHBH�PHH�H��I�AI��   �	A�G�r���f�A��"  A��&  L���
K��A�G�Q���I��(  I��&  H�EH�U I�G@A���  ����I��$  I��"  H�EH�U I�G@A���  �{���HcU Ic��  H��H��H��?H��
 �  H��Hc�I��X  �����H�U I��P  ����I�G H�E I�G@A���  �!���H�E H�UH�EH�U I�G@A���  � ���I�G@    1��u���H�E H�EI�G@A���  �����������f% @f�� @��w fA��"  fA��$  fA��  fA��   �������fA��&  fA��(  ����H�E H�u��f	������I��(  I��&  H��H��������t���H�E H�u��f	�tI��$  I��"  H��H������A��"  A��  �7����U �uI��&  L���������� ��������U �uI��"  L�������������A��"  L��A��  ��H��A�G�7���H�E A��8  H9���  I��@  H��H�E I�G@A���  �~���H�U A��8  H9���  H�MI��@  H��I�G@A���  �I���L���%���A�G����H�m fA;oT�]  1ɀ�.t9��L��H��IG`H�PH�0A���  I���  L��H��H��A���  H)�H����I�wHL��A���  fA��  A�GfA��  �C���A���  ���c!  �Q�A���  Hc�H��I��  H�rH��H�rAƇ�   H����   H�RA���  H�RI���  I�G �h����A�H�I����  H�E H����  Hк    HH�f.�     H�E I�G@A���  �����A�H�u L��H�I����  A���  H�E A�G�s���H�e �I�G@A���  �����H�UH�M H�EH�MH�U�H�E H��?H���H�E I�G@A���  ����AǇ@     IǇ�  �QA ����AǇ@     IǇ�   RA �����H�uH�V�H����  H�} �N��   ��H��tHc�H9��o  ��A"�d  	�A��d  H�������I�H���   �zx(�����H��A��+  �~���fD  AǇ@     IǇ�  �A �]���H�} �R�������H�U �A-  L����C��A�GAǇ@     IǇ�  �RA ����H�U H���H���H����  ���  HO�I��0  �����AǇ@     IǇ�  `RA �����I��0  I9G ��  A�wTfA9�  ��  I���   H��6�>  @ A���   �����I��0  H��I��0  H����  M�G0H��I�W8I�,�fA;��   s�A��  ��L��H��I��   H��IG`H�QH�1H+PH+0A���  ��H��L��H��H��A���  I�W8�v���H�] fA;��   ��  A��  fA;WT��  ��D��I���   D��H��I��H�t$fA��n   �  I���   L�IG`H�QL��H�1H+PH+0A���  H�UL��I���   H��D��H)�A���  A��  fA��  fA��  A���  �����fA��  A�G�:���L���S��A�G�)���fA��l   A�   tfA��n   tE1�fA��p   A��I��0  I;O ��  L�M A��&  D���8@��A��(  D��Lc��%@��Lc�H��:�R  �     A���   �����I��0  H��I��0  H����  M�G0H��I�W8I��fA;��   s�I�H���   �yx(�!  A��+   �  E��u=A��,   t
A��-   u�A���   tfA��(   uI���   ����g���1���A�   L��L��賌��I�W8�H���fA��p   H�] �   tA���   f9������L�D$~H��$�   L��H��$�   H��$�   �@P�����>���1�f��tI���   H�Ӹ   fA+�   fDQ�fA��p   �  E���   D��fA9�w:�����fD  H��$�   A�   D��L��H��$�   ����A��fE9������I���   H9�$�   u�fD9L$~u���I��0  I9G �   L�D$~H��$�   L��H��$�   H��$�   �hO�����f���I��0   I�W83��  D  A���   �����I��0  H��I��0  H����  I�G0H��I�W8H��fA;��   s�H��$�   ��A�   L��H��$�   ����I�W8�I���  ��A+ D�DL��A9��d���A��f����  �   �f.�     I���  H��LH�L��H��f9�s���IG@A���  I�G@�G���H�] ��fA;_T��  H�uI;��  ��  I��H  L��H�D$A��  ��H��I��fA��l   �I  IO`H�QH�1L��A���  L��H��H)�A���  t-L)�H��I���  L��HH�H9L$LL�L��A���  H)�H����I�wHL��A���  A�GfA��  fA��  �����I���  ��A+ D�DL��A9��!���H��A��I���  f��tL�G���H�|� �f.�     I���  H��H�BI���  ��T���H��H�E H9�u�I�G@H�AƇ�   I�G@�~���H�U � @  L���=��A�GAǇ@     IǇ�  �RA �7���L���   A��  H�m I�W8I��H��u&�>   A���   �����H��H��H9��  H���2  I�G0H�J�I�O8H�t��I;��  s�H�<�A���  H��H������t��  L�@ ��uID�A��`  H�H��I9�u���D��H�G�H��H��L��HI�A*�b  H��A��   I�W8�`���H�U ���  ����  I��  I�OHI��  I�OPI��  I�OXI��   I�O`I��(  I�OhI��0  I�OpI��8  I�OxI��@  I���   I�_HM�_PfA��l  M�WXM�O`fA��n  M�GhI�pI���   I�wxI���   M���   M���   M���   M���   I���   I���   I���   I���   M���   M���   M���   M���   I���   I���   I��   fA��p  �?���H�uH�} �@   �=���H�E A�G� ���A���  H�u�SH��H9�����A���  I���  9��  ��H��H�<�H9�r�T  @ H��(H9��C  �JH9�u�z �����A���  A;��  �����H�}  �����A��x  Hc���H��I��  �0I���  H��H�pHcu H�PH�p�2A���  �F�����  H�RL���T���AƇ�   H�E I�0  I��0  I;�8  �����A�G�   ��   �^��� H�U fA9WT��  fA��&  Ƀ��fA��(   t�����IGp A�G�����H�] fA;��   �i  I���   D��L��I��L�H�PH�0A���  H�M��L��I���   H)�A���  fA��p   ����I���   I���   J�T J� J�T!J�!A�G�C���H�E A���   H9������H����F�
  I��   L��H�PH�0A���  H��A�GH�U �����H�u I;��  ��  L��A��  H�E A�G�����H�u I;��  �p  H�UL��A��  A�G����A��x  ����  A���  M���  H��H��I��I9�s%H�U A�AH9�u�6@ A�AH9�t)I��(L9�w�L9�uA;��  �	  ��A���  H�U H���   ��  I���  A�QA�AA���  H��A�9I�AH�E H9�v
��A���  L���l;���������A���  <-�  <�t<,u�A�G�   ��   ����I�O8I�G0AƇ�  A�G    H��H���j  D��GA+G A9������H�rH����  E�������A�x�1��H��H��H��H��H�PH9�u�����I�7H�U H���   ���Hx�    HE���tA��   t����tA��   t����tH���   t���� tA��(   t����(�)���A��)   ����H���� ��@HE���tA��*   t�̀H��H��   ��HE�H��H��   ��HE��������A��.   �����H   �����     H�U fA9��   ��
  H�MfA9��   ��
  ��I���   ��H��H��H�I��I���   H��H�H�H�NH�zH+H��H��H)�H	��z  �����  H)�H��H	���  M��   I��   I�L$H�}I�$H+E H��H��H)�H	��  ����  H)�H��H	��v  L���;7��A�G����H�U I��8  �r���AǇ@      IǇ�  �QA �W���I�H���   �xx#�����I���  H�E I�G@A���  ����H�E fA9GT�o���H�UfA9��   �]�������H��H����I��  I���   IG`L��H�0H�H�PH+1H+QA���  H��A�G����A��x  ����  A���  M���  H�U H��H��I��I9�sA�AH9�u�.A�AH9�t%I��(L9�w�L9�uA;��  �3  ��A���  H����  �  I���  �   A�9fA�IH��A�QI�AA���  I�A     H9�vA���  L���7���������A���  <-�  <�����<,u�����A���  H�M ��H��H9������A���  I���  9���  ��H��H�4�H9�s�PH9�u
��PH9�tH��(H9�w�H9��r����x �h���A���  A;��  �����A��x  Hcу�H��I��  �2I���  H�B   H��H�BH�r�0A���  �V�����  H�PL���{��A�GAƇ�   �����H�}  �   �1���H�} �����!���I�H���   ��	  H�E    I�G@A���  �#���H�}  �����A�   fD  L���6��<�&���A���  <X�z  <Y�c  <u�A��u������H�EH9E ����H�E I�G@A���  ����H�EH9E ����H�E I�G@A���  ����H�EH9E ����H�E I�G@A���  �l���H�EH9E ����H�E I�G@A���  �I���A�G�   ��   ����AƇD   ����H�] I�G@A���  ����H�U H�������H��H�U I�G@A���  �����H�EH9E ����H�EH9E ����H�E I�G@A���  �����H�U fA��  �3���H�U fA��  �"���H�U fA��  ����A�   �f�     <Y����A)������L���g4��<�����A���  <Xu�A����H�U ����
  ���h  I��  I���   I��  I���   I��  I���   I��   I���   I��(  I���   I��0  I���   I��8  I���   I��@  I���   fA��n  �;���H�U ���J  ����  I��  I�OHI��  I�OPI��  I�OXI��   I�O`I��(  I�OhI��0  I�OpI��8  I�OxI��@  I���   fA��l  ����H�U ����  ���Y  I��  I���   I��  I���   I��  I���   I��   I���   I��(  I���   I��0  I���   I��8  I���   I��@  I��   �����AǇ@     IǇ�  `QA ����AƇD  ����I�H���   �xx(�h  I��0  I9G ��  H��7�w  D  A���   �����I��0  H��I��0  H����  M�G0H��I�W8I��fA9�  v���I�0  �0I�W8�H�UH;U �t���H�U I�G@A���  �����L�e fE;��   ��  H�mfA;oT��  ��A��L��H��H��IO`I��   H�QH�1H+PH+0A���  I���   L��H��H��?H�H��A��H��H��H��A���  H����L��I�wHA���  A�G�����H�U I;��  �c  Ic��  HcEH��I���  H��H��?H��0 �  H��H�H��I�G@A���  �����H�U �ʁ��   �`
  ����   ��tA���  9�|AƇe  H�U ��tA��   tAƇe  H�U ��tA��   tAƇe  H�U ��tA���  9�}AƇe   H�U ��tA��   tAƇe   H�U �� �����A��   �����AƇe   ����H�U H�����������  A��h  ����I�H���   �zx(��  H�uH�} E��  ���fA9��  fA9���   f9��E�����I�0  � �f9�s������I�H���   �zx(��  H�}H�u E��  ����fA9���   fA9���   f9��������I�0  �f9�s��r���H�U H�������fA��b  ����1�H�u L��A���  �����H�E �6���1�H�u L��A���  ��H��@����H�E A�G�f���H�M H��~H9���  @ A���   �B���A�G�   ��   ����H�E H���s����=���H�EH)E I�G@A���  ����H�EHE I�G@A���  �h���H�UH����  A�G�   ��   � ���H�UH;U ������F���H�U fA��`  ����H�}  �@��������  �����  �����  ����P  �ˍGA+G f�� ��9�������   H�I��  �H�T��H��f9�s����� L����A�   L��L����u��I�W8�v���H���k�����   �X���A���k�������A���]���A���   t}A�G�   ��   IǇ0     I�W@����A�GI�W@IǇ0     ����A�G�   ��   H�E     �����A��+   �����A��,   �|���A��-   �n���IǇ0     I�W@�����A���   �@���H�E     I�G@A���  ����L���q�������A���   �  fA��  fA��  �k���A�G�   ��   �<���H)к    H��HO��%���A�GI�W@�����A�G�   ��   �	���A���   ��  A�GI�G8    1���L�D$~H��$�   L��H��$�   H��$�   �8��������A��p  f����  E���   fE�������E1��/ H��$�   E1�D��L��H��$�   ��s��A��fE9������I���   H9�$�   u�fD9L$~u���H��L����+��A�G�����I��H  I�OHI��P  I�OPI��X  I�OXI��`  I�O`I��h  I�OhI��p  I�OpI��x  I�OxI���  I���   ����A��+   �`���A��,   �R���A��-   �D����V���fD  H�} �@   �r��H�E A�G�5���I��H  I�OHI��P  I�OPI��X  I�OXI��`  I�O`I��h  I�OhI��p  I�OpI��x  I�OxI���  I���   �����I��H  I���   I��P  I���   I��X  I���   I��`  I���   I��h  I���   I��p  I���   I��x  I���   I���  I��   ����A���   �����A�G�   ��   IǇ0     I�W@����I��H  I���   I��P  I���   I��X  I���   I��`  I���   I��h  I���   I��p  I���   I��x  I���   I���  I���   �t���A��+   �8���A��,   �*���A��-   ��������D  H9�������v����2�F��������H�RL���pm��A�G�W���H)�I��H�E I�G@A���  ����A�G�   ��   �|���A�G�   ��   �j���I��   L��H�PH�0A���  H��A�G�����fA��  fA��  ��   A�G�   �$���A�G�   ��   ����H��H�ЋzH9�����H���-���I�WXL�L$L��I���   I���   H�H�H�RJ�	J�T	D��H�MA��   I���   L�L$I���   J�TJ�L�H�A��  H�QH������A��&  ���"��I�WXA��(  D��H�H�H��f"��IO`H�H�BH�H�RH�H�Q�s���H��H��D�AL9������H���	���I���  I�AA�G����I���  I�A�N���H�u L���p���=���� @  I��$  I��"  �o��������1ۿ @  I��   I��  �P�������H��H������H)�H��I�< I�t H���$��I�G0I�W8H�\��A�G�"���A�G�   ��   I�G8    I�G@    �S���AƇe  �������I����GA+G ��9��!���I���  f�� H�P��H�L� �I���  H��H�BI���  ��T���H��H�E H9�u�AƇ�   I�G@����E�������A�P�H��H�T�H�     H��H9�u������I���   H��A�   fE+�   fDZ�����fA��l   M���  ��   fA��n   ��   M���  I���  IGhI��   L�H�0H�HH�RI9���  ����Mc�Hc�D)�)�H�Hc�I��H��L��H��H��H��?H��?H��0 �  H��
 �  H��H��Hc�Hc�A��H��A�G����f������I���   f������I���   D�TB�A��� ���L�I�G@I�G �F���A�G�   ��   AƇ�   �{���I���   IGXL��H�0H�H�PH+1H+QA��H��A�G�����H�|$(H�t$8�@   L�L$HH�L$@L)���k��H�t$L��@   H+|$0H�D$ ��k��L�d$ H�t$H��I�L���k��H�t$H��L��H�D$�k��L�L$HL�D$I��   M��   LHCM�H�L$@I�A�����A�G�   ����H)�L)�L��H��A��Ic��  H�H��H�H�� �  A�GH��Hc�����H������H��H���x���H������H��H�������    USH��H����   H�oH�T$�P  H�������L$H�Å���   H�h1�L�L$E1��    �    H��ǀ�      ������T$H���  ��uKǃ       H��H�C(    ǃ�      H�C0    Hǃ�      H�    H�C    H��[]� H���4���D$��t
�     1�H��H��[]�@ AWLcٹ/   AVI��AUE��ATUH��SH��H��HL�bI��$�   M��$�   H�$1��H�A��uCE��tfL�[ 1�L�#H�kL�sL�{0Hǃh      Hǃp      H��H[]A\A]A^A_�@ E��u�I��(  D�$L�(L���w��L�kLc$� D��E�����D$.��  ����  ��  ����  ��u��Ѕ�u�H��  H����	  D��H�4$�����~x(�F	  Ɓ*   ��D�l$ �D$H��L��H��D�T$,D�\$H�L$��8�����2���H�4$H�L$D�\$D�T$,�~x(��(  � 	  8D$t2�D$��(  �t$.H��D�\$H�$��=��H�$D�\$���������d  D�ڃ��DEڨ��   1Ҿ   H�       @Hǁ0     H��  H   @H��   1�f��(  H�      Hǁ8  @   ǁ@     ƁD  HǁH  D   HǁP      HǁX      ǁ`  	  f��d  H��h  f��p  �D$.���  H���  H��  H��  �������������3   H�H��   D�\$D�D$,H�D$H���   H��H�D$����H��  H�|$Hǅ       ���H���  H�|$Hǅ      ���H�|$Hǅ�      H���  ���D�\$H��  Hǅ�      D�T$,H��tD�T$,D�\$�N1��D�T$,D�\$H���  D�T$,H��D�\$H�D$ ��1��H�t$Hǅ  ����H���   ����H�t$1�E1�H��  H�|$L�L$8���  H�����   ���  ǅ�       ��  H��x  ǅ      H���  ���  �(   f���   1�Hǅ      f���  Hǅ�       Hǅ�       Hǅ�       Hǅ�       �����L$8D�\$H��   D�T$,����  ��  H�|$E1�1�L�L$8�(   �����D�\$D�T$,H��  �D$8����  H�|$E1�1�L�L$8H���  �   ����D�\$D�T$,H���  �D$8���N  H�|$E1�1�L�L$8���  �   �N���D�\$D�T$,H���  �D$8���  H�t$H���  D�T$/E1�H���D�\$(L�L$<���  �   Hǅ�      Hǅ      �P��)�f�T$,��  1����H���1�H��H�D$H�|$H���  ����D�\$(D�T$/H���  �D$<��uFH�L$H�|$E1�1�L�L$<�   D�T$/D�\$(�r���D�\$(D�T$/H���  �D$<���o  H�|$ D�T$D�\$�0/���D$<D�\$D�T$���D$8�  �D$,� �A L�E D�\$H�t$E1�ƅ|  f���  H��  H�       @H��P  H   @H��X  H��H�      H���  �   fD���  f���  H���   D�T$ E1�H�@L�D$fD��`  H��8  H�L$Hǅh     Hǅp  @   H��ǅx     HD�H��Hǅ�  D   Hǅ�      Hǅ�      ǅ�  	  H���  L����2�����L���H�L$�D$.L�D$D�\$Ɓ`   D�T$ ���  I��X  I��`  ǁ�      H��H�A     HǁH  @   HǁP      HǁX      Hǁ�   @  ǁ�      Hǁ�      Hǁ�      fǁ�    Hǁ�      Hǁ�     H��  H��  Hǁ      Hǁ       Hǁ(      Hǁ0      ��  ǅ      ���  H��  ���   ���  ��  ���  ��  ���  ��  H��  H��(  H��   H��   H��  H��8  H��0  H��0  H��(  H��H  H��@  @ ��  ���!���f����  �t$.��tK�x�H���  H���  1�H��H��D  H�    H�D    H�    H�D    H��H9�u����  ��t-H���  �H�H�BH���
fD  H��H�    H��H9�u�1�E1�A�   D�T$H�       @D�\$H��P  H   @H��X  H�      f��`  H��Hǅh     Hǅp  @   ǅx     ƅ|  Hǅ�  D   Hǅ�      Hǅ�      ǅ�  	  fD���  H���  fD���  �X5��D�\$D�T$������     H��D�T$D�\$�+���D$8D�\$D�T$���g����'���f���tkA��   D���D$ ������*  �   D�l$A������fD  ��.  D8�)  tJD��)  :T$ tH�t$ @��.  8D$���������Ɓ*   D��D�l$ ��    ��   ����:T$ u��{���8D$�w����}���D�T$H��D�\$H���  H���  Hǁ�      ǁx     H�L$A���  H�L$D�\$����  D�T$���������H�L$H�|$E1�1�L�L$<�   ������|$< D�\$(H���  D�T$/�V���H�L$H�|$E1�1�L�L$<�   �����|$< D�\$(H���  D�T$/����H�|$E1�1�1�L�L$<�   D�T$(D�\$�J����|$< D�\$H��   D�T$(������D$,�D$8    fǅ�    f���  �����ff.�     AW�����AVAUI��ATUH��S��H���  H���   �T$H9��  ���  H�}H�G  ���  �G���  I�E H��M�}(L���   L���   H�D$H��p  L��$�   AT�T$���   AXAYA�ƅ���  ǅ�       �D$zǅ�   stibH��H�E0�D$xH��H�E8H�D$|H��H��H�E@H�D$~H��H��H�EH��$�   H��H�EPH��$�   H��H��H�EXH��$�   H��H��H�E`��$�   H��H�Eh����  ���   ���   H�E�@��   A�   ��H��L��L���O����t$1ҹ   L���<p��H�D$x1�1�I��$h  H���   �?��Hc�$�   H�}P Hc�$�  H�UpH�Exu(H��t#HcL$H��H��H��?H��
 �  H��Hc�H�UPH�}h u H��tMc�I��H�H�� �  H��H�H�EhH���  D��[]A\A]A^A_�@ L�]I�C��A����9  H��t�fD  �؃��D$��  A�   ��@u�L�d$xE1���H��L��L���F���A�ƅ�u��t$1�1�L��ǅ�   ltuoǅ�       ǅ�       �o��A�ƅ��  ���   pmocH��$�   ��  H�PH��$�   H���   H�P H���   H�P(H���   H�P0H�@8H���   H���   ���   ����H���<  ��uGH��$�  ��e   �2  ��h  ��t'��  ����  ���  ���   �     H�\$xL��$�   H�D$   H��$�   H���   ��$�   uH�qXH�VH�T$A���   pmoc�s  I���   H�t$8H�L$(H�D$ �h���H�D$ H�L$(Hc�$�   H�|$8L�D$PI�wpH��$�   H+�$�   �xx(I�@M�GHI�wP�r  H��$�   %   H�  u\H�AXD���  ��tJL��   A�fA9��h  ��H�P�   ��    A�H�pfA9��E  H��H9�u�D  H�D$HH)�L��H+|$@I�G0I�8���   tf��   �I  H�t$��Y��f��h  �H����  ���  ���  )�Hc�H��H)�I��I��?I�I��H���   H�PhH��tEH�H�@H��t9H�zH�L$h�   H�L$XH�D$X    �t$L�D$`�Ѕ��4  L�D$`H�L$hI�Ox��$�   u?Hc\$Mc�Hc�L��H��L��H��?M��  �  H��H��?I��H�� �  Mc�H��Hc�I�WPM�G`I�OhH��H��?H�I�W@H��H)�I�WXH�D$xI��$h  1�1�H���   �����D$������I�EXf�x�������      ����f�A���    A�$   �3���������    H��$�   H�t$8H��$�   H�t$@H��$�   H�t$HH��$�   H�t$P�y����    ���   �����@ A���?����     H��$�  H���}�����+   ������k���D  �PPH�@X���   H���   �S����    ���  ���  )�Hc���������x������    �l���@ H��$�  H�t$L)��W��H��$�  1�L��H��$�  H9������H�t$H)�L�D$ �rW��L�D$ ������D  H��H���   1���������H�������1�1�1�1�I���   f�T$6f�L$8f�t$Xf�|$x�f���I��p  �\$L��1�L�D$XH�L$6L�\$����  L�\$1�M��H�L$8��L����P��HcT$H�D$6H�E0    D�t$XH�E8    H��H�EH    L��Ic�D�|$xH�EX    ǅ�   stibH��L��ƅ�   Hǅ�       H��?H�� �  ǅ�       H��H�E@L��H��?I�� �  E1�H��H�EPH�D$8H��H��H��?H�� �  H��H�E`L��H��?I�� �  H��H�Eh�L���1� �T$H��  �rH9������H��H�DH�   ������ ��I�GP����@ ���   ���   �4����    ���   0�D���@ H��H�wH����   H����   ;V rL���   I�xh ��   ��t[H�vA��A�����    AE�A��A��  �ŀuWE��tA�ȃ�A��	H��AE���t$H�pH�pXH��H���I���f�     ��  u(H�p`H�pXH��H���%���D  ��E��u��fD  H�v��    �@ �$   �f.�     �#   �f.�     �   �f.�     ��G�H��H	��FH��H	�H9��H9Ѻ   G���    H��  ��     H���   H�H��   H�FH��  H�FH��  H�FH��  H�F H��   H�F(H��(  H�F01�Ð��0  f�1�� �   �f.�     H��   H��8  H��1��H���     H��P  H��t\D�I�1҉F1�D�E��tA�    H�|�H��H�|H���   L�L�DD���   J�|��H�|H��A9�w�1�� �   �f�L��P  M����   ��u<H��u7A� ��t,�H�I��  I��  1�� H��H��H��H�PH9�u�1�ÐH����   SE���A9�AFم�t*M��  D�S�1��
�    H��H��I��H�HL9�u�A9�v/A��I��  ��A)�I�H��J�T� H�     H��H9�u�H�G��t�̀H�G1�[�D  ��H�G1�[�D  �   �f.�     H��P  H����   �>D�D9�rf1�E��t&L��  E�B�1��H��I��H��H�HL9�u�D��9�v%��A��)�J��L�H�T��H�     H��H9�u�D�1��f.�     D��   ��    �   �f.�     H��S1�H��1�1�H���Ph��`  [�D  ���  ��     AWAVI��AUI��ATA��USH��H��H�o�W8H�H9�vW� ��0��	wLH���SHH��I���S@H�H�PI�M��x.H)�L9�~&�SI�GH1�M�} ����H��[]A\A]A^A_�f�1�E��u��C   H��[]A\A]A^A_� H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ USH��H�GH��p  H��t.H���   H���P�F H�x�2���H��tH���UH��(  H�B@H��1�[]� AWI��AVAUA��ATUSH��H���	  H�oH�L$L��  H���  I�FH�$H���   L�`hH���  H���
  H���  H���
  H���  H���
  H���  H���
  H���  H���
  H���
  M���v  I�$I�|$L������(  ���    �3  �   H��H��$�  A�V0H�D$H��8  H��H��A�V8H�D$IcWI�7H��$ 	  H�$H��$�  �P<�u2H�CH��$�  ƀ0   H�D$� H�$IcWI�7�Pf�     ����   M����   I�$H�z t|H�{@�kM��H�{PH�D$     H��H�D$�PM��H�{XH��H�D$(�>M��1�I�|$D��H��H�L$H�D$0I�$�PH�T$H��H�S@H�T$(H��H�SPH�T$0H��H�SXH���	  []A\A]A^A_�fD  H�$A�WH��I�7�P�:���f.�     H���  ��H��I�H���  ��A�G���    ������ SH��H��0H�L$H�T$ �D$ ������u+H�SH���   H�RhH��tH�zH��D$H�t$ �R�D$H��0[�ff.�     @ AV1�1�AUATI��UH��SH���  L��  H�    H��L��P  L���  I�Fh`B j j H�|$(�H�� A�Ņ���   ��`  Ƅ$�   1�Ƅ$�    ��$�
  H��h  H��$�
  H��p  H��$�
  H��x  H��$�
  H��h  H��$�  ��`  I�$    ��$�  ���  ��~- ��H�|$����H�D$X��tI;$~I�$��9��  �I�FH�|$�PH���  D��[]A\A]A^�ff.�     @ AUATA��USL��H���  ���  H��  H��I����L��P  H��1�1�H�@L���  h`B j j H�|$(�H�� ����   A��`  Ƅ$�   Ƅ$�    ��$�
  I��h  H��$�
  I��p  H��$�
  I��x  H��$�
  I��h  H��$�  A��`  ��$�  E��tKA��D  ��H�    H��A9�t.��H�|$�y�����u�H�|$X��H����I��H��H�C�A9�u�1�H���  []A\A]��    ��t�B�I�D�@ H�    H��H9�u�1���ff.�     �AWAVAUA��ATA��UH��SH��H��P  L���   �D$    H����  E���y  ���t#D9��j  H���   []A\A]A^A_�fD  E��L�L$E1�1�L��8   L���{���H��   �D$���_  L�L$E1�L��1Ҿ�   L���N���H���  �D$���2  L�L$E1�L��1Ҿ    L���!���H��8  �D$���  1�C�$L�L$E1��   L�������H��H��  �D$����   J��H��  H���   H��  H��8  H���  H���  H��0  A��vTA�T$�H��   H���(  fD  H�8H��H�W8H���   H�H���   H��  H���   H�W H��  H9�u�D�# �k������E��tA9�t���z���D�kD��   D�#E��t��tH�{( tU�D$H��[]A\A]A^A_�f.�     H�T$�   L��莩��H�ËD$��u�ǃ�      H��P  �����D  D��   L�L$E1���1�L������H��H�C(�D$��u�A���y���A�L$�H�S0L�D�8���H�s(��H���H�4�H�r�I9�u��I���f�AW�   AVAUATUH��SH��H��  L��P  H��H�t$ H�L$�Sx�t$��   ��x t6��1M��t4A���t-�   9���   �CH�Ĩ  []A\A]A^A_� �   ��1�H���������u�H�CL��P  L�3H�D$�D$��~GL�d$ 1�I�$1�H��I��H�I�D$�H�CI��  L�,��SPI��  I�E H��H��9l$�H�D$L�3H�C1��]���D  H�CL�3H�D$�f.�     AWI���   AVAUATUSH��H��(  H�|$H�L$8L��H��$�   A�Wx�T$8��   ���2  �R  ���I  I��D$    �D$    H��P  H�D$ I�GH�D$(H��$�   H�D$fD  H�L$�   H�t$@L��H�I�H�AH�L$<I�GA�Wx�D$����   �T$<�B��T$����   H�\$�t$8H���F�������   H��P  �D$<LcT$H�l$@E1�M�r��~:fD  H�E 1�L��H��I�H�E�I�GJ�D�N�$�I��A�WPI�$D9l$<̃D$�D$H�D$9D$8�+���H�D$ I�H�D$(I�G1�A�GH��(  []A\A]A^A_�f��D$9D$<�_����   ��ff.�     AWI���   AVAUATUSH��H��  H���   L��H�L$8�D$4    H�t$@H�D$A�Wx�T$8��   ����  ��  ����  I�1�H��H�D$ I�GH�D$(�������D$4���[  �D$8H��P  ���7  H�D$@�D$    H�Ũ   H�D$f.�     H�|$H�L$<�   H��$�   H�I�H�GL��I�GA�Wx�L$<�A����  H�} ��   �H�|$L�L$4E1�Hc�1Ҿ   �[����L$4H�E����   HcL$<H��H��H�M�U ��~gL��$�   E1���    H�EI�u I�ML��I��N�$�    I��H�VJ� I�H�Q�I�WA�WH1�L��H�H�]A�WPL�H�D9t$<��D$H���D$H�D$9D$8������L$4H�D$ I�H�D$(I�GA�OH�Ĉ  []A\A]A^A_�D  �   ��f�     UH��SH��H��H�vH����H�CH    H�s8H���CP    ����H�C8    H��H���C@    H��[]�p���AWAVAUATUSH��H��P  H���o  L���   D�3I��H�s(�kL���6���H�C(    A���T  A�V�H�C0H�T�8�    H�     H��H9�u�H���  L�������H��   L��Hǃ�      �����H��8  L��Hǃ       ����1�Hǃ8      HǄà      HǄ�      HǄ�0      H��A9�w�H��  L���t���Hǃ      Hǃ      ��t]D�}�L�sJ�l�I�6L��I���>���I�F�    I9�u�K�H���   H����   H�u L��H������H�E�    �E� H9�u�I��P  L�������IǅP      H��[]A\A]A^A_�@ H���  L�������H��   L��Hǃ�      ����H��8  L��Hǃ       ����Hǃ8      E�������Hǃ�      Hǃ      Hǃ0      ����� AWI��AVAUATUH��SH��8L��  H�^H���V8M�7L9��  A��PЀ�	vK<[tGI�FH9��2  �Y�F �   L����� ���  ǅ      H��8[]A\A]A^A_�D  I�O H�$<[��  L��A�   A�WH�D$ =   �D$DN�L��A�W8I9s�H��8  I���   H�D$H��tDH�<$�l���H��@  H�<$Hǅ8      �Q���I��   Hǅ@      H��t	I���   ��D��(  Mc�H�<$1�L�L$,E1�L�Ѿ   E���   L�T$谿��H��8  �D$,����   A�GH��8[]A\A]A^A_�f.�     I�FH9�vG�j�F �   L����� ��u/ǅ      �����A�G   H��8[]A\A]A^A_�f�     I�FH9���  �y�F �   L����� ���w  ǅ      �l����     L�T$H�<$L�L$,1�E1��   L���о��H��@  �D$,��� ���I�E H�$D��I���   ��D$,��� ���E1�E��~7H�$D��M���   �    �ރ��   ���F L��A��  A9�u�H�$L��A�W8M�/L9���  D�t$H�l$L���$    D�d$�]�    <]��  ��0��	waE����   L��A�WHL��I��A�W8M�/I9���   I�EH9���  L��A�W8I�/H9��b  �E <du�L�mI9�s
�}e�  E��ubL��A�W@A�G������I���f.�     A�G�   H��8[]A\A]A^A_�f�     I�F�D$A�   I��D$   �����H�EI��H9�v�} /u	�$9L$A�G   �����     A��I��L��M�/A�W@I�H9��w���A�W���k����$9L$~;L)�L��D��H�|$H�ōHA��  A�G���;���I���   Mc��J��� �$�����f.�     �}f������E<>wLH�6  !� PH�������f.�     H�l$M��ǅ      M�7�����fD  I��H�l$M�u�ڃ�߃�[���}�����A�} /�B����$9T$�5��������D  AWA��AVI��AUA��ATUSH��H��8  H�o�D$' H��  H�@H�D$;U rH���   H�xh ��  A��   ��  A������M����  I�F H��8  I�F(H��@  D��H����0  L��ǃ�       ��ǃ�   ltuo�ƃ���1  D���L��P  ��@�t$&L���  H���h`B PQH�D$(H��H��$�   �H�� A�ą���  ��`  D��H�t$'H�T$(��   H�|$x��$  H��h  �L$H��D��H��$  H��p  ��$�   H��$   H��x  H��$(  H��h  H��$  ��`  ��$  �]���A�ą��b  H��$0  ��0  H�|$xL��$P  H�D$8H��$8  @�t$H��$X  H�D$@H��$@  H�t$H�D$HH��$H  H�D$PH�D$�P���   �T$�������   ���  H��$�   �8��H��$�   H��H�CP�8��H��A��H�CpH��(  D�l$�@ �F  H���  H+��  H��H�ChH�Cxǃ�   ltuoM��tfA�~w
���      H�|$8   L���   uH�|$P   �"  H�t$8L���z��HcCPHcT$8H��H�H�� �  HcShH��H�H�CPHcD$PH��H�H�� �  H��H�H�ChL�t$L��L	�tL��L��L���Xx��L{PLsh�|$ u�|$' tj�|$ Hc�@  Hc�8  ��  H��$    ��  HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$XL���w��H�T$XH�D$hH)�H�S@H�C0H�D$pH��H�CH�D$H+L$`H�K8����   H�shH�{0�(T���    A��1�1�M���l���Hǃ8     Hǃ@     �g���@ H��$�   L��(  �|6��H��$�   H��H�C@�g6��H�t$H��H�CPH�D$8I�u8I�EH�D$@I�EH�D$HI�E H�D$PM�}0I�E(A�EH�D$(H��   HcD$0H��  H���   H�@hH��t%H�xH� H�t$(�PHǃ       Hǃ      H��8  D��[]A\A]A^A_��    H�D$H�|$x�P�ՐA�   ���     H��$�   �Pf���1����z�H�@H��H��H�f�     HcH��H��I��I��?J�� �  H��Hc�H�P�HcP�H��I��I��?J�� �  H��Hc�H�P�H9�u�������    H��$�   �5��H��$�   H��H�Ch��4��H��H�Cx����f�     H�D$@HD$H���������ff.�     H���G  USH��H��H��h  H���   H��tH���C���Hǃh      ǃ`      H������H���   H��HǃP      ����H��   H��Hǃ�       �����H��  H��Hǃ       �����H��  H��Hǃ      ����H��  H��Hǃ      ����H���  H��Hǃ      ����H���  H��Hǃ�      �p���H���  H��Hǃ�      �V���H��h  H��Hǃ�      �<���H��p  H��Hǃh      �"���H��x  H��Hǃp      �hD��H��x  H�������H��H  H��Hǃx      �����H��P  H��HǃH      �����H��X  H��HǃP      ����H��8  H��HǃX      ����H��@  H��Hǃ8      �w���H��  H��Hǃ@      �]���H��  Hǃ      H��tH���~���H�C(    H�C0    H��[]��    �ff.�     @ ���  ��~cAUD�h�ATUH��S1�H��L���  �f.�     H�CL9�t'H��I�4�H���h�����u�H����[]A\A]��    H��1�[]A\A]�1��AWI��AVAUATUSH�
H��8H�H�|$H��H�^�F    �V8M�7L9���   I�6  !� PE1�1��xD  <c��   I�F
H9�tv=A�F	<>�(  I��s*f.�     ���F �	   L����� ��tx�     I�W@L����A�G��ucE1�L��A�W8M�7L9�vMA�<eu�I�FH9�tv�A�F<>��  I��s��    ���F �   L����� ��u��     A�GH��8[]A\A]A^A_�D  <FuiI�FH9�t#�e���A�F<>�h  I���N���fD  ���F �   L����� ���,���A���  �t
��A���  I��M�7�����Ѓ�0��	w(L��A�W@A�G���a���L��A�   ������    <RudI�FH9������A�~D�����E�������H�D$I�/1�H�T$(H�t$ L��H���   H�xh ���x�����������   �����fD  <-uI�FH9��_���A�~|t��S���I�W@</�K���I�FH9��>���M�fL��M�'��A�G�������I�H��L)�J�������H9�����A�F��A�|�F A���F H�t$�D$�v   ��I��0M�M�������A� 8D$u�L��L�D$�y���H9D$L�D$u�H�T$L��L������L�D$��u�A���  �Ѓ���A�F(�������t���F �   L����� ���k���H�D$H��P  1�H��t�
��HE�A�v��t^A�~��   A�N�$���F ��߃�[���b�������D  ��߃�[������������D  ��߃�[������������D  L��H�|$A�VA�GA�G�������<��(���A�G    E1�����H�T$(1�H�T$(H�: tރ�	E1�L����L��v	A���   �A���   �H�D$H�   H�D$(1�H�T$(�H�L$H���   H�T$(H��t�H��  ��H�D$1�H�T$(H0  H�D$(�H�D$1�H�T$(H�D$(�n���L�|$(1�H�T$(�]���H�L$H���  H�T$(H��t�H��0  ��9���H�L$H��8  H�T$(H���X���H���  �����f�     AU1�ATI��UH��SH��H��f�H�    H�t$�W��A�ŋD$��uA���  f��vfD�+H��[]A\A]�H�t$H���c���H�D$��u�I�$��f�AW�   AVAUI��ATUSH��L��H��x�D$    H�L$H�t$A�Ux�T$��   ����   ��   ����   1�H�������D$����   �T$L��P  L���   ����   L�|$1��YD  I�t�H��tL�������sH�T$L���ލ��H��I�D��D$��uC��I�7H��H��H��I������� 9l$~<I��8/uH��I�I�_H)Å�u�f��   A�EH��x[]A\A]A^A_��     �D$��f.�     AWAVI��AUATI��USH��hH�F L�.H�^H�D$H��  H��H�D$�VH���B  H�ډ�H�L)�H��H9�O����  A�v����  I���  A��(  H�D$(I��0  H�D$ I���  H�D$8���  �D$3 E1��D$4    �    L��A�V8M�>L9��  I�GH9�v<A�G<>�g  H�6  !� PH��sA�<d�e  <euA�n��  @ L��A�V@M�I9��e  A�V����  A�?/u�I�GL�D$H9��A  1�H�T$XH�t$PL��I��$�   H�xh ����������  A��(  ���6���L�D$I�WD��H�|$ I)�A�HL�D$A���  �D$L����  I��X  Ic�L�D$H��E��B� A�.u?I��X  ���F �   H�<��L$4�t$3�� �����   AD�D��L$4@�t$3Ic�$<  H�L$P����  �UD9���  H9��K  H�|$H�T$LH������I�ǋD$L���/  H�T$PH�t$XL�������H�D$��  L��H�t$P�P H�L$PD��H�|$(Ic�$<  H)�L�H�L$PA���  H�|$L���D$L�K����D$L�r  f�A�d�=���D  E����  I��X  �|$3 E��(  H��  I��`  H�\$8�D$\1��D$X���H�ߋA��@  �D$L���]  I���  I���  �   H�ߋ
H�A��@  �D$L���/  H�\$ �   ���F 1�H��A���  �D$L���  L�|$(�   H�T$X1�L��A���  �D$L����   I��   I��  D��H�ߋ
H�A���  �D$L����   I��   D��L���HI��  H�PA���  ����   A��(  H��h[]A\A]A^A_��    H�T$XD��H�|$(A���  �D$L��uQA���s��� ��߃�[�������A�<d�����A�e�����A�f�����E��������[���f��   A�FH��h[]A\A]A^A_��     L�|$D�mH�T$I���  D��I���D$L��u�I�H�T$D��I��0  ��D$L��u�I�H�T$�   I���  ��D$L�������뀾��F �   H����� �������I��`  L�|$81��L��A��@  �D$L���>���I���  I���  �   L���
H�A��@  �D$L������Hc\$4I��`  �   L����I��X  H��A��@  �D$L�������I���  �   L����I���  H��A��@  �D$L�������I��   I��  ��L�|$ �
H�L��A���  �D$L���{���I��   ��H�\$(�HI��  H��H�PA���  �D$L���I���I��   1�L���HI��  H�PA���  �D$L������I��   1�H�ߋHI��  H�PA���  ���p��������f�     AWI��AVAUATUH��SH��HH��  L�v H��H�D$�V8I�L��I;Gs	�8[�y  A�WH�D$����  I�WI�H9�r H)�H�H��H9�~I���   �T$��  L��A�W@A����  I��X  L��H�D$A�W8A��P  ��u$H�D$L��t$I��X  H� ��D$,���  I�7H�FI9G��  E1��   �    H9���  H�T$,L��躅��I�ŋD$,����  H�T$0H�t$8L������H�D$��  L��H�t$0�P H�L$0��H�|$Hc�<  H)�L�H�L$0A���  L��L���D$,������D$,���q  I�7A��H�FI9G��   �   ���F ��� ����   L��A�W@L��A�WH1�H�T$8H�t$0H��H���   L��H�xh ���r�������   L��A�W@A�O����   L��A�W8I�7H�FI9Gv#���F �   ��� ��uL��A�W@L��A�W8I���  H��tE���L��L��L������A��P  ������Hc�<  H�t$0���~�����H�T$8��H�|$A���  �D$,�����A��P  ��u�D$A��P  H��H[]A\A]A^A_� A�W@L��A�W8I�I;Gs�8]t�A�G   H��H[]A\A]A^A_ø   A�GH��H[]A\A]A^A_�L��H�T$,�(   讃��H��I���  �D$,��u�L��账���D$,���C����fD  L�GL�WI�H9�}PD�A��v<I�HH9���   A����H�<�   �   � H�PI�L�H9�}"H��H9�u�K�D��H���I�H����     I�T �M�L�UH��H��SH)�H)�H��I�I�,��!��H��H)�H��H��H�[]�M�Ѹ   ��f�     AT�   UH���   SH��H��H��0H���Uh���  H�D$H���  H�I��I1�I)�I��   ��   L���  �s!��H�<$L��f���   �`!��H�|$L��H�$�O!��H�|$L��H�D$�=!��H�|$ L��H�D$�+!��H�|$(L��H�D$ �!��H�D$(H�D$H��?H%  ��H   H�D$H�$H���  H���  H���  H�T$H���  H�T$H���  �t&����t0H�D$ H��H���  H�D$(H��H���  H��0[]A\��    �E   H��0[]A\ÿ �F ��2��fD  AWAVAUATUSH��L��  M����   A�D$@I��A��I��1ۅ�u�M@ H�EI���A9\$@v8��H�<�I�D$8H�,�D9m u�H�EL9��H�UH�u L9�}$I�7��A9\$@w�H��1�[]A\A]A^A_�fD  L��H)�H+uH)�����HEI��D  H���   []A\A]A^A_�@ AUATUS�    H��M��II؃�-w��I���$��F 9�`  �9  D  H������H��H��[]A\A]� H����  H����  ��0  �   f���@ H����  H����  ��,  �   f��@ H����  H����  ��*  �   f��x���f�     H���W  H���N  ��(  �   ��J��� L��  H�L$M���+��� L�������H�L$H�hH������H9�����H��L��H���?��������f.�     L��  H�L$M��u������f.�     L��  H�L$M��u�����f.�     L��   H�L$M���k�������fD  L���   H�L$M���K����n���fD  H����  H����  H��   �   H��H���f�     H����  H����  H��  �   H�����f�     �������H���  H����  �н   ��G  f������D  H����  H����  ���  �   ����� H����  H����  ��<  �   ����� H���o  H���f  ���  �   ��b��� H���_  H���U  ���  �   f��8���f�     H���/  H���%  ���  �   f�����f�     H��x  H���������H�L$��,��H��������H�L$I��$h  H���������I��$p  ���jH��tH9�rH�U�H�4�H��������D(� H�������H��H��[]A\A]�D  H����  H���}  ��`  �   ��R��� ��   �;���H�L$9�(  �*���H��@  ��L�,�L�������H�L$I��H�hH������H9������H��L��H���1���B�  ������    H����  H����  ��   �   ����� 9��  �������H���  ���jH��� ���H9������H�U�H���  ����� H�L$9��  �_���H���  ��L�$��%���D  H���_  H���U  ���  �   ��*��� H���7  H���-  ��8  �   ����� L��  H�L$M������������fD  H����  H����  ���  �   ����� �������H��t-H��v'����  ����  ����  H���  f�H��   �r��� H���W  H���N  ���  �   ��J��� H��t�H��v�H��   �   H��(���f�     ������H��t�H��v����1  ���  ���+  H���  �e���D  H����  H����  ��C  �   ����� H����  H����  ��B  �   ����� ��A  9��y���H����  H���v  �н   ��G`  f��V����    H���7  H���.  ���  �   ��*��� H���7  H���-  ���  �   ����� H���z���H���p���H���  �a������C  9������H����  H����  �н   ��G�  f������    H����  H���~  ���  �   ��z��� ���  9��a���H���h  H���^  �н   ��G�  f��>����    ���  9��!���H���(  H���  �н   ��G�  f�������    H����   H����   ��A  �   ������ H����   H����   ���  �   ����� ��@  9������H����   H����   �н   ��GD  f��n����    H��tSH��tN��@  �   ��J��� ��B  9��1���H��t<H��v6�н   ��Gt  f������    H���   [H��]A\A]�D  �   �����fD  �   �����H���  �R���H���  �F���H���  �:���H���  �.���H���  �"���H���  ����fD  H��H�Љ�H���  ��H��H�4��B���1�H���ff.�     H��  H�    H�A    H��tlL�@H�@P����H��H��H	�L��H��H�s�H�L�@I9�w>H��L)�H��H��H��?H�H��H��L��8D�HH��L	�H9�tH9�w�H�p�I9�v�1��fD  HcPHc@H�H�A1��ff.�      H�O����   L�G����   L�W8L�O(����   H�GhHGxHGXHGHL�L�L�H�H�H�GpHGxHGXHGPHG8HG0HGHGH�FH�GpHGxHGhHG`HG8HG0HG(HG H�FH�GpHGxHGhHG`HGXHGPHGHHG@H�F�f�     I�H�H�GHGH�F�@ H��@ K�L�H�H�H�G0HG8HGHGH�FH�G0HG8HG(HG H�F�f.�     USH�� H��P  H��t~H��H��  �UA��H������D9]D��FU��t1�D  H��H��H��9�w�A9�v+A����A)�H��I�J�T�fD  H�  �  H��H9�u�H�� 1�[]��    H�� �   []�@ AVAUATUSH�� H��P  H����   I��H��  �UA��H��E���	���D9eDFuE��t)H�Ũ   1�f�H�4�H��H���`���I�D� H��A9�w�E9�v-A��D��E)�I�D� I�K�T�fD  H�     H��H9�u�H�� 1�[]A\A]A^ÐH�� �   []A\A]A^�ff.�      AVAUATUH��SH��   L���   H��P  H�t$(薾���D$��tH�Đ   []A\A]A^�fD  �D$(H�T$L��H�4@H��H�� �s��I�ƋD$��uD$,�T$(A�F    I�F    A�FI�F A�I�F����   ��L�D$(H�RH��M�TP@ I�PM�HH��L�H�PI�H�@(����H��H�H�H�����H��H�H H�PM��t%���F �   L����� ����   H�@ thgwH��0I��L9�u��SH�t$H��  E1�H�è   �*����D$(��t,J�t�O�,dH��I��I��MnH������I�ED9d$(w�L�u �D$H�Đ   []A\A]A^�fD  ��F �   L����� ��uH�@ htdw�]���f����F �   L����� ���>���H�@ zspo�1���fD  H���  AW�����AVAUATUSD�o�A9�AF�A������   �D$� D�q�1�E�M�L��  �   A�   �    A��1ɸ   E��uS�g�    H�4�A��L��A��H)�E��HD�H��~dH����  H�H��H��H��?H��0 �  H��H�qI9�tH��A9�w�H��H�qI9�u�D  I9�t	I���D$�H�EI9�tH���h���1����D$�������[]A\A]A^A_ø   �ff.�      AWAVAUATUSH��   L��P  M���v  A��A�vI��H�|$D9�DF���%  I���   1��     L�ML�]D�} A9���   I�|� E��E����   I;9��   ��   �   E1�� �    I�H9�toH��H9���   Lc�A�@D9�u�K�D��H�D�H��H��9�w�H�\$H�T$H��P  �������uH�SE����   �΀H�SH�Ę   []A\A]A^A_�I�I���     A��I�D��I+H��H��?H�H���-���f�K��I��I�4�K+4�H)�H)��5��A�v�[���1�H�T$L���m����������H�D$H�PH�D$��H�P1��g����   �]���ff.�     @ AVAUI��ATU�   SH�� ��F�I���t(I��1�I���    I�<��g��H��I��H��9�w�L���L�������H�� []A\A]A^�ff.�     f�U��SH��H��P  ������uH�SH�р΀����HD�H�S[]�ff.�     @ 1�1��f.�     SH���   �P�F H��p  H�x�?��H��tH��tH�H��t	H��[�� 1�[�@ ATI��USH��H�?����H�;L��H����*��H��tH�CPH�S(E1�1�H�s H�8�U[1�]A\�ff.�     f�SH��H��H�?�`���H��1�H��t(H�H�T$H��8  H���   ���uH�SPH�L$H�
H��[��     H�GPH�8 t.SH��H�?�
���H��t
H�SPH�:�PH�CPH�     [�fD  ��    AWAVAUATE1�USH��H����  wk���  ��~aH�t$I��D�x�1�L���  �D  H�CI9�tWH��I�l� A��H��t�A�8E u�H�������H9D$u�H�T$L��H���������u�H��D��[]A\A]A^A_�f�     E1���ff.�     AWI��AVAUATUSH��H��XL�f8H��  �D$    H��tL�������Hǃ      H�T$ �X   L����k���L$ H�Ņ�t$H����   �D$ H��X[]A\A]A^A_��     I�wL����X���D$ ��u�H���  L��  H�EH���  H�EH���  H�EH���  H�E H���  H�E(H���  H�E0I�EHH����   I�OHI�W@H�|$(I�w8��D$ ��t;<uI�GH��vI�W@�z�  �    L����Y��H��L��������%���H���   H�|$(H�l$8H�D$HI�EHH�D$@0HB �PH�|$(�D$ I�EH�P�D$ <t���u�H�EH���  H�EH���  H�EH���  H�E H���  H�EH��H�ChH�EH��H�CpH�EH��  H��H�CxH�E H��  H��H���   H�E(H �  H��f���   H�E0H �  H��f���   �EP������H�K@L��H��  �X���*���D  �JH9������I�G8I�OH�D$$    H�D$H�BeH9���  �Bd�����Bc	���H�DuH�pH9���  �p���0��	�f���i  �@H�H9��Z  L�pL9��Z  �P�����	��EP��L�H9��7  f���!  H�|$��E1�1�L�L$$�   �b����|$$ H��H�EHH���	  �EP�KHD�,�    H���   M�H�D$��~6H�CPH�0f�~��   H����H���H�0H��f�~��   H9�u�M9�sVA�6H��H�T$I���\/��H�T$H�߉A�v��H/��H�T$�BA�F�H������A�F��B�    	Ș�B�M9�w�H�|$ tH�t$H���5���D$$�|$$ H�}Hu3�uP�   ���A ������T$$��u`�D$     �b����D$$   H�}HH��H�|$臮���D$$H�EH    �EP    �D$ �)���H��H�T$�>5��H�T$���D$$����H�}H��    ATI��1�UH��SH��H�� ��R����tH�� []A\� H�T$H�t$H���f�����u�f�|$�t1�H���R����u�H��H���T����u�H�{@H��L�������   H�߅�ED$��U���D$H�� []A\�f.�     AW1��Y   1�AVI��1�AUATUSH��8  H��  M���   IǆX  ����H�\$hM���   Aǆ`      Aǆ<     H���H�L��H�      H��I���  Iǆ�  \  H�EIǆ�   �' �E1ɺ   ���F L��L��$�   HǄ$       HǄ$      HǄ$      HǄ$      fD��$   Ƅ$"   �o����D$X���1  <�  ��$!   �D$X��  �D$PH��$�  H��$�   H��t	H���   ��H��$P  H��t	H���  ��H��$�  H��t	H��0  ��H��$�  H��t	H���  ��H��$  H��t	H��X  ��H��$   H���_��H��$   H������H��$�   H��$  HǄ$       H���˫����$!   HǄ$      ��   H����$�   �D$PH��8  []A\A]A^A_Ð�
   �̷F L���>����D$X�������1�L���(P���D$X�������L�l$`H�t$TL��L�������D$X�������f�|$T���   1�L����O���D$X���}���I�t$H�t$`�y@ H��$   H�������HǄ$       �6����    H��$   L���Ъ���D$XHǄ$       �D$P���/���H��$  1��   D  Ƅ$   H�t$`I�|$( ��  H�D$XL��H����c��D�D$XH��$   E�������H�T$`H��L���QP���D$X�������H�L$`H��$  H��$   �D$P    H�
H�T$pH�T$hH�D$xH��L���j����D$P���y�����$    L��$�   �D$T    L��$�   �x  H��$   H��$  I��H�1��    I��L9��;  A�<$eu�I�T$	H9�v�A�|$eu�A�|$xu�A�|$eu�A�|$cu�I��
H��H�L$hL�d$xL9�r=��  �    H����$�   ��$�   ����  H����$�   H�D$hI9���  �8eu�H�PI9�v��xeu��xxu��xeu��xcu�H��$  H�$   H��H�D$x��$�   L�d$xL�l$h�
   L��L��L)�H��H�L$�}���H�L$H���"  H�ʾ   L��H�D$�Z���L�D$I9�������M9��  A�U �J�����  �� ��  ��u����  H��$   H��L)�H�$  ��$!   H�D$X��  Ƅ$"  H��$  H��$  HǄ$       HǄ$      I�EI9��p  A�E �PЀ�	v��߃�A<�U  A�E�PЀ�	v��߃�A<�:  A�E�PЀ�	v��߃�A<�  A�E�PЀ�	v��߃�A<�  H�EH��L�l$hE1�H��$  H��$  H�L$`�P0H�D$`H��$  H��$  � H��$  H��$  �q�  �U H��$  ��  H��$  �  H��$  �@ H��$  �@ H��$  �@ H��$  H��$  H�T$pH�
H�T$hH�D$x�D$T�D$P���9���H��L�������D$P���"���I��P  A��@  �H���?  �H�   ��9tL���	���I��P  H���  ����  ��t;Ht
ǀ�      ��t�p��uL���˻��I��P  H����  �P��t:���    ��  ��H�RH���f.�     H�����    �  H9�u�A��`  ���;  H��$�   ��$�  �D$8A���  tb��$�  HǄ$�      A��`  H��$�  I��H  H��$�  I��h  H��$�  I��p  H��$   HǄ$       I��x  I���   H�xh ��  H��$�  A��   HǄ$      I��P  H��$   I���  H��$(  I���  H��$�  HǄ$�      I��X  H��$�  HǄ$�      H��I���  ��  A���  �  vAǆ�     A���  �  ����Aǆ�     ����H��$  H��$   H�1I9������@ �   �����fD  L��L�l$`��I��H�l$H�D$H�D$XHǄ$      H��H�D$�*fD  H�t$XL��H�H��$  � I���D$T���{���H��L��L���V����D$T���a���f�|$`�H��$  t�H�l$H���k  �D$P   �9���fD  I�D$L��I$H��$  H��$   Ƅ$!  �H���D$X�������H��$  �>���fD  L�������I��P   �p���f.�     Aǆ`      �e�����$P  ����  H��$X  ��L�t$HE1�H�D$(�D$8H�L$ I��8  ���D$<    H�L$I��@  I��H�D$@H�L$� I�D$L9d$(��   I��H�D$ 1�N�,�H�D$fB�`H�D$J�ࢥF A�D$�D$M��t��D$8��~�E1�L�d$0M��L�|$@� I�D$M9�tnI��K�,�L��H��������u�M��H�D$L�d$0H��   ���F fF�<`H�D$J�,��L$<�� ��D9��A������D$D��D$<�/����    L�d$0����fD  L�t$HAǆ,      �D$<A��0  ��$(  A��(  � ���f.�     H��$   �g����D$P   �Z���@ L�L$PE1�1Ҿ   I���   �5z���L$PI��h  �������Aǆ`      �����f�H�t$L���F���D$T�������H��$  H�T$TL���Z��H��$  �D$T�������HǄ$      L�|$�5 f�|$`�uOH�T$XH�L����F���D$T���Z���H�D$XH�$  L��L��L���(���H��$  H��$  �D$T��t��D$T    �l����D$<    ����I�������   �����H��$  H�T$XL��莮��H��$  H��$  �"���H�pH�T$TL���Y��H��$  �D$T�������H�D$XH��$  �"���f�AVAUATU�պ   SH��H��H�   H���   �׷F �"+����F H��  I��H���   H�x��*��H��  H���{  I��H���   �P�F H�x�*��H��H��p  �����A�Ņ���  ����  ����  ��  Hc��  H�C    H�C H�CH��H��
  ��(   H�St
H
  H�CH��P   tH�K   H��  H�C0    H�K(H���O  H��  H���O  �@ ��t4�1@8���  < ��  <-��  @�� t
@��-�   H����u�H�C0�F H��    H�C    H��  tH�C   H��t:� �F �   H����� ����  H�ƿ��F �   ��� ����  �H���  H���  �C8    H�C@    H��H��H�ChH���  H�{pH����  H���  H��H����  ���   H�sxH��H���   f����  �@A���������A����A������D��f���   )�D)�f���   H��9�f���   H��AN�f���   ���������  ���   f���   ��*  ���   M����   M�f@1�H��1�H�cinu  H�$H�D$I�|$�n{��A�Ņ�t��=�   t��uZ��   �   f�|$����  �	  ����  ��u*�   �D$EBDAI�|$f�L$H��t1�H��1��{����A��H��D��[]A\A]A^�fD  H��  H��tH�C(H��  H��   H���	  H�C0H�C    H�������������    H�K����fD  �BH��H���_����    �BH���K��� H��A�   [D��]A\A]A^�f�A��  ��  fD���   A��  �8���f����&����   �D$CBDAI�|$f�T$����� H��A�   [D��]A\A]A^�f�H�<$����H��f���   �����    @�������H�S0�����fD  1�H��H�C0�F ��H�C�����    �   �D$1talI�|$f�D$�h���@ 1��D$BODAI�<$f�t$�L���H�H���  H  H�G1��f�     H�G    ��    1����   w
H�G���p�ff.�     �1��    ���   w"H�O���    �Q��uH����   u�� ��D  L�H��I���  H��    H��`  t"L�RM��t)�P$I���   E1�� wB A��@ ��   �f.�     �   �f.�     H�H���  H��`  �`ff.�     �H�H���  H��`  �`ff.�     �H��p  H�    H�A    H��tSH�����   H�H�1�[�f�1��ff.�     f�1��G���fD  H���  � H��t��L  ��  t�1��ff.�     @ H���  1�H��t2��L  ��  �   t!9q$v1�H��tH��   ���q�
�D  �ff.�     @ H���  �`fD  H���  �`fD  H���  �`@fD  H���  �`HfD  H���  �` fD  H���  �`(fD  H���  �`0fD  H���  �`8fD  H���  � �    H���  �`8fD  ���t`��t���   #��u���H��f�H�V1�H9Wv8�Fȉ��@ L�FH�O1����   ~FI9�s��   )��V��)Ѓ�lH�� H�V1�H9Wv��F�����F	�H����     I9�sρ��   �F���DlH���    1����   w
����? �F �ff.�     H�WH��t�����   <t1��D  ��+G;G��   D�D�WD��D�BI���A	�E��D9�r�D�J�BH�JE��D�JA��E	�E��D9�s-�Nf�     �H���Q���A���Q�D	���9�r,A��I9�w��l���@ ���2�f�     �G�D��E��D)�D�O�W�G��    H���  �`PfD  H���  H��t�`X��ff.�     @ H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ SH�H��H�w H���   �	���H�C     �C    [��     AUI��ATUSH��H��H�wH��t2�W��t+1�fD  A��L���J�4�趕��H�sJ��    9kw�L��蝕��H�sH�C    H��t6���t0E1� D��L��A��H��H�t.�h���H�sH�D.    D9#w�L���N���H�C    H��[]A\A]�ff.�     USH��H�GH���  H��X  H��t.H���   H���P�F H�x���H��tH���UH��(  H�B@H��1�[]�ff.�     �H���   1�H���H���H  @�~��t�H���P  f�LFH��9�w���I  @�~	��t!1�f.�     H����  f�LF(H��9�w���J  @�~
��t!1�f.�     H���  f�LF<H��9�w���K  @�~��t!1�f.�     H��  f�LFXH��9�w�H���  H�FpH���  �FxH���  �F|H���  f���   H���  f���   ���  @���   ��t1�@ H���   f��F�   H��9�w����  @���   ��t1�@ H���h  f��F�   H��9�w����  ���   Hc��  H���   ���  �F�ff.�     H�H��tXUSH��H��H�8 H�h8tH�w8H���9��H�s0H������H�{H�    1�H���H�C8    H)��K@���H�H��[]��ff.�     @ H�GH=@�F tlH=��F tdUH�����F SH��H��H�H���   H�x�(��1Ҿ��F H�����H��tH� H��tH��H��H��[]��fD  H��1�[]��    ��   �f�USH��H���  �Gt
H��p   uH��8  H��[]�D  H���   H�����F H�x���1Ҿb�F H���)��H��t�H� H��t�H��H��[]���AWAVAUATUH��SH��H��tH�    E1�1�1�E1��   A�   ��t
H��H;ws?D�E��A)�A��D��A��A��tFA��	�|   I�����~CH����t�H��H;wr�E1�L��H�؅�LE�H��[]L��A\A]A^A_û   �f�     E��uM��uE1��p���fD  O��Mc�I��O�B�V���@ E1�A��
�  A���y  A����   E1�M���u���H�N�,O�4)H����  M�I���q  I���  �%  M��M)�M��~DI���   IN�H��L)�H��~,L�� �F I)�M��I���  ~L���
   I��H�H��I��I��L�] ������D$    E1�E1�A�   ��tH��H;w�����D�E��A)�A��D��A��A��	��   I���  O��Mc�O�Z��t�� A�   �A�   ��tH��H;w�g���D�E��A)�A��D��A��A��	�����E��uM��uH����t���fD  I������I���O��Mc�I��O�B��D$   �"����L$��tVM�������I��E��������n���L��J�4���F H�H��H=�  ��   J�4���F L��I������L�u I������M�������E��� ���A��������I���I����w���M����   M)�I��
tiM��uI��N�� �F L��H��I�� �  A����LL��:���L��I�������L�u I���"���L�Ǿ
   �����I��L��L)�H��H�E �����L��H�I��A�	   I��L��J�4� �F H�H��H=�  �����L������I�������L��I��M�H�J�<� �F I���9���D  AUATUH��SH��H��L���  H���   A�}(��   �   �׷F ����H��H����   A�E$����   E1��8 ��  A;�H  sI��P  H�4�H��tH���!�����t`A��E9e$vSI��   D���<Bf���w��U(H����fD  H����F ����1ҾW�F H���c��H��tH�@H��uD  E1�H��D��[]A\A]��    H��H��H��[]A\A]��fD  AT1�USH���O �D$    ����   I��A��H������   H�G�V�1�H�4P� H���f9�B�H�HH9�u��˾   E1�H��L�L$1�L���-e��H��H�E�D$��u)D��H�EH�� �Pf�NH��H���u�] 1�D�e$H��[]A\�@ L�L$E1��   1Ҿ   L��1���d��H�E�D$��t���ff.�     ��? �   t9wt�9Wu�1���t�H����H�wH��H����������H���D  AWAVAUATUSH��X�D$L    ��tH��u�   H��X[]A\A]A^A_�D  L�wI�F� H�D$���   A9��  vƉ��T$(�W I��H��I��  L�G(�t$,�(H�L$ H��L�L$LH�|$�   H�D$�MH��H����c��I�E(�D$L���n�����A�] L�\$��  ��M��1�M��H�D$�D$(��L�L@I��M���LD  I�S�E���A9��  ����I�H(�t$(L�4�    J�1��uI�    H�EH9l$�$  H��H��u�I�@(�    ���     A���  9����������� I���  L�d$ �   1�L�T$L�<� I�?�   H�H�H�wH9�AH�H9�8H��I��A��I��?E��tH��u �   H��tM�$L9�L9�}H1�fD  J�41H��I��HcH��H��H��?H�� �  H���L9��w���L�T$�
���D  L9�t�L�D$8L�\$0PH��L)�H)�H�������L�D$8L�\$0Hc�I�H(� M�ŋD$,�|$(A�E��u!�D$(A�E A�E�D$L����L��H)�H)�뱋\$(A�UL�L$L�   H�|$M�EH��H��H���a��H��I�E�D$L���Z���H�t$ H���9�����    AWI��AVI��AUATUSH��H��HL�?H�0 H�$D�oM�g8�D$8    H�    ��  E��u�D$8H��H[]A\A]A^A_��     1�A�ML�L$8E1��   L��L�T$H�k(�a���T$8H�D$ �Ѕ�u�L�T$I�t- H�t$(M����  H�T$8L���A���T$8L�T$I�ǅ҉��{���H�D$ �KL�K8L�8����  H�D$ 1�1�A�   L�`�zfD  H9k(HFk(M���  H�T L�I�$H9�tAI�|$�L�L�T$H�L$H)�L�L$����I�$H�L$H��L�T$L�L$�  H��I�$�CI��I��L9�r:H�C0J�,�H��H9��w���M����  H�1I��I��L�I�D$��CL9�s�H�D$ �T$8I�M��tM�:H�<$��H���x���H�L$(H��k���f�H�T$�D$<    E���O����GA�mE1�1Ҿ   L�L$<H��L��D$�t_��D�D$<L�T$H��H�C0E��t>fD  L��L�T$蛆���D$<L�T$H�C0    ���D$8�����D�k�����D  �sL��Hs�!+��L�T$���D$<��   �D$L��L�T$H��H����,��L�T$���D$<ueI�G@�|$H�S0H�4(@����   @����   @����   H9�s�H��H��ɉ�H�z�H9�w�L��L�T$�.���|$<L�T$��tUH�s0����@ H��I�1I�$�,����     L�K8H�D$ E1��sL��������H�D$ I��[���f�     D�k�D$8    ����I��6���H9��o����H��H�����H���	���H�J�H9�w��H���1�H9��=����4H�4�H��H9�u��'���H9�������xH��H������	��x�	���H�z�H9�w����������  t@���  wH��`  H��t,H�@(����@ ��  1�;�H  sH��P  H���@ 1��D  H���  ��H��   �4p�f.�     AUATUSH��H���  H��tP��L  ����  tTH��I��I��H��tH��x  H��tBI�E M��tH���  H��tEI�$H��t
H��X  �E 1�H��[]A\A]�D  �   �鐉�H������H��x  �D  ��P  H�������H���  뤐AT1�USH��L���  �D$    M��tGI��$p  H��H��tBH�U H�H�UH�SH�UH�SH�UH�SH�U H�S H�U(H�S(H�U0H�S0H��[]A\�f�H���   H�T$�8   �<��H�ŋD$��u�A��$h  L���?���A��$l  L��H�E �+���A��$t  L��H�E����A��$x  L��H�E����A��$|  L��H�E�����H�E I��$�  H�E(A��$�  �E0I��$�  f�E2I��$�  f�E4�D$I��$p  �����f.�     AU1�ATUSH��L���  �D$    M��tI��$�  H��H��t�f�U H��[]A\A]�fD  H���   H�T$�   �r;��H�ËD$��u�1�A��$H  L��f��"���H��t}���F H��谐��H��tkL�h���F L��蚐��H��tUI9�tPH� $     �,@ �f���w0���f�fA�M �T
�f�I��L9�tA�U �JЀ�	vˀ� v1�f��I��$�  �D$�����    H��r���SH���  �P�F H��X  H���   H�x���H��tH��tH�H��t
H��[��@ 1�[�ff.�     �AWAVAUATUH��SH��H�wXH�?����H�} ����H����   I��H�E H�U(E1�H�u 1�L���  H�EPL�8M���  I�?A�UA��0  ��tv�X�H���RD  L��H��L��H�L$����H�L$H�}(L��H�$H�������L�$H��I�|H��E1�1�L��A�UH���tI��8  L�M H�HhI9�u�H�U(��H��1�[]A\A]A^A_�ff.�     @ AUATUSH��H�GPH�(H��tjH�?L���   H���  ����I��H��t-H�} �P��0  ��t��H�\� H�;H��A�T$H9�u�H��H��L��[]A\A]���f.�     H��[]A\A]�D  AWAVAUATUH��SH��H��(H�?�Gt'H��p  H�T$���   ����   �����H�} H�EXH������H�} �����I��H����   H�E H�U(E1�1�H�u L���  H�EPL�8M���  I�?A�UA��0  ��tw�X�H���SfD  L��H��L��H�L$�E���H�L$H�}(L��H�$H���-���L�$H��I�|H��E1�1�L��A�UH���tI��8  L�M H�HhI9�u�H�U(��H��(1�[]A\A]A^A_��    H�t$H���;���H��([]A\A]A^A_�ff.�     �AWAVAUATUH��SH��  H�?�D$    ����H����   I��H�E H�T$�  H���   L���  �/7��D�t$I��H�D$E��tH��  D��[]A\A]A^A_��     I��h  H�t$ ����H�E L��H�t$ H���   A�$A�ƉD$��u�A��0  ��tr�X�I��H���D  H��H���tVI��8  H�t$ �d���H�E I�H�t$ H���   A�$�D$��t�A���O���@ D�t$�����H�EX�8���D  H�EPH�L$H���f�UH��SH��H���H�t$��"��1҅�u%�;��t1��     �tH��H��H	�9��E H��H��[]�ff.�     @ AW�   AVAUATUSH��(�D$    H����   ���wH��9���   H�G0I��L�?H����   ��L�$�M����   �}���H��H�H�t��D  H��H9�tjH�H��t�I�WH�s H��H9��J  H��H)�M��tSL9�vNL)�H��H�H�C8H����   J�D �I��D$H��([]A\A]A^A_�f�     E1�I�WH�s H��H9�w�I�    �D$H�    H��([]A\A]A^A_� �wH�GH�L$H��wL����H�� ���D$��u�L�kH�;H�T$L���K���I�ċD$���d���M��H�L$�n����@ 9k�b���H�;H�T$L��H�L$������H�L$H��t�������     H�C L��I�t�����D$�������L��H��L���"�������H��H)�H9����������ff.�     �USH��H��(H�W8H��tfH�j8H��8H�L$H�T$������D$��uGH�D$H��H�T$H�p�3��H�ŋD$��uH�T$H��uD�D  H�{p t H��(H��[]�fD  1�H��(H��[]�@ H�{8H�t$�j ��H��(H��[]�H�t$H���#���H�T$�ff.�     �AWAVA��AUI��ATA��USH��H����H��H�n8H�G�    H�G(    H���L�|$)��H@1����H�H�3H������L��L��H�CE��tl�(���|$��u/A���C   E��um�D$H��[]A\A]A^A_�D  �D$   H�s0H���y��H�C0    �D$H��[]A\A]A^A_�f�     ��"���t$��u�D���C   E��t�L��L���("���L$��u��P���w��CA�v���SH��HSD�sL��H�H)�H�S ����D$���a���H�;L��H�s�����T$���F���H���5���H�p�H�s(E��t'H�S8L���4 ���D$������H��[]A\A]A^A_�L���1���D$��ff.�     UH��SH��H��H���   H�@hH��t$H�xH� H���H�$H�HcT$H�U H��[]ÐH���  H��8  �=���H��[]�fD  H��H���   H�@hH��t$H�H�x�T$H��H� H�$�PH����    H���  H��p   u�H��8  ������f�     AWAVAUATI��U��SH��H��h  L�w�T$(M���  A��L  ��  t;I��(  H��t/��t5A;�0  ��  A�   H��h  D��[]A\A]A^A_� �D$(A9E$v؉����   E�I���  H�D$H�@PHǃ8     H�$Hǃ@     M��tII�D$ I�t$XH��8  I�D$(H��@  �����H9�t"I�$H��p  H���    t@����   �� @  �F���E��0  E����  I���  �D$- H�D$@I���  H�D$HI���  H�D$PI���  H�D$XI���  H�D$ I���  H�D$��A��L��L��ǃ�       ��A����A��ǃ�   ltuo�����Ѓ��ǈL$.��A�ȃ���1  A��@�|$/h��B h��B H�D$��0  H��H��$�  �AZA[��   tƄ$	
  ��t$(H�L$`H�T$8%   L���D$��$�  �%���A�ǅ��2���H�$�T$(L��H��$p  �PA�ǅ�����H�L$1�H��$p  H��$�   �Q0H�$H�T$`H��$�   H�t$8�PA��<���  H�T$`H�t$8L���	���E�������I���   H�xh �.  Hǃ       Hǃ      H��$p  ��$  I���   H�@hH��t}H�L�BM��tqH�xH�L$`�t$(H�D$h    H��$�  H�T$`H��$�  H�T$pH��$�  H�T$x1�A��H�T$`H��$�  H�T$pH��$�  H�T$xH��$�  ���$  D�L$E����  H��$�  H��(  H�t$ H�S@H��$�	  H�SPH�T$@H�PH�T$HH�PH�T$PH�P H�T$XH�p0H�t$H�P(H�p8�@�����t$(I��8  ����A��0  ��9�r�B���I���8  M���  �D$- H�P@H�ppL�@hH�T$@H�PHH�t$ H�T$HH�PPH�T$PH�PXH�@xH�T$XH�D$M9�����H��8  L��L��L�D$�~���L�D$H��@  L��H��8  L���`����D$-H��@  ������    H��L���   ��L��H��$x  L���   R�T$8���   A��XZE���0�����$r  ǃ�       ǃ�   stibH��H�C0��$p  H��H�C8H��$t  H��H��H�C@H��$v  H��H��H�CH��$x  H��H�CPH��$z  H��H��H�CXH��$|  H��H��H�C`��$~  H����H�Ch��  ���   ���   I��p  1��T$(L��L�D$`H��$�   ��  �D$`H�CpA���   �}  fA��   �n  I��p  L�D$`�T$(L��H��$�   �   ��  �D$`H�Cx�R���f.�     �T$(�P�D$(���V����)����    H�$ƃ0   H��$�   H�T$`H�t$8�P�D$-A���D$. �#���fD  fA���   ��  I��p  1�E1��T$(f�|$8H�L$81�L��fD�D$`L�D$`��  �D$`H�T$8H�CPH�S@H�CpH��(  �@ A���   tfA��   ��  fA��h  ��/  A���  A���  )�H�H�ChH�Cx�   ǃ�   ltuoǃ�       M��tfA�|$�%   ��H�|$@   ���   L���   uH�|$X   �e  H�t$@L����	��HcCPHcT$@H��H�H�� �  HcT$XH��H�H�CPHcChH��H�H�� �  H��H�H�ChL�t$L�l$ L��L��L	�tL��L�����LkPLsh�|$- u�|$/ tj�|$. Hc�@  Hc�8  ��   H��$�   ��   HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$`L������H�D$`H�T$pH)�H�C@H�S0H�T$xH��H�SH�T$H+L$hH�K8����   H�KPH��H��?H�H��H)�H�CX����fD  ���   f���H����z�H���   H��H��H� HcH��H��I��I��?J�� �  H��Hc�H�P�HcP�H��I��I��?J�� �  H��Hc�H�P�H9�u�������    H��$�	  H�CPH�Cp�q��� �������H�shH�{0���������D  I��p  1�1�L�D$`f�L$8�T$(H�L$8L��f�t$`�   ��  H�D$8�D$   H�C`�D$`H�Ch�H����    H�D$HHD$P��������� I��h  H��������T$(H��I��p  H�D�H��   H�D$`H��  ����@ A���  A���  )�H�H�Ch����� fA��h  �tEA���  A���  )�H�H�Cx������     ���   ���   �����    A�������A���  A���  )�H�H�Cx���� H��tKH��t&��uH�GH9u(�3��� 1��)���f�     �������     �#   �f.�     �%   �f.�     AWAVAUATI��US��H��(H�GL���   ���   H�w% �  ��  �H	�����   H��t�   ���  t^A��$�   ti��tML��D�<L�t$L�l$@ I��$p  ��M��L��   L���H����  �D$H�E�A9�u�D  1�H��([]A\A]A^A_��    ���L��A��A�͉D$A����u"�� E��I�GxIDGp��H��H�E�;\$t�I��$�   D���L��������t�H��([]A\A]A^A_� H��t�   ���  �k���fA��$�   �q������Q���L��D�<L�t$L�l$I��$p  ��M��L��1�L���H����  �D$H�E�A9�u�1�����f�     UH��H��x  SH��H���8���H���  H���ij��H��8  H��Hǃ�      �Oj��H��H  H��Hǃ8      �5j��H��`  H��HǃH      �j��Hǃ`      H��[]�f�     H����  AVAUATUH��SH��p  L���   H��t�PH���  H���4  H���   L�c�v���H��x  �j���H�{8�a���H��8  �U�����0  ��tGE1��     J���8  H��tL�������I��D9�0  w�H��8  L���Oi��Hǃ8      H�Cǃ�       Hǃ       H��(  ǃ      L�h8L���i��H��   L��Hǃ(      ǃ0      ��h��H���  L��Hǃ       ǃ      Hǃ      �����H��h  L������H��@   tH�{H��@  ���ǃH      H��p  L��ƃ8   ǃ<      �hh��H��8  L��Hǃp      �Nh��H��@  L��Hǃ8      �4h��H��P  L��Hǃ@      �h��H��X  L��HǃP      � h��H���  HǃX      H��t#H���  ��H���  L����g��Hǃ�      H���  L���g��H���  L��Hǃ�      �g��Hǅ�      H���  H��tH���PXHǅ�      []A\A]A^�@ ��    �>tkH��I������H��M��u/����H���  H��H��  �H��H�� ���HN�H��� H��H��?H��H1�H)�J;͠�F J�� �F � 1��	���f�     H��H��  �����HO��ff.�     AT��   USH�_ H�S H9W(r}H�31�L�g8H���8���H������H�s1�H��I��$�   ����H���½��H�s1�H��I��$�   �����H��褽��H�s1�H��I��$�   �����H��膽��I��$�   1�[]A\��    �<t1<�t�p����F�V����	��V	Ѓ���H����    H��1�1������H��H���f�AWH��AVAUI��ATUSH��H�wH�$H�W H�GH�W(H�wH9���   I��I���] =�   tyA9���  H�JI�M(L�"���K  ����  ���0  I�T$I��=�   LF�L9$$�|   I�U(M�u A�$H��E�E0L)�H����@�ǃ�@��@��u�A9��o  L�"���  AE4�   � �F =   u��   �9Ct+�S H�� ��u�I��M�u(L9$$w�1�H��[]A\A]A^A_ÐI�E8D�CJ�, ����   ����  ��w~�$ՠ�F �    I�6�   L�������S��tM����  ����  H�E �I���;�����M�u �n���f.�     I�61�L��������S��u�f�E ��@ L���S��t��A����I�m8���\  I�6L��������t���@ I�T$H9$�9  A�D$I�Ԁ������I���o����    9K�SFK����K����A�E1�I�D�H�D$�#f�     <tLL�} �CH�L9t$����I��I�v�L���6���I��C<t<u�D�} �ɐfD�} ��f�     D�} �I�������H�<$I�D$H9��M���A�D$I�L$������tv��<toI�D$H�w�-�     �P�I�ĉ������������H�����s���H9�u�1�������    �E �P����E �H���H���   []A\A]A^A_�I���4���ff.�     �AWAVAUATU1�SH��XH���    H�_H��(  Ɔ!   t
H���    uH��X��[]A\A]A^A_�f�     I��L��H  I��1�H��P  L��HǆH      H���H)����  ���H�H��  Hǆ�     Hǆ�     D��4  ǆ�  ����Hǆ�  \  Hǆ�   �' ��P  L��X  A�}0 ��   I�U A�a   �a   A�    I��H�t$1��   H��L�2E1�H�T$�H�1�D�L$<L��L�L$�   L��L�T$@D�|$H��9���T$H�D$(����   �l$8H�D$0I��$�   H��Iu�����Ņ�uI��$�   H������Ņ���   H�t$(I��$`  AǄ$p      I��$h  H�D$H�8�`���w����A���  I�U A� P  D�XL������ H��L���`���D$H�D$(    ���X���1�1��f.�     H�SHH�s@H�|$�~���H�߉��t�����X���I��$�  A��$H  �H��xVuIǄ$�  �h�:I��$�  �  vIǄ$�     I��$�  �  H�t$(����IǄ$�     �����fD  H��I��$�  � SH�_8H��t6H���  H��t*��!   ��   uH�G H�0�p������  1�[�fD  �   [�f�     SH�_8H��tH�G H�0�:���1�ǃ@    [�@ �   [ÐAT��   USH�o H�UH9W(rBH�u L�g8H�������H�uH��A��$�   �����H�uH��A��$�   �����I��$�   1�[]A\�f�H�W ��   H�J(H9O(s�@ USH��H��H�2H�o8����H�P�H���   H��w'H�S(H+S f��4  1�H����f��6  f�K@f�SBH��[]� AT��   USH�o H�UH9W(s	[]A\�@ H�u H��L�g8� ���H��x+I��$�   H�uH������H��xI��$�   1�[]A\� [�   ]A\�fD  H�G8H���  AWAVAUATUSH��(L���  M���  M��X  ���  I��I��   E��P  H��L���D��������tL��D���H�����������  I�E(L��H�p��[���H��A9E0��  I��(  E��@  �D$    I�u H�xI�E(D��H�X���   H)�H��A9��P  A��p  D�\� A��t  D�9��i  D)�A��p  �+�D$���	  A��D  A��I��H  L��J�4�H�h��������A��@  vND��   )��L$f�     I�u L��H���$D�pH�4��u����E��$�L$�D���4A;�@  r�I��h  I�u ��J��H�pI��h  � �I��h  H�pI��h  ����@�0I��h  H�pI��h  ����@�0I��h  H�pI��h  �0I��h  H�pI��h  �I�u 9\$������D$H��I�E(�D$AƇ!  H��([]A\A]A^A_��     �   H��([]A\A]A^A_�@ M��`  M��h  A�L�L$�   D�\$M��L�$�+4��H��I��`  �D$��u�A��p  D�\$I�u E�t  H��H�I��h  D�M���(���I9�����M�E(H��L)�I9�����L�$H��fD  H�:I9�wI9�vH�H�:H��L9�r�������    �   �f�AW��   AVAUATUSH��hL�w I�V0H9W(�k  L�o8H��E1�H�       �I��������A�E`�    H=�� ��  H=?B ��  H=�� ��  H=�����  H= ʚ;��� �'  ��HL�D����A����	H��H�H��H=�  kMc�N�D<0莲��J�<H��tJ�D<0H9�HL�I9�LO�I��I��0tXK�4>�>��   H���C���H��H=�  �D���J�D<0    H���D  ��Hc�H�4� �F J�L<0�����fD  H�C	H��	wH��L)�H��	vjI�E@   I�EP    I�EH    I�EX   I�Ep    I�Ex    I�Eh   1�H��h[]A\A]A^A_ÐH�D$01�H��J�8�M����
����     H��������1�I�      �I�       ��+fD  I��I)�I9���   H�H�H��H�H��H��0tKH�H��t�H��H+T0H�4� �F H��H��H��y�N�I9���   H)�H�H��H�H��H��0u�@ H�$H��I�}@I�E@H�D$I�EPH�D$I�EHH�D$I�EXH�D$ I�EpH�D$(I�ExH�� �F I�Eh�[���������������fD  H��H�H��H��:����    L��H�H��H��"����    �
   �   �7���f�     �
   A�   �   ���� �d   A�   �   �x��� ��  A�   �   �`���ff.�     ATI��� �F UH��S�\���H��H��tH��[]A\�@ M��t�I�|$H��t徝�F �����H��t�H�[H��H��]A\H�R@���    AUI��ATA��UH��S��H��H���  �(t>H��`   t]H��   �4X1��"���H��tD��H��L���W��H����[]A\A]�f�H���   ���F H�x�K���1ҾW�F H�������H��uH���   ��[]A\A]�D  H� H��t�H��D��L���H��[]A\A]���AWAVI��AUATI�̹   UH��SA�� ������H��   ��H��$�   �T$Hҁ�  L�D$L�D$@H���  H��`��L��H�D$(    E�E1�H�D$H��$�   A��  A��`H�01�L�.H�t$8�   �H�H��D�L$l1�L�L$0L��L�t$p�l.���L$0H�D$X���  D�|$hH�D$`I�~L��1�Iǆ@      H���H)���H  �����H�I�F(  ��H���  ��  I�I�FI�FI���   ��U%�  I�F0  2 ��0A�F<   I�F@   I�FX   Iǆ  "  Aǆ�   ��  Aǆ0  ��  A��@  ����   L�l$(�t$H�L$0H��L���]���A�ǅ��T  �E����   H�}8 ��  E��uA���   ��  ��   H�t$X�+�    H��L���T��D�|$0H�D$X    E�������1�H�D$8H�8�gT��H�Ĉ   D��[]A\A]A^A_�f�H�u L������A�ǅ�u�L�l$(H�u(L��L������A�ǅ��x���H�U(H�T$0H�t$(H�|$8H��3���A�ǋE���.���L��L���j����)���D  H��$�   1�1�L���\���A�ǅ�������t_H��$�   H���   �@t�����   A���  ����   H�l$L��$�   fD  ���U(I���   �Bt��x�A���  ����   I���  H�������H�t$I��   L��H������A�ǅ������1�I��x  ��L�����   H���N���A�ǅ��]���I���  1�1�H������A���B����     H�} L���T��������    I���  A���  �W���H��$�   H���   �E`A���  ��t�L�l$ ��A�U(�E`��x�����H�T$0�_���@ AWAVA��AUI��ATUSH��H��8  H���   ���F �L$H�hL�D$H���5���H���L  I���   �   �׷F I���C����P�F H��H�D$������F H��H�D$ �����H���  I���  �   ���F I���   �����1�H��H�D$(�z���A�ǉ�$�   ����   L�D$�L$D��L��H��A�T$A�ǉ�$�   ����   I��  OTTO��   E����   1�H�ھdaehL��A��@  ��$�   ����  H��L��A�T$@A�ǉ�$�   ��uO�D$1�H�ھ2FFCL��A��@  A�ǉ�$�   ����  Aƅ�  A�   �D$s�^f�     A�   H��8  D��[]A\A]A^A_�D  A�   ���     1�H���f���A�ǉ�$�   ��u��D$s E1��D$I���   H��$�   ��  H��H�D$��	��D��$�   I��E��u�I�{L��I���  E1�H���H�C8H)����  H�D$0L����I�    Iǃ�      L�\$8�H��   H��$�   �H�H���k���L�\$8H�L$0H�߾��F H�D$@I�+L��I�[I�KE�c0I�C�i��L�\$8����$�   �  E���t  A�{(��
  A�{*��
  H��$�   H��L�\$8H��H�D$H�Y���L�\$8��A�C,��$�   ����  A�s*H��Ht$@L�\$8����L�\$8����$�   �
  I��x  E1�I���  Iǃx      H���H��L��Iǃ�      H)�L�\$8��@���H�H���Y���L�\$8H��A�K,I���  I���  �������L�\$8����$�   �  I���   �   �   H��H��H��$�   �����L�\$8����$�   ��  A�CL��$�   �|$ A��H  �f  A�ΉL$8�L$tE��~9��|  A�C E���<  A��AUI��h  H��AS�L�|$PH��% �����$�   D�� 0  M��L�\$H��������$�   AZA[L�\$8�2  I��(  H��L�����L�\$8����$�   �  A��I��8  1�H�މ�$�   �����L�\$8����$�   ��  A��L  ��  u	E����  I���  H�K8Ǆ$�      H�D$X    H�L$8H���  Ǆ$�       H�t$XH�|$8L�\$P�-M����$�    L�\$P��  Ǆ$�       H�t$@H��L�\$8I��  ����L�\$8����$�   �/  L��$�   ��$�   1�H��L������L�\$8����$�   ��  ��$  =   ��  A��0  L�L$H1҉�H�|$0E1���  �.%����$�    L�\$8��  ��$  1��I���8  H��H�  9�w�A��D�d$0I��L��E�D�t$81�A�� ���A�� @  E���>H���8  AUE���SL�D$PL��L��H��������$�   AXAY����  ��$  9�w�I��L��D�d$0D�t$8E��t	����   H�t$@H��L�\$0I��  A��L  �]���L�\$0����$�   ��   H��$�   H���������$�    L�\$0��   A��8  AǃP      ���V  <�>  H��$�   H��L�\$0������$�    L�\$0u?�����  �@��A��H  A��H  I��@  H��L�\$0�����L�\$0��$�   ��$�   ��$�   L��L�\$0膷����$�    L�\$0�4  H��$�   L�\$0�a���D��$�   D��$�   E�������A��L�\$0�D$8�  fD  L�D$�L$D��L��H��A�T$A�ǉ�$�   ���m����D$ ����D  H��$�   H��L�\$8H��H�D$H�{�����$�   L�\$8���g  A�{(��  A�S*<��  ����  H�D$@H��L�\$8H�4����L�\$8����$�   ��  I�{81�1�H��L�\$8�����L�\$8����$�   �~  A�CL��v
I9C`��  I��x  1�1�H��H��L�\$8����L�\$8����$�   ��   1ɺ   H��H��$�   �z���L�\$8����$�   ��   I���   1ɺ   H��H��H��$�   �E���L�\$8����$�   uUI��`  I��X  I��P  H��$�   ����L�\$8����$�   u#A�CLA;��  �:���Ǆ$�      �    H��$�   L�\$0�N�����$�   ��$�   ����  A��E��L�\$0�D$8��  H�D$ H�L$A��L  ��  I��X  H�D$(I��`  I��h  HcD$8I�EA�C$I�E u	H���7���A�EtXI���  A��H��tHE��tCL�\$I���  D��L���P8A�ǉ�$�   �������H��L�\$tL���S8L�\$�    A���   u�|$ ��  uA���   I���  I���  I���  H����  H��H��?H1�H)�H��   ��  I���  H��I���  I���  A��0  ���Q  ��L�l$I��0  M���8  M��M���   �    A���   taI���  A�   H��vI�T$hH��v
H9�HF�I��I�t$@L��H��辣��I�|$pL��H���N���I���  I�|$hL���:���I�D$hM�t$XM����   L��H��?I1�I)�I��   ��   I�D$xH��I��I�|$pI�D$xL9��l  M�e A�|$` �<���I���  I���  I�D$@I���  I�D$HI���  I�D$PI���  I�D$XI���  I�T$xI�D$pI���  I�D$h�N��� I�D$PM�t$PH��?I1�I)��M����    I�|$hL���3���I�|$@L��I�D$h�!���I�|$PL��I�D$@����I�|$HL��I�D$P�����I�|$XL��I�D$H����I�|$pL��I�D$X�ٝ��I�|$xL��I�D$p�ǝ�������f�<��n���1�H�ھ FFCL��A��@  A�ǉ�$�   ���H����D$sE1������|$ �j���f.�     Ǆ$�      �P���L�l$M���|$ A��L  �  A�C I�E ����  �H  A��0  ��I�E I���  �����I���  H��I�EhI��   H��D��I�upH��  H��I�ExI��  H����  I���  fA���   H��fA���   ���@I���   ��fA���   ������)�A��x  D)�����9�I���  L�H��fA���   I���  fA���   H��fA���   ���u  I�E(L��$�   H����  A��t  L��L�\$����I�u(L�\$H��tCH��t>���t7�8��z  �� �d  ��-�[  �� ��  ��-��  ����  H�|$L����F L�\$��C��L�\$I�E0�|$s����  A���   t��H�I	EA��|  1�L��I���   L�\$���6���L�\$H��t1� �F �   H����� ��tRH�ƿ��F �   ��� ��t:I�E0H��t4� �F �   H����� ��tH�ƿ��F �   ��� ��u��A��L  Hc�I�]����  ��  A�]HI�M   ����   I�EPH��z  ��   f�z ��   H��1��(f�     H��y  ��   H��f�y ��   ��9�rځ���  t�|$ u[1�1��@�F L�\$H��$�   L��$�   H�cinu  H��$�   ����L�\$��t*�Ё��   t��t��$�   fD  D��$�   ����I���    Ǆ$�       uA9]HtI�EPH��I���   f�     A��  ��t�I��   �   L��$�   f��$�   H����  Ǆ$�   BODA1�f��$�   1�H��$�   1����F �%��A���#���H��$�   L�\$諭����$�   L�\$����$�   �  A��������     ����  �  A�]H���H������� I���  I���  H��?H1�H)����� I���  H��L�\$�ܘ��L�\$H��I���  I���  �����L�\$H��I���  I���  覘��L�\$H��I���  I���  苘��L�\$H��I���  I���  �p���L�\$H��I���  I���  �U���L�\$H��I���  I���  �:���L�\$�e���A�C I�E �����I�M   ���  �����H����  Ǆ$�   CBDA�   f��$�   �_���A��L  ����L��L�\$葺��L�\$H���p���L��$�   H�|$H��L�\$L����?��L�\$I�E(�Q����PH���w����PH��H���f����t$8L��L�\$�y���L�\$H��I��I�E(��   L��H���1����׃������A�x+������   �\$M�HD)�L��L��A���D  ��tH�����A<�v��t4E1���E��t*�W�Lʃ�t�AH���A�H9�u�����~A�x+t�I�}( �x���A���  L��L�\$�b���L�\$H�������H�|$L��H���>��L�\$I�E(����Ǆ$�   EBDA�   f��$�   �����H���<���H�|$H��L��L�\$�k>��I�](I��H���|M��L��I���qM��L�\$A9�Hc���   ��~B�P�A�N�Hc�Hc��A8<uw��Ic�L�H��H�1�H���D�D�H��D:D�uQH9�u�D��)��ȃ�t@Hc���r�@��?w+H�(     �H��s��H��H�Hcȅ�~��� ��?v�D M�e0����H��H��r�����>����D$t    �����D$��������$�   �*���H��$�   L�\$0Ǆ$�      �m���D��$�   L�\$0E��D��$�   �-�������Aǃ0      I��(   ��   Ǆ$�      ����H�t$8I���  �`�����$�   L�\$P����$�   ������!���H�L$@H��L�\$PH�4�����L�\$P����$�   ��  �   H��L�\$P����L�\$P����$�   ��  H��L��$�   �@���L��H��H�D$h������$�    L�\$P��  f����
  Ǆ$�      �R���A��L  1�1�L�\$0H��$�   I��@  A�C$苲��L�\$0����$�   �����E���<  E�c$E���/  A��L  I��  H�L$PH�K8�D$XI��  H�L$0Ǆ$�       H����  I��  ����  ����  A���   ��  D��H�|$0E1�1�L��$�   H��   L�\$8�h��L�\$8��$�    I��   ��  H� �F ���  @����  ��t�� �@����  �|$X��  t*�|$ t#H�T$0H�|$PD��L�\$8�T���L�\$8��$�   ��$�    �  Ǆ$�       A��L  ��  t"�t$tL��L�\$0聿��L�\$0I��8  �=���1�I��    I��   E�c$Ǆ$�       �=  fAǄ    fAǄ    H��H=   u�H����  I��  �E  I��  H�� � �F H���H)�I��  H�� H)�   ��I��  ���H�H�S8H�|$PD��L�\$0Aǃ      �A���L�\$0����$�   ��   �   �5A;�0  w<I��(  �Qf��t,fA��C
  A��  H��H=  tzA��C
  H�ʅ�u�fAǄC
    fAǄC
    �̋3
 �����F �T(��4��������F f�T(��!���Ǆ$�      ��$�   ��$�   ����M��L�l$0��$�   ��$�   ���?�������H�� I��  � �F H���H)�I��  H�| ��   H)�I��  ���H�����H�t$@H��L�\$0H�I��   ����L�\$0����$�   �W���L��$�   H��L���&���L�\$0��A���   ��$�    �'���L��H���������$�    L�\$0�	���A���   �����  �������Aǃ      �D$8   �D$@    L�l$0M��;l$@��   L��H��������$�    �ЉT$H��   L��H���w�����$�    ��ur��A;�  �T$HvA��  �t$8H��H��<�:A9�v+���   w#��M��   H�L�f��  E�0fD��  ����H��9�rD$@�|$8�L���M��L�l$0�	���M��L�l$0A��     vAǃ     A���   ������L��H��L�\$0������$�    L�\$0���D$@������D$8    L�l$0M�݋L$89L$@�����L��H���j�����$�    ���a���L��H���������$�    �H���H�1�I�T- f��  �I��   H�qf;O��   H��A9�w��   �U��H��L�\$0A��  �A���L�\$0����$�   �����H�s@1��   �2H�HA9�v#�I��   H�L�f��  �<Of��  ��H��9�s�H��L�\$0�]���L�\$0����f��  �D$8�����A���   ��  D��H�|$0E1�1�L��$�   H��   L�\$8���L�\$8��$�    I��   ��  H���y  @���V  ���:����� �@���'���������F f�T(�����H�L$@H��L�\$8H�4I��  �#���L�\$8����$�   �;  L��$�   H��L������L�\$8��A��  ��$�    �  H�|$0E1�1�D��M���   ���L�\$8��$�    I��   ��   f�   A��  ����  ���y  D�t$H�   L�l$8A��L��E9���  L��H��������$�    A��uw��  L��H��tV�������$�    ��uV�ƺ��  A��H)�H9�~D������H��   1�D��A�<A����f�<VE9�v�9�v��z���������$�    ��t�L�l$8D�t$HI��L�|$0I��   L�\$8L����2��L�\$8L��I��(  L�\$0Iǃ       ��2��L�\$0Aǃ      ��$�   Iǃ(      Iǃ      Iǃ       ��$�   ��������l���H� H�xH���H���H���F H�L�H)�H��H)�����H������Ǆ$�      �1���A��Ww�D��H�|$0E1�1�L��$�   H��   L�\$8��
��L�\$8��$�    I��   �����H� �F H�ǉ���~���I��L�l$8D�t$H�l���A��$���H��L�\$8��q���L�\$8����$�   �����D�t$81�M��I��L���L��L�|- L�   ����fA�H��A9�w�H�\$HL��M��D�t$8H������L�\$H������r ������F �T(������H�X H�x���F H���H���H����F H�L�H)�H��H)�����H�����I��D�t$8L��D�d$0����L��H��L�\$P������$�    L�\$PH�D$x��  L��H������L�\$P��A���  ��$�    �r  H�|$8E1�1���M���   �4	����$�    L�\$PH�D$X�+���L�l$P1�I��D�t$`E��M���*H�\$X��L��L��H���������$�    H��  ��A;�$�  r̋D$hH�t$xL��L��$�   H��E��L�l$PD�t$`H�H��$�   ����L��$�   ����$�   �����L��H��L�\$P����L�\$P��$�    fA���  �j���L��H������L�\$P��A���  ��$�    �B���H�|$8E1�1���M���   ���L�\$P��$�    I���  �����D$x    D�d$PL�l$`D�t$hM�ދD$xA;��  �R  �D$xH�|$8E1�M��I���  A���  �   L�,�1������$�    I�E ��   E1��   L��Ik�H��Im ������$�    f��$�   ��   L��H��������$�    f��$�   ��   L��H��I���c�����$�    ��   H��$�   H��H��H��H�EH�U H��$�   H��H�UA���  D9��Z����D$x�����H�D$X    �����M��L��E��L�l$PD�t$`�����Ǆ$�      ����A��H  �����M��D�d$PL�l$`D�t$h����M��H�|$8E1�1�A���  M���   D�d$PL�l$`D�t$hL�\$P�L��L�\$P��$�    I���  �A����D$`    D�d$PM�܋D$`A;�$�  ��   I��$�  �l$`H��H��$�   H�D$hH�D$XH4��������$�   ����   �   H���*�����$�   ����   L��H��H��Hl$h������ЉU ��$�    ��   H�|$8E1�1���M���   �y����$�    H�Eu|1�D�t$hM��M��I�܉�;] sML��L���y���H�M��������$�    u����M��D�d$P�$���M��L��M��D�d$PD�t$h����L��D$`M��M��D�t$h�����M��D�d$P������Hc��   ��x=;�8  }5H��SH��1�H��H��H�@  H���RPH���   H���   [�fD  ��    �ff.�     @ H��(  H�@@    �H��  �  H�T$�H�|$�H�G@H��    H�GHH�  H�GPH�D$�1�3G�G8   ����
�G<��H�GX	  ��1�1�x��[DG`1��D  �؉G`1���     �ff.�     @ H��  H��t1Ҁ8/��H���     H��8  H�H��@  H�FH��H  H�FH��P  H�FH��X  H�F H��`  H�F(H��h  H�F01�Ð��P  f�1�� H��t
H��   H�H��t
H��(  H�H��t��0  �1��f�H��t�1��D  H��t�21��fD  USH��H�GH��`  H��t.H���   H���P�F H�x�´��H��tH���UH��(  H�B@H��1�[]� AWAVAUATUH��SH���	  L��t$I���   M��p  �D$4    H�$I��   H�D$I���   L�phM����  I�I�~H��$   ��D$4����  A��(  H��$   @���5  �V�1���H�L�     H���P�H��H	�H9�u싔$  E1�H�D$    ���  I�I�~H��$   �P�T$4����  H��H��I�X  �H�@Hǅ�
      Hǅ�
      H���
  H��H�����
  H��I�@  H��  H��0  H���
  H��  H���
  H��  H���
  H��   H���
  H��(  H���
  �SH���
  �    �҉��
  I�Hc�H;L$�$  ��x'�D$ H�D$��  L��H�L$(H�t$�P H�L$(�D$ D���   I�t H�t$ E���&  �T$H��E1�)�H�D$H�@�P�D$4M����   ����   I�H�x ��   H�}@�*��H�}PHǄ$      H��H��$   �	��H�}XH��H��$  ��~��I�~1ҋt$H��H��$   H��$  I��P�D$4H��$   H��H�E@H��$  H��H�EPH��$  H��H�EX�f.�     �D$4	   E1�H�<$L���)'��H�ED��1  �D$4H���	  []A\A]A^A_��     E1��� H�D$H�L$(�   H��H��$   �P0L��L�|$H�D$8H��H��A�W8H�D$8H�\$H�L$(H��$ 	  I�GH��$   H)�H�t$ H���P�D$4<������H�EH��H�t$ H��$   A�   ƀ0   H�D$H�@�P�D$4�O����1������f�     )�H�<$Hc�H�T$4H��H�D$�����L$4I�Ņ������H�T$Ic�(  H��H�$   �J4������D  �D$A��,  L��L�D$A�(  I��   ��I�H  H��}���L�D$���D$4��  �4L��L�D$�L����D$4���k  L�D$Ic�(  I�P@@���]  �F�1���H�Df.�     H���J�H��H	�H9�u�A��,  ����   �z�1�@��H��L�8@ H���P�H��H	�L9�u�H�E1�H�48f.�     H���P�I��I	�H9�u�L��H�L$ L�D$�
���Ic�8  H9���   L�D$M9`��   H�L$ I9���   I)�L�D$(H�L$ tyH�<$L��H�T$4L�d$E1������I�ŋD$4���A���H�L$ I��H  L��L�D$(H�H�L$L��������D$4���#�������L���i���Ic�8  H9�w�D$4	   E1�E1������H��1������AWA�   AVAUATUSH��(  L�gA;T$ ��  I��$   A��H����I��H�V H�D$H�F(����  ��H��@  Ǉ�       H��8  ���ʉ�H����0  E1���E1�L��ǃ�   ltuo�ƃ�����1  @�t$%H�D$L��L�x��h��B ����PQH��H��$�   A�H�� A�ǅ���  ��D��H�|$h%   �D$��$�   ����A�ǅ��a  ��0  H�L$H�|$hL��$H  �D$��1  �D$H��$   H�D$(H��$(  H�D$0H��$0  H�D$8H��$8  H�D$@H��$@  H�D$H�A�P���   �������   �D$���c  H��$�   �y��H��$�   H��H�CP�y��H��H�CpH��(  �@ I��$�  I+�$x  ǃ�   ltuoH��fA�}H�ChH�Cxw
���      H�|$(   L���   uH�|$@   ��  H�t$(L���л��HcCPHcT$(H��H�H�� �  HcShH��H�H�CPHcD$@H��H�H�� �  H��H�H�ChL�l$L��L	�tL��L��L��蓹��LkPLsh�|$ u�|$ ��   �|$ Hc�@  Hc�8  ��  H��$�   �Pf��~cD�B�H�@I��I��I�@ HcH��H��I��I��?J��
 �  H��Hc�H�P�HcP�H��I��I��?J��
 �  H��Hc�H�P�L9�u�HcCPH��H��H��?H�� �  H��H�H�CPHcChH��H��H��?H�� �  H��H�H�ChH�t$HL���}���H�T$HH�D$XH)�H�S@H�C0H�D$`H��H+t$P��H�CHH�s8��   H��(  D��[]A\A]A^A_�D  H��8  ��1�1�H��@  Ǉ�       �|���@ H��$�   H��(  �Tw��H��$�   H��H�C@�?w��H��H�CPH�D$(L�u8H�EH�D$0H�EH�D$8H�E H�D$@�EH�E(H�D$H�E0�S���D  H�D$H�|$hH�@�P�8���f�H��$�    ������,���@ H�shH�{0��������fD  H�D$0HD$8������^���ff.�     H����  AUATUSH��H��H��X  L���   H��tw��8  ��~ZE1�f.�     L��H��H�H�EH��t-H�0L������H�uL��H�    ����H�E    H��X  I��D9�8  �L�����HǃX      H��8  L�����H��@  L��Hǃ8      �w��H��H  L��Hǃ@      �]��H��P  L��HǃH      �C��H��X  L��HǃP      �)��H��@  L��HǃX      ���H��  L��Hǃ@      ǃ8      ����H��   L��Hǃ      ����H��(  L��Hǃ       ���H�C(    H��h  L��Hǃ(      H�C0    ���H��p  L��Hǃh      �s��Hǃp      H��[]A\A]�D  ��    AVAUATUSH��0Hc��   ���P  ;�8  �D  H��I��L��@  H��   �   H���Uh���  H�D$H���  H�I��I1�I)�I��   ��   L����  �=u��H�<$L��fA��$�   �(u��H�|$L��H�$�u��H�|$L��H�D$�u��H�|$ L��H�D$��t��H�|$(L��H�D$ ��t��H�D$(H�D$H��?H%  ��H   H�D$H��H��H�$H��L�H��  H�T$H��  H��   H��  H�T$H��  �-z�����5   H�D$ H��H��(  H�D$(H��H��0  H��0[]A\A]A^��     �E   ���    AUATI��USH��H���   H��L���   �D$    �VHH��x1I�UH��H���(\���(H��H��H��H��H9�HB�I��$@   tH��[]A\A]�fD  1�L�L$E1�H�پP  H��������T$I��$@  ��u�A��$8  ��~��K�H�PH�4�H��H��H��T  �    �Bt   H��P  ǂ(���   ǂ����   Hǂl���\  Hǂ��� �' H9�u��U���fD  ���F 醅��fD  SH���   �P�F H��`  H�x����H��tH��tH�H��t	H��[�� 1�[�@ SH��H�?����H�;����H��tH�{PH�S(E1�1�H�s H�?�P1�[�ff.�     �SH��H��H�?�p���I��1�M��t9H�H�JH���   H��H�4�H��H�@  H�T$A���uH�SPH�L$H�
H��[��    H�GPH�8 t.SH��H�?�
���H��t
H�SPH�:�PH�CPH�     [�fD  ��    AWAVAUI��ATUSH��H��8  H��    H�   �T$8�h  I��`   ��  1�H�������A����tH��8  D��[]A\A]A^A_�@ L�t$P1��   I��   L��I���   I���   HǄ$      �H�L��H��H�t$1�H�B1��H��H��$�   �0����   H��H�D$�^�������  H�u@���F �   �H���� ���&  �����D$L   H��$�    tH��$�   I���   �ھ��L����$�   D�D$LE�������D$8������f���  I��0  A�EH    I�E    I�E I�EH��H��  A��h   I�Ut
H  I�EI��P  I�E0�F I�U(H����  I��H  H��t<����t4�
8���  < ��  <-��  �� t	��-�C  H����u� I��`   I�E    tI�E   I��X  H��tB� �F �   H����� ����  H�ƿ��F �   ��� ����  f�     I��p  I��x  A�E8    I�E@    H��H��I�EhI���  I�upH��  H��I�ExI���  H����  A���   H��I���   f���c  �@�������������������D��fA���   )�D)�fA���   9�A��j  N�A���   fA���   �/���苾��L�l$ H��A�	  L��$   谻��H�$    L��I��L�}H��薻��L��H��I)�I9�LG�L����������  O�L<�H��$   C�< I9��;  D��$   �D�@A��s��  H��I9��  A��Su޿��F �	   H����� ��u�H��$   H)�I�D
H�$L�<$H�t$H��L��H)��:������  I���   H��H���P�������  L��$�   H��$�   L��L��$�   L�L�D$XL�D$PL�D$H�\$`Ǆ$  ������$�   L����$�   L��H�\$P��$�   L����$�   L�d$`L�|$PL�D$M�l$�M9��L  �D$h���h  I��	�Df�A�s�e  L����$�   L����$�   H�T$PL9��  �D$hI��L�����!  I��A�?Su�M9�w����F �	   L����� ��u���F �   L��L�l$ ��� ����  �D$L    L��$�   H��$�   �D$h    L�H�C�H�\$`H�$f.�     L�d$PL����$�   H�l$PH9���  H�$H��I9�r�eD  I��I9�sGA�<$%u��F �   L����� ��u�E��8  E��~�I����$  I9�r�f.�     H9���  �    E��8  E���   �D$hD�T$8�D$LE��������������H�|$H�T$L�P   ����D�L$LI��p  E�������H��$   I���   H��$�   H���I  H�BH)�H9�vH��$   H��H�|$H�T$L�3���D�D$LH��I��h  E���B���I���   H��$�   L��$   H���\������t  I�L9���  A�   H��$   L�,$H��E���AfD  �N�1�E���*  ��H��M �   D)�A��@���[  H��H��L9��K  H9��  �
�΃�0��	v��N����K  �N�����  �N�1���     ��F �   H����� ������H��$   H)�I�DH�$�)���f.�     L<$I����  J��<  �	   H��$   I��   ����   H�$	   L��$)  �5����    I�M�6���fD  ��F �   L����� ������L�l$ �   f.�     �D$L�����    �FH��H���?����    �FH���+��� H���   ��F H�x�ӛ��H����  I��`   I��   �s���D  I���   �P�F H�x蛛��I��`  �M����    I���   H�������H�4$H���-���������D  L�l$ �D$L�����f���  ��  fA���   ��  ����@ I��  H�������I�E(�����    A�   �����D  H�E�I9��,��� L����$�   L�d$PL9��h����D$h���t  �} /�����H�EH9������H�EL��H)B��T$����������u�R�A���F ���F H�|$H�z�C   H�\$ H��L�d$0A��L�l$(M��I���@ I��0I�] H����   �A8�u�H������H9D$u؃|$t-�E8Cuȸ   �f�     �TH��:T�u�I9�u�M��H�\$ L�l$(A�W����  A�O����  �Q  ����  I��p  ���G  ��	E1�1�H��$   ��L��L��H��$   �\  ��$�   �D$h���\���L�d$P�r���f�H�\$ L�d$0L�l$(�\���@ A��8  ���)���f�     �D$L   ���� M H�}�����@ H��舳��H�SI��H)���  H��   �   H��$   H��HG���������  H���H���H��$   L)�H��H�����f�1��V���f�     H�2H�0H�rH�pH�rH�pH�rH�pH�r H�p H�r(H�p(H�r0H�p0H�r8H�p8H�r@H�p@H�RHH�PHI��H  E��(  E������E��,  E�������A�������A�������M��p  E��8  I�I+�H  E����  A�A�I��@  H�4�H��H�JxH��L���  �[���   u��������������H���   H9��w������o�����t��H��H)�1�H��H9��U���H��P  L9��^  �9�  v�   �y�  v�A   Hc��   ���x������� �������I�u0�����    A�   �����D  @�� v'@��>��   L�,$��   �����L�l$ �   �����H�6     H��s�H������L�,$I��h  I��p  �D$L    H��$   �+���IǅH      �P���1��
   H�����H���S���H��$   �D$L    �L���I��  �������Hc�$  ����  A;�8  �y  Hi�P  I�@  �����   1��������$�   ����I��   H9������H)�C�1�H��Hc�H��I9�0  �����I���   Ic�E1�1�I��   L��$   �   H�<$H�D$0�w�����$    H�D$I��X  ��  H�D$    1��D$    I�܋D$A9�8  ��  Li\$P  I��@  Lۋ�8  ���=  �C�L$�D$<�E�D$ 9�vL�E���9���  �T$H�<$M����L��$   �   �D$(�������$    I���K  D�T$(D�T$H��@  L��I�H  譮����$   ���  �t$ ��H  L���{�����$   ����  D��H  I�G@1�A�y�@��H����M��E����  L�81�D  H���H�H��H	�I9�u��I�L��9�s�L��菱��I�4$I;t$��  �U�I�D$I�L��H�H��H;�j  H9�u��I��I�GI+�H  H9��K  H)�L$ H�<$E1�H�T$(L��$   1Ҿ   ������$    H��H�D$H�X�  H��$   H�t$(H�<$H��������$    H���  I�4$L��I�H  �T�����$   ����  H�\$H�T$(L��H�CH�0�l�����$   ����  H�K1�I�T�I+�H�H�T�H���P9�v�|$< �+  H�D$�(H�D$H�D$����L��L��A�W�D$h�|���I��P  �B���I��8  �6���L�,$�����I��1��e����D$h�   ��   ����Ǆ$      L��I��X   ��   A��8   ��   I��X  E1�L��H��H�D.H��tH�0H�<$�v��I��X  H�D.H�     H�t.H�<$I���Q��I��X  H�D.    E9�8  �H�<$�/��IǅX      H�<$H�������$   �D$L����1���1��	H�D$H�HH�D$0I�t���  I+4�H�<�H���P 9�w�����I��X  �L���L������I��X   L��Ǆ$   �   �����u���f�     H���H  H��X  �WH�G ��v+�p90s-�J�H��H��H��D  �H��;sH9�u�1��fD  �   �f.�     H�G     �G    ËWE1�A9�sF��L�O D)���B�H��H��A;4t-v#�/D  ��D)���B� H��H��A94tr��A9�r�1�Éȃ�Éȉ�f�D�@����     �D�_D�HD��1�9�sFA��L�W A)�A��A� I��H��E;tHv!�U D��)���H��H��E9
t1r?A��D9�r�E1�D9�s?��t=��H��HW D�
D��D��@ ��u"A���D��A�ȍBD���t���D  1�D�ÍB��D  H�    �   ��t$��H��t9�H  vH��H�X  HcFH�1��ff.�     AVAUATI��USH��H�    H�A    ��t.����H  ����   9�����9�vh�1�H��[]A\A]A^Ð��uD1�1�H��X  H��h  �,0���	�H��t�f�     9kw9ksNH�H��u��@ ��H  ��1�9�w���H��H����u��f�     1�9��x���H��1��fD  L���   H�sL��蕨�����O����s�sL���m������7����SD�[	�   �D�CI�}@��E��A����A�����D����)�tPA��H��
D�rE����   L�R��9�tis*1�E��@��J�|�f.�     �
L�R�9�tAHB�A9�s ���H��
D�rE��u���L�RD	�����OE��tW�L�W�9�u%A�
E��t����A�J	����S
�Hc�I�$L��D$�����D$�;�����L�R��D	��H�����L�W	��ff.�     f�AU1�ATUSH��H�zh �D$    tH��[]A\A]�f.�     L�G�   I9�w��A����A��E��A�C�L- I�L9�r�H��H��D��E1�H�} L�L$1Ҿ   �����H�ǋD$��u�E��H�}hJ��H�UXE���w���A�E�1��@ H���LS���LS��	��ɉ�H�JH9�u݋D$�?���@ AWAVL�wAUATUSH��(H��D$    L9��  I��D�oI���o���   L��M��$�   F�*E;�$�   �   A��1���A��A����������@�����A��A�������@�������@�����A��L�I9���  E���l  ��A�M�H��H�L�I��L���   @ A�M�F��A�N��	��ɉHA��HE����   A�HE�pI�XE�@��A��D	�D	��H@����   �D�sL�C�[��A��D	�	ىH@����   A�H��(I�X��A��A�HD	��ɉH�L9���   �L�sE��tD�C��L�sD	��ɉ@���0���A�M�F�HA��HE���?���A�HI�X��A��A�HD	��ɉH@���E����L�C��A���KD	��ɉH@���J���A�H��(I�X�H�L9��[���D�D$A��$�   H��([]A\A]A^A_�fD  �   H��([]A\A]A^A_�@ A��L�L$�(   H��A���D��D�T$�����I��I��$�   �D$��u�D�T$A��$�   E��$�   ����f�     USH��H��H��X  H��8  H�(H�������H��P  H��Hǃ8      Hǃ@      ǃ4      ����ƃ`   HǃH      HǃP      HǃX      H��[]�H��H��(  H��H��8  H�0H�G�    ��H�G(    H���)���h  1����H�H��X  H��Ƃ`   ��c��1�H���D  AUATI���    UH��SH��H��L�*H�T$�D$    L���P���H�ƋD$���  H�KI9��  D�D�N�S���S��	�H��f�V
�S�V	D�EH+��   L�A��H�~A����   �F   A�   ��tA��D�VA�щ�A��H�I9���   E����   ���{D�KA��H�E����   �K��D	�����A���KD	���	ω~�
�����J	��z�R����	���	ʉVH���   H�    H�2H���   �V��   H��[]A\A]�fD  L������H���   []A\A]��     �F   A�   ����fD  L�������D$�f.�     ��D	ω~�
�R��	ʉV�`��� AT1�USH��H�zp �D$    tH��[]A\�fD  H��H��H�T$I��H)�H�;�u�l���H��H�Cp�D$��uƉ�L��H���@
��H�Cp�( �D$H��[]A\�ff.�     AUI��ATI��UH��S��H��H�1�D$    H��tH������I�$    ����   �S��|  ��   �E �� <_wj�   � �| H���W���_wO9�w�sH�T$L��諴��H���D$��u6H��H��H���	��H��� �D$I�$H��[]A\A]��     �D$1�I�$H��[]A\A]� ��t���h���ff.�     f����F �e��fD  AVAUI��ATM��USH��H���   H��t���  �H��t���  �H��tQ�}���  ��Hc���R���}���  I����Hc���R��M��tM�u M��tI�$[1�]A\A]A^��    �   A�   ��ff.�     �> ��   D�_bH�G`S1�E��A�K�f��~L�GxH��A�TP�9�~\L�OhLc�Hc�H��I��M�I�I�I9tH�WxD�@fD�G`f�B[� �fD  I�YI9Xu�A��A�K�fD�Wbf�     9�~�� [��    �ff.�     @ UH��SH��H���������  ���  9�tH�} H��u6H�}H��uH��1�[]�@ ���  ���  �P��H�EH��1�[]�f��P��H�}H�E H��t���ff.�     ��   @��tvUH��SH��H��H�Wb�OH�ЍT;Ww5H�u H�}H��H��HShH�2H�zH�Sp�1�f�CbH��[]�D  1Ҿ   �T�����u�H�Cb�f�     �ff.�     @ AWI��AVI��H�4
AUL��M��ATUSH��   H�T$����A�ą�tH�Ĉ   D��[]A\A]A^A_�f�     L��L���Ş��A�ą�u�I�F@M�W(J�,(I�:H�XM��t	�8 ��   �D$<    H9���   D�(E����   A����   H�XH9���   �@A�����D$A��E�A�WM�GD9���	  D��I��I�GE���0  A�z�1�1�1��7�L�KL9�rw����KL����	���Hc���I��H�BH9���  H����uH�CH9�r<�3H��@��u�H�CH9�r'D�H��D�� A�w�D$@    �t$H9�sS A�   L����������D  A����  A���d  E1�H�CH9�r���\$E�H������D  ���y��у�?��@�L$D��t_H�XH9�r��P��tNH�XH9��y����@H�H9�s)�h����     H�CH9��S����H�H9��D�����u��    �D$A�WD�9���  D�hL�T$(A���D�\$ A��@�	���M�G D��L�L$@�    �����T$@I�G ���|	  D�\$ L�T$(E�o�|$I��H�|$ I���|$ J�(��	  H�CH9������E�C�I��I��I��   D  L�HL9�������8L���������n  ���U  L�HL9��X����0L�ȉz�r��@�C  H�pH9��6����8�@��	����B���|  H�^H9�����������F	����BH�� A�GL9��  H�CH9�������3H�   ��@��t*H�CH9�������{��A���{D	�����Hc�H�:H�B   �� t)H�xH9������D��@A��D	Ș��H�H�BH���σ�@���+  @�������1������f.�     H�XH9��3���D�XA���S���E���D$    �b���@ 1�����f�     H�pH9������� �B������\$@L��L�T$�����L�T$����  A�G+D$�n���H�|$ ��A�jL��M�O D�d$H�DA��H��H�D$M�H�T$L��L��A�IE�AA����������3  M�O �KM��H�C I��K�)A��)�H�2L�H��   uH�z   ��  ��~n��D�ZLcBHc�H���zH��H��HcH��H��H��H��?H��* �  H��D�Hc�H�P�HcP�I��H��H��?H��* �  H���Hc�H�P�H9�u�I�� L9l$��  E�������     H�^H9��������N����	��N	ȉB�{���fD  I�G�D$    E1�I�GA��thH�SA�   H9��J�������  H�SH9��2����[H�H9�s$�!��� H�SH9������H�H9��������u��D$<    H�D$H    H�T$HE��H�D$@    H�D$@A�G0 H�T$xH�D$pH�؋\$L�`L9�������������D�����x  ���$���F @ A�   H�t$P1��   fD  H�D$pH�F�D����������   ����  ����  H�D$xH�F�A������   A����   M�L$L9�����H�F�H�V�E�$M��A�   H�D$pH�T$xH��H��D��������  ���  ���`���I�T$H9������I�$HD$pI��H�F�D���������J���I�T$H9������A�$��A��A�D$I��D	�A��H��H�F����7����    H�F�H�V�A��A��H�D$pH�T$xE9��E���M�G(���  �$� �F A�   A�+  ����A9�����H�T$p��H�T$@I�WH��H�D$HH�D$@H�T$HH�D$pH�T$x�E9������I�W��H��H�D$@H�D$x��A�   A��  �,���A�w0H�T$@L�������D$<��uL�������L��I�w0�@���I�(�gW��D�d$<�s���L��I�w0L�D$����L�D$A�G0A�PA�@b�DA;@��  A�PA�@`�DA;@��  I�(A�w0H�T$@������D$<�n���fD  I�T$H9������A�$��A��A�D$I��D	�H��H�F��g���fD  I�T$H9������E�$L��E9������M�WI��I��H�F��.���D  I�T$H9������E�$L��A9��q���M�WI��I��H�F��"���D  I�T$H9��J���I�$HD$xI��H�F������@ L�HL9��#����8��A���xL��D	��������     L�HL9�������0��A���pL��D	��������     A�BL�L$<�   D�\$ ���D�T$���D$�J���D�d$<I��I�GE��������D$D�T$A�G�D$ I��I��I�G�����@ �������HcrHcz�Q�H��H��H�f�H0HxH��H9�u��|��� A�������D�d$�����I�G �H���A�   ����A�0 ��   I�PbA�HH�ЍTA;P��   H��I@pH�T$HH��H�D$@H��IphH�VH�H�D$PH�T$XH�FH�VH�D$`H�T$hH�F �  H�V(f��A�D$<    fA�@b������   �   L���$������J����X���A���e���1Ҿ   L��L�D$�������u$L�D$I�@b�L����D$<   ����H���,����D$<����L��L�T$�-���L�T$�9���A������ff.�     AWAVAUATU��SH��XL�o�����M���u  A9�H  �h  H��I��A����	�n  A�� @  �I  H��I�X  ǃ�   ltuoǃ�       A��0  D�EI���   H��X  D�eH�T$L�D$H�4$��P��L�D$H�T$L��ǃH      H�4$H��0  ����A�ą���  H��X  A��H�PH���   H�P H���   H�P(H���   H�P0H���   H�@8H���   �����fA����   w  ���   A���  A���  H�CP    H�Ch    HcE9�tH���B��A���  �A  H�ChL�CPI��L�CpL�SxH�CX    H�C`    E����   ���   H���   Icw(Ic f��~^�J�H��H��H�@ HcH��H��I��I��?J��
 �  H��Hc�H�P�HcP�H��I��I��?J��
 �  H��Hc�H�P�H9�u�Mc�Mc�I��I��H��H��?H�� �  H��H�H�CPH��H��?H�� �  H��H�H�ChH���   H�t$0�k���H�L$0H�D$@H�T$8H)�H�K@H�C0H�D$HH�SHH)�H�C8��    A�   H��XD��[]A\A]A^A_�A��   M��(  ���|������NH�D�I����     I��(I9��U���A9$u�A�GA9D$u�A�D$I���   A�t$��H�<$���������������I��X  ���I�x  �T$H�D$�T�����������T$H�<$��A�t$�'����������A�|$��E1�H�$H��HD$A�t$A��D�L�Y@H�D$A�����|$A����A������A�������A���@��@��   ��@�πH�AHA�Љ|$A�|$I�<H9�rVL��H������D��I9�sNL�d$(I��L�l$ ��L�H��H9���   �E��tD�j��D	���H9��L�l$ L�d$(�D$$�D$�D$��@�D$A�D$1��D$�ty9�r�s ��9�vj�7D������L��L�aE��tL�a�I��	���A9�r�vV�z�@ H�CPL�ShI��������LkD$��H��H��L9��  fD  H�<$�'����T���L�l$ L�d$(�Q���A�T$A�$�D$�z  ��I��	���H�D$A�$A�T$�D$�@  ����E�d$	�A	�H�<$輎��H�|$ �����H�D$A���  A���  Hc@H��9�t��H����=��H�t$A���  HcvA�H�CpH����=��A��0  H�D$L�L�$$L���ۊ�����u���H�t$L��L�$$貌��A�ą��Y���H�4$H�F@H�NHH�PH9������D�D�҃�����  ���V  ���,  L�HL9�������@A������A��H��M��H�D$D��@����@����  @����  1�1�@���[  D��@����@����  @���~  @���P  A��A������E����  A������L�D$�։�H��I��H��I��Mi��   L9���������   ��L�D$H����H��H�s0H��H��ƃ�   ��H�S8L��H��H�����   D�H�S@L��E��H�����   H�SHH�T$ǃ�   stibH��H�sXH�� H�C`    H���H�SPI�W@D���   H�Sh���   A��  @ �0  Hc�H��D�D$H��L�L$H��D�T$�I���D�T$L�L$��A��D�D$�������   ����  ���   ����  ��H���   ���   ��A��D  u������Hc�H�H�$H�SHA���7  E����  A����  I��A��E1�A��   �   �   Hc��'D�0I�D E1�A��I��A��   A��1�E��@�Ń����0  ���  ��tE	�A��t�A��u�D�0A��   H��E1�뼉։�H��H��H��H��H;|$��������I�qH9������A�I�����������I�yH9������A�A�AA�q��	�A�AI������	����I���I�qH9������A�A�AI���+���L�HL9������L�XH�@H�D$�����L�HL9��_���D�X�P�p��A��A	��P��A	��P�@��	�	�H�D$����L�HL9������PD�X��A	��P�@M����	�H��H�D$�\���I�qH9������A�	I����Hc�H�|$����I�qH9������A�9A�I����	�A�yI��	���H�|$�X���I�qH9������A�	A�yI����	�H��H�|$�,���A��A��A	�E������I��H�D$����I��E�A���E�������L9�w������A���   tD�0H�<$�A��������L)�I��A��A��   ��Hc�9�G�1�E1������I�1�A��I��A��   ����t8����9�uE�)I��A�ŀtD	�E�A��t�A��uшA��   H��1���A���   �l�����e���I��E1���E1�E1�A��   �   Hc�A�   �&D�8I�D E1���I��A��   A��1�E��@�Ń���tc��uOE��u��t�A��u�D�8A��   H��E1���E	�A�   ��L9�v�E�I��E��A��E��E1�A��E��u�E��u�E��A�   ��A���   �����D�8����f�     H����  AUATUSH��H��H���   H���   H��  L�hH�G(    H�G0    H���i���H��  H��Hǃ      �O���H��  H��Hǃ      �5���H��   H��Hǃ      ����H��(  H��Hǃ       ǃ�      Hǃ�      ǃ�      �����H��X  H��Hǃ       Hǃ(      ����H��8  H��HǃX      ǃH      HǃP      ����H��h  Hǃ8      ǃ0      H��tD  L�&H���]���L��M��u�Hǃh      H�s@L��Hǃp      ǃ`      �)���H�C@    H��[]A\A]�fD  �ff.�     @ AWAVAUATA��UH��SH��1�H��X袂����tH��X[]A\A]A^A_��    H���   ���F H���T�����uҋ�@  �D$<    ���  �   ���   0RFPu����   w���  9v���   
  u�D��  H��L�������D$@���n���H�t$@H�������ЋD$@���R����ʁ�23  �  H�}�t�I��M)�L9���  k���_H9���  �D$<    H�E���	���E���   I9��������  H��D��@  老���D$@�������H�t$@H��臆���ЋD$@��������   A9������Ak�H��莁���D$@�������H�t$@H���E���D���D$@���w���H�t$@H���x���H�ƋD$@���[���A�ĉ�h  H�����d  �߀���D$@���5���L��H��踂���D$@������H�U@J�4"L�JL9���  ��J����	��J	ȉ�l  �B�J����	��J	ȉ�p  �B�J����	��J	ȉ�t  �B	�J
����	��J	�1ɉ�x  �zL��A��A��t������Ƀ�@��u��A��A��t@�� A������Dك�L�H9��+  E��tI�JH�B@��tH�B�R��	��ɉ��  @��u��HH������	��H�	ʉ��  E��t#�@�� ��   �H��H��	��҉��  @��@t@H�HH9���   �H���H�HH9���   � H�H9��~   ����u��D$@    H�PH9�rf��H��	��ɉ��  �P�x����	��x	����  E��t8H�PH9�r'�@������  � �   �(���H���E����D$@   H�������D$@�D$<�������H�M8���  H��H��h  H��p  D���  H���  H�Ɖ��  Hǃh      H�$H�D$�R~���D$@�������L��H���+����D$@�������H�E@N� L�hH���  M9���  ����P��	��҉��  �P���P��	��҉��  �P���P��	��҉��  �P���P��	�H��H���  �P���P	��	�H��H���  �P
���P��	�H��H���  �P���P��	�H��H���  �P�шT$&�����  �L$'u!L�hM9��  �P�@��	И���  �|$& ��  I�EI9���   A�U A�ME�E����	�D	���  A��N�4(M9���   H��  H�l$L��I��H�L$(L�T$�f����  H��L)���  H�xI9���  �D�`��A	�A��fA����  E��I9���  �HJ� �����H	�f���'  f��u�H�L$(�r�H�$�����D$@��t������D$@   H�����H����|��Hǃ�      H��x  �D$@�D$<���^�����H  L�{H�KH��H��H�C ��t0H��X  �z��u7H��1���     H���r���u��9�u    ��  H�C    ���  @��uH�KH�C��   ��`  H��H��H�� @��HE�H��H����HE�H�C��tH�K@H��  H�C(H����  H��  �����H���  �C8    H���  H�C@    H�C0H���  D��H���   H�ChH���  f���   H�Cx���  H�{pf���   ���@f���   �������)���D)�D��A9�L�f���   ����   ����   ���  f���   ���   ���   �gfff1��@�F H�\$@f���   �����H�T$@����f���   i���  1���f���   H�cinu  H�D$H耳����`  ���t���H�K@�j�����H  H��X  ���2  �r�1�H��H��HƋH9�L�H��H9�u�f���   �C���H���   1҉�L�L$<E1��    H�x8蕭��H��H�C@�D$<��������u�H��(  H��H��H֋G�H�� H��(f�B���f�J���H�B�H�J�H�B�H9�uԉk8���  ����H��  H�C(�����H�P$H9��l����P���P��	���A���  �P���P��	���A���  �P�@��	ИA���  � ���I��  �r������   �#���1������L�T$H�l$L��M�nM9��j���E�L�T$C�M��D�\$L�D��0  I9��B���H�<$1�E1�L��L�L$@�   �M���1҃|$@ L�T$H��8  D�\$t"����A�LV����A�LV	��ɉ�H��A9�w�M�M�M�eM9������A�E D�t$&��@  A�EA����D  A�E����A�E	������  A�E����A�E	������  A�EA�U��	�L��H+E@HD$A��H��P  D���D��H  ���|$' t���|$&�������L$�������@��@�|$����� ���L$&���A��L�I9������H�<$��E1�1�L�L$@�   �����|$@ H��X  �����H��1�D�\$&�n�0H�����p���	����|$�rH����|$ �8�G  H�p�@��	����BE���  ��~L�f�v����	�	��B��H��A9��T���A�4$I�D$E��tA�|$��I�D$	����|$' �2�Z������  �d���I������I�EI9�r~E�u L���  H�\$I��L��E��tiI�}H9�rTA�UE�m I�L9�rB��t�@�F �;tH��H�HH��u�A��뽹��B L��L���х�t�H�\$�D$@����H�\$�   ��I���D$@    H�\$�~����L�f�����F	��������H�p@������fD  H��  ��     H���   H�H��   H�FH��  H�FH��  H�FH��  H�F H��   H�F(H��(  H�F01�Ð��0  f�1�� �   �f.�     H��   H��8  H��1��H���     �ff.�     @ ATI��USH��H�/H�X�Y��H��(  D���;J����uFH��(  H���   H�JH�KH�J H�K H�J(H�K(H�J0H�K0H�J8H�K8H�J@H�K@H�RHH�SH[]A\�ff.�     �ATI��USH��H�/H�X�
Y��H��(  L���+J����uFH��(  H���   H�JH�KH�J H�K H�J(H�K(H�J0H�K0H�J8H�K8H�J@H�K@H�RHH�SH[]A\�ff.�     �H��0  �$?��@ H�GH���    H��(  t+SH��H��H��H�t$�f���H�T$H��0  H��[�@ H���   H��0  1��ff.�     @ USH��H��H�H�t$H��(  �ӡ��H�|$��H�{X�X��H����[]�f.�     H����  USH��H��H���   H��(  H��t��@��H���   H������H��   H��Hǃ�       �����H��  H��Hǃ       �����H��  H��Hǃ      �����H��  H��Hǃ      ����H���  H��Hǃ      ����H���  H��Hǃ�      �{���H���  H��Hǃ�      �a���H��P  H��Hǃ�      �G���H��X  H��HǃP      �-���H��8  H��HǃX      ����H��@  H��Hǃ8      �����H��  H��Hǃ@      �����H��  H��Hǃ      �����H���  H��Hǃ      ����H�C(    Hǃ�      ǃx      H�C0    H��[]��    ��    SH��H����F ��V��H��tH� H�C81�[�fD  �   [Ð���  ����   AW��AVL�<�   I��AUI��ATUS1�H��L���  �.�D  H��L9�t?I�4@:.u�L��������u�I���  �
   1�H�<�K���H��[]A\A]A^A_�@ H��1�[]A\A]A^A_�1��@ AWAVAUATUH��H��SH��H��HH�F H�$H�FI��H�D$�V8H�L9��^  H�PH��8[�N  H���S8L�L;\$�:  A�<]��  �D$ E1�E1�H��H�D$(    L��E1�E���D$    E1�I��<<�p  ��0��	w`�|$ �T  L��L�T$A�RHL�T$H����   L��I��A�R@L�T$A�J����   I�H�T$H)�H�XL9���   J�D0I�H����  A����  M����  L�d$E1�M+"A����  E���K  A����   I��M9�r�L��L�T$A�R8L�T$M�L;\$�@  A�<]����I��I��M��;  L��fD  �C   H��H[]A\A]A^A_�H��    �T$H�<$H��I��L�L$4�   L�T$��L�\$ ��Hc��g����T$4L�T$H��  ����  L9�   L�\$ ��  B�I�UI��B�(I��M9�s1@ L9�   �w  B�H��  I�MI��B�(I��M9�r�A�   ������     B�I�EI��C�(I��M9������L��  I��~�A�@A�P��Љ��D$����Hc�H��   I9���   H�<$�   L�L$4�   L�T$L�\$ �f����T$4L�T$H��  ����  L9�   L�\$ ~6B�I�UI��A�   B�(I��M9��"���I��H��  H9�   ʋT$���\����Pʉ�I9�rV�|$H�p(H��   ��H��H��0�    H�����H�H��   H9������H��ʉ�I9�rM��I)�I9�}��D$4   I�ߺ   L�ӉS�|$ �����H�<$L������H��H[]A\A]A^A_�B�|3� I�F��$���I�������     H��t�|$ �o���L��L�T$L�\$ A�R@L�T$A�r����   L�\$ I�M��I��L�I��I��?I�I���N���H�T$(H�<$I��L��L�L$4�   L�T$ L�\$����T$4L�T$ H�Å�uJL�\$L��L�T$L��A�   H�L$8H��M�A�RXL�t$8L�d$(�D$L�T$�,���@ L���K���I��L�������I��L�����I�������I���D$4   A�B   �����AT1�UH���   SH��H��H��0H���Uh����   H�D$H����   H�H�<$I��I1�I)�I��   trL�����H�|$L��H�$���H�|$L��H�D$�x��H�|$ L��H�D$�f��H�|$(L��H�D$ �T��H�<$H�D$(H�D$H��?H%  ��H   H�D$H�T$H���  H���  H���  H���  H�T$H���  �#����t+H�D$ H��H���  H�D$(H��H���  H��0[]A\�f��E   H��0[]A\ÿ`�F �&0��fD  H��H�Љ�H���  ��H��H�4�����1�H���ff.�     1�@�� wH�6     ��H����D  AWAVI��AUATUSH��8L��  L�n H��H�^�V8I�H9���  � ��0��	��  L��A�VHA�vA��  ����  ����  I�H��H�H)�H��H9�~A��  H9���  I���   ��  I�I���  A��  L��H������j  I�M��   A��  L��L������I  I�I���  L��   H�|$����(  �D$& E1��D$     D�l$D�l$�Af.�     <>ttL��A�V@I�H9���  A�F����  A�</�P  <(�H  L��A�V8M�>L9�v2A�<eu�I�GH9�v�A�nu�A�du�A��Q�����t�D  �D$�|$& A��  �o  I��H  ���F �   H�H����� ���R  I��P  L�|$1��L��A��0  ���,  I���  I���  �   L���
H�A��0  ���  Hc\$ I��P  �   L����I��H  H��A��0  ����   I���  �   L����I���  H��A��0  ����   I��  I��  ��L��
H�A��p  ���~   I��  ��H��HI��  H�PA���  ��uYI��  1�L��HI��  H�PA��p  ��u4I��  1�H��HI��  H�PA���  ��t� ��<t�   A�FH��8[]A\A]A^A_� L��A�V@A�N��u�L��A�V8M�&L9�v�L��1��% <>t,L��A�V@A�V��u�L��A�V8I�H9�s�� </u׃���f�A��  M�&�����<(�9  I�GH9��i���I�W�D$' H)щL$���t$L��A��p  ���E���I��H  J��    H�D$(�D$J��� A�.u?I��H  �   ���F J�<��L$ �� ����DL$�   �L$ �L$&DȈL$&L��A�V8�|$' tL��A�V@I�L��H�T$A�VHM�I9������H�T$�t$H��I)�A�IL�L$A���  �������I���  J��    L�L$I��H�E��B� �D$���D$E9�  �4�������D  I�GH9��0���H��I�W�D$'H)Љ����D$����fD  AWAVI��AUATUH��SH��8L��  H�^H���V8M�>L9���  A��PЀ�	vK<[tGI�GH9��r  �Y�F �   L����� ���V  ǅ      H��8[]A\A]A^A_�D  I�N H�$<[��  L��A�VH�D$ A��=   �>  L��A�V8I9s�H��8  I���   H�D$H��tDH�<$����H��@  H�<$Hǅ8      ����I��  Hǅ@      H��t	I���   ��D��(  Mc�H�<$1�L�L$,E1�L�Ѿ   E���   L�T$�E���H��8  �D$,���  L�T$H�<$L�L$,1�E1��   L������H��@  �D$,����  I�E H�$D��I���   ��D$,����  E1�E��~9H�$D��M���   f�     �ރ��   ���F L��A��  A9�u�H�$L��A�V8M�.I9��^  D�|$�$    H�l$L��D�d$�]�    <]�H  ��0��	waE���_  L��A�VHL��I��A�V8M�.I9��]  I�EH9��  L��A�V8I�.H9���  �E <du�L�mI9�s
�}e��  E����   L��A�V@A�F�������I���fD  I�GH9�vG�j�F �   L����� ��u/ǅ      ����A�F   H��8[]A\A]A^A_�f�     I�GH9�v'�y�F �   L����� ��uǅ      �4���A�F�   H��8[]A\A]A^A_�f�     A�FH��8[]A\A]A^A_�D  I�G�D$A�   L��I�A�V8I9�$���������H�EI��H9�v�} /u	�$9L$A�F   �����     A��I��L��M�.A�V@I�H9������A�V���{���L)�L��D��H�|$H�ōHA��  A�F���T���I���   Mc��$J��� �.��� �}f�O����}�}������>���H�l$M��ǅ      M�>����� I��H�l$M�}��A�} /������$9T$������0���ff.�     f�AW��AVI��AUATA��UH��SH��H�GH���   L�x8H�1�H���  H�<к
   �n���H��0  I��H���&��H�{8��D��H���H�C0    )�H�Ch    �Hp������1��H�D��Hǃ�       Hǃ�       ��Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       Hǃ�       I�vXHǃ�       H��0  ǃ�       Hǃ�       Hǃ       Hǃ      Hǃ       ǃ�       H�Cp    H�Cx    A���   ���=  H��0  H�J0H�M0H�J8H�M8H�J@H�M@H�JHH�MHH�JPH�MPH�JXH�MXH�J`H�M`H�JhH�MhH�JpH�MpH�JxH�Mx���   ���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   H���   ���   ���   ���   ���   ���   ���   H���   H���   H��   H��  H��   H��  H��[]A\A]A^A_�f�     SH�H��H�wXH��(  H���   肹��H��tH�{X��+��H�CX    [�f.�     AWAVAUATUSH��H���  H�   H���   Hǆ(      �׷F �T$�   �L$@L�D$�C����F H�D$H��  H���   H�x��B��H��  H����  H��$�   I��1��H   H��H�T$t�   L���   �H�L����p��D�d$tH��  E����  H��$�  H��t	H���   ��H��$h  H��t	H���  ��H��$  H��t	H��   ��H��$�  H��t	H���  �Ѐ�$8   ��  H��$�   H��tH����D�t$tE����   �D$����   A��A����  ��   Hc��  H�S�CH    H�C    H�C H��H  ��(   H�Ct	H��H  H��  ��H�C0�F H�CH�S(H���>  H��  H���>  � ���0  �
8�t1< �q  <-�i  �� t	��-�
  H������   �
8�u��FH��H���f.�     A�   H���  D��[]A\A]A^A_�D  L���   I�EL��1�1�H��Hǃ      �D$x    �1�L��L��$   HǄ$0      HǄ$(      Ƅ$8   �DZ���D$x����  ��$8   �D$x��  �D$t�����D  H��$(  H��$�   �C���HǄ$(      �(���f�H��  H��tH�C(H���   �C8    ���F H�C@    Ǆ$�   	   H�x�?��H��$�   H��  H��$�   H��   H��$�   �D$@��t��$�   H�D$��$�   H��$�   H���   1�H��(  H��H�x�+�������  H��(  H���   ��'��H��(  H��    H�PhH�ShH�PpH�SpH�PxH�SxH���   H���   ���   f���   ���   f���   ���   f���   ���   f���   ���   f���   ���   H�C    f���   ��*  ���   tH�C   �@tH�K�@ tH�K H�|$ �����M�m@1�H��1�H�cinu  H��$�   H��$�   I�}虑��A�ƅ�t����t=�   �e�����   �   f��$�   ����  v1����  ��uX�   I�}Ǆ$�   EBDAf��$�   �&D  ��u0�   I�}Ǆ$�   CBDAf��$�   H��t1�H��1������A��E������� �FH���k��� A�   ����D  �   L���SY���D$x������H�%!PS-TruI�G@H9�8  �D$x   L���Z��D�\$xE�������1�L���W���D$x�������I�( M�g�u  H�T$xL��L���k��D�T$xH��$(  E�������L��H��L���	X���D$x�������L��$0  H��$(  �D$t    H��$�   I�H��$�   H��L��$�   Ǆ$�       ��$�   L��$�   M9��>  L�l$(M��H�\$ �xD  </��   I�EI9���   M�uH��L��$�   �ҋ�$�   ����   H��$�   I��M)�A�W���wL9��   H����$�   L��$�   M9���  A�E H��$�   <F�x���I�EI9�v���F �   L����� ����    H���ҋ�$�   ��t�L�l$(H�\$ �[����A�������     H��$(  L��蠰���D$xHǄ$(      �D$t������L��$0  1�����D  �   I�}Ǆ$�   1talf��$�   �`���1�I�} Ǆ$�   BODAf��$�   �B����H����H����$�   L��$�   M9���   L���3 H����$�   ��$�   ������H����$�   H��$�   L9�sX�8ku�H�PI9�v¿��F �   H����� ��u�L9�s,H����$�   H�t$xH����$   ��$�   u	L��$�   �L��$�   �;��� L�l$(H�\$ ��$�   �D$t����������  *�  �D$t   �����f�     A��F �|�F 1�E��L�d$8M��I��L�t$0M��� ������  M�.I��0M��t�A�E A8D$u�L��蜾��I9�u�H�|$0L��L��������u�Hc�L�d$8H�IH��H��F �P���X  �@���  H�D$ H�   H�D$xH�4I��	E1�1�H��H��H����F ��H�T$x�  ��$  ��$�   �������r���f�H��$(   ��$�  �D$X���  u�D$t   H��$  ��   HǄ$(      H��P  H��$8  H���  H��$@  H���  H��$�  HǄ$�      H��X  H��$�  HǄ$�      H��H���  �-�����$h  ���,  H��$p  ��L�l$`E1�H�D$8�D$XI��H�L$0H��8  ���D$\    H�L$ H��@  H�D$PH�L$(H�\$h� I�GL;|$8�1  I��H�D$0E1�N�$�H�D$ fF�xH�D$(J����F A�G�D$DM��t�D�D$XE��~�E1�L�|$HM��L�t$P�f.�     I�GM9���   I��K�\� L��H���P�����u�M��H�D$ L�|$HH�߾��F �   fF�4xH�D$(J����� ���=����D$\�L$DD9�OȉL$\�&���fD  L�d$8����fD  H�eTypeFonH9P������xt���������D  L�|$H�����fD  �������H�s0������    L�l$`H�\$hǃ,      �D$\��0  ��$@  ��(  �X���I�GL��IL��H��$(  L��$0  Ƅ$8  �P���D$x������L��$0  ������tN�������H�D$ H0  H�D$x������D$\    �g�����$  �����H��H�|$ �P��$�   �����H�D$ H�  H�D$x����f.�      H�H���   �Pt�W�@u��)ЉG1��+w1�9wv�F�f���O�P�   9�s��)�9Gv���щ�fD  1�1��ÐH��H���   �   H��1�H���H��@ U1�SH��H��H�?H���   ����E\�������UlH�K0)���H�H�C8�Er��H�CHH��1�[]�@ AVAUATUSH��H�6�D$    H����  L���   �   M���@  ;V �7  ���B  ��fA�|$ I�t$�E  ��v   E1�A�   H�V�L)�H9���   I�$�   D�@D��D� ��A	�E��D���   E���  D�h�PA��D	�D��I9���   A�t$lA����H��Ƈ�   A�D$\H�0�wh�����   ��Ǉ�       �G`stibL�H�wL�G H�G    H�G������  @ �9  H�EI��$�   H���   ���   D�pA��D���   t���   ��A��L�I;D$vy��   H��[]A\A]A^�fD  fA�|$ A�T$vI�t$������RA�   A�   �� �   ����@ D�h������    H���#   []A\A]A^�fD  E1�D��L�L$1������I��H���   �D$���e���A�F�J�+I�D  ���   H�H9�v#L���    �2H��@�1Hc��   H�H9�u�I��L9�u�H��(  �@   �D$����ff.�     @ ATUSH���   H��tWH���    H��L���   tH���   H���   �	N��H���   L���z���H��L��Hǅ�       �d���Hǃ�       []A\�@ � �F �&��fD  �FL�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H����t?��uI���   �Hl�   H9�t�@ �   �f.�     1��9���f�     I�@@H�@H�� H��H9�t۸   �D  UH��SH��H��H�7H���IK����tH��[]�fD  H�S���F H���X����u��C���f�� ulH�Sf= tYH��uv\f= uHǃ�       Hǃ�       �CTu:H�3H����J����u�H�sH��H���   H��[]��M��f�     H���   w�H���   []�ff.�     AW��I��AV��AUATU��S��1�)�H��(  L���   D��Hǆ�       H�<$L���   1�L��L���AJ�������D$8�L$���  ��$�   <�e  ��$�   ����  I���   f�{l ��  I�G�KrM�wH��H��I�Wf9Kp�  �{b tI�Of�{fvI�OH��$�   E1�1�L��    I���   H�D$�}����$�   H��I�G@���!  �Cp�{VA�G8   �H   D�cZD�sXf�E�C`��fClfE��Hc�f�E �H   LD�fE��H�}LD�L��� ����{lH�� ��H���Hc�H�EH9��q  H�}�H   L�������H�� H���H�EHǄ$      L��$   �{hMuǄ$  nmra�   f��$  1�H��$   1��@�F ������$�   ��u<�Cu�St8�r%)�H�S��H�I�G H���   H9���  fD  Ǆ$�      I���   L�������I�w@H��芣��I�G@    ��$�   A�G8    H��(  []A\A]A^A_ÐH�T$>� �F L����T���������f�|$>MZ�D$8   ��   L���i����D$8����"T$��$�   ��u�����@ H��I�G����� L��H��$�   ��   �C\��H��I���   ��$�   ���W���H�4$I�   H�    H�FH���   ������$�   ����������������;���Ǆ$�      �����f�     �t$@L���#G���D$8�������H�T$B� �F L����S����������D$B�D$8   f=NE�5  f=PE��  I�H����  I9���  �D$8�������Ǆ$�       ���u������� H�}L��H   �_���H��H�E�v��� L�t$H)�L��H�rH��L���[����$�   H���   �������H��H���   H��H��   �ǯ��H���   �( L���   L������H��M��M��H�H�   L����y��H��H���   ��$�   �������I�W(I�WI�G0�F H�у�����   H�ɺ �F � �F HE�I�W0�~����t$@�D$DL���Hc��E���D$8���b����t$F�D$DL��)�Hc��gG���D$8���?���L���cI��f�D$f��wBD�t$�$�LI��f����e  ���@��   H�ID$@L���%I��L���f��u��H��Ǆ$�      �����H�������I�G0�F �����t$@L����D���D$8����   H��$�   ���F L���Q���D$8����   H��$�   PE  ��   H���  ����H�L  � H#�$�   H9���   f��$�    I�    ��   1�H��$�   D�t$H�D$���'H��$�   H9�$�   ��  ��f;�$�   �}  H�T$���F L����P���D$8��t��\$1��)���Ǆ$�      �����L�l$�\$�l$ �   1�� �����L��\$�T$ �zD��I�L$@I+L$HL��H�DH�D$�G���T$ f�������H�|$ ������Hk�vI;T$�m���I����z  I9��j���H�T$8��   L����W��I���   �D$8������Ik�L��Ht$�9C���D$8���w  �   L���E���D$8���^  L���G���L$I���   L����H���L$H���F���L$I���   L����H��H���   I�D$@�5F��I���   L���V����D$8������\$����H��$�   L��\$�B���D$8���x���H�T$x���F L���RO���D$8���Z���H��$�   f�D$&  L�l$H�D$�\$�l$ ��$�   ��$�   �D$&�9��^  H�L$��L��H�H�t�B���D$8���'  H�T$H�`�F L����N���D$8���	  H�D$P�   ������H��������L��H!�H�D$PH�$�   H��H�D$(�A���D$8����  H��$�   ���F L���jN���D$8����  E1���$�   ��$�   A���9��v  H�L$(��L��H�H�t�FA���D$8���^  H�T$X�`�F L���N���D$8���@  H�\$`��   �����H��������L��H!�H�\$`H�$�   H����@���D$8����   H��$�   ���F L���M���D$8����   1�H�������$�   ��$�   ���9���   �4�    L��Hc�H��|@���D$8����   H�T$h�`�F L���>M���D$8��uz�D$c��V���H�|$Hu�H�t$L��Ht$p�1@���D$8��uMH��$   �@�F L����L���D$8��u0M;7tlI��M����D$8��������A���l���f�D$&����L�l$�\$1ҋl$ �����L�l$�\$�l$ ������|$8 �����Ǆ$�       ����H�|$H�T$8��   �'T��H��I���   �D$8��u�H��$  H��$   L��H�$�   H+�$�   H�H���   ������D$8���0���L�l$�\$�l$ �^���D  H��t;USH��H��H���   ����H�s@H���:���H�C@    �C8    H��[]�@ �f.�     D  H�H  H�G1��H�G    ��    H�O1��Q�y���9�rKD�YD�	D����D�9�w5@��fA9�w)f9�r$��D)��ƃ�D)����H�QD)�H��B�f�1��ff.�     f�H�OD�1��yD�A��E��D�D9���   ATUS�fD  D9�vt�iD�A����E����D�D9�AB�A����A��D��fA9�wD��fA9�sA�ZE��D����D)�A��)�BH�QA����E�D�D)�H��B=��  t�[]D�A\�D��ff.�     H��P  H�H��X  H�1��f�     �   �f.�     �   �f.�     1��ff.�     f��ff.�     @ USH��H��H�/H���|��H���  H��H�C0H���  H��H��H�C8���  ��H�H�CHH��1�[]�f�USH���FH�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H������   ��u H���  H��  �   H9�tH��[]ÐH���   []�@ H��1�H�����H���  H��H�E0H���  H��H��H�E8���  ��H�H�EHH��1�[]�f�     H�C@H�@H�� H��H9�t�H���   []�ff.�     @ AVAUATUSH�.H���\  �   ;U �   H��  ��L���   A��H�RL�4к   A�vE�NE�A�FƇ�   ��0  f���   A�   D)�D���   �����   �����  ~'����  ����  �P?�������   �@ ���o  �P�����   A�V��A��H��D���   H�A��H�0���   ����Mc�H�Hc�Hc�D��H�wH���  �G`stibH��  H�W H��L�GH�G�
��A��  @ ��   Lc��   ���   H��L��L����W������   I�vL���]:������   H���   L��L���;������   H��0  H��H�������   H��H��1��tdH���   ������  ��uJH���   I��v;I��I��J�t�fD  ��HH���H��H��P��P��H��P�H9�u�@ 1�[]A\A]A^�D  [�   ]A\A]A^�f��P�������   �y���@ �P��҉��   �b���D  [�#   ]A\A]A^�f�H���   M������J�<.@ �H��������   ��U	щ��������   ��3	ʉ�������	ʈV�H9�u�H��0  H��H�������H���   I���$���I��I��J�th�     ��HH���H��P�H9�u�1������ H����   SH��H�F 1�H��H;u�2f�H��H�� H9H�t#H��H9�u�   I�    H��[��     H�GH�sH9�wH)�L�$L�D$�8��L�$��t
�S   � H�SL�D$I�H�SI�H��[ø   I�    �f.�     �@�F ����fD  AUATUSH��H��L���   H��  L�������H��(  L��Hǃ      ����H��   Hǃ(      H��t���  ��~b1��fD  H��   H��9��  ~EH�Dm L�$�M��t�I�4$L��苒��A�|$ I�$    t�I�t$L���n���I�D$    � L���X���Hǃ       H��p  L���>���H�s(L��Hǃp      �'���H�C(    H�s0L������H�C0    H�s@L�������H�C@    H��P  L������H��X  L��HǃP      �Α��H���   HǃX      H9��   tH��[]A\A]��     �;6��H��H  H���   H��[]A\A]�f�H��t�V���fD  �ff.�     @ ��~aAVA��AUI��ATI��UH��S1�fD  H�} L����Ѡ����tH��A9�u�[1�]A\A]A^�f�     Hc�H�[[]I�D��A\A]A^�1���     SH��H��   H�Ӌ��  H���t���H�¸   H��t�z H�Bt�   H�C1�[��    �C1��   [�ff.�     SH��H���� ���u ��� �F � �F HD��
B��H��[�@ H�T$���F ��A����u��T$�f��T$�f�S�T$�f�S�T$�f�S�T$�f�S1�f�S
H��[�fD  ATH��UH��SH��H�� H��p  H��h  L�L$L�D$������D$��t
H�� []A\ÐH�t$H����@��H��H�D$�D$��u��� ���uу�H��x  � �F t���F H���A���D$��u�H���  H�H1�H)�H=�  ~H�� ��H���  H���  H���  H�H1�H)�H=�  ~H�� ��H���  H���  H�t$H���  H��I��   ����L!��l����D$���&���H�t$H���  H��L!��I����D$������H�t$H��� ���H��   tYH���  H���  H���  H���  H���  H���  H���  H���  H���  H���  H���  H���  ����H���  L!�H�������D$���u���H�t$H���  H��L!������Y��� AWAVAUATI��UH��SH��H��   H���   1�H�$�2���D$`��tA�   H�Ĉ   D��[]A\A]A^A_ÐH��`  �`�F H���\?���D$`��u�H��`  fcpu�H��h  H��t�H�EH��v�H��H��	wH9�vH��	�	   HF�H��h  H�<$L�L$`E1�1Ҿ    �f��D�t$`I��H��p  E���R���H��h   ��  E1�� H��h  A�WI�� I��H9���  L��@�F H���>���D$`��t�H��p  H�<$�����D$`Hǃp      �D$8�������H�   H�C    M�������H��h  H��p  L�L$`H��L�D$@�   L���   �����D$<���*  L�l$<H��L���=���T$<H�D$@���	  � �����   L��H����  �[=��H�D$�D$<����   H���8��8��H��H�d$`H��H;T$��   H�D$M��   L��A�   H=   LF�E1�1�E1�D���  L��L�|$�}d��I�ǋD$<��ux1�H�|$ �X  H�\$L�t$L��L�l$ I���D  I��H��M9��  H�ھ��F �D$@t���F H���=���D$<��t�H�\$E1���D$<   �E1�E1�L��L���?���L��L���4����D$<�D$8���8���H��h  H��p  H��t/H�>   �4  1��H��H��H�<   �  H��H9�u�   H��H��������D$8��������D$ H��h  H��p  L�L$`L�D$@�   H��L���   �����D$<�������L�l$<H��L���;���|$<H�D$@���|���H�� ���� ����h���H��L��H���H����  ���5  �4���ȋt$<���6���H�|$@H�D$`�� �����  H���������H��H��H��H9�����H����������  M��   L��H����  HG�1�E1�H��H��  �fb���T$<H��  �������H��  L�x��  A�   �^f�     A�fA9G|A�GA�W��9�}%1�E1�E1�E1�fA�G1�fE�OfE�fE�_fA�GI��I��L;�  ��  H�t$@L��H�������D$<I�G    ��t�H��  L��������D$<Hǃ      �D$8�������H��h  H��p  L�L$`H��L�D$@�   ������D$<��������   H���S/���D$<�������H����1��H��H�D$@���
  �1��I��H���0��H�L$@�� ����r���I����  A���  H��  MF�H�P�I9��M���H�UN�d�M���@  A�   �8�    ��6��H��  K�H��H9D$`seL�bI��M9��  H�L$@��L��H��u���8����D  �D$����fD  �{6��H�D$�{��������  �c6��H���m��� L�H�B��    H��L��p  I����  �D$    1�M��E1�1�1�I)�L�|$�    H��I�L �WH��L�AH��H�qH��L�L�PM9�vAL�8L�L�QL�9L�xL�yL�xL�yL�xL�yL�A�   L�PM��H�pL�@H�qL9���   I)�L9Q��   L9��v���L�|$E��t�D$�D$I9��@���H�UI�EH9���  H��H)�I9}�x  1��I�MH9��g  H��H)�I9}�W  �HI�� H��I9�w�I�EH9��;  H)�I9UvI�U�D$8    �h���f��D$`	   �.���H���������H��H��H��H9����������3����������7��H������D�D$<E�������A�   L��H���D$@�  �}4���|$<�������I��u�H�D$@H��h  L�L$`H��H��p  L�D$@�    �D$8    H��0  L���   �����D$<���/  L��H���t6��H��H�D$@�D$<���  �� ����H�����H��  ���F t�`�F H���6���D$<����  ��  ��  f9�����f=� �������  ��  f9������f��� �����D����M��E1�A)�)�1Ҿ   A����L��H�Mc�L��L���C]��H��(  �D$<���P  K�4?H���$+���D$<���  ��   D��  ��  D��  ����  f��fD9�rf9�w@��fD9�rf9�vD��A��D����D�f��   E������D��D)�E�ă�D)����)��Hc�HM@�A�	�D$@�m
  ��	�f���t����H;�  r�   Hk�L��  �   L��(  L��I�4 �fA9�v(�Ef�     �,��1�f�����I��A���fA�F�fD;�  ��  H���D$@u��,����H���l+���D$<�     �D$8���8����|$ �v  H�CH��H����{   H�StH��H�C���  L��   H�C    �<�F �D$<    L���   H�D$@    L����H�D$H    H�D$P    H�D$X    �B���H��t;�x t5H�P����<Ot<Iu#H�C   ���F ���<O�4�F HE�H�D$P�B�F L���������H��t&�x t H�@� ���<BuH�KH�D$H �F @ �N�F L��������H��t$�x tH�P���t���<NtH�T$X�    ��\�F L������1�H��t*�x t$H�x����b  ���<N�W  H�|$@D  1�E1�H�D�`    H��t�X���H�D�`M�tH��H��tH�D�`    H�|�@H��u����    L��M��uH�D$@�F �   H�D$`   L��L���:���t$<H�C0���B���E1�J�t�@J�l�`H��t7H��H9C0t�  H��H��H���Q���H��M���%  I���  H�H��I��I��u��  �D$<�D$8�������H��   ���  �k�F �Q���H��t
�x �|  H�C(    L�t$8H��  H�<$1�M���C8   E1��   �    H�C �Y���T$8H��H�C@���i���H�     A��  H�@    H�@    H�@    H���  H���  H�2H��H��?H1�H)�H=�  �2��1�A��A)�D���  fD�} �F�F L��   D��L���y���H���  H�@H��H��?H��H1�H)�H���� ��  ��  f�E���F L��D���6���H��t'H�PH�xH��?H1�H)�H��� �;  H�E�  ���F L��D�������H���  H�@H��H��?H��H1�H)�H���  ��  H�E�� A��� �w�F L��D������1�H��t*H�@H��H��?H��H1�H)ʹ�  H���  ��1Љ�)Ѻ��F L��D��L$�m����L$H���L  H�@H��H��?H��H1�H)�H���  ��  M����  L�}��  A��  L�}L���H   D�D$�L$������L$D�D$I��H�E�   f����  ����  I��H��L�������D���  L��   H�E���F L��D������H��H��t%���F L��D�������} tH��t
�x �E  D�t$8E������������D  H�������H��H�)�: u�-H��H9�u��������.���������&��I�������D$8    ����H�D$H+D$H��H�4�H�\$L�l$ �v"���D$<���  H�D$����  L��H���D$@�?  ��+��D�\$<E1�E�������H�|$H��H�|$`H)�H9��  �  M��   L��H=  HF�E1�H�T$(H�J1��U��D�T$<I��E�������H�T$(H��H���"���D$<���g���H�L$E1�1�M��   L���GU���|$< �B���H�|$ H��   ��  I�H���F  H;T$(�;  M�GE1�L�|$I��H�l$L��H�\$ L���dH���  H;D$(��  I�4L��L���|��D�D$<I�GE����  H��H;\$��  H�U I��H��H����  H;T$(��  I�4L��L���n|��D�L$<I�E����  �U�A�WH�E����h���I�G뗺   H��H�������D$8���n�������A��fD;�  �,���D��  � ���1�����Hkt$�H���^ ���D$<��������D$<S   E1������I����������L�t$8H�pH�<$L���{���L$8H�C(���l��������,������H�gfffffffH�HH��H��?H��H��H��H)Ș�1�)�f�E������1�)�A��M����   f�����L�����1�)�A��A��Mc�L�}�i���D���  L��   L�}�O���M��u�L�}L�}��   H��H)��e���������D$<    �����L�}�����N �  ����D���  L��   H�E�����D$`   �����D$<   ����L�}L�}f���i���H���Z����   A��  �u���I���   �   �J���D���  L��   f�E�����L�<$H�pL��L���0z���|$8 H��P  �����H�uL��L���z��H��X  �{�����	�����H��(  L���Jy���D$<Hǃ(      ����L�|$H�l$H�\$ �D$<	   �����L�|$H�l$H�\$ ����L�|$H�l$H�\$ �D$<    ����H�U�����AVAULc�ATL��I��UL��SH��H�� ������tWH����  H��L���   ����L��L����@ <��  ����  L��H  L��H��L��L���   �M�������  1����  t	f����   H��X  L��P  H���	  M���   ���߀�I��   �P��߀�S��   �P��߀�O��   H�����F �   H����� ��td���F �   H����� ��u�4�F �   L����� ��t2H�ƿ��F �	   ��� ��uj���F �   L����� ��uRf�H�cinu  H�\$H�D$�Hf.�     �   H��tH�߉D$�*����D$H�� []A\A]A^�f�     H�\$H�D$    H�T$1�1����F �/U��H�� []A\A]A^�f�L��L����F <t���`���H��t?H������H�� �   []A\A]A^�f.�     L���   A��   ��> <�����   �U���f.�     �H����   �1�����   E1ɀ�-��   I����������H�ʃ������� �F 1���r�<D  L9�KH���� �F H��H�P���H�ʃ�@������ �F ��r�H��H��M��HE�� 1��D  H��������H��H��M��HE���     �WA�   H���O���ff.�     f�H���   �1���txE1���-��   ��H�ʃ������� �F 1���r�9 f=�J�� �F H�����B���H�ʃ�@������ �F ��rʉ���fE��E��fD  1��D  ��  ����fE��E���    �WA�   H���c���D  �����H�VH9Wr�����f.�     1��ff.�     f�H�H��  H��  H�RXH�G 1�H�W�H�G     H�G    �ff.�     @ H�OL�O H��H��H��tH��E1��fD  L�@H�H)�I9�s,H9�v,L9�r'H��H��L�H�:H9�t%v�H��H�H)�I9�r�1��f�J�H�����    �B�����D  S�H�_L�W D�HH��H��H����   M��H��1���     H�xL�L)�H9�s,H9�s\H9�wWH��H��L�L�M9�tUs�H��L�L)�H9�r�H9�sPH�������[L�L��G��I9Ӻ    DG���D��fD  H�H����    �B[D�����ÐE1�1�[D��fD  H���   H�H��   H�1��f�     USH��H��H�?H��  �(���H�E@H��H�C0H�EHH��H��H�C8�E��H�CHH��1�[]�f�     AW�   AVAUATUSH��L�6A;V �  �B����E  I��  H��    H��H)�H��H�Q`D���   H���PD�hD�`�hH�p H�H(�@���   ���   ���   �E���fA����   ��   fA����   fA��u�   ƃ�   f���   �    ��A��I��H�{0���   ��A����? H����   ��H�CH���   Hc�ǃ�   stib��L�kPH�C0���   H�S@��H�C8I��  �p
��Hc��5���1�H��[]A\A]A^A_�@ fA���m���ƃ�   �a���f�     A��  ����@ ƃ�   �<���@ ƃ�   �,���@ U1�SH��H�W�D$    H9�sRH��H��H�l�@   H�����t9H9�wAH��H�����w5H��H�L�L$�   L��tI��H��D$��uH�kH��[]�fD  ���������ff.�     �SH��H�H��t'H�3�{p��H�    H�C    H�C    H�C    [�f.�     AUI���   ATUH��SH��L�eH��H���   H���   L���   L�L$�D$    J�"�H��H��H���   �D$��u$H��   H��L��H���2~���(
�D$L��   H��[]A\A]��     �@�F ����fD  I����������ʉ��������� �F ��1���r�L@ L9�w;Hc�H��H���� �F ���H�P��@�������� �F ��r���    H���������    ��ʉ��������� �F ��1���r�DfD  f=�w2Hc�H������ �F ��΍B��@�������� �F ��r�ø������f�     �FL�H�V��t%��H��H�J$H�9��8��8H��H��?H��H��H)ʋH�� H����t?��uI��  H�HHHH@�   H9�tø   �f.�     1��9���f�     I�@@H�@H�� H��H9�t۸   �D  AUATUSH��H��H���   H�7H���n��H���   H�    H��t"H���F���H���   H����m��Hǃ�       H���   H���m��H���    Hǃ�       H���   tQE1��@ I��L;��   s;O�,dI��J�.�xu�H�pH��I���im��H���   J�D.    L;��   r�H��E1��Em��H�{X L�c`Hǃ�       t@�    I�4$H��I��I��8�m��I�t$�H��I�D$�    ��l��I�D$�    L;kXr�E1�H�{p L�cxt:�I�4$H��I��I��8��l��I�t$�H��I�D$�    �l��I�D$�    L;kpr�H�s`H��E1��l��H�C`    H�sxH���l��H�Cx    H���   H�������H���    L���   u�Yf.�     I��I��L;��   s7I�4$H���3l��A�|$I�$    u�I�t$H���l��I�D$    � L���   L��H����k��Hǃ�       H��[]A\A]�H����   USH��H��H���   H��  H��t����H��  H���k��H���   H��Hǃ      �k��H��   H��Hǃ�       �sk��H�s(H��Hǃ       �\k��H�C(    H�s0H���Hk��H�C0    H�s@H���4k��H�C@    H��  H���k��Hǃ      H��[]� ��    AWAVI��AUATI��UH��SH��(L�oH�G    M��t*H�H� ��F H�@��F H�@��F H�@��F H�@ ��F 1�M���s  �U ���g  ��   ���W  H�$    E1��   H�D$    H�D$    H�D$    �)f.�     �ȉ��������H��t���t��+u܀~ u�A�   H��u�I�1�A���F L9��#  fD  ����  �Ѓ�H���������s�  @ �����������rH�����u�I9��P  H9�IC�I�$H�FI�D$H�,�E����   �; ujE1�I;D$�V  H�pL���P�����u<I�t$I�$H��    H�M���,  H��I�t$H� ��F H�DH�     1�H��([]A\A]A^A_Ð� H�kI�t$H9���   1ɀ}  ��M�l$I9��&  �U �������H�1I��I9D$�o����U���������   �������4�у�����   H���fD  ����������o����E  H���E ��u�I�t$H9��_���1��a��� H��L���4���������I�t$A���F ����@ H��I9�tн��F �}���H��H�     H��(1�[]A\A]A^A_�I9�vHH��1����� M�l$I9�v1H��H�������M��tI�$붾   �V���H��H��I��H������1���f�     SH��H��H���   �}���H��tH� H�@H���   [H���@ 1�[�ff.�     �H��  H����   H���    ��   H����   �> ��   SH������H��H��t1�H��tO��t2�   ��t[�fD  H�B�   H�C1�[ø   [��    H�@�   �C1�[��    H�@�   �C1�[��    �   �f.�     AWAVAUATI��UH��SH��H��(H���   L���   H���D$    �[���H��tFH� H�@H���   H�ЋC����  ����  ���F  �D$H��([]A\A]A^A_� L���   H��L�������I��H����  L���   L;��   �^  I�H�IH��H����F H��RvH���   H��8���H���   K�RL�4�H�I��PA�V�P�@A�V���(  ����  ���v  ���F �   H����� ����  �E< ��  H�&     H����  I�����F �   H��L���   ��� ����  �E< ��  H�&     H����  I�FH�C8�D$�����f�H�sL����d��H�C    M�������A�<$ �����H�T$L��L���he���fD  1�M��tA�<$ tL�������H�C�[����M���o  L���   I�JL�L$L�Ҿ   L���'=��H��H���   �D$������H���   H�@H��H�     H�@    H�@    L���   H���   �)����    I�F    M���y���A�<$ �n���H�T$L��L���d��I�F�D$�������L���   �B����     1�M��tA�<$ tL���
���I�F�����H���   I�>L��L���E���D$���M���L���   �)��� L�������I�F������    ��F �   H����� ��u0�E< w(H�&     H��sI�FH�C@�D$������    ��F �   H����� ����   ��F �   H����� ��������E< �����H�&     H�������I�FH���  ��D$��߀�P��  �C0   �Z���@ L��� ���H�C�D$H��([]A\A]A^A_�f�     L��H��L���   �D$    �6���H��ty�D$�D$�������L��H������I������fD  L�L$E1��   1�����@ �E< � ���H�&     H�������I�FH�CH�D$�����    H���   L���   L�L$L���   H�J�d:��H��H���   �D$���\���H���   H��H�@L��I�    I�B    I�B    L�$�,q��L��L�L$E1�L�X1Ҿ   L��L�\$��9��L�$H��I��D$�������L�\$H��L���so��L�$L��L��H���   I�B   I�:H�pS��B���D$�������H���   �D$    ������Mu�C0   ������C������C0    �u����   �k���ff.�     f�AWAVI��AUATUSH��H���   L���   1�H�|$�T$�D$x    L�<$�&���D$x��tH���   []A\A]A^A_�@ L��H�T$|�x   L��H�      �D$|    H��$�   H�       H��$�   �g��I�ǋD$|���@  H��$�   A��  I�WHE1�I�G@I�F�   �   fE�OI�GpH��$�   I�GH    I��I�GP    I�GX    I�~8I�ohI�o`H�T$@1�H�|$ Ǆ$�       H�D$8�(8��D��$�   I��E����   H�\$PE1�E1�   HǄ$�   �C H�D$   �  H�D$(   L�|$HI��H�T$H�|$K�4/L)��%��H�D$0I�M9���  H�|$0 tSM���K	  H�|$��  �t  L�l$L�L$8M���   H�|$ K�\- L��H���m7��D��$�   I��E���  M��H�\$PL�|$HH�|$ L���^����$�   I�o8�D$|����  I�H��H���~  �}0t�Mf�M4I�O@�9��tvH�MXHMptlE�GA�wD����D)�D�ED9�t)�f�}f;Mtf�MA�wf9utf�uA� f9}t��f�}��f�MD����D�D�E
D9�t�f�u
H����  H���   H���'  H���   L���   �   H�JL�L$|�N6���t$|H���   ����  I�G8H���   H���   � I�o8��  @ O�'I�D$E�D��A9���  A��
��	  A����	  M���fD  ��
tI��I�vI9�����C�\7M�7��u�A� A�D��<#��<����tI9�|mM�fH�D$(�   A�A��
�����A���
   �   E����� M����  �D$x<��E���H�������   �3����H�\$�[���fD  L)�L�T$hL��L�D$HD�L$`H��H��$�   H�T$(L�\$X��$�   L�\$XD�L$`�����$�   L�T$hu:L�T$`L�D$HH��L��D�L$XH��$�   H�T$(��$�   L�T$`D�L$X��$�   �������D���D  H��u�D$|   �Af�     � �����   �D$|H��tH������I�o8H�<$H��1��[��I�G8    H�|$@�����L�4$I�w(L���~[��I�G(    L��L���k[���D$|�D$x<��������������D$H��  ��~	f���c  H�   H�C    H�KH����  H���    �  ��F H���S���H��t
�x��  H���    �  �k�F H���)���H���   H�pH����  H�<$H�T$x�U[��H�C(�D$x���G���L��  �D$|    L���   HǄ$�       HǄ$�       HǄ$�       HǄ$�       H�C    M����   I��$�    ��   �<�F L������H��t
�x�[  I��$�    tj�B�F L���[���H��t
�x��  I��$�    tC�N�F L���4���H��t
�x�]  I��$�    t�\�F L������H��t
�x�.  1�E1�E1�JǄ�       H��t�Pi��J���   M�tI��I��tJ���   ���    L��M��uHǄ$�   �F �   HǄ$�      L��H�T$|���H��H�C0�D$|�������E1�L��$�   K�4�N���   H��t5H��H9{0t� H��H��L���<g��H��M����  I����  J�<0I��I��u�� �D$|�D$x���W���H�EP�C8   E1�1�H�<$L�L$x�   �    H��H�C �51��I��H�C@�D$x������I�$    I�D$    I�D$    I�D$    H�E@H���  ��H����  ��  H�EHH���  H����  ��  ���H���    fA�<$��  �F�F H���I���H����  H�@H���� H����	 ��  ��  fA�L$H���    �  ���F H������H���	  H�xH��� H=�	
 ��  I�D$�  H���   H����  ���F H������H��t!H�@H���  H����  �O  I�D$�� H���   H����  �w�F H���y���H���p  H�PH���   E1�H��t#H���  A��  H����  w����1�A��A)�H���!  ���F H���$���H���  H�@I�|$H���i  H��u
I�|$I�|$I�|$H�MPH�<$1�L�L$xE1��   L�e`�5/��H��H��  �D$x������ǃ      H�}PH���X  H��L�M8I�L$1�A������f�H��H��8H��H9��+  H�1f�PH�0L9�w�L9�u׉�  ���    H��M���*���H��J�<1D  �8 u� -H��H9�u�����f.�     L��  H�C(    ����@ I�Ľ   ���� L��K�4'L��L)�E1�H��I���c���]����     H�xH������������������<N�����H��$�   ����H��H��?H��?H% ����H�  f���H�E@������     H�H��?H% ����H�  f���H�EH�����D  H�@H�������� ���<Mt<C�����H�K������    H�@H����������߀�Ot	��I�����H�K� ��F ���<O�4�F HE�H��$�   �\����    H�@H�����������������߀�N����H��$�   �r����    H�@H���7���� ���<B�)���H�KHǄ$�    �F �����    I���7���H���    t=���F H���9���H���    I��t#���F H������M��tH��tA�|$�f  H�BODA   H��$�   1�1����F H��$�   H��$�   �1���SH�D$x������H�SPH�H���   �	����    A� I��M���h����H���  H����  �T  H���  I�|$��  A��  I�|$�H   褪��H��I�D$�   fE���S������K���I��I���x���I�D$�9���fD  H��������   �h���fD  H�E(������    H���   H�U ����H�EH����   H��H��H=�  ��  HF�I�D$����� A�<$H���   �   ����fA�D$����D  E1��w���H�gfffffffH�HH��H��H��H��?H��H)���1�)�fA�T$�=���f.�     �1�)���H�I�D$����@ ������1�)�A��H����  f��������fD  A�D$��H�I�D$�"��� I�o8������    H���N �  H��?H1�H)�����I�D$�����f�M��H�\$PL�|$HǄ$�      �����x�����I�|$ �����H�pH���w���L�4$H�T$xL���Q��H���   �D$x�������I�t$H�T$xL���Q��H��H��   �D$x��������E ���<I��   �E���<S��   �E���<O��   H�����F H���F`����tL���F H���5`����uH���   �4�F � `����t&���F H���`����uvH���   ���F ��_����uaH�cinu  H��$�   H��$�   1�H��$�   1����F �F.���������   A��  �	���I�|$I�|$���T���H�������H��$�   HǄ$�       �I�GH1�H�D$@�7���ff.�     @ H�    L�WM��toH�1�E1�H� D  M9�sJH�N��A���t!I)�f�     H���L�A���u�L�WI��M9�v�� L�WH��M9�r�H=��F t� H��1��ff.�      H�OH��t0H��v1H�H�t��f�     H�PH��H�P�H9�u�H��H�O�fD  H�G    ��    AWAVI�ι   AUM��ATI���&�F UH��L��SH��   ��À� �ۅ���   A�D$< ��   H�&     H����   I�x8H���h  H���    �Z  ��F ����H���C  I�}8H����   H���    ��   ��F �~���H����   �����I!E I���C H�Ĉ   ��[]A\A]A^A_Ð�8�F �   L����À� �ۅ�tl���F �   L����� ����   A�D$< ��   H�&     H����   I�T$��tA�D$ I�T$I�}8L����������j����    A�D$< w�H�&     H���E����q���D  I�}8H�G�4�F H�GHH��H��1���\��I�}8H���F �p������������������I�}8H�G�4�F H�G@H��H��1��\��I�}8H���F �0�����������������A�$M�}8�����  L���	u��  �<	�(  H�����u����  ����   I���   L���^���H����   A�����H�H�RH��H����F H��RvI���   H��8���A���tD�3H��tZ�ytTM�uHH��L��N�F L�������Å������I�EHL��L������H���<���I�}8H��L���=����������fD  �I�4,����   H9�s,�F�<	t< uH��� H9�t�F�< t�<	t�<"��   I�}8H��L����������u���f.�     � A�<$ A�	   tI���   L���A���H�������D�3I�4,H���  �@H����u�i���f.�     H������P���< t�<	t�<"����H��8���f�     �F� �W�����L���P���D  H���A�$ A�	   �{���� A�<$ D���Q����d���ff.�     �AWH��H��AVAUM��ATI��U1�SH��8  M�@8�D$    M��tI���   ���F �   H����À� �ۅ�u]�H�� wTH�&     H��sDI�u@�v��tM��t���|  H��H�pL���������H��8  ��[]A\A]A^A_�fD  M�M A����   �Q�F �	   H�ƻ�   ��� ��u��@	< w�H�&     H��s�M�}hH�T$��   I�E    I�E8    L�������\$���p���I�UhI�E8L���   L��L��H���   I�Eh    �I���ÉD$���9����\�F A���F 1��@ H��I��H��S��  I�<$L��L��H���+���ÉD$��t������D  �   �[�F H������� ����   �H�� ��  H�&     H���r  A����   �����H��I�}HH�¾N�F �����ÉD$������I�EHI�]8H�xH����  �? ��  �����I�UpH���   H��I�EH9���  Hǃ�       �   �+���D  �   �k�F H������� ����   �H�� ��   H�&     H����   A����   �����H��I�}HH�¾N�F ������ÉD$�������M�]HM�M81�I�{H��t
�? t����I�{fA�AE1�H��t�? t�i���A��fE�Q
I�{�����fA�AI�{ �����fA�AA���fE�QfA�AI�M �B���@ �   ���F H������� ����  �H�� �v  H�&     H���b  M�eHH�ѾN�F H��L�������ÉD$�������L������H�t$�#���I��H����  I�E8H��H�0��F��I�]8H�D$1�L�L$E1��   H��H�    H�H�M��H��\$���t���I�E8L��H�8H�D$H�P��T��I�m8H���v  H�] H���i  �; �`  I�E@H���   H��H�D$    H�D$    H�D$     �@H�T$(�E0��U��L�`I���   �  H��L��H�|$0�IT��L��H�T$0�{�F H�|$������Å���  H�|$ �/  H�|$�2���I�M �����     H�pH������ �   ��F H������� ����   �H�� ��   H�&     H����   A����   �9���H��I�}HH�¾N�F �?����ÉD$������M�UHM�M81�I�zH��t
�? t�d���I�zI�A1�H��t
�? t�K���I�zI�A 1�H��t
�? t�2���I�}XI�A(��  �   fA���   I�M ����@ �}�F �   H����� ����   �@< ��   H�&     H����   A����   �R���I�P�4�F H�|$01�I�P@����S��I�}8H�T$0��F �����ÉD$������I�U8�4�F H�|$01�H�JH�JH���S��I�}8H�T$0��F �J����Å������I�$��C ����������fD  �   ����fD  Hǃ�       1�I�E    L�L$E1�1Ҿ   H���L��H���   �\$��tI�E8Hǀ�       �_���f�     I�M I�$��C �D���fD  I�]8H�T$�(   L������H���   �\$������I�E8L��H���   �B���ÉD$�������I�U@I�E8�RH�@8�����P0������   �����I�z �0���f��vfAǁ�    ����H������f���   �   �   E�F�fA���   �����H�D$H�@X���C��-�����H�        �   H��H��u.H�      H��u+H�      H��������E0    �t����E0   �h����E0   �\���H�|$���������f�     AWI��AVI�ι   AUATUL��SH�����F H��H��(M�h8��D$    M���   �� ��u �C���o  �P����#  <�  H�E � ��   �}�F �   H����� ����  �S�� ��  H�&     H����  H�}HL��H�ھN�F �M����D$����  H�EHH�xH����  �? ��  �r���H���������I�EPH��H�EH��H�epH��H9��  I�UPH�UH���X  H���� �  H�U �D$   ��@�af.�     ���F �   H����� ����   �S�� �  H�&     H���  ��  ��  �D$�   ��@H��H����   D�L$�1f�     I�W�H�s����   L��������D$A��E����  H��(D��[]A\A]A^A_�fD  ���F �   H����� ��uw�S�� wnH�&     H��s^%?���H�E0    H�E E1���     ��@�D$�   H��H���I���H�u(L���?��H�E(    �0���H�sI�W��C��� H��@tH�}0��m  �	   ���F H������� ��u4�K	�� w+H�&     H��s��  ��  �D$�   ���� �   ���F H������� ����   ����  H�}0��d  I�uXH��    H)�I�u`L�t��I��A��   ��  H�uA�VH9���  �   ������H��H�E �����D  H�E    I�EP@   �@   L��L�L$E1�1Ҿ8   ����|$I�E`��tPH�U ��@�����@ �K�� �@���H�&     H���,���H���.  �D$�   ����f�     H�M  �9���fD  H�M@�q�����������@ I�uXI�}`���C �8   �L�������D�L$H!E I�ІC �����    H�u(L��L�mH�=��L��H�ھN�F H�E(    L�������D$������L���A���H�t$����H��H���)  H�D$L�L$E1�1Ҿ   L��H�H�����L$H�E(�������H�|$H��H�WH���gK��D�L$H�M @E��������V����    H�}HL��H�ھN�F ������D$���x���L�UHI�z�;���H�E0H����*  �,  H�PH��   �*  H�E0����H�E@�@���   I�UpM�ExI;Uh��  H��    H�M(H)�I��H�H�JI�MpH�PH�E(    H����?����H#E D�L$�H�E ����D  �D$�   ���� �   ���F H��L�D$����� ����   �K�� �  H�&     H����  H�}HL��H�ھN�F �����L�D$���D$�X���H�EHH�xH��t�? t�����I��fE�FH�M    ����I�upH��    H)�I�uxL�t�������   ���F H������� ���h  �K�� �[  H�&     H���G  H�}HL��H�ھN�F ����L�D$��A���D$�����H�EHH�xH��t�? t�B���I��H�E fE�F���  ��H�E ����M�N(M��I��Iv M���  ��ω�@����������F ����  E1��6 A��t�F H���I�҉ω�@����������F ���?  �Hc�I�R��� �F �L9�u�L��A�Nf���7  B�K����������F ��sH�E �   @u
H   @H�E H�ED�L$�����H��������   ���F H������� ����  �K�� ��  H�&     H����  H�}HL��H�ھN�F �����D$���,���H�]HH�{H���X  �? �O  �=���A��H�{fE�^H���=  �? �4  ����A��fE�NH�{����H�{ fA�FA���x���fA�FA���fD9MfE�NfDMMfA�Ff9E fME fD�Mf�E C�f9Ef�E"fMEfD9Uf�ED��fNEfD9UfDMUf�EfD�UH�E    ufE�^H�E@�8 ��  H�M    D�L$�b���H�E0����H�}X��  H�E0H�������I�UXM�E`I;UP�U  H�JI�MXH��    H)�I��H�M(H�BH�
H�E(    �����H�U �D$   ��@����H�E �   @u
H   @H�E A�Nf�������H�E8���   ����H�����F  I9�����������   ���F H������� ����   �K�� ��   H�&     H����   ���Z  A���   A�F��A�N����Hc�I�v(H��=��  ��   H����  ��   fA�N0E1�1�L�L$�   L�������|$ I�F �����H�E    H�M    �?���H�J@L�L$�8   L������T$I��I�E`�������I�EP@I�UXH�E0�p����D$   �[���I�z�+���H�E0������D$�   �<���H�JL�L$�8   L���?���|$ I��I�Ex����I�EhI�Up�����H�u(L���c6������I�UI�U A���@ �׍��D�L$fA�FH�M    ������D$�   ����E1�����E1������1������1������I�UI�U �@ A�~�}���fA9F�=���fA�FH�M    �+���I�MP�D����    ���   ���$��G fD  H���  �1�H���   t^H���  �@ H��0  �H���  ��     f��h  �t.H��h  �fD  H���  �1����   tH���  �D  1��D  1���w�����   ������pG ��!��ff.�      �Wи   ��	v���1���A�����@ D��0  ����������E��tWH��H  1��@ ��H�� D9�t<f9pu�f�x t�f�8tI�8u�f�x t�9�uЉ9��H�� D9�u�f.�     ��   ��x�@ �������     f�xw�f�x	t�:�u��:��     H�H��   H�RH9Qw���     H�w1��f�     1����   wH�W�F��f.�     D�A�PH��HW��BH����u��A�ȁ��   v�1�E1�D��ff.�     f�H�OH�F    �A�����A	���H�1��ff.�     �1�����  wU��H�WH��  ��u�H���N��f	�HD��D  �H�������B�    	�%��  H�H9�HD��H�A������H��1�H��t|�JE�������J	��2�ɉ��r��	���A)��r���r��	���D9�v9��t5B�A�rD�JH�|
����W��f	�tA����	����� 1��ff.�     f��I��L�OD�@A����  ��   fD  D��L�������H��tP�A�����P��	�D���P���P��	���A�9�w0A���   w'A�   L��D������H��u��A���   w7A��두�H���H��	���f��u9A��   u�E1�1�E���    E0�A��   A����  �I���E1�1���f�A9�vcE0�1�E�H�|89�sZB�)��p�����p	���f�H���G������G�f	�t	�����u�A��A9�u�D�A��?����    D)ލ<w띅��(���D���� H�OH�F   �A�����A	���H�1��ff.�     �H�w�F�����F	�f�����G0�����H�G(1���     D�G0L�OA9��  G�\ AUE�P�L��AT��USH���  ��  �fD  f�����   ��A9���   �6I�D������PL�	��҉W<������PH�	��҉W8������PH�	��҉W@������P	�D9�r�H9_8u�f��t7L�'��L�l(I��$8  I�$0  I9��[����G@   1��
�     1�[]H�GH1�A\A]�w4�fD  [�����]A\A]�f��t���H��Ѹ�����f�     AWI��AVAUATUS�_(����  ��   L�7��A�   9_8C_8M��0  I��8  ��A�G4L���p������x}A�G89�B�A�w<9�w�I�WHA�@H��tw��A+G8�H�I�,H9�w��f�     ��9�r�H���B������B�f	�t������t�A�_([A�G,]A\A]A^A_��    �����[]I�G(A\A]A^A_�@ A�N D�>�2fD  ��xL=��  �9���A����  �,���D��)���9������;��9�vʅ�t�A�_([A�W,]A\A]A^A_� E�������������f�     AWA��AVAUATUSL�w�ӉT$�A�VH�t$���A�V��	���  �����|  ����������  �w  H����D$�H��8  H�0  H�\$�H�t$���1�I�|6H�D$�L�wH�H�|$�H�t$�fD  A�|VH�D$�E�DV��A	��<P�DPE����	���9�vE����   ��A9���   H�\$�A�z�4SD�LS��A	�A�2E����	���D��I�\:D��H�\$�!�9T$���   f�����   f���
  H�\$�H9\$��J  �   D  D�A��E��t\L�l$�A;E ��   ���Ä��9  ����  w/��A9�s��    H�BI��H9T$��  H�������D  1�H�T$��
[]A\A]A^A_�@ [1�]A\A]A^A_� f���t�E��t]��D��)��A�DL�H9D$�s��u�D�(D�@1�A��fE	��Y���E�A��L�D$�A;@ sV��A��D!��9����     D�������     E��xsA����  �.���A�=��  �����   )������ 1������f�     f����I���H�BI��H9T$������ 1��|$� ����������fD  D����������������@ AWAVAUATUSH��PH�OD�aD��D�a��A	�A����  �F  D���T$ ���H�t$H�|$�D$����   �D$���  A�T$D�L$1�� A9��  �nD9�sHB�t ��6H�D�8D�@H���D	�D� D��E��D�@A��E	�E��A9�v�A��D9�r�1�|$  ��   A9�s��9t$��   H�|$�������^  H�D$�X(��tV�h,H�D$��hfD  �����<���1�1�A���  말A��f�����  �|$  t4H�|$1��@�����u&H�D$�X(H�\$H���W����k,����  @ 1�H��P��[]A\A]A^A_�D  L�t$M�>M��8  L�|$8M�0  E��L�M��L�L$0�(D�HN�48A�L�t$(��A	���A��E�N�l$D	�L�L$��l$$�l$E�I ��D�L$@A��9�w]D!�f���uTf����  ��I�|>I9�s>E����  �FA��   E1�D$HA���  �D$@��  �A ����������� E��������~�|$Hf����F  D�T$@�|$A��E��D�d$$���  ������H�lD�E �EA��D	�A��D��A9���  D�T$DD�\$L�4f�     G�T �J�lD�m D�UA��E	�E��A9��	  E��H�D A��D�D��D�XL���A	��8E����A���xL�D	�D���A��D��D�PA	�fA���E��EE�E���t���D�\$@D�T$DD�\$LD�t$DD;L$H�  E9���  C�	H�DD�D��D�XH�D���A	�D��D�PL�E����A	��E�҉��P��	��ʉL$J�8�H�L$(�����A	����D$$�L$$��tf��D)ЍAHD$(H9D$0sD��1��D$ �������@��f	��X  fD$D����H�D$8;h �    C��j���A��A���  fD  �L$�|$  ��������H�T$8D��;j �@���1���  =��  �+����L$�   A�)ȁ���  O�����D�L$H�|$E��D�T$@A���  ����E���t����FA��|$E1�D$HA���  �D$@��  ����D�\$@D�T$DD�\$LD�t$DD;L$H�[���D9��X  H�D$(D�\$DA���|$D�T$@D�d$$D9L$��  C�	I��H�D�(�xH���	��(���|$D�x��	���A��9��_  A�|$E��H�L$D�t$DH�lL�l9D�ωt$$E��H�A��H�T$(�<f��u A�E�I���UA�M�����	�	�H��H������9�wCA��A��E��L�E�P�8���xL����H	������	�f���D��EE�D9T$u�H�L$�t$$D�\$@D�t$DH�T$(D9��&���D��D�\$D1��W���D�\$DD�T$@H�D$(�|$D�d$$�q���A������D���(���E1�D;L$Ht9H�D$(D�l$D�������D�������������A���D$   A���  �����|$E��D�T$@D�d$$�Z���A�y�D�d$$E��D�\$DA��D�T$@�|$�@���A�A��|$E��D�d$$A��D�\$DH�D$(D�T$@����H�D$�X(����H��1��t$����  w1�H�t$�G t����H����    �{���H���fD  H�OH�F   �A�����A	���H�1��ff.�     �H�O�A�����A	��Q��)Ɖ��Q	��	�1���9�v�H�L1
������A	�����    ��P1�����  ��   L�OA�yE�A��A	�A��E�AD��E�A	��A	�9�B�E��A��A)�C�M�T	
E9�vcE�
I�JE�RA��fE	�uP����  t8A���H���A��y���f	�u$����  t��A9�u�1�1҉�D  1��D  ����1���A�����     H�OH�F   �A�����A	���H�1��ff.�     �H�O��   H��   ʅ�t6��H�RL���   ��     9�sI9�t��HH���x���9�v�1��)�ω����9��    C��ff.�     L�G�1�A��   �����   Ƀ�M��   ����   �A�AVH�@ATUI���   SL�'������    A�9E�QI��E�A��9�A�B�A�A9�r_��I��E��)���I)�M9�wK��D�u<���t(����A9�r4��I��I)�M9�w'A�)�u�����u�1�[]�A\A^�@ A;D$ r�L9��w���1�1�[]�A\A^�f.�     �1҉�f.�     H�GH�F   �@ȉ�H�1���    H�O1��Q�9�w#)֋Q�9�v�H�L1������A	����ff.�     f�H�G�D�@L�HD��D�@1��Aȃ��tq��9�C�A��A)�C�I�E9�vgE�I�IE�IA��fE	�uU���t;A��@ H���A��y���f	�u$���t��A9�u�1�D��f�     1��D  A����D��A����A��A����H�GH�F
   �@ȉ�H�1���    H�w�F�G( ȉ�H�GH1��f.�     H�G0�����H9���   AUL�_@H��ATUSH�_HL9���   H�OK�[H�/A�����L�L�D  A�1A�IA�Q�A��ɉ�L9��A��IB�H9�r[O�,I)�M9�wO)�A�Չ�A�ukL9�tOH�PD�,H��H9�r.L��H)�L�L9�r E��uCA�   L9�t!H��H��H9�s�@ I��I��L9��o���[]�G( A\A]�@ �G( � D;m s�[]D�o8A\A]H�G0L�_@��    AU1�ATUSH�_D�cA�E����   D�����   I��H��E��E1�� E9���   D�QE9�s)C���I��H�t�D�F�A�A9�s�A��E9�r�1���t6E9�v��A9�t)D���E(H�E0��H�E@H���Q����}( usD�]01�E�] []A\A]�f.�     A���t�A���X����D�ߋv)ǉ�����9��    BƄ�t�D��H�U �E(H�}0��H�}@;B s���t��E8��    �E8D�]0�ff.�     @ H��1҉t$H�t$����H����    H�GH�F   �@ȉ�H�1���    H�w�F�G( ȉ�H�GH1��f.�     H�w0�����H9�wrL�O@L�WHH��M9�saH�WK�IL�H�L���    I��H��M9�t;��QD�Aȉ��H9�A�HB���H9�r�E��t�E;C s�H�w0D�G8L�O@� �G( �ff.�     AU1�ATUSH�_D�cA�E����   D�����   I��H��E��E1�� E9���   D�QE9�s)C���I��H�t�D�F�A�A9�s�A��E9�r�1���t6E9�v��A9�t)D���E(H�E0��H�E@H��������}( u[D�]01�E�] []A\A]�f.�     A���t�A���X�����FȄ�t�D��H�U �E(H�}0��H�}@;B s���t��E8�@ �E8D�]0��    H��1҉t$H�t$�����H����    H�GH�F   �@ȉ�H�1���    H�w�F�G0    ȉ�H�G8    H�G(1��ff.�     @ 1��ff.�     f��    1���    �����H�F   H�1��ff.�     f�D�E1�A��A�E9�v{G�A��B��    H�T��J����	��J	��JD��9�rB�Lf�     C����    H�L�D�Y��A��D	�D�Y�ID	�9�vA��E9�r�1�ÐE��H�L9�s	D�R�h����   �fD  D�E1�A�E9�sfG�A��C��H�L��Q����	��Q	�9�r8�>�    C�
���H�L�D�A��A��D	�D�AD	�9�vA��E9�r�1��D��E�� 9�vD�RE���y����A�����A	����ff.�     f�D�E1�A�E9�vqG�A��C��A�AH�D��HH������	��H�	�D��9�r8�K@ C�
����AH�D�D�@��A��D	�D�@D	�9�vA��E9�r�1��fD  H��E��9�v�D�Q�m���@ AUATI���U��SH��H�_H�{�B���H��t�D�h�Aͅ�uE��u9H��1�[]A\A]�@ �׉�H�������t�I�D$L��H�@H��[]A\A]��H��E���J�<+[]A\A]�(����     ATU����SH�_H�{���������H��t�D�`�A̅�u2�����E��u[��]A\ÐE���J�<#�����1�[]��A\���ډ��f��҉�H�<�����   ��t����     L�H��I��x  I���   H�@H��tI�Q E1��`YD ��D  �   �f.�     H�H��x  �` H�H��x  �` H�GH�@`H��t�����   �f.�     AUATUH���  SH����   I�@H����   A�A9X��   H�pI�p�0��A���pD	����2H�pI�p�p�@��	����1�O 9
skf���t��0  9�sZ[�   ]A\A�@A]�A�A����A�Af	�t5E�Q��E�IA�0��D��Hc���D	�H��%�� H�H;u ��   [1�]A\A]�fD  �]L�eA�@    �����t�E1�� D�XA9��A��E)�D����D���D�D�@E�Mc�M�E�A��E��E�QE	�E��D9�w��<����X���    HE������    H���  H����   ��  �   9���   �HqD��0  �D�I���VL����	¸   ��A�E9�U��    H��H  H�HAH�4�H9�s+ �H��H���J��H��J��H��J��H��J�H9�w�1��D  �   �f�AWH��H  AVAUATUH��P  S��X  HŅ���  H�HH��
H9���  A���D��\  E1�I��A�   I	�f.�     D�AD��D�A��A	�E��I�L9�LF�E����   �QH�qM��I)���Q��	��ҍR�H�I9�}H��������*I��I��?D)�D�y�AA��A	�fA�� �uRD��`  uy��tE�Aȉ�I9���   �B�H�@H�TA��    �ȉ�I9���   H��H9�u��     Eۃ�tI�@L��H9�����[D��]A\A]A^A_�f.�     E1�D9�v�F�2A��C�I�H��ɉ�I9�t=v)�kf�     C���I�H��ʉ�I9�twUA��E9�r��x����     �P�@��	ИA�A��DE��R���f��F�����F	И��D��A���     D�qD���W���E1�[]D��A\A]A^A_� H�L�HI9���   D�L�GfE�D�PfE�PfD�PfE�PfD�PfE�PD�PfE�P��t6L�HI9�wMf�PfA�P
f�PfA�P�@fA�@1��G L��fD  1�A�@
    fA�@1��G L���    �   �f.�     L�WH�GE�ZD�H����  AWAVAUATUSA�	D9���   E����   D��   C�A;��   �_"A�ٍ{��A��Hc�H�H9���   IcjA��A��D��E�Mc�MJ��A����   E��tl�S�Lc�A� �  ����A����I���,�f�     J�<L�ȃ��P  H���V�H��H9�u�K���H����tD��H����"M�A��u�1�[]A\A]A^A_�D  [�   ]A\A]A^A_��     E��tэS�A� �  1�����A���؍�I��L�ʉD$�N�&����    H���F�D��	�������@:H����L9�uދD$�K�!D�:��tf��I�rE��E�A��D��D�E!�D	�A��A��E	�D�:��~��D����@zI�A���&���N�&L��1����v�����I��D�:��u����D��L����D	�����    �   �f���L��H������ AWAVAUATUSL�OH��H�GE�QH�T$��P���  D�
E9��	  E���   D�8�   G�E;��  D�w"D��D��A�փ���Hc�H�H9��  E���t  E���k  IcAA�˺   ��A��)�D��A��D����   H�D$�E��D�|$�E��E�Mc�MYD9�N�1�E1��ى\$����)�����D��)ى|$��L$��   )ىL$�f�E����   D9l$��L  D9D$��1  H9t$��F  DD$���D��I�[�����L$�"T$�AA�ʃ��)  A��H��D��D����A��I��N�&H���~�H��	�������@z�L9�u���A��L�E��L��E��~F� �  D���;��E9�}kL��L;L$�s
A�	H��	�D��D����A��D!�	׺   @�;D)�A�L\$�A������1�[]A\A]A^A_� E��L��I��A���:���� D����E)���!�L��	�@�;�f�     [�   ]A\A]A^A_�f��D+D$������f��E��H���������H��	�����I������f.�     ��G �x��fD  AWH��AVAUATUH���nrekSH��H��(H�L$��@  A�����  H�t$A��   H����  H��H  H���ʴ��A������  H��H  H�|$A�    H��P  �AH�L�A�����A	�f�� DF�E��f���k  H�A
H9��^  �A�Q�q�I	����	�	�D��f���6  A�   E1�1�1�I��������*A�   �S�    ��A9��  E��H�FA��H9��  �F�VD�F��	��V��D	�I��D��f����   ��L�H9�HF�A��u���f��u�M�pL9�r�A�@����A�@	�H��L)���I�֍@�Hc�I9�}L��I��?I���D)�D	���K���A�PM�pʉT$�P���t5E�@A�D��D9D$r� ���E�A�E��I9�����L��I��H��u�E	������f�     E1�1�1�f�     ��X  ��\  D��`  H��(D��[]A\A]A^A_�ff.�     SH��(  H��H���   �I���Hǃ0      Hǃ8      [ÐD��   H��(  I��I�L9�r�3 H�� I9�v'H;0u�L�HM��t�H��tL�	H�pH���%���D  ��   �f.�     AWAVAUI��ATI��UH��SH��8L���   �    ���   ��  ���  H��h  ��    �t$H�L$M����   H����   H�����A�   I��H����   �t$����   H�L$�A
D�AH�\H�Q��A�����AE��D�A		�A�E	���fD9�t[��H�t��,��
H�����J���	��B���A���B�D	���f9�t%���H�H9�u�A�   H��8D��[]A\A]A^A_Å�t��H�D�L�<C�CD�K��A	�A��D�L$tv�3M���  Ή�L9�sdL��L�T$H)�L9�vTI��x  H��H�H�D$���A����u6�CD�L$ȉ�D�ȃ�f���Z  L�T$��  f����  D  H��
L9��c���A�   �6����     L��h  H�L$(� FDBH���   HǇh      I�F    H��I�F    I�F    I�F     H�D$�p������P  H�t$(H���A  H�|$L���������,  I��h  H�T$(H�I��p  �1D�I�A���qA����A	��A	�ȉ�f����   H����   H�p�A��H��H9���   H�pH9���   A��H)�L�I���  ��    H�QA���  H�<M��x  fE��t2�F�L�L�D  �BH����A���B�D	������H�L9�u�I9�rAƅ�  �����f�     H�|$L���s���Iǅh      I�F    I�F    I�F    I�F     A�   �{���D  A�$   A�T$�d���fD  ��D�D$I9�� ���HD$1�L��H��H�D$�9��D�D$H�������H�D$A�$   I�D$����@ A�$   A�T$�����ff.�      ATI�����F UH��SH��H�� H�T$�������tH�� []A\� H�⾢�F H��������u��|$u�<$tH�� �   []A\ÐH�T$I�$H�T$H�U �ff.�     �AUH��ATUH��SH����tLL���  L���  �xtmvH�L$H��H����@  �Å�uH�D$H��I�E �Ѫ��I�$H����[]A\A]�L���  L���  �xtmh�ff.�     AWA��A��AVAUI��ATM��USH��H���  H��8L���  H���  H���  H���  H���  E��uH���  H��H���@&f��t.��H���   H�D9���   B��    H�H�FH9��P  1�1�fA�E fA�$M��tTA�$�D$(A�E �D$,E��uVI�H��tH�T$(D��H����I�FH��tH�T$,D��H���ЋD$(fA�$�D$,fA�E H��8[]A\A]A^A_�f.�     I�FH��tH�T$(D��H����I�F H��u���    D������H�$Mc�I�I�@H9��9���L��H��D�L$L�D$H�L$����D�L$���D$$����H�L$H�t$$H���|����t$$D�L$fA�$�������D��L�D$H�$)�H�L$�t L�H�FH9���   1�fA�M ����� H��D�$H�L$�����D�$���D$$�����H�L$H�t$$H�������D�D$$D�$fA�$E���f���H�L$H�t$$H���Ԭ���|$$D�$fA�E ���M����:���f.�     H��D�L$H�$����H�$D�L$���D$$�K���H�t$$H��D�$�y���D�$fA�E �����ff.�     UH��1�E1�S�   H���_H�oH��L�L$�K�����T$��u]��ti�U H�u��t]�{�H�HA�?   L�L=�f�     H���V�H����t�z���`H��ACЈQ�I9�u�� H��[]ÐH��1�[]��    H����ff.�     ATH��1�E1�U�   SH���_H�oH��L�L$f��D��A�L$�J����T$����   f����   �u H�M���u��	���f��trA�t$�H�xA�?   L�Tu�#@ H���q�H�����q���	���f��t�r�I����`ACшW�L9�u�A�  H��[]A\��    H��1�[]A\�D  I���� USH���G0�D$    9�r1�H��[]�f�H��I��L�G8��H�S@L�L$�¾   L��H���Y���H�C8�D$��uĉk0��     AUATI��USH���Ʌ���   D�i�H��H�F1�J�|�D  �0H���L1H9�u��qL��H�]�Q�����uYI�D$8J�|�H����sH������	��s�	��s�H�t�fD  �
H����H9�u�H9�u��    H��[]A\A]�H��1�[]A\A]þ   �������u�I�t$8H����ff.�     @ ATI��UH��S�ˍs������uVI�D$8��t]�S�H�MI��H�t�	H� ��yH��I������	��y�	�A�P�H9�uډ�H���    []A\Ð[1�]A\�f�     H����ff.�     AWI��I����AVAUATUSH��L�wI�~�����H����  D�(�@A�D��ȉ�	���  I�4>L��E����  E��M����q  I�A�m I�EA��˅��S  �U�I��I�t�1��    �H���T
H9�u����+  ���X  �tL��L���q������)  A�UM�UI�G8E1�A�MA�vI�~	A�   ������	�A�ME�m	�A�NF�*��	�A�vA�   	� Ic�A9�rFH��L�<09�vA�A��L�|0A��D9���   ��wH������	��w�	�Ic�A9�s�H�4��@ D���D�zH��A9�u�A��C�tE�A9��?  A�E�BA��I��E�j�A����D	�E�B�D	�F�*�Q�����u5H��L��L��L��[]A\A]A^A_�����H��1�[]A\A]A^A_��    L��L��H��L��[]A\A]A^A_�L���@ A9���   Ic�H���fD  ���rH��A9�u�C�TA��Hc�L�<�A9�sdE)�O�\�@ A�2A�RI������	�A�R�E�J�	�Ic�H���VB�<
�
�    ���1��H��9�u�G�DM9�u�Mc�N�<�A�    H��[]A\A]A^A_�Hc�L�<�A9�w�A��A�A9�sNIc�H�4��S�D)�L�D�I�D  ��OH��H������	��O�	ʉV�I9�u�D)�A�Ic�L�<��Mc�N�<��x���AWH��AVA��H��AUATI��USH��L�o(H�oA�u��������   M�|$8E����   A�E�H�]
M��H��H�DPH��fD  ��utH9�tP�CH���S��ʅ�t��D��I|$�T$������T$��t��C��S�I������	��S�	�A�E�H9�u�A�E     H��L��[]A\A]A^A_�D  ��D��I|$�������u�����    E1��� M���ff.�     ATH��I��USH�o(H�_�u������ubI�D$8��ti�U�H�K
H��L�D�f.�     ��yH��H������	��y�	��V�I9�uۉ�H���    []A\�f.�     [1�]A\�f�     H����ff.�     AVH��1�AUATUH��SH��H��L�f8�psag��@  �D$��tH��[]A\A]A^�D  �   H��胠���D$��u�H���S���H��f���  �D���H��f���  �ա��f���  v1�f���  H���   []A\A]A^�D���  E1�1�L��L�L$�   L������H���  �D$���Y���J�4�    H�������D$���=���H���  E��t4A�E�L�d�f.�     H��H��蔡��H��f�E�舡��f�E�L9�u�H�������D$�����ff.�      AWAVAUATUH��SH��(D��0  L���   �D$    L��H  fE���  I������L��1�E1�Ic�Mc�D�D$A�   �D  ��H�� fA9��   f9pu�f�x t��f���  f����   f����   f��u����t�Hf���f��	u��Hf��
w�M��I��A��  t��HHc�f���f��	A���v���fD  A�����   ���t
E��x<E��u7I��L��A� �C L�����t7H�{ ��   L��H��A��H�D$� H��L��Cf��vf��
t1�1�H�U H��([]A\A]A^A_�f�A���C ��     Lc�������     f�x u9Lc����������uC�|$���   A���t�I��L��A���C L����N���f��L$f�x DʉL$�{��� Lc\$E�������E����KL��`  1�E1�L�L$�   L���c����T$H�C��uH�sL���[����D$��t(H�CH��L������1�H�C    1�f�C�D$������SH�sL���[����D$��������Lc\$�|��� USH��H���  H��t.H���   H���   H�s藜��H��H��H��[]����fD  H��[]�f�     USH��H���  H��t.H���   H���   H�s�G���H��H��H��[]����fD  H��[]�f�     AUATUSH��H�����   t"H���  L���   H=   t$H= P ��   ƃ�   H��[]A\A]�fD  H��  L���A���1�f��   Hǃ      f��   H��  t71�f.�     D��L���J�4������H��  J��    f9�  w�L�������1�Hǃ      f��  �\���@ H��  L������1�Hǃ      f��   �0����     AUATI��USH��H���   H��H  H�hH��tXD��<  I��I�L9�s.f�     H�sH��H�� �@���H�C�    I9�w�I��$H  H��H��� ���IǄ$H      I��$X  H��tSA��$P  H�@L�,�L9�s'f�H�sH��H�������H�C�    I9�w�I��$X  H��H�������IǄ$X      AǄ$P      1�fA��$8  IǄ$<      H��[]A\A]�fD  H����  ATUSL��p  H��H���   M��t>I��$�   H��t��I��$�   H��tH����I��$�   H��tH����H��A��$�   ���   H���   ��  H��H  ����H��  H��HǃP      HǃX      ǃ`      �����H��(  H��Hǃ      Hǃ      ����1�Hǃ(      H���   f��   H��0  �������   Hǃ8      Hǃ�      Hǃ�      ��  H���  H���G���1�Hǃ�      f���  M��tH��A�T$hH�s(H������H�C(    H�s0H������H�C0    H�s@H�������H�C@    H��@  H��������C8    H���  H��Hǃ@      ����H���  H��Hǃ�      ����H��   H��Hǃ�      ����H��(  H��Hǃ       �l���H��8  H��Hǃ(      �R���H��H  H��Hǃ8      �8���HǃH      Hǃp      []A\�D  H��h   tH��h  肗��H���   Hǃp      Hǃx      Hǃ�      �����D  H��   H�������H��(  H��Hǃ       ����ƃ�   Hǃ(      �:����ff.�     @ SH��H�8H�3�p���H�    H�C    H�C0    [��    H�G@�G0    H��t H�w8H��tSH��H���+���H�C8    [Ð�ff.�     @ SH�H��H�w H���   �����H�C     �C    [��     AWAVAUATUSH��(H���   L���   H�D$    ��  H��H��H���RLOCH�L$��@  �D$��ukH�t$H��w@E1�L�l$�D$   L��H������L��L���b����D$H��([]A\A]A^A_��    L�l$H��L���(����D$��tE1�� L�l$E1��fD  H�T$�(   L��L�|$�a���I�ƋD$���z���A�����A�W	�fA�f���U���A�OH�t$��A�O��	�fA�NA�Wʉ�H9��)�����H���IH)��Hc�H9�����A�A�O��ɉ�A��A�D	�fA�~H9������H��I������ I)�L9������H�|$I�v H�H�I�~I�VI�NL���  �����fD  H��(�   []A\A]A^A_�ff.�     �AWH��AVAUATUH���LAPCSH��H��8L���   H�D$     H�L$(��@  �D$��uqH�t$(H��wFE1�L�d$ �D$   L��H������L��L�������D$Hǃ�      H��8[]A\A]A^A_�f�L�d$ H��L���P����D$��tE1�� L�d$ E1��fD  H�T$�(   L��L�|$ 艦���T$I�Ņ��t���A�A�W��	�fA�E f���O���A�A�WL�D$(��	�f��0  A�OA�W��	�f��  A�wD��A�WG�\��M��	�fA�uA�Wʉ�M9������I9������L��    A���� L�$M��I)�L9$�����f9������H�t$ I��M�}H�I��I�Uf����  A�AI9������C�H�I�D�D�zD�RA�E����   E��D�T$M9��X���M)�L�$L9��H���E1�1��ɾ   L�L$L�������|$ �+���D��  H�t$ H��L�$D�T$M�I�I�L9�s"I��A�K�H������A�K�	�f�J�I9�w�H��(  L�D$(A�E����   E��D�$M9��������  M)�H� ���� L9������E1�1��Ⱦ   L�L$L��������|$ �x�����  H�t$ H��D�$H�I�H�H9�s$I��A��H����A��A��D	�f�y�H9�w�H��   L�D$(A�E��u]��0  I��M�E ��L�L$E1�M�]1Ҿ   L��L���  �B���H��H  �D$�������1�H������������������E��M9��������0  M)�H� ���� L9������E1�1��Ⱦ   L�L$L��������|$ �t�����0  L�\$ H��H�M�H�H9�s"I��A�w�H����A�w���	�f�q�H9�w�H��8  L�D$(��0  ���� I��H��H��tE��   H��(  H��H�H9�r��   �D  L�HM��uWH�� H9�v�H;0u����    H���   L�HM��t9I�H��tH���   L���Ɏ��f�     M�1��f.�     LPM��u�H���   L��L��镎��D  L�W8LWHA��d��  AWAVA��AUA��ATE��UH��S��H��HH�w@H���E  I�BL�PH�D$(E�D��E�Z��A	�I�BH�D$(A�BE������A�B	���9�L��wD9�sHf�     H��H����   D�D��D�X��A	��PE�ۉ��P��	���9�r�A9�w�H�PH�T$(�@L��L)�ȉ�H9���   L�H�HL9���   H�PH�T$(����P��	�H�pH�t$(�xD�PH�L$(@�|$D�@f��wE���$��G D)ۍ�    H�H�AL9�w%H�QH�T$(�H�D$(�Iʉ�ɉ�H9��,  �A���%�   ��H��H[]A\A]A^A_� H��H�   []A\A]A^A_�@ �   �H�PD�L$D�T$D�D$I9�r�H�P�   H��D�XH�T$(H�t$(L���h�����u�H�T$(H�BH�D$(I)ǋ2L���H����H9��^���H���U���H�BD��D�D$D�T$H�D$(�Bɉ�D�L$�����B1�	���9�u6�L  �     L�\$(I�CH�D$(A�����A�C	���9��O  H��H9�u������f�     H�PL9������H�HH�T$(L9������L���pH)�H��Ή�H��H9������H�������H�xH�|$(�x�@��	���9���  1��4D  H�zH�|$(�z��A���zD	�L�ZH����9��Z  L��H��H9�u��#���D)ۍH�H�qL9�����H�AH�D$(����QH�t$(��	��A�I����	���H9������H9������H��D�L$�   D�T$H)������A�D��H�H;M0�����L�}HU(H�L���ۉ���������H�T$8H��L���������y���D�T$�D$D�L$A��A	�H�D$8E��H�fA��H�D$0w!�   D��H��� ��  � ��  fA����  B�$�xG H�PD�L$D�T$D�D$I9������H�P�@�   H�t$(H�T$(H��L���D$������������D$��D�D$D)�D�T$D�L$ȉ�H��H�������   H�t$8L���D$萊���D$����H�D$0H��H9��  H�D$0A��D �}! �
  E����   E��E��D��H��H�t$0H��A���A���C ��H�UA���C �
�B�P�����у���9�s�H��H+D$09¸��C LD��A���C �I��1�H��L�\$(�Q���Q��	�H�yH�|$(�y���I��	���H9����������@ H��H�����D�L$1�H��H�t$0H���U���D�L$���M��������D�L$�   �Ҹ   ����1������}  t3H�MH�U�1�A�2H��B�}"�w�@����   @���$�G �   �r������B�Bf�B HcrH��H�������L�T$E��u�H�E H���   �x������/����E!L�T$�k����B�Bf�B 밃��B��f�B �B뜃��B��f�B �B뇃��B��f�B �B�o����   ������     AWL�~�   AVAUATUSH��I9��  D�6E��D�FA��E	�E��F��    M�L9���   H�WA��H���Bf�D$�Bf�D$�Bf�D$�B
f�D$
�Bf�D$�Bf�D$fE����   A�@�A�iL�t��	@ M9�t9A�7A�WI��E1�A��H�߉�A�w�A�O�D���	�D����������t�H�Sf�L$fD�|$f�J�L$fD�zf�Jf�L$
f�J
f�L$f�J�L$f�JH�K�q�	f�rf�
H��[]A\A]A^A_�1��D  AWI��AVAUATUSH��H��XL���   ���   H�T$0D���   H�L$���   �t$���   M����  H�\$0�Ɖ͋��   D���   9�N��A�D9�E�։t$���   DM�D)�A��D+��   ��D9�E��DN�9�M�A��9ǉ\$ ��A	�D9���A�u	D9��?  �\$ D+t$H�T$LI���   D����D)�F�$�    �ƉD$$A�������H��H�D$(�D$L����  H�T$0D�d$8E1�+��   ���   ��L���   ���   D��A�̉t$<+t$����Hc�H�H�H���tE�l$<H�l$0 ���   L��H��A����    �d���H��Hc��   H�I�D9��   wˋl$<H�\$0H�t$(H����N���L$ H��(  ���   D���   L���   ���   �L$���   �L$$���   �Hǃ�   stibH�\$���   ���   D���   �|$��  ��  �T$I��H  L��A�9A�qA�QE�IH�\$+D$��H���   H�H�\$�\$ )ˋL$8�D$8    ��Hc�H�I�E���Q  A��A������D$@�ǉD$ @�ƉD$$�D$(H�D$E1�E1����   ����   �    H�\$D��E�Ժ�   M�D�L$ A�jE�Z��D$A�ZL�A�<$L�M��u �E�;I��H��')�D������M��I��I��I��'��H��'A��D�H��'A�<$�|$$I��I����H��'H��'I��H��'�@�u �t$(��I��H��'��A��A���A�H�D$D9��   �)���H�\$�D$8Hc��   HD$H�D$0Hc��   IŋD$89��   �����1�H��X[]A\A]A^A_�A��P   u6I��(  H���%  A��@  A������r��   D��D��D������A��Q  A��R  A��S  E��T  �����L�t$0A���   ��L��A���   A��A���   �   A���   E���   ��AƆ�   H��fA���   �����D$L���/���I���   H��1��@���A���   H�T$A���   M���   �D$8A���   ���   �\$�D$ D���   ���   ����1�1�1��:���H�\$0�|$�t$ ���   �\$8�����A�����1�1�1����� AWAVAUATUH��SH��H��H��@  H���t  HcW8A�   H9�vu�4���8  ���D  ��vw���6  H��(  A�   �t�΍FH;��  w7L���   ��H��  L�����A�ą�u�   L���s���A�ą���  H��D��[]A\A]A^A_�fD  H��(  H�vH��H�T�B,f�E H���B-f�ED�JA��A��Ic�H�u�J��Hc�H�E D�R����   E����   H��H)�H��H����   H�E(�J�B�  @ E1��R����R  ��H�H�E0�1����R  �}�  @ H�E�v1��H�E�%���D  A�   ����D  ��<  A�   H9�����������fD  A	��]����B��D��8  ��A��Hc�Ic�H�uH�E �4���fD  I��A���?  L)�L�E(H�u �)���D  H��H�H��H�M ����fD  L�������L��A��赁��L��E���I���D��R  fD�} I��fD�}H���  L��L���0��H���  L��L��H�E�i0�����  L��L��H�E ���  )����  �Hc��>0�����  L��L��H�E(�(0����R  �} �  @ H�E0�0����R  �}�  @ H�E��/��H�E����D  L��H�E     H�����?  H�uH��������    H��1��L��fD  AWH��AVAUATUH���CLBCSH��H��(HǇ(      HǇ0      H�L$HǇ8      ��@  ���`  ǃ8     H�|$wN�   H��(   tL��(  L��H��D$�~���D$Hǃ0      ǃ8      H��([]A\A]A^A_ÐH����|��I�ŋ�8  ���g  ���n  ���U  �   H����}�����w���H�����H��A�����H��A���2���H��I���7��fE����  A���fA���0���I����  �#���H�D$J��   H9�vL�p�I��H���/|��H��H�p��s{���������B�4�   H��(  H��H��0  �}~���������D��<  ��8  �>   H�L$H��CLBEH����@  ��uǃ8     H�|$���������� H�L$H��colbH����@  ��t�H�L$H��xibsH����@  ���G���ǃ8     H�|$�,����u���D  L��(  H�t$H��L���}��������H��(  H�L$H��0  ��RȉƁ�  ���H��   t%��  =   t�   �����fD  ����  �,  ��H�@H��H��H9�sH���������H��H��H��H����<  ��8  Hǃ�      Hǃ�      ��u@H�D$L���  H���  H����   1��w����    Hǃ�      Hǃ�      ��t^H�L$H��TDBCH����@  ��t\H�L$H��TDBEH����@  ��tBH�L$H��tadbH����@  ��t(H���  �u���@ ǃ<      1�������    H����y��H���  H�D$H���  �9����   ����fD  �   �m���fD  U1�H��H��S�TLCPH��H����@  ��tH��[]�f�     H��H���  H���G []�v���fD  AWH��AVI��AUATUSH��H��(L�f8H��`  �emanH�L$��@  �D$��tH��([]A\A]A^A_��    H����x��I��8  ��G H��H�������D$��u�A��<  �I��L�lH�D$H�H��H�D$��   I9�w�fA��8  �6  L�L$E1�1Ҿ    L��跫��I��H  �D$���^���A��<  H�ߍ4@���y���D$���=���E��<  M��H  E���:  @ L����G H��D�$�D���D�$���D$uHA�Wf��t>A��@  H�IGI�GL9�r'H�H;D$wfA��8  ��  I�� f.�     A��u�M��H  E��<  M)�I��D��D��D�ʾ    L�L$L���ʪ��A��<  H��I��H  �4z��A��<  fA��0  �D$�V���@ L��H���v���D$���;���H�t$H���{��D���D$L��E��P  ������L�L$E1�1Ҿ   L���C���I��X  �D$�������A��P  H�ߍ4�    �x���D$�������B��   M��X  I�A��P  H�@I��H�$I9�sM@ L����G H��������D$A��@  H�IGI�GL9�rA�H�H;D$v1�fA�I��L9<$w�H���y��H�uH���u��A��<  �D$���� A�Gf���T���- �  A;�P  �P���I��X  H�@H��f�8 �)����2���1�M��1��G���fD  U1�H��H��S�tsopH��H����@  ��tH��[]�f�     H��H���  H��`G []�Ɓ��fD  AUH��1�ATI���pxamUSH��H����@  �Ņ�tH����[]A\A]�D  L���  �@G L��L���q����Ņ�u�Hǃ�      1�H���  ��  Hǃ�      Hǃ�      f���  ~�L�� G L���$�����u@f���  ?w�@   f���  f���  ��b��������1�f���  �O���f�     ���?���f�     U1�H��SH��H����H��@  H��tD�aehvH���  �Ѕ�u$H�ھ�
G H��蒀����uH�C(    H�C0    H��[]��    �aehh�Ѕ�u�H�Ð  �ff.�     �H���   H��0  H��8  H�D$H�H�D$8H�D$8H�4$H���|  H�D$8H��H9��j  H�D$8H��H�D$8H�D$8H�T$8�@��R���f	��>  H�D$8H��H�D$8H�D$8H�L$8�@������A�	����D$,�D$,����  H�D$8H��H9$��  H�|$�4f.�     �D$,���D$,�D$,����  H�D$8H��H9$��  H�D$8H�|$H��H�D$8H�D$8H�L$8�@������A�	�f�D$lH�D$8H��H�D$8H�D$8H�L$8�@������A�H�|$`�D$h    	�f�D$nH�D$8H��H�D$8H�D$8H�T$8H�L$8�@�H�t$8�R�����	��V�	��Q���	��%���H��8  ��H�V�H�t$H9��
���HD$H�D$@H�D$@H�L$@� �����A	����D$0H�D$H�G H�D$HH�8 u&�   �     H�D$HH��H�D$HH�D$HH�8 tdH�D$HH� H�D$PH�T$P�D$09BPu��D$4    H�$H�|$p1�H�t$@�7��H�D$H�|$p���  ��$�   �B�����t>��$�   ��tSH�D$H�9���f�     1�H���   �fD  �   H���   � H�D$PH�t$pH�|$@�PX�D$4��     H�t$@H�|$PH�L$XH�T$`�ש����u��T$4H�D$X�P �D  AWI��AVAUATUH��SH��   H��p  ���
  �A�E1�E1�   H��I�T ��H=spgiDD�I��L9�tI� H=fpgiu�I��A�   L9�u�I���   H�xh �Q  1�H��xibsL��A��@  A�   ����  H���   H���O  H��L���ЉD$D���;  E���D$A�    �/  1�H��CLBCL��A��@  1�H��L���D$�TDBCA��@  D�D$E���  ���  A��R  �P�   f���?��  H��L���SHH��L���D$D�S@H��L���D$D�S`H��L���D$D�SX�|$ �D$�D$D��   1�H��L���S8�D$D����  1�H��L�����   �D$D<���	  ���k  �   H��L���S8�D$D���/  �   H��L�����   �D$D���  AƇ�  H��L���SP�D$D��tA�����fE��h  H���   H��tH��L���ЉD$DH���   H��tH��L����H��L���D$D���   �D$DH��L�����   H��L���D$D�SxH��L��I�o(�D$D�SpI�G(    fA��h  ��D$DA���  I�G0    I�G ��  A���  ��  E���  H��   L��� ����D$D���A  E����  I�0 �9	  A��8  I�G�W���v
I���   t��@H��D�D$H��A��HD�H��H��E��uI���     t	H  H��I��   tH��A���   tH�� A��\  ��tH��@A���  ��  A��   I��(  H��H�H9��q  H���D  H�� H9��;  H�:fylgu�H�z t�H���fD  H�� H9��  H�:ravgu�H�z t�H��   ��  �    �D$ E1�H��L���S0�D$D�������H�Ĉ   []A\A]A^A_ÐE1�������     H��   L�������D$D��u�I�G(E��u	H����  H���	  I�o0�   L��H���I����D$D��u�A��I�G0u	H����  H���E���H��   L�������D$D���)����Q���@ A��   I��(  H��H�H9���  H���@ H�� H9�vH�8fylgu�H�x �j���H�� H9�w�H���D  H�� H9�vAH�8 FFCu�H�x t��9���f.�     �D$ ����H�y ����H�� H9��Z  H�92FFCu���<������I��  eurt��  I���   �D$D�   H�Ph��   H���f���H�H�z �X���E1��D$D    fE���  ����� H�x u!H�� H9�vH�82FFCu���<����������H��   I�wA���-  A���  H�Ѓ�H�H��H����HE�I	GL������A�OH���*  M�OP1�E1� I�<�   � 
G D�G�O��    H��H=�
G �0  �9�u�P���tA9�u݋@�G=cinut=bmysuA�   H��A9wH�E����  E��<  E���  I���   A��R  H�@8H�D$f���  fA��h  ��   A��D�fEE�j  E��H�|$E1�L�L$DL��1Ҿ    L�t$0����I�G@�D$D�������H�|$L�L$DE1�L��1Ҿ   ����H�D$8�D$D���������E1��D$,    H�D$    f�����D$$A�D$�L�d$HH�D$A�ŉD$(L��A��H���
�    I��L�m@L��L��H�����   �D$D��uzH�L$�t$HA��H��H��I�H�D$pH��fA�E �D$(��D$$�����fA�E��I�E�D$J��Hc�I�UI�U��t!��t�D$,H�|$8�D$,D�4�H�D$fD  I�FL9t$�Y���H�T$0L�D$8L�L$DI��H�L$H�|$�   軛���T$,��tNH��@  H�E�\$,H��H�E�]8�6�    �G    �����1�H��xibsL��A��@  ��A������I�G���  H��I�GI��x  fA��h  �I�GhI��z  I�GpI��|  I�GxI��~  I���   A��R  fA���   ��  A���  ���  A���  A���  fA���   fA��  )�fA���   fA���   H�  ����  I���   u;I���  �A  A���  A���  ��fA���   ���fA���   fA���   A���  A���   fA���   ��  A��  A��  fA���   A��   ��fA���   f���f��)�fA���   �   E1�E1��#���fA��h  ������A���  1�f����H��H���� HE�����L�d$H1�1��@G H�cinu  L��L�|$HH�D$P������t�Ѓ�t���   �]����D$D    ������*����D$D�?���H��   L��������D$D���#���I�( ���������fD  A�   �   �����A���  A���  fA���   fA��  )�fA���   fA���   ����H��   L���i����D$D�������I�G0�&���H��   L���D����D$D�����������I���   �D$D�   H�Ph��   H��������Z���I�W0�   L��������D$D�������8���A���   ����A���  A���  fA���   fA��  )�fA���   fA���   ����I�W0�|���H��   L�������D$D�������I�G(�����D$D    E1��K���f�     AWH�GAVI��AUI��ATUSH��(H�VHH9��-  A�E����A�E	�I�VHD��K�L% H�L$H9�w^f=vXI�]E1�I��  �D  ����A9�DB�L9�tAH���C������C�	�A�vP���vШt̾   L����)��뽾   L����)���F�,�   J�+H��H�D$I�FHH9���  E1��A��L���C�sL�k��f	���   ���CA�vPD�[D�C�D$�C�$��vF�3���s��	�f��� w���   )�9�s#�   L��D�D$D�\$�C)��D�D$D�\$D����fD	�t2��I�t5�H9t$w�|- H�H9t$s�	   L���)��A�vP��uA�GE9��,���H��(1�[]A\A]A^A_�D�D- M�M9�s��l$�$��	�L������     I9�vCH���E������E�f	�t����A9FXwھ   L��L�$�T$�u(��L�$�T$I9�w�H������H)�I�I��O�lE�U����   L���A(��������   L���/(���e���f.�     AWH�GI��AVI��AUATUSH��xH�VHH9��#  A�_I�VH��A�_��	�����L�H9�sA�FP����  I�^HD)����|  A�G����A�G	�A�VP��A��A���v���  B��   9���  A�FP��v^A�GE�oE�O
E�G����A�G		�D��E�o����A	�D	���  ����D9�w���D9��  �   L���'����%��  I�TH�T$H�H�,H�T$H�H�D$XA�FP��v'A��$����I�L������A	�f����m  E���,  A�D$�E1�E1�E1ۉD$dI��L��H�D$0���D$`    H�D$hL�|$��   fD  E��E9�w(E��t#�rP����  E9��  D9��v  �L$`����@  ����  �4  �JP��LÅ��k  H9\$Xw��H�t$Ht$hD)�L	H�H9�vH�׾   �D$@H�T$8��%��H�T$8�D$@�JP���_  I�L$E��A��I��L9d$0�>  I��H�D$H�|$I�h�]��M�F�4`F�|`H�D$B�4g��A��	�E	�F�|`B�D`��@�t$ B�tgE��A��A	�@�t$(A��A9������H�׾   D�T$TL�D$HD�\$P�L$D�D$@H�T$8�,%��D�T$TL�D$HD�\$P�L$D�D$@H�T$8���� f��������JP��wD;L$d�+  H�׾   �D$(H�T$ ��$���D$(H�T$ ������    D;L$d�E  H9\$X�������H�rHD)�L	H�H9�������JP�������fD  A9�������H�D�|$ �D$ D)�L�tK�L$(A��H�l$(L��H��I��A	�E��D��I���	@ M9�t;I��A�F�����A�F�f	�t����9EXwپ   H���$��M9�u��    H��D$ H�l$(�����    �L$`����fD  H�׾   L�D$H�L$D�D$@H�T$8D�d$P�#��H�T$8�D$@�L$DD�L$PL�D$H�@����D$`    �D$`H��x[]A\A]A^A_�D  E!�fA����x�������D  �   L���K#������fD  �   L���3#��A�G����A�G	�A�VP��A��A���v �t�   L����"���i���f.�     �   L����"���]���fD  �   L����"�������fD  E!�fA�������������D  E��A��A�D D9��l���D��A����	��   ��9��Q����Y��� �   L���L$D�D$D�L$�U"���L$D�D$D�L$����D9��������� �   L���#"��I�^HD)��R����    AVAUATI��UH��SH�FHH�_
H9���   A�D$E�l$H�MH����A�D$	�D��E�l$	��A	���L�E��H9�rfC�T6
��9�wZ�EP��tEfE��t?A�F�M�dD�f�L9�t-H���C������C�	���9EXw�   H���c!��L9�u�[1�]A\A]A^� �   H���C!��뗐�   H���3!���=���ff.�      AWL��   AVAUI��ATUSH��H��H�FHL9��H  I�UH�CH)��9��<  =   �1  I�UH��   �����H�kL)�ȉǉD$������9��  �T$���$  �$    1�A��   �A�A�GI��E�O���A��9��"  �$��t9�w�   L��D�L$�U ��D�L$A�UP����   D��A�UX)�9�r�A�D)�D9�w�   L��L$� ���L$����  ����   ��u*�p�ډ��������  �t D������tz�SA9�tJ�Ӊډ������t ��D������u��   L������fD  �   L���������fD  �$D��$9D$�����H��1�[]A\A]A^A_� �   L���[���t���fD  �   L��T$D�L$�:���T$D�L$����@ A��  ��uO��u�f�     �SA9��t����Ӊډ��������  �t D������tԾ   L��������D  �   L��L$����L$�f�     �   L���������fD  �   L����������fD  AVAUI��ATI��USH�FHH�_H9���   A�EI�T$HE�u�L)��A�D��H9�rH��vH��H��H9�s�   L���#��A�D$P��tE��u([1�]A\A]A^�f.�     �   L������H��t�H���C������C�	���A9D$Xw���fD  �   L������U���fD  AWAVI��AUATL�gUH��SH��(H�FHL9��3  �E�]I�VH�ˉ���H)�H�$H9�r H��vH���������H��H��H��H9�s�   L���@������   1�E1��l�M��t$I9�w�   L��L�D$�D$���L�D$�D$A�VP��t-��A�VX)�9�r
��)�9�r�   L��L�D$����L�D$I��L��L9,$tUA�$A�l$I��A�D$���A��A��M9��p����   L��H�T$L�D$�D$���H�T$L�D$�D$�B���f�H��(1�[]A\A]A^A_��    �   L���K������fD  AWI��AVAUL�oATUH��SH��H�FHL9���   �E�]I�WH�ˉ���H)�H�$H9�r H��vH���������H��H��H��H9�s�   L����������   1�E1��8�M��tH9�w�   L�����A�WP��tD���A;GXsFI��H��L94$tSA�m A�]I��E�e��ˉ��H9�v��   L��H�T$�Z��H�T$� �   L��I���?��H��L94$u�H��1�[]A\A]A^A_�D  �   L����������ff.�      AWL�
AVAUATUSH��H��HH�FHH�|$(L9���  H�|$(H�CHD�w�oH)�A�D���A��H�t$H9�r"H��	vH�V�H���.�袋.H��H��H��L9�s�   H��������  H�D$   K��I�DD
HD$(H�D$ �*@ I�D$H�D$E����   ���`  L9|$ ��  E�'A�GI��H�L$��A��A	�A�G�A	�A�G�A�o���A�ŉ�M��H�D$L9��,  H9��#  L;d$s��   H������I�D$H�D$E���w���Ll$(H�CHM�uI9���  H�CHE�e L)�A�D��H��H�<$H9��T  H�<$ �4���E1�L�|$0E1��l$<M��L���f�M9�rRM�}I��L94$v_F�d�B�D�A����A	�B�D�A	�B�D�N�, I���� v��   H�����M9�s��   H��M�}I������L94$w��l$<L�|$0�������L�l$H�CHLl$(M�eI9��z  H�SHA�m H���������L)�͉�H��H�4$H��H9��5  H�<$ �M���E1�L�|$0E1�M���Ef.�     L9���   �CPL�z��tA��@��A	�E��D;kX��   I��L94$��   A�$A�T$I������	�A�T$�E�l$�A�l$�	Љ�=�� v��   H��H�T$����H�T$L9��z����   H��H�T$����H�T$�^���D  �   H����������fD  �   H��I�����L94$�X���D  L�|$0L9|$ �F���H��H1�[]A\A]A^A_��    �   H���S�������fD  �   H���;���t���fD  �   H���#������fD  �   H������`���fD  �   H����������ff.�      H��tKM��tF��   H��t,D�ȸ�   A9�v1��H��H�(  H�H�H�FH�H�FI� 1���     �   �f.�     �=��  w'�G u;G(t$�   ���f��   ��|��fD  1��D  UH��SH���K{���C,��t�S(�U []�ff.�     �( t�H9G0t�   �8����     UH��S����1��( t
H�W0�G8�U []Ð�( t�H9G0t�   �����     UH��S�v���1��( t
H�W0�G8�U []ÐUH��H��H��8  S�pamcH��H����@  ��tH��[]�@ H��8  H��0  H����Q����t�Hǃ8      H��[]�@ AW�tsopAVAUATUSH��H��XH���   H�L$HH����@  A�ǅ�tH��XD��[]A\A]A^A_�@ H����N���    H��L�l$HI��L���  �tN��A�ǅ�u�I��   t$A�   I�� P �a  ƃ�  ��     H�t$DH��L�u8��R��D�|$Df�D$E��u�A�   f;��  w�D��E1�L�L$D1�L���   L��蓁��D�D$DH�D$E����  K�4?H���tO��A�ǉD$D����  �D$f���6  H�t$��L�d$ H�\$0H�DFH�t$(H��H�D$I��H��H���Q��f�C�L9�u�H�T$(H��L�d$ H�\$0H�T$ �P��H�T$ H�|$1� �
�ȁ�  ~D�Ɓ�  f-D9�O�H��H9�u�f�t$��L��L�L$DE1�1Ҿ   觀���|$DH�D$ ���  f�|$ ��  K�,D�|$<E1�I��H�\$0H���   fD  H��D$(�M��H��L)�H9���   D�l$(A�ML�L$DE1�1Ҿ   L���,����L$DK�����  E��H��H��L���[M���D$D����  K��I��B�( fD9d$��  H��E���L��H9��2  H�t$DH���uP���t$D���V  D��L9��D���H��A���aL��A)Ÿ    DH��I���H�t$DH��L�m8�P��D�|$DA��E���}���A�   f;��  �j���D��A�F�=  �W���E��L�L$DE1�1�L�Ѿ   L��L�T$�%��H���D$D��utL�T$H��H��H�L$L��L�T$�ML��H�L$��A�ǉD$DuGE���0  H�L�T$I9�|(H��x#�   @ A9��  H�H�H��I9�s��D$D   H��L������D�|$D�����H�D$     H�t$ L���ʥ��H�t$L��轥��D�|$D�r���H�\$0�D$H�T$ ��H����L�d�fD  H�u L��H��耥��H�E�    L9�u��H���M��E1�1�1�L�L$D�   L��� ~���|$D H�D$ �i���f�D$  �D$f��   �D$f��  H�D$H��  H�D$ H��  �����fD��   H��  ����H�D$0L��D�d$D�|$<H�D$(A��1�L�L$DE1��   �   L��H�\� �c}���T$DH���u1A���  fE9�r�H�l$ H�\$(fD�d$�M���D�|$<H�\$0�>���H�l$ H�\$(fD�d$����f�AUATUSH��L��x  M���  H��H��A��1�A�T$ H�E H���  H=   tkH=   tH= P �   H��1�[]A\A]�f����   ��   ��   A9�s�H��  D���<pf��vlH��  H�������H�E �D  A��  w�D��A�T$ H�E H��1�[]A\A]�fD  ���   tg��   A9��h���H��  D���<D�A�T$ H�E H��1�[]A\A]�H���x������M����,��� H���   []A\A]��     H���H�����t�� ���ff.�     @ H��t���  9�v���� �   �f��#   �f.�     AUATUSH��H�G H��xT�����H9�~cA�����I��H��1�D  ���  9�v$H�T$��H���&�����uH�t$L��������t
��D9�r�1�H����[]A\A]�f.�     A��H��u���fD  H��H�D$    H��t&���  1�9�sH�T$����H�D$H���D  1�H��ÐATUSH��H��tS���  A�   9�sH��H�T$���s���A�ą�tH��D��[]A\�H�t$��H��葢��H��D��[]A\�D  H��A�#   D��[]A\�ff.�      AWAVAUI��H��ATUSH��H��XL�v8��F��H�t$H��H�D$(�P��H�D$�D$��tH��X[]A\A]A^A_�f�H�T$��G H���R���D$��u�H�D$H=OTTO�]  �L$ I��fE��   E1�1�L��I��  L�L$�    �y��I��(  �D$��u�H�D$(H��H�p�wE���D$���j����t$ H��H���JG���D$���M����l$ f����  1�E1��3f�     I��xtmh�s  I��xtmv�f  A��fD9|$ �f  H���^I��H��I���SI��H��H�$�GI��H��I���<I��H�SI9�w�L)�H9�w�I��(  f��t-L;7t��M�H����H��H���     H�� L;2t�H9�u���H�$��H��H�L�7H�OL�gH�G�W���D  H�D$(H��H��H��H�$�PD���D$���C���f�|$  �x  E1��D$    1�E1��D$    �4fD  H��GNIS��   H��ATEM�   DD� ��f;l$ ��   H�T$0��G H���P���D$����   H�t$@H�CH9�w�H�L$HH)�H�T$0H9�vH��xtmht	H��xtmvu�A��H��daehtH��dehb�h���H��5��   H��H���jC���D$���]���H�t$H���QM���D$���D�����H�߃���Hc�H4$�-C���D$��� ����D$   ����@ �D$   ���� ��f�l$ fE��t2�D$��u��   D�|$������D$    H�D$A������@ �   ����fD  H�Ѓ�������D  fA��   H��� F���D$������   �|���ff.�     f�UH��1�H��SH��H��H����@  ��t
H��[]� H��H��0  H��@G []�O��ff.�      �dehb�f�     �daeh�f�     AUH��1�ATI���2/SOUSH��H����@  �Ņ�tH����[]A\A]�D  L��h  ��G L��L���N���Ņ�uѸ����f��h   Hǃ�      Hǃ�      Hǃ�      ǃ�      f���  t�L�꾀G L���:N����uNf��h  �n���L��`G L���N����u,f��h  �L���H��L��L��PG []A\A]��M��@ ���'����AWI��AVAUI��ATUSH���   H���   L��p  �T$@H�_M����  �   �׷F �+'��I���   I��x  ��  I���   �P  I�G8L�t$Iǅ�       H�D$Iǅ       Iǅ      f�     L���A��H�t$XL��H���HJ��H�D$X����  H��FFOw�d  H��L���!@���D$X����  H�T$h��	G L��I�_8�D$\    ��L���D$\����  H�D$pH=FFOw�j  H=fctt�^  H�D$xI;G�O  ��$�   f���>  H��H��,   H9��)  H��H��$�   H��H9��  ��H�l$�  H��$�    H��$�   �  H�$�   ��   H��$�    uH��$�    ��   H�T$\H����S��H�ŋD$\����   H�$    E1�E1�L��H���>���H�4$H���2���D�\$\E����  �D$X    @ M���   �l���@ L�t$H��   �&  Iǅ�   fcttH��fctt�i  I���   ��	G L���jK���D$X��uI��  H���r  f��   H���   []A\A]A^A_�f�     H�������H��$�    �������fD  H�T$\�P   H���R��I�ƋD$\���/  ��$�   �Ѕ���  1��f�     ����qu��   ����A��A����H�t$p��)�H��f��@�u H�t$pH��@�uH�t$pH��@�uH�t$p@�u��$�   @�u��$�   D�ML�L$\@�u�0   D�EE1�@�}H��f�U
1҈M	��$�   �Aq��H�$    I�ËD$\���1�����$�   E1�1�H��L�L$\�   L�\$ �q��D�d$\L�\$ H�$E���������$�   L��H�4�H����>��L�\$ ���D$\�����1�M��f��$�    ��  H�\$ H�\$H�l$(H�,$L�l$0I��L�\$�!H����$�   N�d� I��I��0D9��O  L����@��L��I�$��@��L��I�D$�@��L��I�D$�@��L��I�D$�@��I�D$ I�$H9�w�L��H�\$ H�l$(L�l$0�?���D$\   L�\$����D  H��H���=���L����;��L��H���*����D$\�D$X�������j���D  ���F H���"��I��H���w  I��p  H� I���   I��@  �����f.�     H��fctt�����H��OTTOt:H��eurtt1H��1pytt(�dbk�H9�tH H9�t�   H��   ������Iǅ�   fcttH�|$H�T$X�   Iǅ      Iǅ     �O��H��I��  �D$X�������H��D$`    f.�     �\$@I��  ��A����A1�A)�A�ǅ��[  Hcи   H9��?���H��    I��  I���   H�4H���:���D$`������H��L��A���   �D$`�������A��H�L$hH��L��M���   D�<$�ravfA��@  ��uH�|$h�  1�A���  E1�E1�f�|$1ɨ�?  E1�E1�1�L��L���<���L��L���1���1�H�ھfylgL��A��@  ��t91�H�ھ2FFCL��A��@  ��t!1�H�ھ FFCL��A��@  ���]  D  ��9$��   �D$@1���6  I��  I�mI�E HcD$@I�E�D$`�����D  ��H�H9���	  1����� ���F H�����1Ҿ��F H�����I���  �������F H������1Ҿ��F H���t��I���  �R����     ��H���^���@ H�$    E1������A��1�D$H�D$`H�D$�D$H�T$L��E1�D�L$(��H�L$ H�H��H�D$0�1M���t$`I�ǅ��{���H�T$H�t$0L���M���L$`D�L$(I�ƅ�H�L$ �P���H��D�L$ H�L$��8��H�L$�T$D�L$ Hȅ�H�D$L�X�t|�D$M��A��f�l$ fD�L$FH�̓�L�|$(I�D�L�d$8M��L�l$HI��M��fD  L��L��   H���8��I��I�D$`M9�u��l$ L�|$(L�d$8D�L$FL�l$HE��D�L$H�L$E1�Ic�L�L��ŉD$�D$H�D$f����  f�l$H�l$0L�d$ M��L�l$(E��� Ld$A��D9l$�n  L��L��H��H����7��H��L��L���D$`聡����u��l$L�d$ L�l$(����f�     I�GH��H9��  H�|$L�L$XE1�1Ҿ   ��j��I��  �D$X���X���I��  L��H�4�    �8���D$X���5���1�I��   ~(@ I��  L��H�,�H����:��H�E I9�  �L����9���D$X�D$`���t���������    1�1������    �����A�   E1ɸ   ���J���fD  H�D$`H��H��H�D$�@��D�T$`I��E�������H�t$H���;��D�L$`��E��������   H��H�L$�6��H�L$���D$`�����H�t$H��H�L$�:��D�D$`H�L$A��E���\���H�t$H��H�L$�:���|$` H�L$A���7���H�t$H��D�L$H�L$�m:���|$` H�L$��D�L$�	���H�t$H��D�L$ H�L$�?:���|$` H�L$f�D$D�L$ A���  tf�D$  E1�E1�1������fD  I��   �����fA�������A�V�f���?weA���t$��   �|$9�t��9������f���~w;�|$��������Hc�H�Hc�H�H;T$hw��A�   A���  ���� A�   �>���D  �   �����fD  �   �����fD  H�\$ H�l$(L�\$L�l$0L��L�\$ �7��H�<$�p�C ��$�   �   �t�����$�   L�\$ I��H��H�L$(H��H��fE��H��,   H�L$��  H�<$H�7H�~H9���   H�FL�d$xL9���   L��H)�H9���   H�VL��$�   L9���   L�$A��L�|$ I�HO�L�M��I��H�L$�S�    H9�rSH��H��H�N(������H�H�M9�tgI�0H9~u-H�FI9�r$L��H)�H9�wH�VI��L9�wM��I)�I9�s���D$\   ����� �
   �k����l$L�d$ L�l$(������H�L$L�|$ H��$�   H��tH9�u�H�$�   H;|$xw�H��$�   H��t"H�W���H9�u�H�$�   H��H;D$x�u���H�D$H9�$�   �b���H9|$x�W���H�T$(H�L$I��H��L�L$\�   L�\$ H��H���f���|$\ L�\$ H�������f��$�    L�`�D$(    ��  L�\$L�l$ M��M��I�$I��L��H��A�E�I�$H��A�E�I�$H��A�E�I�$A�E�I�D$ H��A�E�I�D$ H��A�E�I�D$ H��A�E�I�D$ A�E�I�D$(H��A�E�I�D$(H��A�E�I�D$(H��A�E�I�D$(A�E�I�D$H��A�E�I�D$H��A�E�I�D$H��A�E�I�D$A�E�I�t$�1���D$\���(  I�t$L����2���D$\���  I�|$(M�D$I�D$I�O@H�I9���   H��H�T$`H��H�D$`�7W �D$\����   H�D$`I9D$��   L���4��I�D$ID$(�tD  �D  H���u�D$(��$�   I��0�L$(9��y���L�\$L�l$ H��$�   H��L��L�\$��/��I�G8I�uI�F0 D I���   I�F8H��
�������M���   L�\$I�e���������L��H���y����I���H���'���L�\$L�l$ �����L�\$L�l$ �����H������D  ATH�GI��UH��SH�VHH9���   A�D$H�MH����A�D$	���L�H9�rSf=vM�EP��t:I�\$I��  ��     L9�tH���C�;EXr�   H�������L9�u�[1�]A\�D  �   H�������뤾   H�������j���ff.�     @ AWAVAUATUSH��x��8  ����  H��A�Ճ��  ����  H��@  ��H��$�   �     H��(  D�t�A�D;o �U  H���  E��L9��`  B��   L)�H9��L  �D$   M��H���  A��L��I�tL��>.���Ņ��9  �   L���0���Ņ��"  L���u2��L��I���j2��L��H���o1��A9��  ��   A��E)�A����   H���  ��L)�H9���   H���  E��L��L�L��-���Ņ���   D��L���/���Ņ���   L���\1��L���T1��L����1��= gpjte��   =epud��   �l$�  L���!1��L��D���0��D;k �  H���  L9�vL)�B��   H9������ �   ��L���x0���     �   H��x��[]A\A]A^A_�f.�     =lbgrt�=ffitt½   L���50���� H���   ��   t�H��@  L���   A��M�ϋ�H���  L��D$�,���Ņ�u�H���   L�d$ D�d$H�\$H���   H��$�   H�D$(1�f�D$8H���  H�L$0H��(  H�D$@H���  H�L$`H�D$HH��0  H�H�T$hK�dH��H�r7H9������H�t�ʉ�H�T$P�Nɉ�H�L$X�v.@�t$:H9������H)�H��H9������E��E1�1�1�A��D��H�|$A���՝���Ņ������A��  P �����A������H���   H�|$L� �� �   H�T$L��L���: �Ņ�t,H�t$L���� �G���f��   �i����   �1���@ �D$2H�t$(A�G�D$ H���   A�G�D$0fA�G�L���H���   H��(  �H�������   �����ff.�     AWI��AVAUATE1�UH��SH��H��(�BH�t$H�T$H�pH�<$�D$    �3?���T$����   H�sL��I���x*���D$��uY�sL���T,���D$��uE�CM�w@��t��M��M�l� A�I��I��A�G�M9�tcA�>�Յ�u�H�|$�-��L�4$L��E1�L���E���1�H�sL��H�C    f�C�+���H�C    H��(L��[]A\A]A^A_�M��fD  A�E  H�|$�)-�����    AWI��AVAUE1�ATUH��SH��H��(H�t$�rH�T$H�<$f���D$    �����>���T$����   H�sL��I���S)���D$��ul�sL���/+���D$��uX�CM�w@f������   A�> u4�A�M��M�d�A�FI��I��A�G�M9�tjA�> uA�~�Յ�u�H�|$�O,��L�4$L��E1�L������1�H�sL��f�CH�C    ����H�C    H��(L��[]A\A]A^A_�M��fD  A�$ H�|$��+����ff.�     @ AWAVAUATUSH��HL���  M��tH��HL��[]A\A]A^A_�@ H���   H��tH�G  ���   �G���   H�L$0H�T$(�   H���dN����t��D$(���uG�D$0���t/Hc�H��`  �p�C H���   H��H��H�H  H�������I��L���  �]��� Hc�H��`  �p�C H���   H��H��H�H  H�������H��u��D  H���   L���   H���  ��  H�T$L�D$ 1�H��H�t$�SPH�EH�T$ �  ��!  �E��  H��L��p  %�  H�X�H�BI��$   H��H؋pH�D$(    �� ������~  ��  ����  H�T$0H���p��H�|$0H�T$ H����   賑�����  L����H�tH�T$�8;���L$I�ą������H���  H��躏�����  L�� -H�L$0H�p���t/fD  �Ѓ�0��	v��߃�A��w�H��H�����u�� H�^H�t$0L��M���X����:   �D$L�bL�������tH�T$��  �:���T$���!���H���  H���������  I��HËD$����  H�D$1�H�|$0A������    I�L$H9��  �_H�D$H�A�ʅ���   L�[y�C-��L�[A����E����  H��f�     ��H��A�������)��A0�шC���u�H9���  L��H����B�H��H���A�H9�u�H)�L�E��tQ�.C��L�[�D L�S��I�K��A�Ճ�0�Q�%��  ��  ���L9��  I����fD  �C0H��I�D$ H��H���� t#�ʃ�0��	v�у�߃�A��w�I�D$ H��H��H���� t#�ʃ�0��	v�у�߃�A��w�I�D$ H��H��H���� t#�ʃ�0��	v�у�߃�A��w�I�D$ H����< t�Ѓ�0��	�9  ��߃�A<�+  H�D$H����I��0H�D$;t$�<���M��L)�H�������ۍCI���A����A����Mc�M���K  ��    ��Hc�A��[H�Hcɿ�[��[H��I��A��[M�L f�i��#H��iQ��J�8��i������iғ��1�iA����D1����������VD�i��J�81�iA������D�D���5͖�����G��i���#D1����D���;�2I9��v���H�؃��$�	G f�     �H��H�D$�����L��H)�H��t4��0��  L���	fD  H��H�C��@ �{�0t������f.�     =�B ŀ�1��  = � ��  ��t�A�U/�S��    ��H�T$(H����L�|$(M����  L��M���*���I�\�G���1�A�@1�i������i���#A1�A�P����A�P
��1�A�@	��1�A�@1�i��J�8��i����A1�A�P����A�P��1�A�@��1�A�@1�i������i��J�81�A�P����A�P��1�A�@��1�A� 1�i���#��i����1�1�1�A1�D1ۍ>D���Aʉ�ˉ�����1�1�i�k��i�k�녉ȉ�����1�1�i�5���D����i�5���A1�Ai�k�녉ȉ�����A��1�A��D1�i�5�����1׉���1��>1��i�k��A��A��D1�i�5���A��A��D1�L�D$0�ƉD$0���t$4���  I�x�D$8L�T$<H���F�-�F	... H�F�     ��H��������`G �HH9�u�H��L9������H�����1�����1�����1�����1��`���1��c���1�A�@��1������1��U���1�����1������1������A�P����fD  L��I��H)�H��������1�  ��0����A�U/A�R������fD  L������H�L$H�T$�   H����E������   HcD$���tgH��H��`  ���C H�H  H���   H������I��H��t9L���A�����[vA�D$[ �[   L���  ���  �����D  L���`���HcD$����C���H��H��`  ���C H�H  H���   H������I��H��u������    =� ����������     A�B�0�����fD  H�L$H�T$�   H����D����� ���H�L$H�T$�   H����D��������������A��[A��[��[��[�\���H�D$ I��$   HXH���P���f�     AWAVAUATUS�H�|$����g  ��  �C�L�~I��H�@M��L��L�\�0�    H�M H�E�H��� H��H9~7L�H�zH��L�J L�RL�PL�R L�PL�R(H�xH�x�H�L�HH9�u�H��I9�u�L�&D�k�1�   ��     D9���   D��D9�v��D�OH�@H��L)�L9�~�9���   A��K�RH�Ɖ����L�H�@I��1� HH�    H��H9�u��H�H��K�RH��D9�s�D��D��D��H�@L�$�D9�w� �    I�8 t#��I���H�@H��H�I�HH�HI�HH�HI��M9�u�H�D$��[]A\A]A^A_�@ �GD��A��9��>���1�A���o����   ��ff.�      H��t
H��@;  H�H��t
H���  H�Ð��AWHi��	  AVAUHi�P9  ATL�4USIcFXH�<M�N`LcPH��H�P�����L�|$�I�����fHH�\$�����I��H�H�� �  �    H��H�H�� HN�H�T$�I9��  ���  H��   H�t$��D$��H��H��    H)�L�$֐�T$�H�D$�E1�L�l$����   �    �P0I������   A�IA;Nh�����8�tzI�1H�H�hH��I��H)�I)�H��L��H��?H��?I��I1�I)�H��L1�H)�I9�~
L�XL��H��H)�H��HH�Hc�H�T$�H��H��?H��
 �  H��Hc�L9�}I��M��H��8L9��U���M��tM�y(I��XL9L$�����[]A\A]A^A_�f�H�FP�N4H��   �V0H�GH�FXD�B�A�щ�  H�GH���9  H�GH���9  H�G 1�A����A���A���uE��A��uBA��A����AD�H�V@H���  �ʃ��~  t���ʉ�  1���  �@ A��t̃��ff.�     f���t\�F�L�GA�b   H�@L�T� H�� I�0H��H��H)�H)�HH�L9�}H��I��I��M9�u�H�H H���H9�~H��/H9�HO��H�J H��H���H��/H9�HL��f�     �F4H��   ��  H�FH�GH�FH�GH�F H�GH�F(H�G 1��ff.�     f�����ff.�     ����ff.�     H��t
H�� K  H�H��t
H���  H�Ð��AWHi��	  AVAUE1�ATH�USL�@PHc@HL��I��M�t�F�H�@L�,�H��   �hH�   I��I��LD�Hi�p  H��M9��/  Hi��	  L��I��)g>îH��D  H��PI9���   D�^D;[hu�H�~L���fD  H��PI9�v��QH�AD�u�H9�}�D�I�QfD9NfDNNf9VfMVM��H��I)�M9��H)�I��M��t<H��
A� }  H�I��H-   H='  E1�H��~H��I��H��I��f�     H��H�I��L�H9F0~H�F0H�N H9A0�M���H�A0H�q �@���I�@ H��tL9@ tI�@     H�@ I�@(I��PM9�w�[]A\A]A^A_�ff.�     f�H�VPL�VH��   �F4�N0H�WH�VXD�A�A�ɉ�  H�WH���I  H�WH���I  H�W 1�A����A���A���uI��A��t`����tFA��t
A�Bt ��H�N@H���  �y  u����  1���  �f�A��t҃���u���A�Bt��fD  ��u�����fD  H�T      H�G<	  H�G�   f�G H��  �  H�G$H��    H�G,H�  H�G41���     �ff.�     @ AWAVAUATUSH��   H�D$�L��$�   f��     H��I9�u�L�_0H�_ I)�L�W(H�GN�,L��L)�M9�L�_8A��HL�K�,M��M)�L9�MO�)�A)�D9�A��A��@A��E��  ���  �L$�)���$�   A�݉L$�A)ͅ��  H��$�   Mc�Lc�Hc�H��$�   H�h��$�   ��H��H��L�tRD  H�E D�]H�T$�I��H��H��?L�� �  �EI��I�A)�H��M�I)��    I� ��?���G A��T��H��A9�}�H��PH�T$�I9�u�HcD$�D+d$�E�H)��f�     tCH��A9�|(�D��A�9Gh}�GhH�H���OlH�wXH�G`A9�}�H�Ĩ   []A\A]A^A_�9Ol~���Hc��ff.�     @ AWAVI��AUATUSH��H��XH�GL�g�G,    L�o�D$L    H�D$H�G H�/�G<    H�D$��GH    �GX    Ǉ0
      Ǉ@
      ���?  H�@ ��  A�F�P����`��  H�{0 ��  �C,A�L���Ch   �C<ǃP
  ����������u�Ch����ǃP
     H�D$L�cL�kH�CH�D$Hǃ(      H�C HcC,Hǃ0      ���u  L�{0H��M�FH��M�^M�NI�H��   M�H�$H�@K�<�L�\$H�����   L�����	�D$4I9��  1ɉ�L�D$ L��L�D$L�|$(Mc�Mc�L�t$H��A��L�t$H�\$8�y��������f��N�P�^)�Hc�H��H��?H1�H)��H)�Hc�H��H��?H1�H)�H�H9�}f� H�pHH�F@H��H9���  H��PI��I��H9$��  �@�@I�I�Sf�HHc�I��f�PHc�I��H��H��?H�� �  H��Hc�L�H�H H�HH��H��?H��
 �  H��Hc�L�H�P(H�PL��H��HT$H�
H�Rf�Of�WA���������   f�������W89������L�G@H��8  I9��c  ��L�L$L�   H������I���@E��H�C@�D$L����   A�FD�{8�P����`�|����s(9��|���L�C0H��x  I9��  ����L�L$L�P   ���H��A����D��H�C0�D$L��u-D�{(A�F�1���H�S@HcC<�l$4H��I��H��H9�ww�D$LH��X[]A\A]A^A_�H�\$A��H���D9��O���H�\$ Ic�L�SK�<�H��H|$(H���-���H�\$8L�D$ L�|$(H�S@HcC<H��I��H��H9��A  1�H��@ H��H��I��H��H��L�H�B�A�@���H9�r؋D$4L�|$I���������I��D�d �Mc�f�I�H�KHD�A�yH9���   �sD�K��)�H�H�H1�H)�D��D)�Hc�I��I��?L1�L)�H�I9�J�\  D  D�N��D�VD)�H�H�H1�H)�D��D)�Hc�I��I��?L1�L)�H�L9�}H��E��D��H�qHH9�u�H�A0    H��H��1�H�A8    E1�A����    f�
H9���   D�BD�RH�R@�zD)�Hc�I��zD)�M��Hc�I��?H�L��I��L1�I��?L)�M��I1�M)�N�I9�|�I��I)�I��M��L�P0I��L�R8M��I��I9���  A�   L9�}L��L��A�����L��    �   I)�L��H�H9�DM�D�HH�@@D��H9�tfD  @�p@�pH�@@H9�u�@�rH��E1�H)�H��I��H�p0H��H�q81�H9�����I��M9�����L�|$L;<$�H���L��H�4$I����������D  H��PH9���   ���u�f�xu�H�x8H�H0�XH�<�H��H��H����L�8L�E�CD)�E�BA)�D1�x��XE�C��D)�E�BA)�D1�x���H)�H��Pf�P�H��H��I��I�S0H��I�R8H9��m���H���������H�$�%A�WA�O8�t[�tfD  I��PL9��[���A��u�tσ�fA���fD  L9�}H��A������Z���D  L��L��A�   �D�����u�I�G0A�wL�$�I�G8I��L��O�,'A�GI��A�MA�UO�4L�$A�~)�)�Hc�Hc�)�A�~Hc�)�Hc������L�$���C���L��L)�H��H��I�F0H��I�E8A��:���H��E�ȉ������H��8  �G8   H�G@A�F�P����`������]���H�G@    E1�����H�C0    E1������H��x  �C(`   H�S0�1��� AWI����$I�AVAUATUSH��  H�H��$�   H�G@H��H��$�   Ic@<H��H��$�   I��   �PH�����
   ����H��$�   H��H�D$h1��H���HǄ$�    }  H��$�   Hi��	  L��Ph�xh�@H    I�@0��1�)�IcP,�|$PH��H��H���  H9�v!fD  H�HH��PH�H�H�H�H�H�H9�r�H��$�   H9�$�   ��  Hi�$�   �	  L�D$XE1�I�| pH�D$`H�|$x�|$P�|$H��$�   H� H�PHH�D$�B����1�)�;D$P�  E1��D$ 1�1�H�D$H ���H�\$H�� ���E1�H�D$@ }  E1�1�A� }  H�D$8 ���H��� }  H�D$0 }  H�D$( ���H�D$  }  fD�L$f�L$V� }  f�t$TH��D  H9\$t<��uLD�cE��E��A��E��E1�E)�D;L$P�:  H9[H�0  H�[@H9\$uĀ|$ ��  �D$��t�H�[@L�K0D�L9�IO�L9�IL�L�K8L9�~E��L��L9�}	fD�T$L��A��uM9�MO�L9�IL�D�KD;L$u�   H9\$�B���M��tM�OHM9K@��  L�I�[HI��fE�KI��I)�I��fE�KD�L$E	�A��tI��M)�L;L$h}A�D�|$A��fA�K1�A)�fA�sfE�K
fD�|$VM��E1�H�|$HL�D$@fD�t$TH�t$8H�L$0H�T$(H�D$ �����    Ǆ$�       H�L$XHL$`HcAH����   H�QPH����  �pL���qHI��I�H��$�   M��I�[@I�[HI�H��$�   E�kD�3H�K8H�SHI�CH��$�   I�CH��$�   I�CH��$�   I�C H��$�   I�C(H��$�   I�C0H��$�   I�C8I�C�LE�H�C0A����   H9���  fD�t$H��H��H�� ���D�d$A� }  �����@ HcQL9���   ������x  ����D�TD9���  Ic�A������u  L�t$XLt$`D�T$L��$�   M�FPL;D$x�7  H��$�   �P   �;����$�   I�FP���8  IcFHD�T$�PL��E�VLI��A�VHM^P����D  H9��G  H��I��fD�t$H��H��D�d$���� H�D$x�AL   H�APHcAH�PL��I���QHLYP�=���D  L�T$ L9�M��L�T$(LN�L9�LM�O�d L�T$pM)�L��I��D�SH��E8Q��   L�T$8L+T$0M��I��?M1�M)�I��I)�L�T$ M��I��?M1�M)�L9L$ �.  L�\$pI�_HfE�gfA�oL�\$(L�l$ L�\$XL�T$`1�C�lHE1�������    A�H�� ���A� }  fA�C1�fA�KH��fA�S
H��fA�KE1�fD�t$D�d$�����fA�CH��I���� H�D$0H9�~	D�t$TH��H�D$8H9�}�t$Vf�t$H��H�D$@�T$I�_HfE�gI9�fA�oLO�H�D$HH9�HL�D	�A����  H��L)�H;T$h��   ��A���H�T$p)�fA�OfA�G
L��fA�w�����@ �D$I�[HfE�cD	�fA�k�tH��L)�H;D$h}A���fA�KH�T$p)�fA�sfA�C
I�H�|$HI�I�CL�D$@I�GI�CfD�t$TI�GI�CH�t$8I�GI�C H�L$0I�G I�C(H�T$(I�G(I�C0I�G0I�C8I�G8I�C@I�G@I�CHI�GH�D$f�D$VL��L�l$ �(���f�     ��������     �@   H��  []A\A]A^A_�f�     ����A�����{���H��$�   H��$�   H9�$�   ����Hi�$�   �	  HD$XH�PPHc@HL��I��I�L9�r7�~    H9�~
H)�H��fJ
H�O@H�I8H9�~
H)�H��fJ
H��PL9�sLH�r@H�zHH�N8H�G8H�vHH�v8H9�|�H9�}
H)�H��fr
H�O@H�I8H9�}�H)�H��fB
H��PL9�r�1�����fD  H��$�   E1�1ҾP   ��6����$�   I�FP��t�������H�t$xH�xH���H�H�H���  H���  H)�H)��  �����H�IcFHD�T$��$�   �PL��E�VLI��A�VHM^P���������f����H�D$�@����1�)�;D$P�����H�t$�|$P H9������H�RH�B����1�)�9�t�H�B@H�D$����H9����� H�HH��PH�H�H�H�H�H�H9�r������AWAVM��AUA��ATI��U��S��H��(�G�D$    ���  L�GE1�M����  Hc�H��H�JI��L9���   �   @ 9�@��@����   9���   H�B�H�J�H��XH�BXH�BH���   H�J@H�B`H�BH���   H�JHH�BhH�BH���   H�JPH�BpH�B H���   H�BxH�B(H���   H�B0H���   L9�v�r�@���i���9�@��@���i���A�D$��A�D$D��I�H��([]A\A]A^A_��     E9l$ �<����� HcW9�}L�GE1������@ ��]t��   ��L����D�|D9�}Ic�A��]tqM�T$I��$�  I9�toL�L$M�оX   �*4��D�L$1�I��I�D$D��E���U���E�|$A�D$�o���L���  �G   L�G�X����@   1��#����]tA�]t����1�L�L$E1��X   L�T$�3��1�H��I�D$�D$�������L�T$H�yH���I�L��H�I��$�	  H��  H)�H)΁�   ���H�M�D$D�L$�I����     ��AWHi��	  AVAUATUH�SH��(H�h`Hc@XH��H�PH����E�L�D A���A��L9��%  HcG,H�_0L�<�I��I�L9��	  H���.�袋.H��A��H��H��f��3��D����   ���   A���   H�CL�cH�u L9���   I�x�I9���   H���  ��   H����  L9���  �X   1�� L�HXI9�~L��H��L�T H�t H9��I9���  L�\�I�C A�;M�KH���  A)�H�Mc�I��H��H��?H��0 �  H��L�E��u&H�C fD	+H��PI9�����H��([]A\A]A^A_�f�H�C(��f.�     HEH+E�fD  H�CL�c�����f�I+@�I@��fD  I��1�L9�}KJ�4H��H��H�FL�T� M�
M9�|)�B�    H�7H��L��N�HN�T� M�
M9�}+H��H9�|�H��H�GH��L�T �����H��L���    M9�~cH�xI���|����    A�2H�L$H�T$)�I�zL�\$Hc�L�$L)�蘰��L�\$H�L$H�T$L�$M�KA�;I�C ����@ I�B����I��1��]���ff.�     f�AWAVAUATUSH���҉�L�~L�n LD~LDnHi�P9  H�L9��9  �m  Hi�P9  L�4A���  M���9  M���9  M�~PM�nX���J  Ic�H��   E1��D  A��H��8E9��  �   H��c0�Hc�H��H��H��?H��
 �  H�KH��Hc�)�Hc�H��H�L�H��H�{H�{H��H��?H��2 �  H��Hc�L�H�S H�S(H�H�� �  H��H�H��0H��`�j���H�� L��H���H�{�&���H�SH��H)�xBHc�H��H�H�� �  H��Hc�1�H��~H�B H���H�s�K0H)�H�s(����fD  H)�Hc�H��H��H��?H�� �  H��H�H��+1���    L9��9  �����H��[]A\A]A^A_�@ H�� H���H���ff.�     U1�H��SH��H��H�H�GH�FH�GH�FH�GH�FH�G H�F H�G(H�F(H�G0�����H��H��H�ߺ   []������     �ff.�      AW��I��AVAUATUSH��XH��   H�$Hi��	  H�U �RH�\HH�L�`PH�\$H�� -G HcPHH��@X    L�,�H�GI��H�\$ M����  H�_H�ƿ@   耭���D$ I��H�޿    �k���Hc�   H�D$Hi$0I  H�t$(Hc��  H��H��H�H�� �  H��H�H��HN��%���H��M9��5  Hi$�	  L�T$K�4vL��M��D$L�d$M��I��D$4L��M��I���f�H��PI9��3  H�S
H��L9�|�H�SL9��D�KA��t�H�{( t	�H�L9�|�A�GX�s��~C��I�W`H��H�HL�D�X����)�Hc�H��H�߅�HH�H9�}
D:J�  H��XI9�u�L�D$ �L$4A��L�L$HH�|$L�T$8L�\$����L�\$L�T$8����  H�D$HH�xH�     H���H�@P    H)��HX1����H�H�T$HH�ZHH�ZP�C�BH�Cf�H�D$(H��H��?H�� �  H��H�BH�BH�[H��PI9������f�Hi$�	  L�d$M�I�s`McSX�D  I��PM9�vA�|$u�E��~�A�B�E�D$H��H��H�HL�L�X�fD  H��XI9�t��D��)�Hc�H��H�߅�HH�H9�}�H�BHI�D$H�BPL�`L�bPI��PMcSXI�s`M9�w�D  K��H��I�BH�,�H9�w�x  �    H��XH9�v/H�JHH��t�H�� H�PH�@H9�u�H��XH9�w�f.�     L�^H1�E1�L���   �    H�x(A��H�H H����   H�WH9�A��H����A!�H���6  H�y �+  H�V0E1�E���$  H��t:D��>D)�Lc�M��I�م��yMH�D�HA)�Ic�I��I��E��IH�I9�~H�QE����   H�V8�JH�@I9�t>� �M���H�x(��H�H H���N���H��t�H�y t�H�V0E1��n���f�     E����   A9���   �FH�~8 tH�~0 tH�F8    H��XH9������1�H��X[]A\A]A^A_�fD  H�BHH�CH�BPH�XH�ZP�W����    H�V0�@����    E���0���H�V8H��A�   �����D  �F �m����YE1��\$H���l���Hi$�	  M�McSXI�s`�����ff.�     AWAVAUA��ATUSH����L�~L�f LD~LDfIi�0I  H�L9�pI  ��  Ii�0I  A��H��Ic�H�L��pI  L��xI  ��,K  ��t/��pK  H���K  ��t��   f��
H��H����   ��9�u�Ii�0I  H�L�xPL�`XE���'  L�{L�c(Ii�0I  1�H�3H��hH�ǋ@`��t=@ �Ѓ�H�@H��H�HcH��I��I��?J��  �  H��H�H�AH�A9W`w�Mi�0I  I�Ic��  H��H�H�� �  H����'A���  A����   H��[]A\A]A^A_�1�fD  H��H�K@Hc��HK  �IH��H�H�� �  H�CH��H���   Hc��@9�@�ƃ���@��t	�4   ��u�(   H�H���H9������A����  L�{PL�cXL�{L�c ����� L9�xI  �G����O���fD  ��,K  ���;�����H��0K  A�@   A�    L��I������I������I��J��xK  �>@ E1�H��~H��/M��MO�H�� ��H����r@H�BL)�H�B(H��HH9���   H�
L�rHc�D)�H��Hc�H��H��H��?H��0 �  Ic�I��H��I��?H��J��1 �  H�H��L�I��Hc�H�BI��?L�q0H�BJ��> �  H��Hc�L�H�r H�r(�r@����r@I��`�f���H���0���H����~   E1��2���fD  L��@K  J���K  L���@ H��HH9�������y0������u�L���f�     H��HH9�tϋP0��u��t�H�YH9�H�H9X|؃���y0�H���M��ML�����H��L���%�����,K  �sH��t9��H��`K  H��L��ӨK  f�H�QH�9H��H9�HL�H9�HL�H��HI9�u߉�Hc�D)�Hc�H��H��H��?H�� �  H����Hc��ޅ�Hc�HI�H�ƀ���uHc�I��L���I  L���I  �\���ff.�     U1�H��SH��H���F(�G0H�H�G�F,�G4�z���H��H��H�ߺ   []�d���@ USH��H�/H���	  H�wPH�GpH��H�GH    H9�tH���~K��H�CP    H�s`H��  H�CX    H9�tH���VK��H�C`    H��8
  H��X
  Hǃ0
      H9�tH���(K��Hǃ8
      H��H
  H���  Hǃ@
      H9�tH����J��HǃH
      H�s@H��8  H9�tH����J��H�C@    H�s0H��x  H�C8    H9�tH���J��H�C0    H�C(    H�    H��[]�ff.�      H��twATUH��SH�1�L���   �     H�t H��t6H��@*G �@H���.G H�@ H��t
H����H�t L���)J��H�D     H��H���  u�[H��L��]A\�J��� ��)G �ִ��fD  @���&  SE1ۉ�H����   ��uB����   ���9  H���9  H�ʉ�����H��?�  �@   H��[H��E��HE��@ ��Hi�P9  D�D`��tTH�|hH��D���=�����H����   �@   H��?~�H�B H����@ H��A�   ��u��c���D  D���9  E��t"��Hi�P9  H�DpH��H)�H��'H��N��   H��5~DH��H���   �I���H�ʃ�?H��	�9���H���H����   H�A
�"���D  H���@ �6   [H)�H��H�H��H��E��HE�� H��H�������� H��/~2H���"���H�BH�������� H��0�0   HL�����fD  H�B@H������@ H��*H��6H��HB�����ff.�     AWI��AVI��AUI��ATUS�@   H����  ���T$u+�F�q  A�G�f  A���7   �1   HE�@ M�gI�mD��H��   ��L��H)�����H��I�,H��H��?H�H��H��?H��H�L�H��H)�H�4
H��H����?��?�\  H���S  A�@   M��I)�H9���   H��?'H9��/  L9��&  I)�L9��  H9��  H�Ѓ� �  A�@   I)�L��I��I��H��L)�M)�H)�M)�I)�I9�IN�I)�L9�IM�H��H��?I��I��I��?I1�I)�L��H1�L)�I9�HOƋt$��u|H��~gH���   H�4
fD  I9�~jI�MI�wH��[]A\A]A^A_�@ 1�A����H�\;����D  1�H9�~�L9�}tD�D$H��H��E��utH���H������HL�H�H�4
I9��I�uI�OH��[]A\A]A^A_�f�1��q���f�     I��A��?M9��X���L9�������J���f�L�������     H)�H�4
�,���@ Hc�H�<�H��H�H9�w�; � H��PH��H��H9�v$H�F H�H�F(H�B��u֨�������f��ff.�     @ @����   ��A��Hi�0I  ��>�   ��   U1�SH��H��yH�۽   ����   Hi�0I  D�T`A����   A���O  H��O�@   HN�E����   Hi�0I  H��H�DpH��H)�H)�HH�H��'��  H���   �v  H����  M����  H�FH���   �@��	�  ����   H�K H���H��[H�؅�]HE�H���fD  H���@ H�|hH��D������A����   �@   H��?~�H�H H����f�     A��u2�D$uD���I  ������    H���   �H���w����    ���I  H���I  H�ډ������@   H��?�J���H�HH����=���D  H��8�8   HL�����fD  H��/~BH���U���H�HH��H���H��H)�H)�HH�H�������H�K@H��H��0HM������f�H�H@H�������@ H��H�ك�?H��	�����H��H����� ��   H�J
����@ H��0�0   HM�����fD  H���o���M���f���H�FH���   �@��	v;���I���H�gfffffff�   )�I��H��H��H��H��?H��H)�I��H���}*L������   )�I��I���������H��I��H��I��L)������H��6H��6HL������@ UH��A��D�ESH�ZH�BH��   H�I��  API��D�JH)�D��I)�����ZH�H�][]��    UH��SH��H��H��H���i�����tH��[]�fD  H�MH�U�D$H�s0�{,� ����D$H��[]�D  AW��I��AVAUATI��UD��SH��XH�D$Hi��	  H�H�XP�hH�l�������  Hc�H�4�H��H�H9�sV��H�S@L�KH����
�L9�t4H�R@�:A��	�A����u��H�R@�
��A	�tA��I9�u���H��PH9�w�E����  I�wHiD$�	  ��   L�H�XPHcPHD�hhI��   H�,�D�pHH���9���H�D��H��H�T$H��H9�r�  D  H��PH9���   D�ZE9�u�H��fD  H9���   �qD���   D�A�rA)���   �q�yf9rfNrf9zfMzH��H��H)�H9t$lL�R0Mc�J�<�    N��    O�4L9�}M)�L9�|H;r8~L�B0H�r8H�J L�Q0N��    O�4L9�}M)�L9�|H;q8~L�A0H�q8H�Q  H��PH9��3���H��PH9�����H���f�     H��PH9��+  L�A M��t�I9H u�E�PD�IfE9�~�L�i0L9�~�N�4�    H���fD  H��PH9�v��rH9�t�fA9�|�H�z H��t�H9W u�fD;W�ufA9�t�H�r0I9�}�L9�}�H�r8H�4vH9q8�
  H���D  L9���  H��PH9�v�L�^ I9�u�H�F     L�F(���    E����  E9���  �@H�x8 tH�x0 tH�@8    H��XH9���  1�H��X[]A\A]A^A_�fD  I�w�q����    H�S H��t)H9Z t#H�J0H�C     H9�
H��H9K0}H�R H�S(H��PH9�w�HiD$�	  I��   I�\HL�H�\$(HcPHI��@X    H��H�\$0H�XPH��H�<H�|$ E����  I�wHiD$P9  L���  Hc�H��H�D$8Ic�H��H�H�� �  H�����y  1�H;\$ ����HiD$�	  H�D$fD  D�k����  H�D$���  I�t`�A�H��H�PL�FX1�I��H�D$�*�     H��H��f.�     L��L;D$��   I��XD8nu���C)�Hc�I��I�م�L��IH�L9�HN�H9�~�L�[ M��t�L�VH1�M��M���f.�     A)�Ic�L9�}�M�IM9�t$M�Q M��t�A�BE�SfA9C�D)�H��� L9�HL�HL�L��L;D$�]����    H���  H�BHH�CH�BPH�XH�ZPH�D$H��PIcLXH9\$ �����HiD$�	  H��H�QI�D`H�,�H��H9�r���� H��XH9�v/H�rHH��t�H�� H�QH�IH9�u�H��XH9�w�f.�     H�XHH����   H��E1�E1��{�     H�q(A��H��txH9FtrH�P8A�   H��t3D�
�8D)�Lc�M��I�څ��~MH�D�QfA9�~fA)�Ic�I9�~H�VE��tBH�P8�JH�IH9�������u�H�q(A��H��u�H�q H��t�H�P0E1��f�     H�P0��f.�     D)�Hc���     �@ �E����    �sL�D$01�A��H�|$(L�L$H�������=���H�L$H1�H�yH�    H���H�AP    H)���X���H�H�T$HH�ZHH�ZP�C�BH�Cf�H�D$8H��H��?H�� �  H��H�BH�BH�[�����f.�     H�F     H�N(�P����    I�w�T����    �   莒��I��HiD$�	  IcLXH;\$ �n�������D  I�@     H�A     �C��� AWAVAUATI��USH��H��L�j8H�i8I9�H��L��I��H��H��H��L�q0H�z0M��H��I)�L)�I9�tL9�uWI9�s�<�     L�H��PH�C�L9�w$H�C8H9�~�H�L9�H��IL�H��PH�C�L9�v�H��[]A\A]A^A_�D  L��L)�H�L$H)�蕑��I9�r�H�H�L$��    L�H�S0H��PI9�r�H�S8H9�~�L9�|
H���D  )�Hc�H��H��H��?H��2 �  H��Hc�L��@ AWAVAUATUSH��8HcG,L�G0L�O@�t$$L��HcG<I��M�M�<�����   L��M9���   H�P(H��PH�P�H�P�H�P�I9�w�A�   M9�s4M�1M�fHM9���   @ I��M9�wo�D$$����   M9�sfD  I�@0I��PI�@�M9�w�H��8[]A\A]A^A_�M9��s  L��@ H�P H��PH�P�H�P�H�P�I9�w�A�   M9�sL@ M�1M�fHM9��x���A�L��D��t�Jf.�     �D��u8H��PI9�s��J���M9��r����I�@0I��PI�@�M9�w��[���f.�     H��H�xPL9�s�PPD���'  H��H�xPL9�r�I9��  �PPD����   H����VPD����   H��H�nPI9�s�H9���   L9�s6H��H��L��L�D$(L�L$L�T$H�D$�����L�D$(L�L$L�T$H�D$I9��z���H�s�L9��m���H��H��L��L�D$L�L$L�T$����L�L$L�D$L�T$I��M9�������8���H��H��f�     H9���   H��H��L�D$L�L$L�T$�]���H��L�T$L�L$L�D$�����fD  I9������H9��K���fD  H�C0H+C8u����f�     I�V8I��PH�I�V�I9�r�H��PI9�������    H�S8H��PH�H�S�I9�s�I��M9�������k���f�H���;���A�   M9�������u���A�   M9�������a���AW��AVAUATI��USH��(H���  �  ��Z跍��I��1�I���  �/  �E$D�E(D�}<M���1  A��Ic;   Mc�L��L��H��?I�� �  H��Hc�A���Ƀ�)Ή����   ��   B����)����-�V  D�����ǉ���H9���   D�M,�U0�M4D�u8E�ʉT$�m@A��L9��[  ����H9���   D����H9��&  A)�H���ӌ��E���  D)�A)�Ic�A��Hc�Ic��ҋ��D��H��H��褌��H�| �D  A��H��D��艌��H��L���~��� �  ��H��([]A\A]A^A_��    �   A�  K �  K ����� ��L��H�މL$D)ʉT$�0����L$HcT$�������<���D�|$A)�Ic�E)�A��Ic�� ���D��H��H������H�| �b����     Hc�H��H��H��?H��1 �  H��Hc�����fD  ��H�މ�請��H������ D��H��L�T$)L$D�D$D�L$�T$�|���HcT$D�L$D�D$�L$��L�T$����D�|$A)�D�D$Ic�E)�Ic��a���D�D$H��H��A��D���*���H�| ����AWAVAUATI��UH��SH��8H�G H���   H�4$H�T$(H��    �����I�ǋD$(��t H�$L�9H��8[]A\A]A^A_�f.�     H�U H���   1�I�/I��   M���  I�WI�_fA���  IǇ�      IǇ�      IǇ�      IǇ�      IǇ�      H�D$��t$��H��I��W  @ ��?  H��f�H�H9�u�cinuH����������  E1�A��(G ��9G H�D$ HG A�p9G �7f.�     I��M���c  A�EH�� -G H�D$L�pL��N�,�H*G M��t΃x
u�E�E��twL��H��L�D$�`���L�D$���D$,t3����    A�VI9�w:I;GsH�C�f%�?f=�?ufD�"@ L��H�T$,H���P���I���D$,��u�I��E�E��u�H�D$L�@E�0E���4���@ L��H��L�D$�а��L�D$���D$,t;����    A�PI9�wLI;Gs!H�C��Ɓ��?  D9�u��@f��    L��H�T$,H��L�D$賰��L�D$I�ƋD$,��u�I��E�0E���s���I��M�������fD  A�0   f.�     L��H���%�����t��I;Gsf�C �I��I��:u�I���  �p���?  t:I�GH��~1H�<Cf.�     ���f���?f���?u	f% �	�f�H��H9�u�H�t$H���`���A�G    1������AWAVAUATUSH���3  H�GH�|$8H��$H  H��$H  H��L$1���  �H��   H��$�   D�D$ �H�H��$�   H�^H��$�   H��$H  H���   H���   H��(  H�VPH�L$(H�	H�L$0�   �H�D����H�B��H��t9Jt;H�FH�~(�JH�BH�F H�z H�~0H�BH�z(H�~8H�z0H�~@H�vHH�z8H�r@H��$�   L���   H�B H��$�   ��$�   H��$�   H��$�   L��$�   M����  �|$A�   Ǆ$�       H�|$PI;|$�%  H�?H�D$I�D$D�xA���?  N��@*G O�|� A�CL���.G M���H  H��$�   H�\$@M��L��L�|$XM��H�D$H�l$H�   fD  H�CL�} L�e@H����   I�4$H���Љ�$�   ����   H�C H��tH����H��L���j-����$�   ����*  I�T$H�\$D�,A���?  N�<�@*G K�|�  A�WH���.G u.I�$H�sH�T$L���   L���l���H�ŋ�$�   ���J���A��H��$H  HǄ$�       HǄ$�       HǄ$�       ����H���3  D��[]A\A]A^A_ÐM��I��H�\$@H�l$HO�l� M��I��@L��$�   L�,��.G I�EH���e  H��$�   L����I�E0H��tL��H��$H  ��A�ƅ��P����T$ �t$H�߃����(  �����A�ƅ��,�����$�   �U  H�D$(�P��$�   ����  H�\$0H�����   ltuo��  H��$�   A�   H�D$IcwH�EXH+E@H�M`H�H+MHH��Hc�H��H��?H��0 �  H��H�H�D$pIcGH��H��H��?H�� �  H��H�H�D$x���x  H��$(  H���O  H�t$H���B���H��$�   H��$�   H��$�   H�H?H��$�   H���H���H���H��$�   H��?H��$�   H)�H���H��$�   H��$�   H�M0H��H�U@HT$pH)�H�EHHD$xH���H�����$�   H�M8H�UXH�E`t%H�E�@�g  H��$�   H�\$PH9X�0  H�EPH��tH��$8  H+�$(  IcOHcUhH�� ǅ�   ltuoH���H��H�EPH��H��?H��
 �  H��H�H�� H���H�Eh�@����    H�\$@H�l$HA��L�|$X���~��������H��$�   I�GH��$�   I�GH��$�   I�GH��$�   I�G H��$�   I�G(H��$�   I�G0�[��� H���   �xp t�����H�D$8�x! �����H���   �  �L��$�   H�D$h    H�D$8H���   L�L$@H�@PH�D$p    H�D$D�`A���  f�D$���   ��H��H�D$H襁��f���    HǄ$�      H�D$ HǄ$�       HǄ$�       HǄ$�      �����I��@H���.G H�@(H�������H�T$hH�t$pL����fD;d$H�L$hL�L$@uH����  I;��  ��  H���   ���   L�L$@H��$�   ����H�t$��HcVH�H�t$ H��H�H�� �  H��Hc��À��L�L$@H�T$hH�t$ �  I���  ���VH��I���  fA���  fD;d$��  H�L$pH���   ���   L�L$H��$�   �}���L�d$H�t$ ��Hc�IcD$ H��H��H��   H�H�� �  H��Hc��"���L�L$H�T$p �  H�t$HI���  ��A�T$H��H��L�L$fA���  H)�I���  ����L�L$I���  H�\$8I���  L�L$I���  H���   H�������L�L$H��I���  H��$�   H��$�   H�����������@ H�D$(L�HH�xH�p H�H(H�P8H�@0H��$   H��$�   H��$  H��$�   H��L��$�   H��$  H��$  H��$   L��$�   H��$�   H��$�   H�D$覀�����  H�\$0��$�   H�����   ltuotQA�   ����fD  H�T$8H��$�   H������A�ƅ��9���L��$�   Hǃ�    �D L���   ��������tH��$   H��$  H���   � ���HcUPHc�$P  H��$X  H��$h  H��H��$(  H��$0  H��H��$@  H��?H�� �  H��H�H�f���    H��$8  �  M�M8M��t%L��H��H��$H  �|$A�х��j���H��$8  ��$�   �  Hc�$�  ���m  ��$`  �_  H��$�  H�4�H�rL�QL�IH�TѨL�ZH+BL��L)�J�4I��H�W�HL�H��H�VHL�H�O H�V H���H���H��$(  H��$8  M��~I9�H��@H��$(  H��~I9�|H��@H��$8  H)�H)�H��$�   H��  ��$�   H��  H�D$����fD  H�@f�<X �����A�8 �����fD  IcWHcEPHǅ      Hǅ      H��H�H�� �  H��H������H��1�H����������fD  L��$�   H��L���ս��L��H�|$p訽���c��� H��$(  H��$p  H��$x  H�H�� H�H���H�� H��$(  H���H)�H��$8  H)�H��  H��  H��$�   ��$�   H�D$����@ H�t$H��$  ���������f�     H��$(  H�P H�N H���H��$(  �f�H�L$pH�������I;��  ���������H��t[UH��SH��H��H���   H�D$H��tH�E 1�H��[]ÐH�t$������u�Hǃ�    �D H�D$H���   ��f�     �#   �f.�     SI���   ��G I��H��H����� ����   ��G �   L����� ������   ��G �   L����� ������   ��G �   L����� ����   ��G �   L����� ������   ���F �   L����� ������   �բF �   L����� ������   A�Q!��f�     A�QH��@*G �R�H��[�f�     H�;L��H�t$�p�����u�H�T$H�RH�SH��[�f�     A�Q�H��[�@ A�Q ���    H�;L��H�t$� �����u�H�T$�R�S��    A�Q$�A�Q(�SA�Q,�SA�Q0�SA�Q4�SA�Q8�SA�Q<�SA�Q@�S�=���@ �   �/���ff.�      AVH��AUATI�ԉʹ   UH����G SH��0��À� �ۅ�u@��u\A�4$1�1ɸ�9G �D  H��H��@*G H��t7�H9�u�x
u�U�*D  ��G �   H����À� �ۅ�u��t`�   H��0��[]A\A]A^�@ �   ��G H������� ��tO��G �   H����À� �ۅ�us����  A�$�E 릐A�$�EH��0��[]A\A]A^�f.�     �   ���x���I�<$H��H�t$�����Å��]���A�T$H�D$�P�K���fD  ���F �   H����À� �ۅ��8  ����  L�l$M�u�
   H�t$L���-��A�E H�D$�8,�����L9������I��L�`M9�u�L��
   H�t$�c-���ǉD$,H�D$� ������I9������L�d$A�$A�D$��������������A�L$A�t$���v������n���9��f���9��^���E�T$A���  �L���9��D���E�L$E�D$A���  A��A���  A��E��������  �����U$D�U(�E,D�M0�M4D�E8�u<�}@������    �բF �   H����À� �ۅ�u8��uQA�$�E!�����1��
   L���L,��H��t'H��������E �����   ����A�|$������E  �|���1��
   L���,��H���E!�a���ff.�     �AWAVAUATUSH�Ӻ   �H��HL�fH�FH�WhH�VPD�vHH�L$L�gXD�N,H�G`H�$H�V0D�t$L�#H�E����  �JA����  A��L�Bh��O��I��N��
�   �A�9�O�9�L�I��PM9�u�9���  Hc�Mc�Lc�H�T$I��M��L�T$ I��I��?N��
 �  M��I��I��?J�O�� �  M��I��I��I��H�L�I���I���L�OL�H?M�{ I���H�GL�OI��I���L9�L�_ LL�L9�M�Q LO�M)�L�W8M)�L�(L�O0L�G@I��@�0  H�W(M��A�   H�G0L�GHL�WPM��M)�M9���  L�HO�M9���  L�OPO�@M��M�SMI�I��M9�~L�WHM��O��M��M�SMI�I��M9�}L�WPM��L�\$Mc�H�\$0H��H�t$(L�\$8M9���   )�Hc�H�|$�    H�K I��H9�~I��I)�H��M�, �։�)�)�H9�L�I9��   D)�D�4H�t$I���s��H��G��M��I�4E�H��Hc�H�D$H��H��?H�� �  H��H��H)D$P�t$藩��XZL9{P|?H�H�CL�C@L��H��L)�H)�M9��O���H�s(I��H9��X���H)�I)�H���J����H�KXH�s`H�\$(��D)�Hc�H�D$H��H�H�� �  H�D$ H��H��H�H��(  H�H�� �  H��H�H��0  H�D$0H�H�D$8H�0H��H[]A\A]A^A_�f.�     D��)�D�4
�����f�L�OP�$����    L�H�����    L+O(L�WPL�OHI���   ~A�   �����E1�I��`A��N��   �����     AWI��H��AVL��AUATUSH���   H�T$H�L$�����D$���U  A��  ��4  ��T  E1�I�XM��E��H�|$ E��tA����  H�D$ �	  A��E��u�u�H�|$��G0�  H�D$ �D$0    H�XHc H��H�\$8H�PH��H�,H�D$XH9��#  E1�D�d$(M���:�     L�i���CL�kH��tH�z( ��  M��LD�H��XH9���   �C�u�H�K(H�S0H��u�H��t�H�B(H��t�L�h�JI��L�jI��   A��  I�L$H+J�T$0�\���A�L$I�M�l$�@ 1�L���~�����tJ�D$�D$H���   []A\A]A^A_þ   L���S�����u�H�t$�   L���m���A��  �}����H�t$1�L���Q���A��  ��^����D�d$(E1�E1�L�|$@H�\$8E1�D�L$4M��D��D�d$TI��D��H�D$H    ���D$P�AI��   A��  A���T$0H�KI+M�m���IED�sH�CL�T$(H��XL9���   D�sA��u�L�k0M����  @��tI�B?H;C��  I;E�z  I�}( L�T$(�z���I9���  �D$P��  H�|$@ ��  E1�1�L��H��L������H�D$H�K�   M�UH�\$@H��XA�ML9��_���fD  L��D�d$TD�L$4M��E����  H�D$XH=  ��H=   ���Ƅ���  ����  E���=  H�D$8�     �P��u#H�p8H��tH�H��H+NA��HN�PH�HH��XH9�w�E����  L�l$8M��L���D  H��XH9��c  H���Cu�H��XI9�w��@u	H��XI9�v�H���
@ �Au2H��XH9�w�I9�w�H�SH+PHPH�S�f��D$4�:���fD  I9���  H�CH+AHAH�C�r���f����   H�D$ �D$0   H�XHc H��H�\$8H�PH��H�,H�D$XH9��<����A��  ���H9�sl�    H�CHH�K����   H+K@ H�P@L�@H�fD  ��HJ f�2L9�tH�R@�2E��t��HJ(f�2L9�u�H�@H;CHu�H��XH9�r�L��D��L�\$(����L�\$(D��L�������A��L�\$(��   H�D$I�s0A�{,H�HH�P�����/���D  H�@H;CHt�H�KH�P@L�@H��     ��H�J f�2L9�t�H�R@H�K�2E��t��H�J(f�2��D  L��H�T$`H�|$pL�\$(H�L$h�t���L�\$(L�D$hHc|$`IcC,I�S0H�4�H��H�H9�s1D  H�BH��PH��H��H��?H�� �  H��L�H�B�H9�w�A��  �=���M��H�D$ H�XHc H��H�PH�,�E���<���A��  ���9���D  D�D$0H�L$HL��H��L�������i��� I��   A��  A���   �T$0H�KI+M����IED�sI��H�C����@ E�������H�D$ H�XHc H��H�PH�,�����H=  ��H=   @�Ƅ�u	@���F���H�\$8E1�f.�     H�D$8H�HX��u[H�D$8H���  L��  H���   H�GM�PI)�H��H+QM��I)�L)�IH�H9Y0��   E��t+H;l$8��������� H��H���   H��L��`  �f�H�D$ H�XHc H��H�PH�,����� ��0f9�u%H�@H�C������     I��H���Y���D  �;L�p��H�q)�)�Hc�L)�Hc��0i��I�L�s����@ H�GXH9G0�B���I�@0I�XXH9��1���H���'���H�WH�H+QH��I�PI�HH)�H��t*H)P@��tH�|$8H)��  H)��  A�H�H�����@��tH�D$8H)��  H)��  A�H����ff.�     f��;���ff.�     AWI��H��AVAUATUS��L��H���   H�T$8H�L$�5����D$����  A��  ���  ���  E1�M��tA����  A���J  I��M��u�A��  H�|$��W0��  �u�IcGXI�`�D$O E1��D$    H��I��H�|$@H�PH��I�H�D$PL9��R  �D$H    H�\$@L�t$XL�l$ M��M��D  D�cA����   H�k0H���4  H�}( �i  �EH��L�sE1�L�UI��   E�̈D$8A��  PM)�T$L��L�T$8�+���M��ZYL�T$(D�\$0��  A���+  H�uH)�H�sA��D�c�MH;\$@vM�|$O H�CH�S��  H9�����t0H�C0H��t'H�@H)�H��H��?H1�H)�H����
  f�     H��XH;\$ ����M���D$HL�t$XM��M��L�l$ ����	�M���  ���o
  �T$Hi��	  L�H�BPHcRHH��H��H�H9�vKf�     H�xH��t0H�P@H�pHH�f�
H�z(H9�tfD  H�R@H�z(f�
H9�u�H��PH9�r��\$L����蠳����L���v���A�������H�D$8I�w0A�,H�HH�P�R����D$H���   []A\A]A^A_�@ H�D$1�L���h`�֦�����>  �D$���     H�D$�   L�����I  訦����u�L�t$��L���   I���I  �i����   L���������u�I�F@H�@�DX@�����Ic�@
  I��H
  H�t$H��H�PH���I  H��H�D$H9�������FH�����Hc�������H��H�H�� �  H��Hcظ    H�� HN�H�D$(��,K  �D$ ��H��H���xK  �    �t$ ���N	  H�D$L�\$(E1�E1�H��0K  � H��HH9��	  �A@�t��WA��A��A;�P
  ��D8�uE��t�H�7L�H��M��I)�L)�IH�Hc�H��I��I��?J��2 �  H��Hc�L9�}	I��E��I���G�{���H���r������j���L9���A8��[���H�AH��H)�H)�HH�Hc�H��H��H��?H�� �  H��H�L9��%���L�aI��E������fD  A��  �����Ii��	  E1��D$   M��I�t`IcDXH��I��H�t$@H��H�PH��H�D$PI�I��   H� �@H�� -G �@�D$OL9�r~����D  H���  H�}( t(�M����  ���H�E(    �MH�S(H��t3�C��H�R�CH�SH��H��   L�������M M��LD�H��XL9���  �C�u�H�S(H�k0H���s���H��t�H�E(H��t�H�S(H�@�MH�EH��u�H��H���H�D$1ɉ�L��H�Ph�[���1�L�������������A��  ����������D  �t$H��H��L��������K�E���D  L��M+wMwH��L�H��_�  H�J �    �&   A�   H���H��AHL�LL�H��H)�H��I��H��I)�H)�IH�L�I��I)�H)�IH�H9�H��HM�H��?H�H��H��H��H��H�H)�H�KH�E�H����     �D$H����fD  H��@��  H��_��  I�� I���L�sA���t$H��H��D�cL��I�������N���fD  ��  H�R���CH�S�5���D  H9��������D  M�F H��H��I��H��I���I�4H)�H)�HH�K�| H���I��I)�L�I)�H)�IH�H9�}I�< M��L�KH�}�a����M��   �     H�D$PH=  ��  H=   ��  ���k  L;l$@��  L�d$@�l$OL�� �rH�ZX@���  H�K�H���)  H�{�H�AI��I)�H)�IH�H��O�
  LAL�C�I�Ѓ�@�s�M9�sKH�C�H��`���@����  H9�����t-H�C�H��t$H�@H)�H��H��?H1�H)�H��~
H�S�fD  I9��  �T$Hi��	  L�H�BPHcRHH��H��H�M�������H9��F���@ H�xH��t0H�P@H�pHH�f�
H�z H9�tfD  H�R@H�z f�
H9�u�H��PH9�r������f�     I9��p���H�������    M����   H�C�I��L�C�H�� H���H�C������ L�C�I9��"  L9��  I9��  L9��  H�QH�xL�HH9���  L�K���@�s�M9�������    �C�g���H�C�H�S@���M  H9������H���H�C�H���;���H�@H+�`���H��H��?H1�H)�H������H�S������    H9����4���D  H��P���I9�w#��h���t�f�     �@u	H��XI9�v�I9�v'H���Ct�����fD  �A�����H��XI9�w�L�C�H�C�I+CH��H���ICH�C�����@ �    �    L��H��I�I�N H���H��H)�H��I��L��M)�H)�IH�H�H��L)�I)�LH�L9�HM�H��H��?H�H��H)�H�H�SH�E�����D  H9�������D  M�������     IcWHI�GPH��H��H��k����     H�|$P  �1  H�D$@H�xXL���  H��  I�HH�^H)�H��H+GI��I)�H)�IH�H������I�@H�NH�H+G�~H)�H�FH�F0��H����  H)HH�|$P   uH�\$@H)��  H)��  @�~�H������     L;l$@���������H�S�7����    ���H�C(    �CH�E(�W���f�     H�C�H�qH)�L�\$0L�D$(H)�L)�L�L$ H���x[��L�L$ �s�L�D$(L�\$0I�L�K��
���f�     H�|$@L���   H��`  ������     M��tL�g(E��t�OH��XH9|$����������f.�     H�T$`L��H�|$pH�L$h�����IcG,I�W0L�D$hHc|$`H�4�H��H�H9������ H�BH��PH��H��H��?H�� �  H��L�H�B�H9�w�����H�|$P   uH�D$@H)��  H)��  @�~�E����T$Hi��	  L�H�BPHcRHH��H��H������   �&   ����� 1��ff.�     f�1��ff.�     f��ff.�     @ ATI��UH��S�< u�    H���< t���H�_H��v"H���   ��   �W��H�_H����?H	�E1��f�     H�{D����x4H�����u�M����   H�E     H��[A�$    ]A\�f�     I���   vWI���   I����   A��A�   E��H��I�H��L��D�A�H��A��?I	�L9�u�A�B�H�\�y���f.�     D���H��H��A��?I	��T���D  H���   H��vs��A�   D��H�D  �GH��H����?H	�H9�u�A�@�H�\����� H�F@H��H�8�)�����H�E H��[A�$   ]A\� A��A�   �$�����A�   �fD  AV1���  AUATI��USH��H�쀥  H���   �C`    ǃ�9      H�l$H���H�H�H�T$�@H�� -G H�@ f.�     �����  �� u	H���8 t�H��$�2  H�T$H��H��������$�2  w�H�t$H��t��   L���������f  M��$�   fA���    �O  1�H��$�2  ��r  �;���CHH��I���   HǄ$�2     ��$�2  H��$�2  HǄ$�2     L��$�2  H��$8  Ǆ$0      ��������   L�shI��E1�D��H���D$    �R�������   1�H��D��1�����IcUHI�EPH�<�H��H�H9�sFMc�D�D$E1�Mi�P9  �H�P H��tH9B @��H9���@ ��!  H��PH9�w�E��tD�D$���QL��H�|$I��P9  ����$�2  I���	  ���a����D$A������A��tA�   �0���D  �S`����   �CHH��H��H��
H��H���  H�gfffffffH��H��ƃ�   H��?H��H)��9  H���  ��ub�CHH��H��H��
H��H��@;  H��H�gfffffffH��H��ƃH;   H��?H��H)�H��8;  �Q���H�Ā�  []A\A]A^�H�Kh�b���H���9  ��R�p)�Hc�I��I�ۅ�IH�A�������D��A��A��H�4vI�4�H�T3h����AWAVAUATUSH��h  H�H�t$�@L�<��HG ���HG =�  ��  I���    A�GH���PG I���9  �D$    I�EPA�   HD�1�H�D$���u�L  @ H���< t�<|�m  H��H�L$$H�T$(L�������|$$H��w�H�t$(H��t�L�t$�   L������I���   f���   ~���u����   f����  H���   ��L���   1ɺ����L�FM�@1� �6�~9�}JE�_E��A��A����   Hc�H��L�fE��t8�     L���xL9�}��L�ك�H��9�u�Hc�L��M9�t0I��� L���xL9�~��L�ك�H��9�u�Hc�L��M9�u�E���d  ���H�L�0�������� �D$	���   I��A�=�  �Z���H��h  []A\A]A^A_��     H��E1��d���@ fE��t:f.�     H��H��I�|9��xH9�}��H��H��9�}ލ~�"���fD  H��H��I�|9��xH9�~��H��H��9�}ލ~�������v]H�|$0D�]�A�   E1�I��I���     L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��M9�u�H�D$�|$���  D�c�6  �D$H��$�  A�   E1�I��D�X�I��f.�     L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��M9�u�H�D$D���  �D$H��    H�|$H)���H����  ����   H��H��H���  H���  A�W��H9�t?@��@��f9�t2H�H�|$H��H��?H�H��    H)�H��H��H���  H���  H��    H�|$H)�f��unǄ��      ������D$H����  �@�D$�D���H�|$�D$D���  ���$������H�L�0H��    H)�H��H���  H���  H���1���Ǆ��     �R���H�4׉���H���  H�L�0H���  ����1�������    H�0 1 2 3 AVE1�AUE1�ATUH��SH��0H�D$H�\$H�4 5 6 7 H�D$    H�D$$�D$,8 9 �
D  �; t_H��H�L$H�T$H�������|$H��w�H�E@L�d$H�L$�  H�8D���^���M��t�H�D$E��tL9�u#�; I��A�   u��   �E8H��0[]A\A]A^�1��E8H��0[]A\A]A^�D  ATUH��S���   H��L���   �cinu�GHH���(w����tL��H���~��[1�]A\�f�H��H������H��H������H���������ATUH��S���   H��L���   �cinu�GHH����v����t$Hǃ�       L��H���N~��[1�]A\��    H��H������H���]�����ff.�     AV1���  AUATI��USH��H��@�  H���   �C`    ǃ�I      H�l$H���H�H�H�T$�@H�� -G H�@ f.�     �����  �� u	H���8 t�H��$�2  H�T$H��H���?�����$�2  w�H�t$H��t��   L���>������f  M��$�   fA���    �O  1�H��$�2  ���  ����CHH��I���   HǄ$�2     ��$�2  H��$�2  HǄ$�2     L��$�2  H��$8  Ǆ$0      臆������   L�shI��E1�D��H���D$    �Ҏ������   1�H��D��1�蛁��IcUHI�EPH�<�H��H�H9�sFMc�D�D$E1�Mi�0I  �H�P H��tH9B @��H9���@ ��!  H��PH9�w�E��tD�D$���QL��H�|$I��0I  ����$�2  I���	  ����{���D$A��ȶ��A��tA�   �0���D  �S`����   �CHH��H��H��
H��H���  H�gfffffffH��H��ƃ�   H��?H��H)��I  H���  ��ub�CHH��H��H��
H��H�� K  H��H�gfffffffH��H��ƃ(K   H��?H��H)�H��K  �Ѩ��H��@�  []A\A]A^�H�Kh�b���H���I  ��R�p)�Hc�I��I�ۅ�IH�A�������D��A��A��H�4vI�4�H�T3h����AWAVAUATUSH��8  �GHH�H�t$��$I��$�K��H��$�   ��H���HG H�|$��H�\$ ����H�D$p���HG =�  ��   �D$h    H���PG 1�E1��D$L    I��I��L�� A�����  < u
I��A�; t�H�t$L��H��$�   H��$�   �������$�   I�Å�t�H�D$ �D$K L�\$0�@f�$��f��H�E1�H�D$�D$H�D$H�D$   ��fD  A��D9�$�   ��  H��$�   H��t�L�t$�   L��臹��I���   f���   ~���u�H�D$ ���   �pf�t$Hf���   H���   ����E1��D$    L���   1�A������$    L�HH�l$(M�4Q���    �0D9�~dIc�D��f���}   ��    H9�|"I9�LO�H��9�|(H��A��H��I�T��y�H9�H��D��HL�H��9�}�D9�t�t$A��D�$D�^L��M9�tHI���f�H9�"H9�HL�H��9�|�H��A��H��I�T��y�I9�H��D��LO���f.�     H�l$(1�E���@  �D$H�%  H;|$�r����D$KA��H�|$D9�$�   �i����    H�|$L�\$0H��   ������H�����������|$K �D  �D$hH��Ę  �@�D$hA��������f.�     I�܋D$h�\$LL��	��o  H�D$ H�D$ � =�  ����H�D$��,K  ���B  H�D$H�P@H�BH�RH��~,H��$�   H�P�3����?  9�u�A   f�H��H9�u�   H��8  []A\A]A^A_�fD  H;|$�M��������Ic¹����H�\$@D��L���   H�,$L�l$8H��D�d$PD�|$A�I���H�T$(I��<ADʉ�A����    A9�tq��9��N�AM�Lc�L��H��L�H�BH)�I��I��?L1�L)�H��~$H�H��H��L)�I��I��?L1�L)�H9���  C���<u���E��y�A��A9�u�L�l$8�\$8H�\$@D�d$@D�d$PL�l$XE��D�,$�L$`D�|$D�d$l�L$8H�\$PD�d$@�A9�tpA��E9�A�sAN�Hc�I��I��M�I�AH)�H�H1�H)�H��~&I�H+T$(H��H��H��H��?H1�H)�H9��  A���<u�A���y���A9�u�H�\$PL�l$X�L$8D�d$@HcL$`D�d$l�D$HtWH�D$���QD�XHD����Hc�H��I� ��A��Hc�H��L�|$PI+H�H1�H)�I9�~���T$+$)ȃ�9��!  HcD$8��x+HcT$@��x"H��H��I�I+ H��H�H1�H)�H;D$p0A���<t�   �D$H�p��������Hc�A�6��<u�1��U����D$LH�L$H���   �@�D$L�8����L$8H�\$PD��L�l$XHcL$`D�d$@D�d$l�����L�l$8��\$8H�\$@D�d$@D�d$P����1�1��������vb�D$hH��$�  A�   E1�I��D�X�I��fD  L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��M9�u�H�D$�|$LD��,K  E�k�a  �D$LH��$   A�   E1�I���X�H��f.�     L��I�IL��L)���H��H�H9�~H��H�P�H�H9�u�I��I��I��L9�u�H�D$D��,K  �D$L�L$hH�\$��H���   K�ۅ��  H��H��H��HK  H��0K  H�D$ �@H9�t=�@��H9�@��@8�t+H�H�\$H��H��?H�K��H��H��H��HK  H��0K  1�H�\$�K����H���L��`K  H��hK  ��pK  �tK�ۃ��pK  �tH�\$K�ۃ��pK  ������H�\$K�ۃ��pK  ����H�\$�t$LD��,K  ��������D$h��H��Ę  K��H��H��HK  H��H��0K  ����H�4ËD$hH��0K  ��H��Ę  H��HK  �����D�Ћl$L�|$(�L$X�$�	A9��	����P�9���M�Hc�H��I�L9�t�HcL$XA9������H;T$(��L��$�   �D$lA��A��D�؉�$�   �4$H�D$`1�D��$�   D�d$�D$X    �D$(    L��$�   H�\$x�   Lc�M��I��M�I�BI�L)�I��I��?L1�L)�L�H��L)�I��I��?L1�L)�H��~L��I��I9���   G�>A��A���l  L9�A��D:T$luH9T$P��  �   9�tgIcՄ�u&Hc�A���<�K  �D$X����A���D$(����A9�EN�H��L�L�J��H��L)�I��I��?L1�L)�H;D$`����1�9�u�H�\$xL��$�   ��$�   D��$�   �-���H�T$D�m�L��$�   I��L��H��0K  K�LH�H��H��HH9�u�L��A�   E1�����   H�KM��E��H��M)�D�I@A���-f.�     H�:E��t-H�1H9�~.J��H�P�H�I9�tH��H��B@u�H�zE��u�H�qH9��A��D9�v9I��I��H���D�T$(�l$XE��������l$(�y����l$XA��l$(����M��"H�HH�PI�@�@@t.H�@H9�~H�I��M9�tI� �@@u�H��H�I�@�@@u�H� ��1������L�L$PH��H�\$xD�T$X�T$(D�l$`H�<�    L��$�   L��$�   D��$�   9l$�EN$Hc�H��H��H��I�D H+D$PI��I��?L1�L)�H��~I�L)�I��I��?L1�L)�H9�~1A�6��<u��H�A��9�u��L$@��H�|$P�T$8HcL$`�5����T$8D�T$@94$}�v�HcL$`H�|$P�����t$HcL$`H�|$P����f�AWAVAUATE1�UH��SH��H��HH���   H�$���   �cinu�GHH���Wf����t#H�4$H����m��H��HD��[]A\A]A^A_�D  H��H������H��H������A�ą���   �D$<8 9 E1�H�0 1 2 3 L�t$,H�D$,H�4 5 6 7 H�D$    H�D$4H�D$    �D  A�> tdL��H�L$H�T$ H��������|$I��w�H�E@L�|$ H�L$�  H�8D���E���M��t�H�D$E��tH9D$uA�> H�D$A�   u��   �E8������1���A�����������USL��H��H�.H��tH�G@�  ��H�8�ܵ��H��tH�    H��H��[]�fD  D�A9�vx��H�vH��HG�P��ubD�G��USH�_�PH�@     E��t,D�D�PA�P�H�l�H��E�H�2�D9�-NA9�%H�p E9�vA�P�WJ��[]�fD  ��    H��H9�u���ff.�     f���Hi��  H�7�B����   L�D7Lc��  IcI��H��H��?H��
 �  H��Hc�H�Q I�HH���I�PI�P��tg��H�@M�T�0��     I�HHcH��I��H��H��?H��0 �  H��H�H��H)�H)�HH�H��HN�H��H�B�H�� H���H�B�L9�u��ff.�      AWI��AVAUATUL��SH��H9��  u	H9��  tI���  L��1�I���  �����I9�(  uI9�0  ��  I��(  L�߾   I��0  �����I��8  H���I��  H��H��H)�H��I��X  H��H9�A��l  A��`  ��~RLc�Hc�I��H��H��?H�� �  H���� ~0L)�L���#D  H��I��H)�H��?I�� �  H���� ~��u�A��d  1�Hc�M��@  M��P  M��H	  @ �H�G����   ��H�RH��H�|8f.�     HcPH��0H��I��I��?J��" �  H��Hc�H�H�P�HcP�H��I��I��?J��" �  Lc`�H��Hc�L��H�H�P�HcP�M��H��I��?I��I��?J��2 �  H��Hc�H�P�K��, �  H��Hc�H�T H���H�P�H9��\�������ttL�׃�� �����L��ID�����f�     []A\A]A^A_�D  I��X  H���S㥛� H��    H��H��?H��H��H)�H9�A��l  �<���fD  1�Hc�M��P  M��H	  D�P����   A��@  L��I��H  ����   D���H�_H�t@A�@�H��H�@H�H��H�l8�E��tD�	D��+GH�I��I��?L1�L)�H�H��I��I��?J��0 �  I��H����?=�   D  D��A+H�I��I��?L1�L)�H�H��I��I��?J��8 �  H����?~MI��0I9�u�H��0H9��o���A�������D��D�P������A��8  L��I��@  �������� I�F(H��0H�A�I�F H�A�I�FH�A�I�FH�A�H9������f�     H���   ��     H���   ��     H���   ��     �G    �G   �G    �G(    �G8    �GH    �GX    �Gh    ��    �G    �G   �G    �G(    �G8    �GH    �GX    �Gh    ��    L�GH�G     H��H�wHǇ�       H�(��H���)����   1����H�L�BHǂ�   0E Hǂ�   PE Hǂ�   P)E Hǂ�   PE Hǂ�   @,E Hǂ�   (E Hǂ�   PNE Hǂ�   `$E Hǂ�   0NE H���   Hǂ�   �E Hǂ�   @,E Hǂ�   p(E Hǂ   �RE Hǂ  `RE Hǂ  0NE H���   �UH��SH��H��H�w(H�������H�C(    H�sH���C     H�C0    ����H�C    H�sH������H�    H�C    H�C    H��[]� AUI��ATUH��SH���GH�_��tK��H�D@L�$�f�     H�sH��H���0���H�C�    �C�    �C�    �C�    L9�u�I�]H��H�������I�E     I�E    H��[]A\A]�@ D�H�GE��t(A�K�H�LIH��H�@ �`�H��0�@�����H9�u����   �F�UE1�1�SH�\@H�O1�H��1��H�    A����E��t.L�WI�E�BA��uA��E�BA9�vA���N��fD  H��0H9�t��u�D�
�@   H��A��   �fD  �o��~pI�ɍ]�I������E1��     I�qI��>;:/J��    O��D  H�T�H��9:|H�TI�t H��u�I�BI��I��I9�tI���fD  []��G    �ff.�     f����`  A�   AWA��Mc�AV��   AUE��ATUSD��D�AD�A�݉D$��A�H�D�	�\$�L�$G�L�T��WfD  E9���  D�Z!E9�tTE��t	E9��o  ��@t"�L$���   �L$���   H�z( ��   H��HL9�t`�J��u�D�Z H�B0E9�u�I���u���     I��M9�t�I�+I��Hc] I)�M9�}�H)�L9�}݁�  H�j(H��H�J�L9�u�[]A\A]A^A_�@ ��t�I��I�+I��Hc] I)�M9�}H)�L9��  I��M9�u�H�z( �N���I���f�     I��M9��3���I�Hc+H��H9�|�KHc�H9��H�Z(�����������I��D  I�+I��Hc] I)�Hc]M��I)�M9�}L)�L9���   I��M9�u�H�z( ������q����    �������I��� I��M9������I�+I��Hc] I)�Hc]M��I)�M9�}�L)�L9�}ρ�  H�j(�J�e���D  ��  H�j(�J�N���fD  ��������;��� ��    ��  H�j(�J����ff.�      AWI��1�AVI�΍6AUI��ATM��E1�U���   SH��L��H��(L�L$�w���H�C�D$��tH��([]A\A]A^A_�@ ��L�L$E1�1�H���0   L��H�$�8���H�C�D$��u��    A�ML�L$1�E1�L�������t$H�C(����u�H�SH�<$�+�C    I�H���C     H�SH�SH�C0    ���  �E�H�t@H��H�D  �H��0H���BЋA��BԋA��B�H9�u�M����   A�M�~L�s8����   ��H�D@I��H�D$D  E�7M�o1�E1�1�E��u�I ������u$A��E9�t5��u�A�U ��   I���@   ��t�D��H��A���$�����$E9�u�I��L;|$u��+;kt8��tE1�D��H��A���q���A9�u�D$H��([]A\A]A^A_�f�     �t$���J���D  M���<���A�M�~L�s8���������"���ff.�     f�AUI��ATUSH��H����WL�G�i9�r0��H�@I�T��1��    �B    �+I�U H��[]A\A]�D  D�aH��L�L$�   A����D$    D������1�I��H�C�D$��u�D�c�@ D�GE����   ATU��SH��H���t�   �CH��[]A\��    �G(L�'��tH�O0H�@H���p�H�{(H�T$L��������u��CX��tH�S`H�@H�h�H�{XH�T$L���������u�H��[]A\�fD  �ff.�     @ AT��U��SH����D$    D�@1�A��A9�r	H��[]A\ÍZH��D��L����I��H���   ��L�L$H������I�$�D$��u����] H��[]A\�ff.�     �ATUH��S��97v#�؉ٺ�   ����HE��1�[]A\�D  D�fH��H�wD��H��9�����u�D�e �ff.�     @ AWI��E1�AVM��AUI��ATA��U��SH��8����   M��tA�����A�M M�E���N  L��1��fD  ��H��9�tE9*u�D9bu�A�E��tdH�@I�EH�|��L�ډ�������uM��tA�H��8[]A\A]A^A_Ð��A�ED�yA9�sqD��E�} H�@I�D��(D�`D�PA�E��u�I�}L��H�T$(L�\$�����H�|$(L�\$��t�H��8[]A\A]A^A_�@ ���tsA�   E1�����D  �D$(    v�����L�L$(�   ���L��D�T$�L$L�\$����I��I�E�D$(���+����L$D�T$L�\$A�M�3���@ ��A�   E1�����1��
����     AU�   ATI��U�j�SH��H����E�H��H����H�H�vH��L�lf�     I�$�SE1�L��3������uH��H9�u�H��[]A\A]�@ A�D$H��[]A\A]�ATA��UH��SH��H��H�:��*��H�{H��H�$�*��H��H�D$�E��uH��   D��H���3���H��[]A\�f.�     AWAVAUATUSH��  H�<$�t$����   A��H��E1�fD  A��A�   EN�E1�C�\6��\$�@ I��N|� L��� *��H��J�D�I�D$L9�u�D�d$H�D$A��I��J�L$(�    H�P�H)H��H9�u�H�$�P��u�t$H�L$D��H���a���E)�E���e���H��  []A\A]A^A_� H��H��tHH�?�F    ǆ�      ǆ8      ǆ@      ǆH	      ǆP      �����    �ff.�     @ �D�P�E���o  AWIc�AVI��AUATL�$@UI����   S��   H��8H�t$fD  M�^E�j�D��K�#I��L�HD� K�#f�D9D��F
H�B����  A�1@�0uiL���@ D�>D�8uW��H��H����w��t�6@"0@�Ɖ������х�u-��H�����u�E��E���m���1�H��8[]A\A]A^A_�@ D��A��9�wsӉ�E���    E9>v�D��H�RM��E�E��tKH�@M��E�E9���   I�SA��I�pA��t%A�y�1��f.�     H���H�HH9�u�A�     A�@    A�����D)�A����~[��E�HI�HI�pH�@L��Mc�H��D�L$H�L$�a���D�L$H�L$I��K�I���     D�HH�H�@    A���A�E��E���R��������D  L������H�L$I�sI�{D��D�T$,L�D$ L�\$D�L$�7����������L�\$L�D$ D�L$D�T$,I�S�    E9vD�щ�D�Ѓ��������� I�SA��E9�u�����1��ff.�     @ �G��t	��     ATUS�G(L�'��tH�O0H�@H���p���H��H�8L���2�����u.�CX��tH�S`H�@H�h�H�{hL��[]A\�����     []A\�ff.�     AWAVAUATU�)SA�����   ��A�����L�t��   @ D��2D�Z��   ��M�H��E1�D)߅�u��   �     ��   I��0��tlE9~�p�I��H�4vH��L��f�     A����L�>H��0H�@H��L�L�8L�~8L�xL�~@L�xL�~HL�xL�~PL�x L�~XL�x(D��E��u�E�A�yE��tQ��H��1�I9��7����)A�[]A\A]A^A_��    D��L�I)���tA��A��A�   �B���E�XA�x ��� A�A��x9�}�A�y�fD  9�~���q�y�f.�     AVM��AUA��ATUS�D$0D�˅���  L��  H��	  A�$    L��I��1��E     �I���D��L��   �9���E�$�u I�L$E��tME��H���D�XԉP�D�H�A����xH��0A��vD�E��A)�A9�|�D�:��fD  �P���P�E��t�H�}��tJA��H���# E��D+A9�~D�X�D��D�D�@؉P�A��D� �PH��0A��w�D�D�@؉P�E��t�A�   E��uA��H��A����   A�   E��t�)Y�QA����   A�B�L�T@I��I����H��0�A�A؋QL9�t2D�I<E��A)�D����D���9�|ӍA)�H��0�A�D�I�QL9�u΍H��A�BA��A���u���[]A\A]A^�f.�     I��H��  �\����I����ff.�     AWAVAUI��ATUH���p  SH��H��(H�T$�ʄ��I�ċD$���A  ���   M�,$I��$�  A��$�  ���   H���   ��t!�O�H��M�    �H��H���J�H9�u����   ��I�T$(A��$�  A�D$���   H���   ��t"�O�H��M�   @ �H��H���J�H9�u�H����L�UD�M|A�|$L�}(�M	L��j �uM��L�mXI��$8  L�u<H��L�T$H�D$����H�D$M��L���M�u
�$   D�M|H�������D�EXH�MZ1Ҿ   L�T$E��t����fA+zf9�L���H��A9�w�D�E	E��t&H�M*1�@ ���fA+f9�L���H��A9�w�D�E
E��t&H�M>1�@ ���fA+~f9�L���H��A9�w�D�EE��t'H�MZ1�@ ���fA+D} f9�L���H��A9�w�H����  ��!��H9EpHNEpI��$X  �ExA��$`  �E|IǄ$�      IǄ$�      IǄ$(      IǄ$0      A��$h  �D$L�#H��([]A\A]A^A_��     �G��5  AWI��AVAUATI��USH��H��8�7Hc�Liǘ  H�|$Hc�H�$H��M�Mc��  I��I��I��?J��	 �  H��Hc�I��  H�L$HcK�L$(I��I��I��?J�� �  H��Hc����  A���    ��  H�<$���    ��  H�k�D$   H�D$     L�k M��t[A�E�  �T$(���A�U��AU )�I�UHc�I��H��IUH��H��H��?H��> �  H��Hc�H�H��H��H)�H�T$H�4$���    ttH��@��  HiT$�  H��I�TH��H)�H)�HH�H��'�6   H��/~;H��H���   ��  H���?H��	~H��H���@�� ��  H��5H�i6@ L�|$H�kI�O I�T/ H���H���H��L)�L)�H)�H��I��H��?I��?H1�H)�L��H1�L�L)�H9�HO�E1�H�K�T$��tYH�SH�KH��?�j  H�� H��H���A���"  A��t,A����  H�sH��H��@�a  H�� H���H)�H�K���CH��8[]A\A]A^A_�fD  ����  H�$���    ��  H�$���    �  H�k�D$   �L$(E��$8  D�A��$l  �L$,I��$@  E����  Mc�$L  Mc�E��$h  M��M)�M��L�T$ E��A��Mc�M9���  E��$H  E�E9��m  E�A��D$ O�@I��O��p  �(f.�     HcAM��I)�M9�|�AD�A9��"  H��0L9�uًD$ E1�H�D$     A��$@  I��H�IH��I��  E��tnE��$h  LcAE��I)�A��Mc�M9�|QD�IE)�D9���  A��I��N��    M)�I��I��LcAI)�M9�|D�IE)�D9��T  H��0L9�u�1�A����   A����   H�T$ H�{H)�H�S�������    H�k�D$    �i����    H�t$��H�k�CH�sH��8[]A\A]A^A_�fD  A����   A�������A����   H�C@   �    H�� H���H�� ����@ H�k�D$    ������    H�$L��L�������C�3�D$(�C�����A�������H�T$ H)�H�S�����D  H�{������    �@   L�|$ H�sI)�L�{����fD  �@   H�s����f��|$,��uMc�$d  1�M9������A��H�y�����     �D$ L�D$ D�D$,E��uMMc�$d  L;L$ }>H�D$     E1������D  H��~:H�T$H��H�@   H���H�T$�����@ H�IA�   H�L$ ����@ L�T$I�R H���H��~@I�4*M��H��H�N I)�H���L)�IH�I��I��I)�I)�L��IH�H9�HN�H�L$�V���H�T$�L���H�� H����?���H�i
�6���fD  AW1�I��E1�AVAUATUSH���  H�H�|$8H��$�   L�L$x�L$@�   �H�H�NH�T$ �H   1�H��H�\$0H��$  �К��H��$   �D$x�D$��tlH��$  H��$p  H������H��$(  H������H��$   H�������H��$  H��HǄ$       �����D$H���  []A\A]A^A_�f�I�H��L�L$xE1�1Ҿ   �5����|$xH��$  �|$���a���E�GA�?L��$   D��$�   ��$�   ����   I�W�O�L�JI�I1��f�H��L�ʉ�L9�t|I���2����)�H��M�̉PL�tԉ�I�BH��I�L̸I�
����  ��H�T�	M��L��f.�     H�JHH�I�H�RHH��H�AL9�u�M�SH��L�ʉ�L9�u�I�GL��1�E���y  L�d$I����   �    D�[D�߃��|$H��Hc�L�H��L�iL�L�1L��H+rL��H+:I��H��I��?H��?L��I��H1�I1�L)�I)�L�II��M9��\  ���D�BH�D�C H��L�H�H�HL)�L)�H��I��H��?I��?I��I1�I)�L��H1�L)�L�@I��M9���   H����  �D$�C!����   A����   �    ��$�   ��H��H9���   H�|$H���H�9��8��8�H�CH)�H)�H��H��H��H��I�w�������C   A�   �D$   �����@ D�l$�C!E��u"A���x����C"�����k���D�[�    A��D�[�S��� O�II��L9�~�H����  D�t$�C!E��u�A���"�����K�@A�   H��H9������A��E�B�����@ H�D$ L��$  I�W��$�   H��$   H��$   ��t?�q�H��H��H�fD  H�
H��H��H�@�    H�@�    H�H�H�J�H�H�H9�u��D$    ��u�  @ �D$�D$;�$�   �r  �D$H��H�$  �xv�L�L��fD  H�[I9�t�H�k0I+i0L�s8H��M+q8L	�t�H�l$L��H�\$L���D  L��L�e L9�t�L�m0M+l$0L�}8L��M+|$8L	�t�H�|$L��L��L��� ����t�M��M��H�\$�D$(H�l$HL��H�l$L�l$f.�     E1�H�C0H�K8I��I��E���f.�     H�U0H�E8H��I��H��I�n�   H9l$DD�H�U0I��I)�H�E8L��H��H)�H	�t�H�t$H��L��L��������t��|$(M��E��I��L��1��
  H�\$HL��H��L�d$�D$(E���U����x���H�D$8L�D$0H��$(  �pH�H(H�P �n����D$�D$x���R���H�D$8L�D$0H��$p  �pHH�HXH�PP�<����D$���$���L��$   H�D$ I��$(  Hc�@  M��$�  Hc�H�|$`H��L�t$XH�H�� �  H��Hc�H�s H���H����  H9��x  H���X��L��H��H9���  H��H��$   E1�1��T����D$WL��$   �|$@A�  fD��$�  �G���������(  Ƅ$�   ����$�  ����$�  H��$(  H�D$H�D$ �D$    HH  H�D$hH��$  D��$�   L��$   D��$�   H�PE����
  A�y�L��D�\$H��H��H��f�     H��H�H0H��HH�p�H9�t0H�rH�
�@    H�@(    E��t�H��H�p0H��HH�H�H9�u�E��t#H��$  E1ۋ{����  A��H��E9�r�E1�E9�s$D��H��I�z@��@�+   A��E9�r�H�|$L��H�_��t<��D�l$H�l@H��HݐH��D��L��H��0H��$�   ����H9�u�H��$   H�D$�    H�@8L�`D�8HcD$H�D$(D�hHi��  H���  �2���   D��$�   H��$   ��OƉD$0A����  E����  A�G�E9t$D��D�l$8H�@AFT$I�l$L�|$I�D�0I����H��D��L9��\  D9uE��DFeA9�v�E��u L��A)։�H��H��H�U�@���I�wA�D��D�L$8D�D$0H���s���D��$�   H��$   두H�H����     H�r0H9p0uH� H9�u��y���f�     H�hH��H��fD  H�RH9��#���H�r0H�O0H9�t�H;H0~H9�|H�H���� H9�~� �O@H�H9�t��O@H�H9�u���@ �D$W ����fD  Ƅ$�  �   ��$�  ������    H��� H�p8H�J8H9��  H� H9�u�����f��  E���  A�F�I��H�D�	H��H��fD  H�x( t�P��u���PH��HH9�u�HiD$(�  H�$   �|$L���  ��  K�D�	Mc�H�,��$f�     LiL�k@�� �CH��HH9���   H�K(H��t�CL�i��u���u�HcH�{0H)�H����  HcQH�qH9���  )�L�Hc�I��H��H��?H��
 �  H��Hc�H�H�S@�L��H��?L�t$XH�ףp=
ףH��L�H��H)�L������L��$   H��$   HiD$(�  M���  ��$�   H��L�4�L9���  H��1�f��P�������H��HI9�w����  L��$  H�l$x���=  H��E1��D  H��HI9�vM�At�D��H�D� H9�s*H�P�H�q0H9r0�@ H�P�H;r0}H�H��H9�r�H�H��HA��I9�w�A�D$�I��H�D� H�D$0�;fD  �S ��t:S!uH�   @   H�s��  fD  H��HI9���   D�CD����u�C�u�L�M H�{0I�A0E���,  H9��#  H�E�@ H�0H��H9~0
�эQD9�u�H�D$0H�0D��L�V0I9�}�N  �p�H��H�t� L�V0I9��1  �Ѕ�u��H�L� H�A0H9��F  I�Q0I�q@H9��>  H�s@��  @ H�D$xH9�tH��L���۴��HiD$(�  L��$   M���  HiD$(�  L��$  M���  ��$�   ��t~D�P�Mc�I��I��M�@ A�GI�H��H�4�H9�sKH��1�1�D  �@ t
H��HD؃�H��HH9�w�I�܃�w��  f��A ��   I��I�L$H9�u�I��M9�u�H��$  ��$�   H��$   D�\$L�HL�P1���u0�  �L���tL׹    �7	�H��H��;�$�   ��  �ǋJL�B@H��H����L�E��t�L�F��t�L׹@   �7�fD  H��D  H�m�E t�I�t$0L�E0L�]@I�|$@L9���   L)�L)�I��H��H��L��L�T$HL�L$@L�\$8L�D$0H�T$(���L�\$8L�D$0I�L$L�T$HL�L$@H�T$(L��L��H�L�:�<�    L9�|{D)�Hc�I��I��I��?J�� �  H��Hc�L�H�Q@H�IH9�t9H�Q0H)�H���Hc�I��I��I��?J�� �  H��Hc�H�H�Q@H�IH9�u�I��H9��S����X����Hc�H����    L��H)�I)�M����  �   �E���@ u.HcC0L�K@I��H��H��?H�� �  H��H�I)�f.�     H9�t$HcB0I��H��H��?H�� �  H��H�L�H�B@H��HH9�w������f�     �|$W ��   H�D$H�|$������D$   L��$   �����    L�t$H A�NM�vL9�u�K�����f�     Hc�I��H��H��?H�� �  H��Hc�I�L�k@�����)�Ic�Hc�H��H��H��?H�� �  H��H�IA@H�C@A�� D�C�i��������C�}���H�T$`H�t$XE1�1�H��$   ��������D�l$8L�|$I�G8L��H�@H�P�0�����I�wA�D��D�D$0H��E���)���D��$�   H��$   �����/��IŋCL�k@����H���	 H;H8uH�@H9�u��$���H9�}H;H8����@�π�z�	���M�����������H;H8�������   �z�����E������������D  I��   E1�1�L��軈���t$xH�Ņ����������A9�u7D)�Ic�Hc�H��H�H�� �  H��H�HF@H�C@����H�A@H�C@����L�L� ����D��H��L�D$ L�L$hH�D�	H�,��fD  H��HH9�������G ����t�G!����u��Gu�A��8  H�w0I��@  ����   Ic�L  I��E��h  I)�L��E��A��Mc�L9�|`��H�RH��M��p  � HcPH��H)�L9�|9�PD�Hc�H9�"A��l   uIc�d  H9�|H�P �O0H�W@H��0L9�u�A��@  I��H�@H��I�T�E������E��h  HcJE��H)�A��Mc�I9������A��I��J��    I)�I��I��@ HcJH)�L9�������BD)�H�H9�|"A��l   uIc�d  H9�~H�B(�O0H�G@H��0L9�u�����H�D$ L��$  H��$   �����D�L$�C!�E�������A����E��������D�T$�C!�E�������A����$�������H�I@H)�H)�D�\$@H)�H�L$8�3��H�L$8D�CD�\$@H�H�K@�[���I��I���'���ff.�      f�~ tf�> u1�������ff.�     �G����  AWAVAUATUSH��H��8���  ���   L�/I��E�H�l$$��H�vH��H�D$L�tI��H��I�?I���=��L��I��L��H��H��L��H���!������.  H��H�D$0I��H9�u�H�D$D�t$,D�d$(�l$$H�H�z@�B8H�|$����   ��   ��A��E����A��A��D��A��D���A����A��H�D@Mc�A��D����Mc���Hc�L�<����    �9�vH�OB�	D����   D9�vH�OB�D����   D9�vH�G�0���|   H��H�|$L9�u�H�D$H�T$L��H�|8�������u0��xH�|$L���������uE��y_E��xH�|$�9 �   �CH��8[]A\A]A^A_�f�     ��    ��y�E��y$E��x�L��D���O�����t��f�     H�|$L��D���0�����t��f.�     USH��H�PH��H�GX    H�o�HǇ�       H������H�{@H������H�s8H������H�C0    H���   H��H�C8    �]���H�{pH���Q���H�shH��赪��H�C`    H�Ch    �C     H�C    H��[]�ff.�     @ AWAVM��AUI��ATA��UH��S��H���G��tH�WH�@H��D�@�L�}H�T$L��L���i�����tH��[]A\A]A^A_�fD  �E����   H�@H�EH�l��H�uH�}L����f�����u�D��D�῀   �] ����H�u��Iչ�   ��t�@ �E�M A��A��A!�	�A��AD����u	I����   ��u	H����   ��u�H��[]A\A]A^A_�fD  H�T$L��L������H�l$���S���H��[]A\A]A^A_�ff.�     ��G��u)AVAUATUSD�gD�oHC�,9�t[]A\A]A^��     ��    L�7H��H��E1�1�H�D��H��M���h�����uE1�H�{HM��D��D��H���L�����t��C[]A\A]A^�ff.�     ��G��u)AVAUATUS�GD�gHF� D9�t[]A\A]A^��     ��    L�7I�͉�H��A��H���D��M��L���������u1�H�{HM��A��D��L��������t��C[]A\A]A^�f.�     �H���    H�O0��   H9O(��   H���   H�@(    H�@     H�HH�@    H�@8    ��   ��u5A��A����E��AE�f�HH���    t.�   ���   f�Gz1��@ ��tT��(H���    ��f�Hu�H���   ���    �G8b   �   � H���   H���   H��@H�O0�7���D  ����f�H�y����H�G0H���   H��H+JxttOH��H�J @��t�rA����A�� ����AD�f�JH�H@H���   H�O0H�@     H�HH�B8H��f�GxH9G(v�G{ 1��fD  �G8b   �   � �G8c   �   �ff.�     HcG<L�_ I��M��H��D��I)���x/I�S�Lc�L9�~OA�B�H���    H��I�T�L9�~2����y�H�G(H��H�G(H;G0vjA�BA��Hc�Mc҉G<1�K�4�� 1�L9�}ALc���I��H��K�O�D�I)�Hc��	 H�Hc�H�H����L9�u��f.�     ��    �G8b   �   �ff.�     H�OH�G H�H�G@H�H�H��H�H��H��H��H�O0H�OH�G H�G(H�WH�WH�GHH�H�H��H�H��H��H��H�O8H�G(H�W�ff.�     �H�w H�G0H�OH�H�G`H�H�H�H��H��H�H�wPH��H��H�w@H��H�H�H��H��H�WH��H��H�wH�w(H�G0H�G8H�O H�OH�GhH�H�H�H��H��H�H�wXH��H��H�wHH��H�H��H�H��H��H��H�wH�O(H�G8�AWI��AVAULc�ATI��USH��H��(L�g@H�w0M�t$O�,I�QI9���   L9���   �H��H�����Hc�I!�M9�MN�H9���   �{z t�H���   H��H�B(�Cz L9���   �L��L��H)�H��L��H�D�H��H9C(wR�,  @ J�/L�RL)�I��HcCI9���   H�L$H�t$H�T$A��H�T$H�t$H�L$H��L9�r2L9�-�C{ H�GH9�|�u�C{H�H��H�F�HcCH�H�L9�s�L�c@�
@ L��H��I�H�s01�L�c@H��([]A\A]A^A_�fD  Lcǃ�I�D�H!�H��f��������{{ ��   H��H��I�I�, H��{z ����������@ L�H�H��H�L)�H��L)�H��H�I��L�H�F�HcCH�����fD  H�s0�   �C8b   H��([]A\A]A^A_�f�     H�N��C{ �v��� ATH��UH��SH�_@H�[H�[H�[(��uH�[8L��H��D�ezH��H��I������E��t�}z uH���   H�Z(H�[[]A\�D  AUI��ATL��(  UL��SH��H��H�GXL�g@H��8  H��H  H�G`H��@  H��P  L��H��(  L��0  �> H9���   H9���   H9���   H�� H�{@I9���   H�G(H�WH�oL�/H9�}�H9���   H9���   ���   ��tX�sA�   �V�Hc�H!�HcSH9�A��E�Ʌ�tD��H����������   D��D��H����������   A����   H�KhL�Cp��UE H�߾   �y�������   H�{@I9��H���L�kX1�H�k`H��[]A\A]��    ����H�C@H�x H�{@����f����   �4�����t/HcsA�   H��H�t0���Hc�H!�H)�HcCH9�A���$���f�H�KhL�Cp��UE H�߾   ��������]���H���   []A\A]�ff.�      AUATM��UH��(  SH��H��H�GXH�o@L�l$0H��H  H��X  H�G`H��P  H��`  H��8  L��@  L��(  L��0  H����   �     H��L��L9�~	I��L��M��H9���   L9���   I9��  ���   �  ���,  HcsA�   H��H�t0���Hc�H!�H)�HcCH9�A��E�Ʌ�tD��H���������  D��D��H����������   A����   H�KhL�Cp�`VE H�߾   ��������   H�{@H9�wDH�G8H�W(L�GL�oL�'I9�����L��H�������    �{���H�C@H�x0H�{@H9�v�L�cX1�L�k`H��[]A\A]�D  H��0H�{@�fD  ���^����sA�   �V�Hc�H!�HcSH9�A������D  H�KhL�Cp�`VE H�߾   �������7���H���   []A\A]�ff.�      H�H����   H�АH�pH�H��H��f��H�H�h H���H�LH�HH�@H��u�H�BH��H��u�G�    H�JH�RH��t;H�BH��t&H�0H92~�H�H�HH�JH��H�PH�H�BH��u�� ��    �ff.�     @ Hc��   ����f���   ���H�H��H���   �ff.�     LcWA�pL��M�L�����H�I!�H!�f��tH��LcGH)�L)�L9�L9�tH9�IE��H��H����   �wHI��L��L9���   M��A�    IH�H9��ƃ�H�I�ɾ�   ��H������H���   ����I��A����H���   �Ɖ�L�D)�HOP�����~;A	�D���t$��H��H�|H��f�H��� �H9�u�Hc�H�L@q��    D!�	�@�1��    AUATUSHc_H��L�T���H�I��I!�I!�M9�D���I��L��M��x'�GHL9�~L�Ѓ���   H��H��   HGP��[]A\A]��    L�L9�u�A�h���f��tf����   f��t#f��u�M9H8��   M9A8��   L��f��tH�T
�H��H��?H�HcWH��H�H!ƋH��x��H��H��H���WHH9�|_L��M��I�҉�I��M���&����WHL9�����L��A��H��HWPH��   D���2��   ������������� L��� L9�t�M��I��� I�x  �<���@�������I��LcgI)�M9���������� H��I9p(������ �����I��HcwI)�I9����������f�     H���   H��   ��ff.�     @ LcGI��I)�L��M9�}��I�T�H�H!�H!�H9�t
�f�     �H��H��x싇�   H9�v�Hc��   ����f��H��H����H)к�   HGP���Lc_AVAUL��ATM�T���UH�SH��I!�H!�I9�Z���I��L��M��x8���   L9�v-Hc��   ���f��H��H�҉�H)�H�GPHк�   ��[]A\A]A^�f.�     I�M9�u�E�`H��E��A��fA��tfE����   fA��t%fA��u�M9H8��   M9A8��   I��fA��tH�T
�I��I��?I�HcWI��I�I!��M��x��L��H��H�ы��   H9�rrH��L��I�҉�H��H���������   H9������Hc��   ��L�OPA��   f��H��H�҉��A��H)�E������� ��� I���y����     M9�t�L��M��� I�x  �&���A�������I��LcoI)�M9��	������� I9h(����A�� �����I��LcGI)�M9����������@ �ff.�     @ �ff.�     @ 1��ff.�     f�H��H��1�H�hH�@1�H�@p�P1�H���ff.�     @ H��H�hH�@H�@p�`ff.�      H��H�?�U���D  AWM��AVI)�AUATUSH��8M9�A��H;T$p��A��|  M���s  I��M��M��I��H��I��I��I)�L9���  �H��H��H��I�ŋG��!�L;t$p�I  H�|$pH��1�I�����P  E9�L�T$ L�D$�L$D�L$�   A�t$L��L��L�\$(A��)�Hc�����L�\$(D�L$HŋL$I�D$0L�D$L�T$ ��A�D${A�|$z tI��$�   Ic�H�J(A�D$z E)�E��E�MIc�H��I9D$(�!  Ic|$D�L$M���.  L��L��L�\$�����L�\$D�L$H��IcD$I��H�I���   L)�M�D$0H��E���*  K�t�D  I��I�h�H�H�xL)�H�L9�u�I�t$0H��81�[]A\A]A^A_��    A�t$L��H���N�I��D!�������A�|${ I�D$0�����H��I�D$0�����D  H�t$L��L��H)�L��H�L$L�\$�����L�D$A�$L�\$L�T$I�, I��1��+����    A�D$8b   H��8�   []A\A]A^A_� M)�L��L��L�D$�����L�D$D�L$H��H��IcD$I��H�I��H����������� L�������AUATI��UH��SH��H�����   ���>  ����   ��uUH�W`H9�|hH�ChH��L�KpI��D�kzH�sXH��L��H��I��I��H��P�����ZYE��t�{z uH���   H�Z(��uLL�cX1�H�k`H��[]A\A]��    HcO1�H��H�L
���H�H!�H)�HcWH9�@���������(  H���   []A\A]�H�G`H9���   ~��O�Q�Hc�H!�HcS�   H��H9������k�����u����   ����   H�S`H���spH�sXH��L�KhI��L������^_���1����x����     H�W`H9�~ËG1���H�H!�HcGH9�@����������B����G��H�H#G`�\����HcOH��H�L���Hc�H!�H)�HcGH9��¾   H�����������@��������f��������H�S`�F���fD  HcWH�O`H��H�T���H�H!�HcWH)�H9��D  AWAVI��AUATUSH��X��x  @�t$@ ���T  H�IcNI�^ E1�I��E1�H��:  H��I�VpH��8  H�S�Iǆ�       H��fE�VzfA���    I�V(I�F8    I�FhI�FI�F0I���   H�@fE�^x��  H�D$    1�f�H�|$I���   ��Aǆ�       Iǆ�       IcN�4zH�?H��H�D$(I���   H��I��I��I�H�IcVH�(L�`I�} H��L��H��I�UH)�I)�H)�H)ʀ|$ tH��L��I��H��H��H��M���   L����t��A��   ������G  ��u9A�0�����R  H�I�H��L��H��?H��?H�I�H��I��H��H��I�nXM�f`I9��3  H�l$L�d$ �SL�xH�k���2  ��uMIcVH�pIcNH��H�PH)�H)ʀ|$ t	H��H��H��L�����������  H��M9���   L��뚐H�P I9��{  �S�����k  Ic~H�pL�x0H�PH�H L�@(H��McVH��H��L��L)�L)�L)�M)Ѐ|$ �   M9���
  L�X0L��H�x8H��L��I��H��H��M)�H��I��M)�H��L��AS����AXAY���%  H��M9��B���H�l$L�d$ L��H��L����������  ��    Ic^H�pH�PIcNH��H��H)�H)ʀ|$ t	H��H��H��M9��Q	  M��I���O����`  H�L��I��I��?I�H�D5 H��I��H��?H�H���������uyM9��`  H��IcNIc^H��I��I�/I��A�E H���I�_H)�H)ˀ|$ t	H��H��H��<�x���I��I��L��L��L��M���q������'���f�     A�~8b�W	  Ic�x  A�F8    I��H����:  ��8  A��։׉����������  f9���  f��<  ����fD��>  f��:  A��x  �������H��X1�[]A\A]A^A_� M9��7  L�H0L��H�x8M)�L)�I������@ A�F8   �   H��X[]A\A]A^A_�@ I��I��H������f�     I��L�d$ H�l$M��H��H��L��L���O����������I���   H�\$(I�V`I�v0�A�FM���   �H���Hc�H!�u6I;Vh|0I;Vp*I���   H��t�fA3y��uH��I�v0�     Ic~I9q��   A�A��   H9�@��@��L���������L���I���   H��tI�A8H�D$A���   H�|$9������E�fxI���   fA��@��H����@ �u<�|  @ D�l���L��������������A�u������������H�[fA��teH�C 1�fA��tH�SH��H�SH�S(�Cu��rA��)�H������HCHc�H�K(�D  Hc���H�L
�H�H!�H)�H9�@������f�I�F(I9F0�R���I���   H����   A�I�FhE1�E1�H�D$8    H�D$@    H��A��f�D$6I�FpH�D$H    H��A��f�D$41�fD  H�r(�J H�z��fD9�}A��A��fD9�~A��A��H�    H����  H�8 ~�  @ H�8 H�HH�@H��u�H�BH�H��tIH�D$8H����    I�V(I�F0Iǆ�       H9��d���A��x  ��A��x  �n���fD  E��tfD�D$6E��tfD�L$4A�N<����  H�T$6H�t$4L��A��   H�D$8H���\  �L$4��D  �P()ʉP0H�@H��u�A�N<����  ��I�v H����H�H9�u��A�N<1�f�T$f�     ����  H�D$8D�l$H��u�    H��H����   D)h0H�pu�H�T$8H��t%H9�u��  fD  H9��?  H��H�JH��u�H��@�^  H�T$@H���h  H9
~�^  fD  H9
H�zH�RH��u�H�PH�H��H���w���H�|$@�a���H�|$H�W���A�F<I�V �H���H�A�N<L�$�D��)�f�D$fA9��#  A�\$�D��)�A�o�ۍ+�D$L�l$HH�\$@M����   1�H��uJ��   @ L�H9���   @ �D$ M��I��D��L��A��  �D$ H�[M�mH����   M��tH�I�M H9�~	H��H��H��McFH��H)�L��I9�|���N�L�Hc�H��L!�H!�H9�t�H9�t�H9��r����s��f��t�H���I�M M�m�C0   H�[H��u��    f���?  L��A��A��  9l$�  A�N<D��H�T$@H��u�MD  H��H��t@H�z  H�zu�H�D$@H��t�H9�u	��  �H��H�pH��t�H9�u�H��H�8H��H��u�H�T$HH��u�����H��H���t���H�z  H�zu�H�D$HH��t�H9�u�m  D  H��H�pH��t�H9�u�H��H�8�fD  H�T$HH���"  H9
~�  �     H9
�����H�zH�RH��u�H�PH�����fD  H�|$@�������H�|$H����������@ H�\$@L�l$HH��uB����@ �C0��t!�C0    M��I��H�I�M D��L��A��  H�[M�mH���p���M��u��f���D  H��H�2�����@ H�L$8�a���fD  f;l$6�����D  L����A��  f9l$6}��k����    H�|$@H�PH������    H�|$HH�PH������    H�D$H����fD  H�D$@�3���fD  H�T$8�Z���fD  H�l$L�d$ H��I���P��� A�F8   H��X�   []A\A]A^A_�@ I��H�l$H��L�d$ L��H��I��L��H��H��I��L��H��ATL��I���G���^_������������     I��H�l$H��L�d$ L��� Aǆx      �   A�F8   �p��� �l$4�����   �Y���@ H�VH����  H����  �Bf����  H�:f����  L�BM����  H�z �x  A�|x��ȸ   ��9��Y  �   �F�J  H�H���D  �p���1  ����'  H�x �$  H��G  H�
H��$�   H�JH��$�   H�JH��$�   H�JH��$�   H�H�R H��$�   H�HH��$�   H��$�   H�HH��$�   H�HH��$�   H�@ H��$�   H��$�  H�D$H��$�G  H�D$ ������  �$   �@   �   H�      H�L$�   �t$�L$�T$��y  Ƅ$   ��	1ҋ�$�   HǄ$   @^E ��f��$8  Hc�$�   HǄ$  p^E ����$!  �A�f��$:  ��$�   HǄ$  �_E f�D$HH��$�   HǄ$  @aE Ǆ$x      H�D$P��~��H��H�H�D$P1�H���l�������   ��$!   ��   ��$   ��   1�H��   HǄ$   PaE f��$8  ��$�   HǄ$  `aE HǄ$  �aE ��HǄ$  �cE Ǆ$x      f��$:  �����H�ĈG  � 1��D  �   �f.�     �`   �f.�     1�H�ĈG  �fD  ������ �JDш�$   �s���@ H�       �   �@   �$   H�L$�    �)���fD  UH��SH��H��H�    �   H�T$�;���T$��uH�(H�H����[]��    H�    H�B    H�B    H�B    �G 9��   t�D  H���   H���A���AWAVL���   AUATUSH��H��   L��G �D$    9��   tF�D$   H�D$    E1�E1�H��(  �@�V  M��ua�D$H�Ĉ   []A\A]A^A_� �   ��u�H��(  H��I���@�G  L��   H���w�����t3�D$b   �f�     H�t$L��L��H��H�������     ���   L�L$E1�1�Hc��   L���Y��H���   �D$���(���H��(  D���   D+��   �H���   A��Mc�����H�H�D$M��tI�$Ml$H�H�D$L�d$M	���   H���   L�t$(H�}hH�t$ H�D$ �D$0    �Up�D$�������ǃ�   stib�����     H���   L�����H��(  Hǃ�       �`�����fD  H���   L���a��H��(  Hǃ�       �`�����fD  H�t$L��L���@���C���ff.�     ATA�   US�G 9��   u6H��H��H��tH���   H������E1�H��tH�UH�u H���   ����D��[]A\�f.�      �ff.�     @ 1��ff.�     f�H��H�GH��1�H�hHǀX  ����Hǀ`      Hǀh      Hǀp      Hǀx     Hǀ�      H�B1�H�@p�P1�H���f�     H��H�hH�@H�@p�`ff.�      H��H�?�~��D  A��A��	���   ��   D�ȹ�  %�  )�A��   E�Hc�  A������   D�QL���   H�ID��  I�I�A��  
f�1fD�At�f�S��H��H���   L�ʾ
   �����   ǃ      [��    ����   A1�Hc�  A���   AN�A�����w������   Hc�Hc�H)�H��   H��A��wPE��B�$ŠfG D  �H��D�H��D�H�GD�H�xD�H�GD�H�xD�� H���� H���� Ic�������ff.�     f��GDH�Wh+GP�O@H�H��H�H��t;|�tNH�PH�@H��t9~�H���   H;wx}=L�FH�4vL���   L�GpI�4���OX�N�O\H�F�NH�2� �WXP�W\P�AQ�   �����    SH��H�<$�t$�����@   ��u7�L$��t�
 H�$��hG H���   �����T$�Å�uH�$�@`��tH����[�fD  ��	 H�$�@`��u�H�<$�����H����[�ff.�     @ AWAVAUATUSH��@  �GTD�wPA���D$E)�Mc�I��Uv(H���������I�PTH��H��H��I�D�H��1�H��I��N�,�   H���������I�U�H��H��H��$�   H�whH��H�RH��H�Gp��  H)�H�GxD;t$�%  I��I�E�D�D$H��H�$I���   E1�H�D$L��E��I�ƋD$D�|$$H�l$ E�,�D$D�l$D9�DN�D��E��A��D�l$ �@���@��  ����  D�D�eH�D$ H���] H9��e  D�m D�eA�   I�~hH�$1�D��D)�蠉��E�fPD��L��Iǆ�       A�F`   E�nT�������u�E�fPE;fT��   L�l$D��D��I�Vh)�Hc�H��H��tu�E1�fD  �S��	A�D��+Kt
A9FH��   H�[�pH��t)�E��t�9�}�)�D��D��L��A���������    E��tE�FLD��D��L��A)��v���A��  ��~I���   L��D��A���   Aǆ      A��E;fT}2A�FP�9���f�     ��A�   D��L��������Q���fD  H��H�D$ H9������D�|$D9|$~)I�~hA�   � ��� �   H�Ę@  []A\A]A^A_�1���D  H����  �N�   ���  H�VH���  �Bf����   L�fE����   L�JM����   H�z ��   G�DA����   A��D9���   H��(  H�:H�H��$�   H�zH��$�   H�zH��$�   H�zH��$�   H�R H��$�   ���}   H�FH��tUH��$�   H�F8Ǆ$      H�VPH��$�   H�F@�T$L���D$HH�FH�D$P��H�VX�T$T9�~�D$P9D$T��   1�H��(  �D  1��D  �   �f�H��t{�P��tՋ0��t�H�xH��te�@��xD�F�D��Lǉ�$�   ��H��$�   HǄ$�       HǄ$�       Ǆ$  �����D$H    �D$P    �T$L�t$T�Q���f��   �Y���fD  H���X����F��� �   �f.�     SH��H���G`��uH�X uR�KHH�CX    �SD�A�9�NƉC@�   9ST~9SP~�C`H��[�f�     1�9sL���C`H��[��    �T$�t$�����T$�t$뗐AWAVI��AUATI��USH��HH���   H��H�t$H��H�Ɖ��|$H��9�N�A9VT��  A�VPA��9��N  9���  H�L$I���   M��I)�I��H��H)���I��H��I��D�D$D��M����  M���z  H�D$0    Mc�Hc�M��I��I)�;l$tH�������� H�I��H�D$0H�D$(    9�tH�������� H�I��H�D$(I��I��L�d$8A��L�\$D��L�T$ L��A�F\H+T$A�vXM���G  H�L$ H�<H���~  H����  H�T$()�A��A�F\H��I��L|$H��8��ݽ   )މ�A�vXD��D��L�������D;d$u�D;l$�{���A��L�d$8�8�I���   L�T$D��I��I����I��D�T$D��E9���  9��y  �D$A��D)�AV\���A^XH�D$M���   I���   H��H[]A\A]A^A_�fD  M���_  L�d$E��D�l$A�   @ D��A����L��D)�AF\D�����AFX�$���E1�E9�u�L�d$�i���f�H��~;H�|$0A��I��L+|$ H��8��)�����A�F\޻   A�vX�����fD  H�L$ H�<H��~BH�|$A�   A��A)�1�L)�H�|$(D�I��A�F\H��8�A��މ�A�vX�y���@ H�|$ L��6���H�T$0��   A��I��H��H��8A��A)��A��D�A�F\�1�A�vX�-����     L�\$M��I)�I)��)���D  �t$��L���
����u���D  D�|$ E)F\A��A����D��D��L��E�EFX�����A�   E9�u�����D  H��H��H�OH�7H��H��    H������1�H����    ATI��USH�H�_L��H�,�    H��H��H��H��H���`���I��$�   1�I��$�   []A\�f�     UH��SH��H��H�    �   H�T$�N+���T$��uH�(H�H����[]��    H�    H�B    H�B    H�B    �G 9��   t�D  H���   H���	���AWAVL���   AUATUH��SH��H���   H��(  L�W�D$l    � �@��9��   t6�D$l   1�E1�E1��u>H��uu�D$lH���   []A\A]A^A_��    A��D9�tp�D$l   1�E1�E1��t�H���   L��H�L$��p��H��(  H�L$Hǃ�       �`�H��t��     L��L��L��H��H������r����    I�˅��m  L��D��H��L�T$L�\$�M���L�\$L�T$��t'�D$lb   H��(  �@1�E1�E1������D  ���   E1�1�L��Hc��   L�L$lL�T$L�\$��H���L$lL�T$H���   H��(  ��u����   ���   D���   �H����L�\$��A��Lc�Hc�A��I̀��   Mc�u��VUUU����)�Lc�I�M��tM#MkL��L	���   H���   L�t$xH�D$pǄ$�      A����   A���@  H�L$H�}hH�t$pL�T$�UpH�L$L�T$�D$l����   ǃ�   stib�����D  H���   L��L�T$H�L$�o��L�\$L�T$Hǃ�       H��(  �`��U���f.�     L��L��L��H�L$L�T$����H�L$L�T$�!���f�     H��(  �@���`���fD  ���   L�;L��H�L$L�T$�D$$���   I��`  I��X  �D$���   H��H�މD$(�a��H�}hH�t$p�UpL�T$H�L$���D$lu��D$�����L��H�L$0I��X  I+�h  L�T$�����H��   �T$8I��`  I+�p  H�D$����H�}hH�t$p�UpH���   H+T$��L�T$H�L$0�D$lH���   �����D$8I��h  L��L�T$I+�x  H�L$@�H�H�D$0H���   I��p  I+��  �~��H�}hH�t$p�UpH�T$0H)��   ���D$lL�T$��  H��(  H�L$@�@�������fD  �����L�;L��H�L$D���   L�T$I��`  C�	D�L$�D$$D�H�މ��   �����   �ꉓ�   I��X  ����H�}hH�t$p�UpLcL$L�T$���D$lH�L$�����I��h  L��   L��I+�X  I��`  H�L$I+�p  L�T$L�L$���H�}hH�t$p�UpH���   L�L$L�T$H�L$�D$lL)ʅ�H���   �����LcD$$I��p  L��H�L$I+��  L�T$L�L�D$H���   I��x  I+�h  ���H�}hH�t$p�UpL�D$L)��   ��L�T$H�L$�D$l�������   �VUUUM+��  M�x  �����ꋃ�   �@)�L�ቃ�   ���   L	��I���HcD$(H�T$lL��M+�x  M+��  L�T$(H��H�D$�$���T$lL��L�T$(L	�H�Ņ�������D$$1�1҅���   A�   A�   L�T$HH�L$XA)�A)�L�t$@D�t$8L�d$PE��E��L�l$8A��H�\$(H��D  H�D$(H���   H߃|$vIH�D$0H�L$H��L�L�1� ��
A�4A�@�t A�4A�H��H��@�t A9�w�H�T$H��A����x��H\$D9l$$u�L�t$@L�T$HL�l$8L�d$PH�L$XH�\$(L��H��H�L$L�T$�9j���D$lL�T$H�L$�����fD  ���    D�E1��}���ff.�     f�A�   �e���D  A�   �U���D  AVH��I��AUH��H��ATN�$�    USH��  L���   L���   H��$@  L�$$H�L$H�,�    �GTL�D$I��H�l$I��H�t$ H�T$(L�T$0L�\$8A9�|L��H��9���  �GPI��A9�}+M��I��D9�~I��I��D9�~M��I��D9���   I��L��f.�     H��    H��H)�J�gL�H��H��?H1�H)�H=�   ��   J��    L��H)�H�oL�H��H��?H1�H)�H=�   ��   H��    H��H)�H��L�J�PH��H��?H1�H)�H=�   oH��    H��H)�H��H�J�XH��H��?H1�H)�H=�   BH��L��L�������L9���   H�K�L�C�I��M��H�s�H�S�H��0H�kL�#����D  I�L�1I�2L�L��M�H��L�H��H��I��H��H�{L��I�I�H��H��L�S`H��0H�{�I�<H��I��H�H�H��H�s H��I��H�I��I��H��H�KH��L�#L�[8H�S(L�CL�K�H�{�H�k�l���@ H��H��9�����L��H��9�����L���   H���   H��  []A\A]A^�ff.�     �H���rH��L�
L�FH�H�WH�7H���-���1�H���fD  ATI��H��    H��    UM��SI��H��  L���   �_TL���   H�L$H��    H�$L�D$H�L$L�\$ L�L$(A9�|H��H��9�L��H��9��D  D  �_PA9�}H��9�~L��H��9��   �L�H��A�   H)�H��H��H��?H1�H)�H��K�H)�H�H1�H)�H9�HM�H��@~H��E�H��@�H��H��D  E��A��E!�A����   L�S H�{L�K(H�K�@ H��H�I�4:I�	L�S@L�KHH�H��H�H��H�CH�CH��H��H�{0H�H��H�s H�H��H��H��H�K8A��H�CH�C H�S(u�H���'���A���e���H��  []A\ÐH�SH�3H��H�� �����A���;�����H���   L���   H��  []A\��    H��H��L�FH�WH�H�7H������1�H���ff.�     �ATA�   US�G 9��   u6H��H��H��tH���   H������E1�H��tH�UH�u H���   ����D��[]A\�f.�      AWH��AVAUATUSH���   H�L$�L��$   H�D$�    H�D$�    H�D$�    H�D$�    H�$    H�D$    H�D$    H�D$    �T$�H��$  L�D$�A��L�L$�N�� H���H��D��L9�u�D�T$�A9��i  ��D$��   fD  �l��������   H��H��u��D$�   �   �   D�L$�D9�v	�L$�D�L$�L�\$�   �A���uYI����u����    D)Ӊ\$���  �D$�E1Ƀ���D$$    �D$�    �D$�    �   @ �D$��   ��� �t$�;t$�s�t$�A��\$��9��  ��+D���m  D�Q���J�T��I�J�L���fD  +H�����B  �H9�u���+\���\$��)  �D�����D$$    ��1�1��f�     H��T��H�H�T�(H9�u�L��$(  1�f�����t�L� �qA���t� H��L9�u�HcD$�E��H�D$`    A��H�ËD� �D$     ;\$��  E1�H��$(  �D$�    H������A�   H��1�H�D$�HcD$�H�D��H�D$��D$����D$�1�H�|$����|$��|$��O�D����|$ċL$�����  �|$��l$�G�D)�D)��J�D��L�\�`L��B�\� A��L)�A��H��D��A��I��A)�@�2D�|$�D�JD�zE��D)�D)�Ic�E�D;D$���   D����D�R����9D$�s�t$�9�A����DG�A9�wEE�u A����  ��   L��$  A�M O�4�Mc�N�t�`E���P���H�t$�L�6�fD  �wA9�v/L�|$�+D$��A�9�w�@ I��A��9�s
��)�A9�w��D��E�u ��A����  �}���fD  �����H���   []A\A]A^A_ÐD�D$������H�|$�E)�H;�$(  v4H��$(  H��$(  �?�|$�;|$���   ��   �`   �    E��L$�D��A�ڋl$�D)���D��A��D��D9�vfD  A���O��A�2E�BA�j9�w�|$ĉ���tfD  1����u�1�D��D��Hc������!�;L� t+��D��Hc�D  D)�D��Hc�H�����!�;|�$u�A�˃l$�����f�     H�D$�H�     1��    ������    H�|$��L$�+L$��<��|$��|$��wPH�|$��<��|$������D$��|$�H�D$�;|$��-����t$Ѕ�t�|$�u1��q���������g������+\���\$��P����D���D$$    ���G�������ff.�      UH��SH��H��H��tH�GhH���P���wH�sH�}P�UH���uH�sH�}P�UHH�C@�    �C,    H�CXH�CPH�C`H�C0    H��t1�1�1���H�ChH�E`H��[]�H��tGH�W8H��t>H���zH��H�G(    �H�G    ��H�G0    H�z ���1��;���1�H��ø�����ff.�      H��tsH�w8H��tjH�GHH��taUSH��H��H�n H��t51�H��H�������H�u@H�{P�SHH�u8H�{P�SHH��H�{P�SHH�CHH�s8H�{P��H�C8    H��1�[]� ������f�AWD��H��AV��AUATUSH�D$�H����  ����  I��f����  ��  ��F�)ǉ|$����  ���D$����D$�H��H��L�H�D$� A�E�rI��E�j�E�b�L�A�j�A�Z�I�E�Z�E�J�M�L�E�B�A�z�M�L�A�R�E�z�L�L�H�H�I�4E�Z�H�H�t$�H\$�I�A�r�L��E�Z�H�L$�H\$�I�A�J�M�I�M�M�L�M�H�L�H�H�H�H�I�H�L�HT$�L;T$��.����D$��|$���)ǉ���   H���/�  H�|$�I��L��H)�H��H�H���/�  H��Hi���  I)�H��H��H)�H��H�H��Hi���  H)׋T$�H�|$����u���H�D$�[]A\H��A]A^L	�A_�fD  L�T$�H�|$��H�L$�H��H�tH�� H���x�I�L�H9�u�H�|$�Hc�H�L$�L�T�5���[�   ]A\A]A^A_�ff.�      ATUH��SH�_L�g8H��tiH�{�#���H�CX    H��L��H�C`    H�Ch    H�C    H�C0    �C     �C8    H�C    H�    H�C    �Z��H�E    H�}( t[]A\��    H�u L���Z��[H�E     ]A\��    �kZ��ff.�     �[Z��ff.�     �҉�H��H��H�T$���H���D  �҉�H��H��H�T$�z��H���D  U1�SH��H��������D$��tH��[]Ð�   H�t$H��������D$��uހ|$�   uҀ|$�uˀ|$u��D$�u��   H�������D$�D$�uj�t%H�l$f�H��H�������D$��u���u��D$�t0H�l$f�     H��H������D$���O�����u��D$�uF�D$�9���H�l$H��H���������D$������H�������D$�������D$�Y����   H������������f�AWAVAUATUH��SH��H��L�PH�GXL�fL9�sH�GH�M L)�9�F���thE1���u`)�A��Lu(�M H�K`H��tH�{h��L����H�ChH�E`L��L��L��M��f��M�L9sHt&L�eD��L�sPH��[]A\A]A^A_�@ A��� H�SXH�K@�E I9�txH)�9�G�A��)�O�<N�4��tA����    DD�E H�C`LE(H��t#L�D$H��H�{hH�$��L�D$H�$H�ChH�E`L��L��H��M���f���[���f�     H�KXI��M��E1�1��ff.�     @ H����  AVAUATU��SH�G@H��H�G0    H���%  H�PH�{H �  �(   �   ��I��H�C8H���r  H�@     ����   �@    �E����7  A�D$��H�{PA�l$A�   A�@�E �p   �   A����    LE��S@H��H����   H�{P��  �   �S@H�{PH�E8H����   D��   �S@H�E@H����   L�L�u`1�H��H�EHH���E     ����I�l$ H���.���1�[]A\A]A^� ���@   �/���f�H�CH@�E ����� H�G@p�E �p�E H�GP    1������@ H���SHI�D$     H���)���������f�H�u8H�{P�SHH�{PH���SHI�D$     ��H�������������b��������ø�����R���ff.�      H���w  H�O8H���j  AWAVAUATUSH��hH�/H���L  E1�������A�ă9G�d����   �H���$� kG �    ����������   H��W�H�C�SH�pH�3� �   H��H�AD������   H���H�C�SH�pH�3� �   H��HAD����t\H���H�C�SH�pH�3� �   H��HAD����t/H���H�C�SH�PH�� HAH�AH�C`�   �   H��h[]A\A]A^A_��    �GA���������  ��H�C�CH�H�PH�� HAH�AH;A�  �   H�C0�iG �A   H��h�����[]A\A]A^A_�@ �W����  H�E��H�GH��W�u ���q��<��  �   H�G0�hG �A   렋W��������*���H��z��q�{H�PH�C��H�� ��B�A�������)����������)�9��R  �   H�C0iG �A   �0����W��������� �   �����H�G04iG �A    H��h[]A\A]A^A_��    �W��������z���H���H�C�SH�pH�3� �
   H��HAD�����I����B�H�H�C�CH�rH�3��   H��HQ�=���@ �W������fD  �W������l��� �W��������� ������S�������H���H�C�SH�pH�3� �	   H��H�AD���*����   @ �   ����fD  A�� �[  �   H�+D��L�Q D�sM�ZXM�BPM�z0E�j,M9�s%M)�A��A�D�$$M��A�҃�	�_  �$�pkG �E�BHE)���M��L��M�|$0H��H+�����E�l$,H��L��HCD�sH�+M�\$X�������m  I�t$H�{P�SHM�\$XM�D$PH�+D�sM�|$0E�l$,M9��+  M)�A��A�T$(����  A�$    E1�A���#  E���6  �E D��A��L�MA��E1�H��I	�D����A�D$(D��������l  ����  ���i  A��A�$   I��L��D���I��A)�A��w@E����  D���f�     E����  H���E�A��H����I	ǃ�v�A��E1�L��H��H��L1�f����  E��E�l$E����  A�t$(����  D��M��E1�D�$$A�   �[  M��D�$$M�z0H��H+E�j,HCD�sH�+M�ZX�����H��L������D  �����
  ���o
  D���A���E�L$A�T$���������э�  D9���  A�t$D9�v>E����  D����     E����
  H���E�A��H����I	�9�w�A��E1�I�D$ D��#��lG H�ȋxD�@���  I�D$A�QD��E)�A�T$I��B�<�E�L$�M���A�D$A�t$D����
��9���   H���w!E���   �E A��H�UE1�H����I	Ǎ~I�D$�4� lG ��A�|$D��I�����<�A�D$A�t$��
��9���  H��H���v��f��VI�D$A�T$�� lG ��    A�t$��v�M�D$8I�D$M�L$ I�L$D�T$<H�{P�   �   L�\$0A�D$   L�D$(L�L$ H�L$H�D$�D$X    �S@H�L$L�L$ H��H�D$L�D$(L�\$0D�T$<�0  D�T$ �   �   L�\$�t$H�D$`PAPE1�QH�|$01�� ���H�� L�\$D�T$ ����  H�SHH�{P�����  A�|$ ��  �D$ H�t$D�T$L�\$�ҋD$ L�\$D�T$����  A�D$    E1�A�$   �v���M��D�$$M�z0H��H+�   E�j,H��L��HCD�sH�+M�ZX�$������������������D$�t$(L�\$0A��}G H�|$ �t$�`~G ��H�<�H�T$TR1��t$(H�D$`PL�L$x�!���H�� L�\$0���(  �|$H H�SHH�{PD�T$<u�|$  �P  D�T$0H�t$L�\$(��H�L$PH�{P�0   D�D$HD�L$D�   H�D$XH�L$ D�D$D�L$H�D$�S@D�L$D�D$H��H�L$ L�\$(D�T$0�s  H�|$D�HD�@I�t$H�x(H�{PD�T$L�\$�     H�H I�D$�SHA�$   D�T$L�\$I�t$PH��M�D$M�|$0E�l$,H+D�sHCH�+M�\$XL9��m  L)ރ�L��A� I��M��I����	��
  �$��kG A�$   I��A��L��A��w:E���p  D��� E���  H���E�A��H����I	ǃ�v�A��E1�D��D��%�?  ��A�D$����  ��������  D�T$��  H�{P�   L�\$�S@L�\$D�T$H��I�D$�   A��I��1�A�D$    A�$   D������A�$   E1�E1�E����  E��uRM9\$H��	  M�\$XD��H��L������M�\$XI�L$PI9���
  I��I�T$HM)�A��I9��e  E����  A�L$H��L��D�D$D9�AG�D9�AG�A�ɉL$L��L�L$�LX���L$L�L$D�D$I��L�A)�M�A)�A)L$�����A�$E1������D��M��D�$$M�ZXL��H��L�$�����L�$M�ZXM;ZP��  A�   �\���E1�D��#��lG H��I�D$H���B��A)�I���
�ȅ��O  �BA�$   L��A�D$��u_M9XH�g  I�HXD��L��L��L�L$L�D$�>���L�D$L�L$I�HXI�PPH9��+  H��I�xHH)΃�H9���  ���  A�D$L�Y��E1҈A�T$I�D$ A�$   A�T$I�D$D9��$���E��u�
  @ E���$  H���E�D��A��A��H��I	�A9�r������A�T$A9�s4E��u�	  E����  H���E�D��A��A��H��I	�A9�r�E1�D��#��lG H��I�D$H���B��A)��I���	  ��A�D$�BA�$   A�D$A�T$D9�v9E��u�:	  D  E���\  H���E�D��A��A��H��I	�D9�w�E1҉Љ�A)�A�$   �<��lG D!�I���AD$A�D$�A�D$L��I�P@H)�H9�sI�@HH)�f�     H�H9�r�A�L$����   �r���fD  M;XH�&  M�XXL��D��L��L�L$L�D$�:���L�D$L�L$I�xXI�PPH9���  H��I�HHH)���H9���  ����  �L�_��H���I;XH�U  A�l$A�    ��������m���L����A�T$�����M��L��M�|$0H��H+�   E�l$,H��L��HCD�sH�+M�\$X���������L��L��M��I��A��vA��A��H��M�\$XD��H��L��L�D$�M���M�\$XM;\$PL�D$��  A�    �t������  ��A�D$�BA�$   A�D$A�T$D9�v<E��u�5  �     E���T  H���E�D��A��A��H��I	�D9�w�E1҉Љ�A)�A�T$�<��lG I�D$(A�$   A�T$D!�I�D$I��A|$�����L������ �������H�K8H�މ$H�y H�Q����H�K8�A��t]�   �$�����    H�C8�    �@    �����f.�     ����;qvu�   H�G0	iG �A   ���� �   D���_���f.�     M��D�$$A��1�M�z0H��H+H��E�j,L��HC�C    H�+M�ZX��������@ �   D������I�X@����M��H��H+�����M�z0H��L��D�$$E�j,HCD�sH�+M�ZX�U����P���������A�t$HD)�����E�D$HE)������I�@PI�x@H9��������  H)��p����
���I������A��D��M��D�$$����I�|$8I�t$  L�\$0D�T$<�   H�|$H�{PH�t$ �   �L$(I�D$     �D$D	   �D$H   �D$�D$L    �S@L�\$0H��H�D$��  PA��~G �`G H�T$TR�  �t$(H�D$\P�t$0H�|$@L�L$p����H�� L�\$0���}  �|$D ����M��D�$$H�C0�jG �����H�{PH�t$�D$L�\$L�$�SHL�$L�\$�D$����D$�!  I�rH�{PL�\$L�$�SHL�$L�\$�D$A�	   M�z0H��H+H��E�j,L��HS��D�sH�+M�ZX��������M��L��E1�M�|$0H��H+D��E�l$,H��L��HC�C    H�+M�\$X�Y����������������I�HH��)��+�������  �G��D$   �D$�D$A�4 D9�v@E������D���f.�     E������H���E�A��H����I	�9�r�A��E1�D��L��D�D$A)�H��I�t$I��D��I��D��#��lG �L$�D�9��3  ��u	E���%  1҃�uA�A����I�t$A��A�AB��9�u�A�L$A���}���M��1�D�$$A�   �l���D��)��-���I�x@H9��h  ��  H)��r�����������r���M�x0H��I+�����E�h,L��L��M��IAL��E�qI�)M�XX������?���I�T$PI�D$@H9��8����  H)�D�B�I��E���f��������    A�$    E1��Y����D$   �D$   �^���L�L$H�{P�0   �   L�\$D�T$�S@L�\$L�L$H����  �	  I��A��L���     D�T$f�xH�@ �mG H�@(�lG I�D$A�$   �%���M��I��A��L��D�$$H+A�	   H�C0DiG M�z0E�j,D�sHCL������   D���]���I�T$HA��E)��U���A��H���*���L�d$H�t$D�$$H�C0`jG L�$��L�$L�T$I�rH�{PL�\$L�$�SHL�$�����L�\$A�	   ������)��E���M�|$0H��H+H��E�l$,L��HS��D�sH�+M�\$X�!����{���I��������@��  A�D$�BH��I�D$A�$�P���M�\$@L9���  I��L)�M)�A��L9�DF��t���H������M��L���.���E��A)������H�{PH�t$L�d$H�C08jG D�$$L�$�SHL�$L�T$�����M�x0H��I+L��E�h,M��L��IQ��E�qI�)I�xXL���N��������@u3A�L$�BH��I�D$A�$����M���H��D�$$L����������L��L��M��I��� ��  �   �|���I�PPI�@@H9������H��I)�H��H)ƃ�H9�AF��������e���M��H��H+D�$$M�z0E�j,HCD�sH�+M�ZX�����H��L����������M��D�$$A�	   H�C0jG �9���L�d$H�{PD�$$L�$�SHL�T$H��L�$H+A�	   H�C0tiG M�z0E�j,D�sHCH�+����I�������I�x@H9�������  H)�H���r������I�xH��)������M��D�$$A�	   H�C0WiG ����M��D�$$����������M��D�$$���uH�C0�jG �������������n���M��D�$$���tc���uOH�C0�iG H�{P��H�SH�D$H�t$L�\$L�$��L�$L�\$�D$�W���M��D�$$H�C0�jG �������H�{PH�SH���t���H�{PH�SHH�C0�iG ��	   I�A0�iG �3�����H��)������M�x0H��I+L��E�h,L��M��L��IQ��E�qI�)I�HX������"���M��L��D�$$H+I�B    M�z0E�j,D�sHCL������M��D�$$�����L��L��M��� 	   I�A0�iG ����ff.�      AUH���  L�oATL���   USH��H��H���   H�G0�G8   �JD  �   L��H����H����   ��HEL�c�S 1�L���+�������   ��uv�C8����   �S ��u�H�+H�E(H�uH��u�H�EH)�H=   ��   H��t<��Hu ����sW���   ��t��>A�<$���{����t�fA�t��k��� H���   H���   �U   H��[]A\A]�f.�     H�I�$��H�|�I�|�H���   L��H���H)�H)�����H�����@ H�C0H���   H;��   t#H��1�[]A\A]��    �   �   �/����U   �r����>A�<$�t�A�t����� AVAUI��ATI��UH��SH���   H��H9���   H9���   M����   E1��    H���   H���   H)�L9�r*M�L��L���G��L��   L��L��   []A\A]A^�f�L��H��I�I��_G��H��   H��I)�H��   ������t�[L��]A\A]A^�fD  H���   H�?��������   E1�[]L��A\A]A^�f.�     H)�D  H���   H���   H��H)�H9�rH�H�H���   H���   ����fD  H�H���   H���   H)������H��������u�H���   뙐H�{�����H���   �C     H�CH���  H�C0H���   H���   H���   1��C8    Hǃ�       �p���ff.�     �H��7����    H���  H���v  AWAVAUATUH��SH��H��H��L�f8�����D$���8  H�{H��1�H�    H���H�T$��   H�CH    H)���P���H�L�c8L�������L$I�Ņ���   H�XH��H�(H�C8Iǅ�       I�EI���   I���   I���   ��������  H���n���I�}�����I�EXP�E I���   H�E8I�E`0�E I�EhI���  A�E     I�E�.������6  I�} �+  �D$    L�kH�EH��L�uH�p��K�����tG�D$A����L�{H�C    H�    H�C(��E H�C0��E H��[]A\A]A^A_� �(   �f�H�t$H���S����T$L��H��I�ǅ�uR�����I�G�H=��  �+  H�T$L��L���]���H�ŋD$��t:1��n��� �D$L��L����5���D$�v�������A�����D$�?���@ L��H��1�L������I��L9�t*1�1�1�L�������H��L���5��1������D$   �I�}����I�EX    L��L��I�E`    I�Eh    I�E    I�E0    A�E     A�E8    I�E    I�E     I�E    �5��L�s�D$H�C    H�C    H�+H�C(    H�C0��E �����D$M���X���A�����M���f.�     H��A��H����A���   H����   USH��H��xH�H�t$�/   H�|$PH��H�$D�D$�D$ H�D$@P�E H�D$H0�E �������uC�   H�������Ń�tOH���_�����t3���tf���t)1������H��x��[]��    �   H��x[]�@ H��x�
   []�@ H�D$(H��H��������@ �   �f.�     �@   �f�     S1�H��H���q�����tH��[��    �   H�t$H��������u݀|$tH���   [��     �|$��   E�H��[�ff.�     f�USH��H���G �o<�w@�WD���
  �9{�&  9�r5f����k<���G  9k0�0  �   ��H���   �SD����   �C���  �S<H���   H�s������S<HC(�C    H9�H�����҉S��    9���   )ʃ��SH����   ��   �   1�1��K�D���H����M�L�B��vL�B�R��   )���M�	Ѕ�t�������A���!ʉ���	�H��[]�D  9�� ����C<	   �	   �CD   �C  ����@ 9���������L= �   ����)�H�P�Z���@ �s8�V������S������ H���   �Ox1�H9�rUH��SH��H�lH���   H��L�GpL���   I9�t_H��H��   vH��   tl�   �   H��L�L$�   L���
��H�Cp�D$��uAH���   1�H��[]��    ��    H��   �   H�Gp    HG�1�E1�H��랸������ff.�     @ H�G    �G  H�G(    �Gx    �G<	   H�    �fD  H�    H��H�1�HǇ�       H��H���H)����   ���H�H���   H�F8H�BX    H�B`    H���   H���   �Bh    H�BpHǂ�   @   H�B    �B  H�B(    �Bx    �B<	   H�    �fD  H����   H����   AVAUATUH��SH��H��H�� L�f8�0����D$��upH�{H��1�H�    H���H�T$�  H�CH    H)���P���H�L�c8L���
���I�ŋD$��t?H�C���H�C    H�    H�C(��E H�C0`�E H�� []A\A]A^� �(   �f�H�C8I�]H��M�uI�m I�EI���  I��   I���  Iǅ�      �d�����tL��L��D$�/���D$� H��L���D$�9���L�k�D$�M���ff.�     �UH���   SH��H��H�wp�G  H���   H�G    H�G(    �Gx    �G<	   H�    H9�tH���.��H�Cp    H�sXH���{.��H�{H�    1�Hǃ�       H���H)����   ���H�H��[]�f�     ATUSH�_H��t:L�g8H��H�{�C���H�C    H��H�    L��H�C    �.��H�E    []A\�@ AWAVAUATU1�SH��H��(�GPD�wLD�oH�$H��t�I��I�ԃ�t\����   ����   �$D�kHD�sL�CPH��(H��[]A\A]A^A_�@ =   �}  �K4����  �C@    E1�E1��C H���	�����y��   �D  ���CxM��tH�Sp�A�/H��I9��x����Cx��uՋC@;C8s"D�[hD9���  H�SXfD�,BH�S`D�4�C@�   D�,$��    H���   �   ��������   H���   �   H�t$�����H��H����   �D$����������щC4�S0H��H�⍲ ����s8��wg���C<	   H�������   ��
���C@�   CЉSD�����=�   w*M��tA�I���!  �   A��A���$    �����$    �1��   �W��� ��=�   �@  �$�KxH��H;��   �}  H�sp��A�։Cx��   ����f��C@�   �$   ���  H�{X uD�H���D  H�{`��   ��H�sp�CxH���H�CX�P���   �w���H���	����KxH��H;��   r�H�߉T$������������Kx�T$H����    H���   E����   D����B��L$L�CXL��L�L$�   L�\$����T$H�CX��������T$L�\$H�<PJ�4XL��H�{`��8���L$�C@�Kh������ ���;K@��   �$�F����SxH��H;��   seH�Kp���CxD�4D��A���   ������y���f�     H�߉T$�����T$��x�KxH���d����   �D$   �%���A�������H���_�����������SxH���A��A���$    �Q����$�L���D  AWAVAUI��ATI��UH��SH��H�_H���  H9���   H���  H��H���   H)�H��H)�H9�wvH��H���  H)�H�H���  M���\  H��   H���  E1�L���   H)�K�|= L9��=  L��M��7��L��  L��  H��L��[]A\A]A^A_�f�H�;1����������   H�C0    H���  �C8 H�C@    ǃ�       �CT	   H�C    Hǃ�      H��   H���  1��    H9��0���H���  H��   H)�H)�H9�HF�H�H�H���  H���  H)������I��L�{A���  �6�    1��   L���q���H=�  v/H���     H��   �����I9�u�1�L��L���?���L9�sZE1������f�H��I�I)��b6��H��  L��H�{L���  �   ����H���  H�,H��   H���j������� L��  �5���@ ��G�H��H	��FH��H	�H9��H9Ѻ   G���    L�E1�I9�sUH�B�I��H��"wHAUATUSA��Cը�ugM�HL9�tQA�H�Aը�tE��-������H�I��L9�wOD  L�� L���@ E�����L�LE�L��H�؄�LE�[L��]A\A]� ������M��1�H�I���� ��   ����   ����   E1�E1�H� 6     �=f�A�   I��L9�v�A�	I��A�    I��A����!ECń��f���E���]�������G ���N���L��M9��A���I9��u8��M��M��D  A�6  E1�E1�I���l��������L�E1�����f.�     AT�
   I��USH��H�H�|$H�\$�n���H�L$H9�t9H9�rI�$H��[]A\�f��9#u�H�YH��H�|$H�\$�5���H�L$H9�u�H��1�[]A\�H�H9�sWH�6     �@ H��sAH��H9�s8��� v��%u+H9�w��D  ���tր�
t�H��H9�u�H��H9�r�H��ff.�     f�H�H9���   �E1��@ <(��   <)��   H9�sC�H��H�Q<\u�H9�t0�AD�@�A��Lw2E��B�$��G fD  H�QH9�r��    �   H���    H9�v�HЀ�w�1ɐ��H����w�H9�������D�@�A��v��y���f�     A���_����    A���N���1��H�ʸ   ��     H��H�I��I�� H��H�T$L9�s7L��H�|$�u���H�T$L9�s �
�ȃ�߃�A<v̍A�<	vŸ   ��>uH��1�I�H���ff.�     f�SH��H��H�H�T$H9��  I��E1��<�    <%��   <(uLL��H�|$�_���H�T$����H��H�T$L9�sA��t=�<<tLv�<{��   <}uA����   @ H�T$�   1�H��H�T$L9�r�E�۹   E�H�H��[�f�L��H�|$�����H�T$������    I9�w� f�     �<t<
tH��I9�u�L�ҹ   1��H���D  A���o���H��1�H�H��[�1��ff.�     �UH��SH��H�_H�H�|$H��H�D$�����H�T$1�H9���   �
�q����   ��   ��{��  ��(��  ��<�  ��>��   ��/�?  �� wH�6     H����   H�     � PH�rI�6     �ȃ�߃�[������>wH��H���	Є���   H��H�t$H9��H  �H���� w�I��H�rs�1��fD  H��H�T$H9�vH9U �   D�H9�sH�] �EH��[]� H�\$�EH�] H��[]�D  H�JH�L$H9���   �z>t/H�ʸ   �fD  H�T$1���    H�JH9�v�z<uH��H�T$�l��� H��H�|$����H�T$�R����H�rH�t$H9�si�JH������fD  H��H�|$�����H�T$����f�     H��H�|$�s���H�T$�����f�     H�ʸ   ����� 1������H��������H�w������    AUATUH��SH��H���F    H�    H�F    H�w����H�L�gH�D$L9�sX���[��   ��{��   ��(tNH�E �8/�����D@�E�M����SH����?  H�EH���     H��t@H�H��[]A\A]�D  �E   L��H�|$H�E �p�����uHH�T$H�UH��H��u�H�E     �E    �f.�     �E   L��H�|$H�E ������t�H�UH�D$�v���fD  H�PH�E L���E   H�H�T$����H�H�D$L9�st�wA�   ��t7�eD  ��]t;H�H���P���H�sH���D���H�H�D$L9�s7�K��u0���[u�A����f�A��u�H�PH�UH�������f.�     H�U������    AWAVI��AUATI��UH��S��H��8�����H�t$�����|$tH��8[]A\A]A^A_ÐI�D$M�,$H�$H�[M�<�H�D$H�PH�D$I�$H��I�D$H9�sL���9fD  M��tI9�vH�D$ H�H�D$(H�CH�D$0H�CH��I�D$I9$sH�t$ L���p����D$0��u�L)�H��ië����E H�$M�,$I�D$H��8[]A\A]A^A_�1����     H�w�����H�w�n���ff.�      AVI��AUATUH��SH�wH������L�H�GI9�s-I��E��t2A�9<��   I��L9���   H�    I��M�
[1�]A\A]A^�f�H�T- D)�H9�HF�H����   1�E1�   1�I�6     1��fD  I��s�}H��H9�sOL�I���7@�� v�@��x>������G ��w/��	���t�A��A��}�   D��H��I��H9�r�@ Lσ�t��E�eA�L�#I�:E���9���I��M9J�%���A�9>����[�   ]A\A]A^ÐH�T- D)�H9�HF�H��� ���H�    L��H�    L������ff.�     f��G    H�wH�WH�7H�O H�G(��E H�G00�E H�G8 �E H�G@��E H�GH �E H�GPP F H�GX �E H�G` �E H�Gh �E H�Gp0�E H�Gx �E HǇ�   0�E HǇ�   ��E �ff.�     �ff.�     @ H�GH��t:H�W H�
H���   H�JH���   H�JH���   H�JH���   H�R H���   �ff.�     �H�G(H��t7H�D�@f��~0H�pH���LN���A��9���   fA���? ��    1�f��u�fA��~�M��H�xHc�M��H��I��H�J�|�L�L9t$f��~��p�~���9�t9H�@f�|P���    H�H9~u�H�pB�|�u�A��fD�@��    ��f�xf��D  ��f�ÐH�GH��t:H�W H�
H���   H�JH���   H�JH���   H�JH���   H�R H���   �ff.�     �L�G(���    I�@t-H��
H��H��
I@H��Ix��H�W��H�7�A�@��fA�@��     H�G(H��t7H�D�@f��~0H�pH���LN���A��9���   fA���? ��    1�f��u�fA��~�M��H�xHc�M��H��I��H�J�|�L�L9t$f��~��p�~���9�t9H�@f�|P���    H�H9~u�H�pB�|�u�A��fD�@��    ��f�xf��D  ��f�ÐH�GH��t:H�W H�
H���   H�JH���   H�JH���   H�JH���   H�R H���   �ff.�     �H�7H9�sF��H9�HF�H��t8��E1�1ɐH�A���A��A1��i�m�  D�A�II���X  ��H9�r�É���1ǉ���1�����1��f.�     �G(    H�G0    H�G     H�G    �H�H��  ���  H���  �O(H�G0H�B(H�G H�B0H�G1��ff.�     @ H�H��  ���  H���  �O(H�G0H�B(H�G H�B8H�G1��ff.�     @ H���,  ��0  H��8  )щWH�G 1��O�ff.�     H�G    H�G     �ff.�     @ �W1�9�wW9�v
H�G ���p�D  �D�O�PD9�AB�DOD9�sEH� ���G��u*��H��H�<W�D  D�H��E��u����A9�w�1҉�@ D����1�1���ff.�     �H���  ��H���f�L�H��I��  I���   H�@H��tA���  E1��0�E ��f��   �f.�     H�H��  �` H�H��  �` ��L���   H���  Ǉ�       H�L���  H��x
  H���  H���  H���  H9�vwM��A������L�^<��   <s[<vc<��   <u_L�¸�   L)�H���B  Ǉ�      I�@�HG@I�@�H�GX    H�GP1��D  <s�H��w��   �fD  <s�<t�<v���<���   ��u���L�����- <v�<�u�H�NH9�r��Fȍ� }  �� �  w���H��L��L)�H���  �I��H�I�@�L���  H9������t����     L9��c����~�Y���L�¸�   L)�H��U� L�^L9��7����v<�w���   ���DlL���F���fD  ���   ���1D��)Ɖ�L���%���D  �Ǉ�      I�@�HG@I�@�HGHI�@�H�GPI�@�H�GX1��f.�     D�G E����   � ��   �G$A����PH��H��9t8��D9�r��tC��H��H��D�D8D9���   ��H��H��H�L8�D  H�� D�A A9�~{���Ѕ�u�O8���W<�G$    )�H�9�K1�H��Hct@H��H��H��?H�� �  H����fD  HcGHc�H��H��H��?H�� �  H��ÐHcw�f.�     �щG$H��D)�H���T<Hc���     AVI��ATUSH�����t�I�����   1��	@ I��1�E�Y E��E����  A�y8A�r9���   I�IX1�� H�� �y�9���   ��D9�u�I�y� t
A���   A�C�H��A�D<A9B|[E�A E9��  D��H��H��A�D<����  A9B1A�p�A���   w$D��E��D)���   D  �   �F9B�<���H��[]A\A^�1�f�9�t��t9z}��H��H��A�D	u�I�y� tjA�udA�Ä��x  rH�$�����������H�$�J��A+r�����Icq��Hc�H��H��H��?H��1 �  ��H���)�A�r�BD�؅��X  E�A E1�E9������A�p�E�Ą�tE��A��A���   �'���D��D��D)�tN��A)�)�@ ��A�0��H��H��H��H��L�L�L�qL�pL�qL�pL�qL�pH�I H�H 9�u�H��I�
H��I�9H�HI�JH�HI�JH�HI�JH�H A�D$A�A �������A�CH�
A��H��H��L�H�HH�JH�HH�JH�HH�RH�P E�a H��[]A\A^�A�p�9B�	����?���H�$�5���H�$A�BD�������I�y� tE�A�������A�r�G���E1�����A������D  L�SD����)�)�L�T$A��4   ��   A��A)�D��A��E)�E��A�    A�    ���H   t~����L�_��������)�AC ��xwE���  C� 9���   �Hc�I  D9���   Hi�3�  H�H�� �  H��A�Hc�I  Hi��L  H�H�� �  H��A�[��    A�����X���fD  ��E��xiC� 9���   �Hc�I  D9�|jHi�3�  H�H�� �  H��A�Hc�I  Hi�3� H�H�� �  H��A�[�fD  A�    A�    [�A��C� 9�|M�Hc�I  A9�~W��A���I  A�[��    A��C� 9�|��Hc�I  A9��Hi��L������� A�    ��I  �A�[�@ Hi��L���<���@ �ﾭ�H9Gt�@ USH��H��H�o8H�7H������H�    H�s(H������H�C(    H�s0H������H�C0    H�C    H��[]�f.�     USH��H�GH�/H��t:H�W H�
H���   H�JH���   H�JH���   H�JH���   H�R H���   H���  H��t&H��H���  ��H���  H���=��Hǃ�      H��[]�ff.�     SH��H�wH�?���H�C    [�fD  SH�H��H�w H���   ����H�C     �C    [��     ATUSH��L�'M��t#H�o8H�wH��H�T$H�������T$H���tH��[]A\�@ H�SL��H������H�C(HcS H�3H��L)�H9�s!f.�     H�H��tH�H�H��H9�w�H�CL��H��H�C�6��H��[]A\�ff.�     f�AUI��ATI��UH���    SH��H��H��H�T$�X���H�D$��u)L�bL�"L�j�B   H�+H�SH�C    H�C    H��[]A\A]�f�     AUE1�ATLc�   UH��L��SH��H��H�W81�H��L�L$�/����T$H�C(��t#H��H���h��H�C(    �D$H��[]A\A]ÐL�L$E1�L��1Ҿ   H�������H�C0�D$��uZ�ﾭ�D�c H�K�C$    H�    H�C    H�C    H�C@��E H�CH��E H�CP� F H�CX��E H��[]A\A]�@ H�C(�T����    H��������AT1�USH��H��H�O�D$    H��H9�s%H�S1�H��t�
��u�@   H��[]A\�D  H��H�W0L�G8I��H�?L�L$�   H��������|$H�C8��u�L�c�   H�k0L9c(v�H�CH��t�0��u� �   L�c(H��1�[]A\�f�     UH��SH��H��H�(H;{t*H�SH��H��H{8�&��H�C(H��[]�f.�     H�s H�H���������t�H�{(��    AVAUATUSH�o(���    H�Eu��f�E[]A\A]A^�fD  H��I��HEA��I��H��I��Lm�`��L��H��I�E �`��H��E��I�E������E��f�E[]A\A]A^�f�     AWAVAUATUSH��8H�/H�l$(H9��Q  �E I��I��I���PՁ��   �  E1�<.�
  L��H�|$(L�D$����H�L$(H��H9��  H=�  A�   L�D$�8  L9�s	�9.�g  A�   1�H�QL9�s����<E�#  H��1�H	�I�H����   E���f  @����   M���^  H������G  H�gfffffff�8 I���.  L��I��?H��H��L)�I��I����  H������  H��H�H��H������H�l� H���fD  H�MH�L$(H9�t�U�rՁ��   u 1�H��8H��[]A\A]A^A_�@ <-A�ǀ�.�f  L9���   E1�1�A�   1������fD  ��E1�L9�����������@ L��H�|$(H�T$(H�T$L�D$D�L$�����H�L$(H�T$H9��l���H��D�L$L�D$H	�H=�  �o  I�H���C��� ����H��H��E��HE��+���H��fD  E1�1�H�MH�L$(L9��'����U�� �o  �B�<�B�@��<��@�� ����������H�EA�   1��P@ I��H��H�D$(I9��������� �  �r�H��@���r�@��@��@��@�������������H����G ��	��   I������H������H�L� H�,JH��u	M���z���O�$�M��r���ttH�����������     O�$�M�H	�����I��tJH��H��H��H��H��I�����~�H��H��H��H����f��   H=�������I�1��
���D  H���|���L��H���]��H��i���H�L$(�����H��1�H	������H��A�   1�1������H���X���H���A���ff.�     AWAVAUATUSH��8L�?D�D$E1�H�|$�T$L�|$ I9���   A�H��I��<[��   �}   <{��   I��L�|$ I9���   E1��nf.�     A8/��   M��tD9t$~rM��O�D� H�D$(H��HcT$IE�H�|$ I���E���H�T$ I�$I9���   D�D$A��@��t]I��H9�sTH��H�|$ D�t$E���g���L�|$ I9��y���H�D$L�8H��8D��[]A\A]A^A_��    �]   �-���fD  I���� 1��*���f�     I���f.�     A������E1�� H��A��H�wI��A�������H�wL��D��H���w����    AWAVAUA��ATUSH��H��   H�t$H�t$xH�|$0H�T$�������$�   ����   H�T$x�KL��$�   H�T$p�L$ ���O  �D$    �D$$   ����  B��    D�d$H�D$8C�D- �D$@D�D$XA�E��D$D@ H�t$H�L$D��H�|$p�YH�L��������D$ ��w�$�H�G �    �   H�ĸ   []A\A]A^A_�f�     H�D$0H�L$8E1�1�L�L$l�   H�@ H��H�D$H�����H�ŋD$l��u�1�A�   ��E1�D��L��H�L� H�|$p��������  D9���  L��H�|$pD��H���A��u��D$DE1�H�D$(E����   L�t$PL�t$D�d$\M��D�|$X�@ I��J�|� K����X��H�C�D% H�|� ��X��H�C�D$@D�H�|� ��X��H�CC�'H�|� ��X��H�CI�D$L;d$(u�L�t$PD�d$\H�|$HH���O���mD  E1��   H�|$pH��$�   �.����������H��$�   �hX��H�H��$�   �XX��H�CH��$�   �GX��H�CH��$�   �6X��H�Cf��D$$A��D$A9�����1��9���@ H�|$p����H�t$�V��tc���O  ���6  H�뱐H�T$pH�BI9�v	�:t��  H�J1�I9�v�:fu�za�-  �    H�t$H�T$p�V��u�f��]���D  �   H�|$p�����n���@ H�D$pL9��2���H�T$0��$�   H�J L��H)�A�׃���   ���W���H���j�D�z�H�D$pH�3H��tH��H�L$(�����H�    H�L$(H��D��H�T$l����H���D$l������H�t$pH��H�������( H����� 1�H�|$p�\��������    ��y���f�     ��i���f�     E�������H��D�l$$I�^�H�T$pI���D$   ����D  H���j�H�D$p�(����    1��zr������zu������ze�����H���   �r���f.�     L�|$0H��I�^�H��$�   M�'I�oI�L��I�_�%�����$�   M�'I�o�D$    �D$$   �z���E�������H�D$p�D$    �/���@ H�|$HH���D$l   �;����D$l�����zl������zs������ze�����H������ff.�     AWI��AVAUATA��UH��SH��H��H  H�H�D$H�FH�D$H�F�D$   H�D$ H�FH�D$(H�F H�D$0H�F(H�D$8�F��
��   ����   H�L$�    H�t$@L��������D$����   �S 9���   �{M�7M�ot�S$��uH�\$@��"�   ��D$,D$(H���D$���D$��~tH�E1�D��H��H�t$L��I�H�CI�G������t�M�7M�oH��H  []A\A]A^A_� �ЉT$�r���D  H�M ��D$�q����D$   �"��� 1��@ ��   묐AWE1�AVI��AUATI��USH��(�t$H�w�����H�L�oH�\$I9���   �<[��   <{��   �D$}H��H�\$I9���   L��E1��^D  �D$8��   M��tD9|$~W1�L��H�|$�����H�T$H��M��HE�f�H�D$H9�t{A���|$ tHH��I9�v?L��H�|$����H�\$I9�w�I�H��(D��[]A\A]A^A_� �D$]�O���fD  H���� �D$ �I���fD  H���f.�     A�������     E1��ff.�     H��A��H�w����H�wIc�H��� ���H�    I��H�1�H�G`    L��H���L�V0H)�L�N8��p���H�H�~@H�NPH�F`L�M�L�^M�XL�^M�XL�^M�XL�^ M�X L�^(M�P0M�X(M�H8I�x@I�HHI�@P��t;A�@X ���   A�@Y���   A�@Z���   A�@[A�P\I�@`p F I�@h��E ����   A�@X���   A�@Y���   A�@Z���   A�@[�f�ATUH��SH��H��H�    H�B    H�B    H�B    H�H���   H�xh t9H�L$H����x  ��uH�$H�L$H�H�SH�KH�SH��[]A\�fD  L��  I��$    tG���   w?I��$h  ���A�L$$��t*I��$   1�H�Wf;u�(@ H��f;B�t��9�u�   ��     ��x�H�}�R��� SH�Ћ\$H�    H�G    H�G    H�G    H;V(rL�V1�M��tE�E����   @ H�FHF8D�XD�PD��D)ց�  ����   ��  ��tM����   ����   �   E�ھ   ��0  D�OH�WE�HE�D�G�8 t/�@���G[�7�@ ����   DG�    D�GD�OH�WMc�Mc�[M��L��H��?I��  �  H���GÄ�t��   �   E�D�OD�GH�W�8 t��@��     A��   ����@ �   E�Ӿ   ��   �   �1�����t�   �   ��    �   �   �	����     H�|$�H�zH��1�H���H�T$�H)�H�    ���  Hǂ�      ���H�H��P  ��HǂH      Hǂ      H���)���   ���H��~@��H  ��t�     H�LFH���P  H��9�w��~	1�@��I  ��tf�     H�LF(H����  H��9�w��~
1�@��J  ��tf�     H�LF<H���  H��9�w��~1�@��K  ��tf�     H�LFXH��  H��9�w�H�FpH���  HcFxH���  HcF|H���  ���   H���  ���   H���  ���   1�@���  ��t"f�     H��F�   H���   H��9�w����   1�@���  ��t H��F�   H���h  H��9�w����   H�L$����  �F���  H���   ���  H���   H��  H���  H�D$�H���   �Vt���t.���  ��t.@ ����1Љ���1Љ���1�x�Vt�D  ���  ��u1H�T$�H�D$�1�H�T$�1Љ���
1�����1�9¸�s  EƉ��  �ff.�     �U1�SH��H��H�G�    H��HǇ�      H���H)����  ���H�����   H��������H���  H��(  H���
  H���  ���
  ��h  H���
  H��`  ��h  ��l  H��`  H���  ���
  ��@  H���
  H��P  H���
  H���  H���
  H���  H���  H���  ���  ���  ���
  ���  []�f.�     H��1������H���   H��  H�  H��(  H���  H��   ���  ��D  H���  H��X  ���  ��L  ���  ��@  H���  H��P  ���  ��H  H���  H��0  ���  ��8  ���  ��l  H���  H��x  H���  H���  []�ff.�     SH�_(H��tn���    t=H��W�G`�D;Gw8H�f��~�sH�K�V�f�TA����f�1�[�f�f�1�[��     1��   ������t�[�fD  �   [ÐS���    H�_(tbH��W�G`�D;Gw-H�f��~�sH�K�V�f�TA����f�1�[��    1��   �D�����u�H�f�����D  f�1�[��     AUATUSH��H��Ƈ�   H���   Ǉ�       H�wH�OH�H��t\H��(  I��H��E��H�8H�GH�{H�C H�G`H�C(�W��I�EPH� Hǃ�       H���   E��tH��(  H�@@H���   H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    Hǃ�   @	F Hǃ�   @�E Hǃ�   @1F Hǃ�    �E Hǃ�   `1F Hǃ�   @F Hǃ�   �1F Hǃ�   ��E H��[]A\A]�ff.�     �AU�   ATUSH��H��f���   H���   H�wH�OH�H��tuH��(  E��I��H��H�8H�GH�{H�C H�G`H�C(�V��Hǃ�       Hǃ�       E��t.M��t)I�D$PH� H��tH� H���   H��(  H�@@H���   H�C0    H�C8    H�C@    H�CH    H�CP    H�CX    Hǃ�   p
F Hǃ�   p�E Hǃ�   �4F Hǃ�   ��E Hǃ�    5F Hǃ�   �F Hǃ�   p5F Hǃ�   �E H��[]A\A]��     H���  ���   ��   AUHc�ATUSH��H��H�P0�<r�P(I�ŋ�h  ��tUH��`  D�`�1��fD  H�CI9�t7H��H�|� H��t�A�E 8u�L��������u�H����[]A\A]��     H�������[]A\A]ø�����f.�     AW1�AVI��AUI��ATM��UL��SH��H��H��H��H�T$D�|$P�   H�G�    HǇ�      H���H)����  ���H�H���   �׷F �z��H����   H���
  L��L��H��H�T$E���M���I�E L���
  H��`  ���
  �D$XHǃx  `F ��h  H�D$`Hǃ�  ��E H��p  1�Hǃ�  ��E Hǃ�  rF H��[]A\A]A^A_�f�H���   []A\A]A^A_�ff.�     �AV�A   1�AUI��ATI��US�/��G ������IKHc�H�<���G ��XHc�@8�u��    L��L��D�s�������t�؃�I�H�<���G H��@:/t�A�K   [D��]A\A]A^�ff.�     H�OH�f�     H9�w������G   �fD  H��H��B��� t؃�	tӃ�t��
u	�G   Ð��;u�G   Ã�t��ff.�     f��W��YH�������G��JH�H�H�B�H9�w
�F   �f�H�JH���� t��	t��t��
t��;t��t�H���� 1��D  �F   ��F   ��     �WH���������W1���?H�H�~H�B�@ H9�w�F   � H��H��J���t��
t��u���@ ��    �F   ��     AWAVI��AUA��ATU1�SH�^H��(L�g�K�L�����   �_���H�D$H��t?M�<$I)ǃ{�I�O�wT�S��$Ր�G f.�     1�H����   ���H��A9�u�H��(��[]A\A]A^A_�D  H�4H�|$�r������H��A9�t΋K�L����r����Q���H�D$�m����    M�FM����   I�V H��H��A�Љ�f�H�41�H�|$� ���H�� I�>H�T$L��H�L$�����T$H�L$H����o���H�t$H��H���?���H�B�D8� �Q����H�ƿ�G ��� �������D  �    �%���D  H��t;H�D�Gf��~4H�OH���TQ���A��9���   fA���C�    ��    1�f��u�fA��~�M��H�wHc�M��H��I��H�J�t�L�L9t$f��~��O�q���9�t9H�Wf�tB���    H�vH9qu�H�OB�|	�u�A��fD�G��    ��f�wf��D  ��f�ÐSH�_8H�{(�����CX [�ff.�     �ATUH��SH�GH���  ��0  ����   H��h  H���  H���   ���  H���  1����  ���  t�k   ���  v��l�  �%k��� �  ���  H��   H���  H��  H���  H���  1�[]A\�fD  H��h  I���H��8  �P�и   ;�0  s�Hc�H���    H���8  �@���M���7���I�L$PH�	H�D�H���   �����    I��UMc�H��Ic��H  I��Ic�SIc��H  H��D��L��H��L��H��H��?I��  �  H��?H��H��
 �  H��H����C���Hc�I�H�HcqDHcQLH��H��H��H��?I��H��> �  A���H  I��?H���J�� �  HcQHHcIPH��H���H��Hc�H�u H��H��?H��H�� �  A���H  H��?[H��]�H��1 �  H���H�I��f.�     AWAVI��AUATUH��SH��H��   H�H�4$D�D$D�L$0H�D$E��uH�� ��  H�$A�~ L�h(�  I�H�C     H��$�   I�FH��$�   I�FH��$�   I�FH��$�   I�F H��$�   I�F(H��$�   M9n�-  H�D$��A   ��  M����  L�t$ A�����1�L��$�   L�t$�0f.�     H��A���H��u
I��A�����H��L9���   E�'t�H��D�KL��H��jD�D$H�t$H�|$P����D�D$H�t$L��D�KH�|$p�$    �����D�\$PAYAZA��u�D$`�D$����  H�T$`H�t$@H������D����A �N���fD  I�H��t�(��u�    A�~ �����H�L$�y t
�     �C H�ĸ   []A\A]A^A_�f��|$0 L�t$ ��   A�����L��L�t$1�L��$�   E��I��M��D�|$�.�     H��A���H��u
I��A�����H��L9���  E�.t�H��D�KH��E��jH�L$ H�t$H�|$P�����H�L$ H�t$E��D�KH�|$p�$    ����H�T$pH�t$PH�������XZ�v���fD  �K ��t)�{8��"�A�H���t8��xH�CH�@(    �   f��CH�T$`H�t$@H��H�D$T    H�D$D    �D$XH�D$L    �D$\    �D$@1   H�D$`    H�D$h    H�D$p    H�D$x    �X����K H�CH�@(    ���   L�t$1�f.�     L�mI��L��H���D3A��A��tM��H�� L�m��  H��   A�    A�    H��D�D<L��H��A��D�L<)���DE�A���   )�AD�A9�AN�9�Nǃ�����I9���  M��A�� �  I��B9L<��  H��tH�M�A� ���A)�H��E�D9L<�  A��9�}�D3(�  D��H��D�H���t<E����  L��H��Dt<H���&  L��I��H��I��H�I܋p8A�T$89�t)֋x<A+|$<Hc�Hc��K;��A�D$@�C L��H��L9������L�kL�t$M�](M����   M�eI�{�I�m8L��I��H��     H��H��I9�w$I�EH��H��tD�8E��u� �   f.�     H�
D�BH��H�AH��H��H�H�D�J<E�E�� �  D9P<|D�J<�@tH��H��DD<L)�H��u��|$0 �f  �CA�F	 �4����     H��t6H�M�H��H��H�L�4�u8A�F89�t)Ƌ}<A+~<Hc�Hc��):��A�F@E�������������    D��H��tHH�M�A� ���I��A)�I��E�F9L<~*H��A�H��D�D<E���{���L��H��T<�k���f�9�O�A������ H���a����G���f�A��<  A��L  ���j���D�T$pD�L$PD��L�|$(D�D$D�\$4I���  ��D�T$<E��E��D�L$8A��
�=fD  ��t$D�A)�E9�D�HF�E9���  �     ��H��9���  �x u�E��t�D�E��A)�E9��D�PA�E9��A��@   L�|$(D�\$4�L$t��  ��H��A����  ��)�E���  �D$t�D$���D$`�����H�M(L�H��`�'���H�qA�  I�NH��fE�^I�vH��t,I�F H�0H��tf�� �H��H9�u��ٸ��������A D6H�$L�h(�|���fD  L�t$�K H�CH�@(    ���s���@ D�S E�������H�S(1�H�<$��    D�@� �C H�� H9��c����2H��@�� u�H�BH;G(r#L�G1�M��tE�E��uA� �   �2�    H�GHG8��
D�Bu�D�@��     L�|$(�V���fD  I��H��x  H�T$`H��H�D$`    H�D$h    H�D$p    H�D$x    �����I��X  H�t$`H������������@ H�A�   H��$�   HǄ$�       HǄ$�       H��$�   H��HǄ$�       HǄ$�       HǄ$�       ���������fD  E1�1��D3(�����)�H�{H�t$`L�d$`�T$h����H��H���t<������    �|$0 �K �����5���A��@   L�|$(D�\$4�L$Tt=��H��A����  D�D$��A���D$T)�D�\$@E��������L$t�
�W���@ �� �  D+L$8f1�E;�H  |���H��A����  ��   9�O�럋t$<�� �  f1�D)�A;�H  �������H��A����  ��   9�L������A��T$TD�\$@�u���f�     H�H��t���u� U   1��f�     H�GH��t���u� �   �f.�     �O H�WH�GH��H9�t�0H���@�   H�G�f.�     �ff.�      �O H�WH�GH��H9�t�0H���@�    H�G�f.�     �k���ff.�     H�GH;Gt>H�P�H�W�P��@���t������D���    ��    ��)�����    H�W1�H��t�
��u���   �H�WH�GH)�H��9�s5��H��P� ��t������D�Ð��    ��)�����    H�W1�H��t�
��u���   �H�WH��H+GH��9�w��H��H)�H�W��    H�GH��t���u�� �   �f�H��tKUSH��H��H�/H�wxH���3���H�Cx    H���   H������Hǃ�       H��[]�f.�     �ff.�     @ AWAVAUATLc�USH��8E����  H���   D9g �J  H�A��H�]I��L�u J�/H9��  M��M)��9  L9�H������LF� H��H��H��   H�� ���H9�w�H�E8H�T$,H�މL$L�L$H��H�D$諓��L�L$�L$H��H�E �D$,����   M����   H�UL���L$L�L$�a���H�E(HcU H�} L�L$H�4ЋL$L)�H9�sH�H��tH�H�H��H9�w�H�|$L���L$L�L$�����L�u L�L$�L$K�I���H�]H�}LE�H�E(I�L��L��N�4�H�E0H} B�������Lm1�H��8[]A\A]A^A_� I��� I�����������@ H��8�   []A\A]A^A_�@ L�u H��8[]A\A]A^A_�D  AWM��I��AVI��AUATI��USH��(L�JL+JI���l$`D��E�̓�@��u��utI���8   uSA9�vD ��L��������s��ŉl$�����H�t$L���D$ H�D$    ŉl$����A9�w�I�D$I�D$A�H��([]A\A]A^A_�f�A�? u�H��1��p���I�H��   H��  ���A��a���f�AWL���I  AVAUI��ATL���I  USH��H��xD��|I  H�t$H�L$L�D$D�$A��tL���I  L���I  I�I�M I�WI�}H9�uH9�t{I�,$M�T$D�D$D�L$)�D)�A)�A)�������A��A����A��A��H�Hc�Mc�Mc�I��I��H��I��H��?I��?H��0 �  J��2 �  H��H��)���  E1�1�H��XI  H��`I  H�D$ H�T$(A���U  E1�A����   H�D$ �<$ M�MH�L$8M�E H�T$0H�$��  H��H��8  �T���H�$H��XI  H9|$0��  H��XI  H��`I  �D$`   H�SH�t$ H��H�|$(H���RH�D$0H�T$8H��XI  H��`I  E����   H��x[]A\A]A^A_ÐA�   E1�L�t$D���I  H�L$8H�T$0D���I  H��D�\$L���D$`   ����H�L$HL��H��D���I  D���I  H�T$@����H�T$PL��H��D���I  D���I  H�L$X�\���H�CH�t$ H���PH�D$PH�T$XD�\$H��XI  H��`I  E�������I�m M�eH��x[]A\A]A^A_��    )�D)�Hc���������Hc�Hc�L��L��L��L��H��?H��?I�� �  I�� �  H��H��)�Hc���-��I�7M�$H�M�L$��D)�Hc�H��H��H��?H��
 �  I�WH����B�,D)�Hc�Hc�H��H��H��?H�� �  H��F�$Mc�I9�u����1�)�9�$I  HO�I9�u����1�)�9�$I  LO�I�E H9D$u���)�)�H�9�$I  HO�I�MH9L$uD��A��E)�)�AH�9�$I  LO��H��D��|I  �������Hc�)�H)�H�H��HH�Hc� I  H9�������L��������Hc�D)�H)�Hc�H��HH�H9������I�/M�gH��XI  H��`I  H�D$ H�T$(A���;  A��A�   D�$�o��������A�   E1�H�D$ �<$ �D$`   H�L$8L���I  D�\$H�T$0L���I  H�D$��   H�t$H�������D�\$H�D$H�t$0H9t$ ��   H�SD�\$H��H���RH�D$0H�T$8D�\$H��XI  H��`I  �r����H�t$H������H�$H��XI  H9|$0�?���H��`I  H9t$8�-����m���fD  H��8  H���Q���H�D$D�\$H�t$0H9t$ �`���H�t$8H9t$(�P���������D�$A�   �����SH��H��H���   H�@hH��t8H�xH� H�����u!H�$HcT$H�    H�CH�CH�H�C1�H��[ÐH���  H���  ��H��Hc���fD  S��pI  H��Ƈ�H  ��hI  �  ��xI   u1�ƃ�H  f���H  ƃxI   [�f�H��8I  L��@I  H�sH��H��(I  A�   ������    ATA��U��S���H   H��u{Ic�HcՀ{( ƃ�H  H��hI  H�� I  H��HI  H��pI  H��PI  t
�y	 H�kt$H�kH���H  E1�H���H  D��I  H������H��8  H��  �H�[]A\�������{���fD  ATI��UH��SH��H��PH��XI  H��`I  �( �D$@   H�$H�T$tZH�T$H�L$A��E��H�sH���>���H�CH��H���H�D$H�T$L��(I  H��0I  H��XI  H��`I  H��P[]A\� ��pI  ��hI  �����ff.�     f�AWAVLc�AULc�ATM��UL��SH��(H�� I  H��PI  H��HI  �x	 ��   ���H   ��   A�   H�D$D��A��H��PL�L$�+����L$�D$��HI  ��PI  �A��΀��H   Mc�Hc�Hc�Hc�H�t$H�T$ X��   ��xI   ��   H�D$H�T$ƃxI  ǃ|I     H���I  H���I  L���I  H���I  E��uAL��HI  L��PI  H��([]A\A]A^A_�@ E1�I9��0���L9��'�����f�     H�� I  H�{E1�H���H  H���H  D��I  �����fD  H�sE1�L��I��H�T$H��������4���������ƃ�H   ƃ�H  L��8I  H��@I  � ���f.�     AWA��AVMc�AUA��ATA�̉�UD��A��SH��H��H��PI  ��HI  H�D$$PL�L$(蟾��H�D$4��D��PD��$�   D��L�L$8������D��D��D)���H�OD�\$8������D��E�E�D)�Mc�Mc����֋�HI  )Ћ�PI  A �D$4�L$0�AǋD$<�F�)Hc�Hc�Mc���$�   ���H   Mc�H�t$@Hc�H�H�T$HYAX��   ��xI   ��   H�t$0H�|$8ƃxI  H�� I  L���I  ǃ|I     H���I  H���I  L���I  L���I  H���I  L���I  H���I  �y	 ��   Lc�$�   L��HI  L��PI  H��H[]A\A]A^A_�D  H�D$L�\$L�T$�����L�T$��xI   ƃ�H   ƃ�H  H�D$L��8I  L�\$L��@I  �&���L��H�sE1�M��H�T$0H��H�D$L�\$L�T$����H�D$L�\$L�T$������    H���H  H���H  H�{E1�D��I  ������ ���f.�     AWAVAUATI��UH��SH��H��XA�x	D��A��E�H�$D�\$A��	E1�1��D$�I�BM9�t4D�\�I��C�< F�\� t�H��D�v�'���D��A�I�BF�\� M9�u�E���
  D�l$DE����   A�$D�|$@D���D��D)�)E Hщ�D)�)ǉ�H��H�9���   �����A�$F�4(�T$H���D$<PD�L$@D�D$<�L$8�T$4�t$0H�|$����D�L$E��D���T$L�t$HD�4$H�|$����H�CH�C�D$A�$D�u H��h[]A\A]A^A_� �C���D�u D��D$�{��� A�x
 u9A�$A�x �D$HuL�D$HD�u D�|$@�D$�L���@ D�m ������    D�T$@H��D�N�����D�A�x D�ΉD$Ht�H�������D�|$@E�t �D$H�D$�����ff.�     @ H��G�Wb��;Gw1���     1��)���f�     ��t��f.�     1��ff.�     f�ATI��UH���   SH��H��������tH��[]A\��     L��H��H�߹   �D$�Y����D$H��[]A\�ff.�     ����   u1��@ ATI��UH��SH��Ǉ�      �T�����t[]A\� L��H��H��[]A\�V���fD  H�?�G�Wb��;Gw1��f�     1��)���f�     H�O(�Y H�At%H��
H��H��
HAH��HyH�7H�W� �A��f�A�@ AUATUSH��H�o(�GXH����   �Y I��I��H��tvH��W�G`�D;GwqH�E f��~�uH�M�V�f�TA��E ��f�E H�{�   ������uL��L��H�߉D$�8����D$H��[]A\A]�f�     f�E �f�     1��   �$������{�����f.�     H���   []A\A]�ATI��UH��SH�_8�{X uH�VH�6H�����������   H�{�   �w�������   H�C(�{Y H�Pu ��f�PH��f�Bf�@[]A\��    H�uH�}H��H��HPHHH��
H��
H�9H�q��KYH�S(f�@����   H�BH�u(H�} H��H��
HBH��H��
HJH�9H�q� �KYH�C(f�B���n���H�PH�u8H�}0H��H��
HPH��H��
HHH�9H�q��;���@ I�T$0�
���-����[]A\�H������f.�     H��G�Wb��;Gw1���     1�鉠��f�     ��t��f.�     1��ff.�     f�ATI��UH���   SH��������uDA��$�    I�t$(H�Vt(H�NH��
H��H��
H��H~H�H�/H�_��V��f�V[]A\�ff.�     ����    t1��@ ATI��UH��SH��Ƈ�   �'�����t[]A\�fD  L��H��H��[]A\�F���fD  AWI��AVAUATE��USH��(H�D$`E��u*�E��A��E�A��A�E�H��([]A\A]A^A_�fD  D�Hc�Hc��Hc����0D�@H�у�D�HH��H��?L��
 �  �   I��A��)�A�̓�A)�D��-��   D�ɉ�����9���   D�P�PD�pD�$A��D�P�@A���D$D9��V  D����9���   D��Ic�H��D�L$)�D�T$�D$�J��D�T$HcT$D�L$D��������   A)�D+4$Ic�Ic��;���<$H��I����Hc����A�| A�?�    �4Hc�Hc���������D  IcՉ�H����H��H��?H��
 �  H��9�����A��H��Ic������A�� D����9�}VE)�Hc�H��D�$���D�$E��t;�t$A)�Ic�Ic�D)�A��Hc����Ic�H��I���Q��A�| A�?�L���@ �|$H����Hc��.����A��,���@ ��Hc�D�\$)�H��D�L$D�T$D�D$�T$�L$�����L$�T$D�D$D�T$��D�L$D�\$�i����4$A)�Hc�D�$Ic�D)�Hc�����D�$H��I��A��Ic����A�| A�?���� AV��AUATUSH�GH���<p�S �k(��t<L�c0I��D�m�1��f�H�CI9�t7H��I�<܉�H��t�A�8u�L���i�����u�[��]A\A]A^�f.�     1�[��]A\A]A^� ���   w�s��� 1��ff.�     f�ATI��US��X���   w4H����    ����   t��H���+�����t�A�$[]A\�fD  1�1�A�$[]A\�ff.�     L�GI��A�xL���j���A�@    L�������H��u%A�xt�M��u	��     1�I��f.�     M��t�H��H��II��ff.�      AWAVAUATUSH��   H�oH����  H�t$(H��L�/A�   �\���H����   H�|$(��   H�ƿ�G �   ��� ����   A��   H�t$(H������H��tYH�t$(H��������1w܉��$���G �     H�C�   H�t$@H���D$@   H�D$�������,  @ A��   H�u8L�������H�E8    H�uHL���E@    ����H�EH    �EP    �E  H�Ę   D��[]A\A]A^A_� E1��� �   H�t$@H���D$@   �6�����u�H�D$HH�E0���� �   H�t$@H���D$@   �������S���H�D$HH�E(������    I�      � A�   H�t$0H�������H������H�t$0H�����������7������$�P�G f��   H�t$@H���D$@   �����������D�T$H�fD  1�H���v���A��H��t>E����%fD  H�t$@H���S������*  ���!  H�t$@H���4���H��u�A��   ����@ �   H�t$@H���D$@   ��������C����D$H�E ������   H�t$@H���D$@   �D$P   �D$`   �D$p   �����������H�D$HH�EH�D$XH�EH�D$hH�EH�D$xH�E �g���@ �   H�t$@H���D$@   �^�����������D$H�����2���A�   ����@ H�C�   H�t$@H���D$@   H�D$�������\����D$H���P���H�T$�BP��  E1��;D  H�t$8H��������H�A����7����L��H�� @ ��  L���^  H�t$8H������H��u������ A�   ����D  �D$H�������H�T$�B@�  A�����H�t$8H���k���H�������H�t$8H���U�����tv��8t9��Kt����������s���H�D$A��D�`@�9����E1�������     H�L$A��D;a@�=���Ic�H�t$@H��H��H�A8�D$@   �D$P   H�к   �D$`   H�L$�D$p   Ǆ$�      ������������D$HH�L$�H�D$XH�AH�D$hH�AH�D$xH�AH��$�   H�A �����H�;1҉�L�L$@E1��(   �#���H�T$D�d$@H�B8E��������}���H�;1҉�L�L$@E1��   ����H�T$D�d$@H�BHE�������H���H�D$D�D$D9`P�.���L��   H�t$@H��H��HHH�D$@   H�L$�D$P   �D$`   �D$p   ������������T$HH�L$D�D$��T$X�Q�T$hA��%tN�QA��"uA��u<�D$x�AI������������H�D$Ic����E �   D�`PH�xH�����P���1����A    �Q��     ATI��1�E��UH���  E��SH��H��H�G�    H��HǇ�      H���H)����  ���H�L��H������H��@  ���   H���   H���  1����  ���  t�k   ���  v��l�  �%k��� �  ���  H�D$ D���  H���  H�D$(H���  []A\�f�     H��`wjH�B�  H�WH��f�OH�GH��tGH��tBI��1��H�PH�V� A�D H��I;Hs!H�FH;Fr�H������A�D H��I;Hr��@ H�H��t�0��u��    �ff.�     AUATI��UH��SH��H�_8�{X uH�VH�6H��������uH�{�   L�mH�m������tI�T$0�
��u�H��[]A\A]ÐH��L��H��H��[]A\A]�����     H�GH;Gt6�x�t H�W1�H��t �
��u��   ��     H�P��@�H�W�@ H�W1�H��t��2��u���   ��     AWAVI��AUATUSH��H�wI��H��Hd  H���   L�'�8H�T$PH��$�  L��$�  H�D$@H��   H�L$X�   D��$�d  �|$LH��  H��1��H�D�D$pL�ߺ�I  D�L$|H�t$hH��$   HǄ$�       Ǆ$�       HǄ$�       HǄ$�       HǄ$�       L��$  HǄ$(      HǄ$0      HǄ$8  
   HǄ$@      HǄ$H      H��$`  H��$�  H��$�   1�HǄ$P      L��$X  HǄ$h     HǄ$p      HǄ$x  
   HǄ$�      HǄ$�      HǄ$�      L��$�  HǄ$�     HǄ$�      HǄ$�  
   HǄ$�      HǄ$�      HǄ$�      HǄ$�       HǄ$�       HǄ$�       HǄ$�       HǄ$�       �J���H�T$P�|$LH��$�  H���H  A��   L��$�  H��$�J  H��$�2  H��$�  A�F,H��$�  H��$�J  H��$�J  H��$�2  H��$�  H�T$X��$Hc  A�F4��$�J  ��$Lc  H���$�2  H�R��$�  L��$c  L��$c  HǄ$c     HǄ$(c  
   ��$�J  L��$�J  ��$�2  L��$�2  ��$�  L��$�  ��$Pc  H��$Xc  I��8  H��$�c  A��  H��$`c  H��$X  ��$jc  A��0  H��$pc  H��$�  ��H��$xc  H��$�   ��H��$�c  A��,  ��$�c  1�)ȉщ�$�c  ��Ƅ$kc  1�D��$�c  Ǆ$�c  �  )�H�L$@9�L�H��$�d  �A�~ ��$�c  H��   ��$�   H��   ���A�~ ��  H��  D���  D�l$`L��(   H��$X  Ǆ$X      �/n����$X  I�ǅ�uL� H�D$hI�G�   E1�L��1�L��$X  L���H�����$X  I�G���  �T$`I�GH��$0  A�W �R  HǄ$@     A�V����  ��H��$P  �D$0    ���D$ -1�D$xH�H�L$H�H�C�D$(    H�AH�{H���D$? H�yH�K�D$  �D$t    L�t$H�HE�f�    H9���   �|$0ۃ���E��t_�|$? u�؃��<t�C�<�R  f.�     �L$(��t�C�<v���    G��D$(�|$  t��������!ȃ��D$ ����   �l$�   ���Z  ���$��G E����  �    I�GH�L$H�II�GH9��?���H�\$H�AH�C���t	���.���H�D$�x �    E�����f��D$0���4  L�t$A�   E�nH��$@c  H��$c  HǄ$ c      HǄ$0c      HǄ$8c      茲��H��$�  H��$�  HǄ$@c      HǄ$�      HǄ$�      HǄ$�      �G���H��$�  H��$X  HǄ$�      HǄ$p      HǄ$�      HǄ$�      ����H��$P  H��$  HǄ$�      HǄ$0      HǄ$@      HǄ$H      轱��HǄ$P      M��t"I�I�wH��蝱��I�G    L��H��花��H��Hd  []A\A]A^A_��     A�0   �D$`0   �n���D  �������I�GI�GH�D$H�H�Y���f�     H�L$H�QH9��.  H�BH�A�2H9��:  H�L$H�PH�Q� ��L��	��������=  D  I�GI�oH)�H������)�9���   I�GH�D$H�H�������L�������$�d  A��A�ƍED��A��L��������D$|D��A�������uF��{����u��A��m���H��E��D��ATF�,D��D��E��H��$�  �g���D��$�   D��$�d  ^_9���  ��D��$�d  D�M)�E����r����M���D  I�GI�oH)�H������)�9�������D�M)���   f.�     D�\$|E��L���������$�d  D��A�������uA������u��F�����H��E��D��F�, D��D��AUH��$�  ����D��$�   D��$�d  AXAY9���  ��D�M)��s�����L���9���D$|A��A�ÍED��A���Y����I�oI+oH��A�����  E1�D  D��L��A�]�����A�uD$|������t$|�$�d  H��$�  ��$�d  �3���A�EA��D9�r�9���
  �    L���������sD$|A�������s�$�d  A���}����sF�4�q����sF��e����s��F�,0�V���H��E��D��B�, D��D��UH��$�  �T���D��$�   ��$�d  AZA[D9��p����S
   I�GI+GH����v��$�    �  H�\$@Ƅ$�   ��8   tML�t$E1��  fD  I�GI+GH�����k  H�\$@Ƅ$�   ��8   u�L���5����$�d  L���&������  D$|�ƉD$|����  I�GH�T$H�L$D�b�RH�yH�I���� I�GI�OH)�H����v��$�    �����H�D$H��D��L��j L��$�d  H���   L��$�   H��$�  �����]A\H�D$@��8   ����H��$�  H�$�  ����  H�\$1��  H��$X  �H�L�t$H��$�   HǄ$�       ��   H��$X  HǄ$�       L����$q  �D$LHǄ$       ��$t  H��$�J  H��$`  H��$c  H��$h  H�D$hHǄ$      H��$�   HǄ$      ����H��$�   E1�E1�H��$�  H��$X  H��$X  �2���I�GD�c�SI�~I�N����f�     H�D$�x �q���H�D$H�xh �����H�X`H���   ���   ���   H���  H���P��t-H�D$H��H���   ���   ���   H���  �P ���	  L���������9D$`��  L�t$A�   A�F���H����G���@ H�D$�x �����H�\$�{a ����L���������E  H�T$���   I�G�q���fD  �|$? �i  E���`  ��$�d  �t$|H��$�  �����H�D$h�\$0HǄ$�       HǄ$�      HǄ$�      HǄ$�       HǄ$�       HǄ$�       HǄ$�       H��$�   Ƅ$�   ��ttH��$(  Hc�D�S�H��$P  H�A�L��$@  H��L��$   H��L)�H��H��    I��I9�wI��M��tE�E��uA� �   �H��H)�H9�u�L�T$H�\$H�T$�D$0    I�G�D$?H�KH�{H�KD�b�R�X��� I�OI�GH)�H�������Å���   E1��2@ D$|��$�d  �D$|��H��$�  A��������A9���   D��L���'�����u��$�d  �t$|��$�d  �D  I�OI�GH)�H���Å�t[1퐉�L��������uD$|��������t$|�$�d  H��$�  ��$�d  �&���9�r�H�D$I�OD�`�PH�D$H�xH�D$I�OH�H����fD  I�GI+GH����v��$�    �`  H�\$@Ƅ$�   ��8   �l���L����������  �$�d  ��$�d  ��������t$|H��$�  �0������� E���/  ��$�    �����1�H�\$H��L��D��PL��$�d  H���   L��$�   H��$�  ����AYAZH�D$@��8   �����H�L$I�GD�c�SH�yH�I�T����    E����  ��$�    �)���1�H�\$H��L��D��PL��$�d  H���   L��$�   H��$h  �s��� I�GM�WI)�I����D��A�ƃ��A)ʉL$HA9���   �-����    D��L��E1��������D$|D��$�d  A�������B�D�ƉL$d�������F�(�����L$dB� ��A����  H��D��A��D��SH��$�  ������$�   E�≜$�d  ZYD9d$H�  D�L$HA�jE�BA�ZE�bE)�E���S���D��L��D�\$|A�   �5������$�d  A���$���B�D�ƉL$d������F�(�	����L$dD�Í,A���P���D��������L$dB� E�b�7���@ HcD$0�������H��H;�$@  r$H��$   1�H��tD�*E��u��   �    H��$(  L��H�$P  H�D$�
���H�T$�z t/H�T$@H���  H��t���W��H�¸����H��t
��     ��H�\$H�    H�C    H�C    H�C    �k  H�|$@�H  ;�@  �����H��P  ��H��H�K�\ ��  H���  H����  �<�H�H�{�  f�E���w�����$hc   �(  H�L$I�GƄ$�   H�I�\����    I�GI+GH��A�Ń��  �   �\$H�D  ��L���u��S����u�D$|A���D����u��$�d  A���2����u�F�4�&����u�F������u�F�$0����H��D��E��B� D��D��SH��$�  �����ED��$�   ��$�d  A^ZD9��n����\$H���  I�GI�GH�D$D�`�PH�D$H�xH�H����f�     H�L$H�AH9��f  H�|$�T�����A���Q����  �$��G  I�GH�T$H�L$D�b�RH�yI�GH�D$H�H�<���@ �   H��$  �F��������������f�     �À���$  H�t$H�V�����  ��	�����H9��7  H�|$�����tlL������������D  ���D$0H�H;�$@  r-H��$   1�H��t�)��uH�T$��   D�b�RD  H��$(  H�$P  H�xH�HH�D$�]���D  ��$�    �����1�L���0���H��$�d  D$x��j���D  H�PH�Q�A������D  H�L$H���������H�yH�AH9������H�|$����������H�D$@H�@@� �����H�D$@H�@@�@�H����    H�T$@�L  ;�D  �Y���H��X  ����H��H�KH�KH�<�H�{H�D$�D$0D�`�P�j���f.�     L�������H�\$@H�H�SHH�H�B    �����H�K@��Hc�H��{[ Ƅ$�   �2���H�L$�|$? �Q��  D$|H�L$I�GD�aH�L$H�yH�I����fD  ��u���L�����������D  D�������L$dE�b�,�������$�d  H��$�  ���������    L��L��E1�A�@   �\����:����    ����*  �������H9���  H�\$H�BH�C�������L��)��D����g�����H�<�H�D$H�xH�D$H�H����1�L�������H��$�d  D$x�����1�L�������H��$�d  D$x������A�   A���G H��$�  H��$�d  L��H�t$|���������H�BH�F������E1�A� �G ��E1�H�t$|L��A��G H��$�  H��$�d  ����������E1�A� �G �D�aH�L$I�GH�yH�I�����H9��o  H�L$H�BH�A�
H�\$H�SH�CH9��-  H�zH�{�2H9���  H�\$H�WH�SD�H9���  H�\$H�BH�C�����H�\$	�A��D	�	ƀ{ �7  �� }  �   L��=�  �D$ CD$ ����H�D$D�c�SH�xH�H�r���1�����1�����H�D$�x �����A��%�����H�T$D�bE���x  �\$(����  A����  H�L$I�G�D$(    �RH�yH�I�����H�\$H��$�   H���[���H�T$I�GH�{H�KD�b�R����L���������uD$|�����t$|�$�d  H��$�  ��$�d  ����������H��$�  �$���H�D$D�`�PH�D$H�x����H�D$M�_A�   M+_D���   I��D��E)�B�,A�����   �\$HL�t$@ I���   D��L��H�X����A���   A��vKD��E��A)�@ L��H��D�V�����HcS�H�D��H��H�H�� �  H��A�C�A;��   r�E��I�WI�GH)�H��A9�wFD��H��D� �@    A��A9��`����\$HD��L��)������H�D$�@a����f�     L���H�����H�|$��������H�\$@�    D���  E��I��  H�\$��Hc�H�H�KH�<�H�{�����H�|$�Ӿ���.���H�\$H�������H�SA��H�C�����H�\$H��褾��H�{��H�C�����H�|$苾��������L���,���I�WI+WH�������������  1�9�s��)�L���k�����L�����������I�GI+GH��L�t$�����u��$�    ��  H�D$@E1�Ƅ$�   ��8   �������$hc   ��  E1�fA�~ �����I�GI+GH����������|$p A�   �����L���]���A���U������^�����$�d  �R���H�|$@H��$X  D�ƉD$|�I���A�Ņ��a���L��$�   A�   L��AT��$�d  PD��$�   H�L$hH�T$`H��$h  H��$p  �<���L�l$PH��$x  H��H+�$p  I�}A���  ��L��H��$h  �ǟ��Y^A�Ņ������ATE1�A�   L��j H�L$hH�T$`H��$h  �����H�D$PH��$x  H��H+�$p  H�x���  XZ����f.�     ��w	���$� �G H�L$H�T$I�GH�y�RH�I�Q������D$tH�D$�PH�D$H�xH�H�s�����!w����$���G H��$�  ������9���A��L�t$�	���1�L���,����l$x�H��$�d  �(�����E���l���L��1������   A��������   A�������   A���ݼ��I�OI�WH)�H������   A�D���A    D)؉A�   L��襼��I�OI�WH)�H������   E)��A$    A)�D�I H�D$@A��H�@@uu� H��$�  H�\$�SH���   �T$HL��ASPL��$�d  �|$XL��$�   �o����|$? �����L��輻����$�d  谻���D$|H�D$@ǀ�      �����@H��$X  ������e����ܺ���%���E���Q����D$t���>����|$( �����l$(HcD$(����   �8���E������L��� ���A������Lc�I�GA���\  D���$��G E���,���H�D$@H��   ���  ����1��҉���1�����1��r���  L��艺��H�D$�D$(    �D$t   D�`�PH�D$H�xH�H�
���A�������苺��A��胺��A���{������t���E9�LƉ��H�\$@H���   ����A���u����8������h���9��  �\���H�T$@H�H���  H�4��L���H�\$@H���   �2���A���(��������Hc�������9��  �����߹��H�T$@H�H���  H��H�D$�D$(    �D$t    D�`�PH�D$H�xH�H����A�������菹��Hc�臹���������Hc��7���������A��������a���Hc��Y���H�H��H�H�� �  H���o���A���^����1������*���)����P���A���?���������������3���H�\$@A��L���  ����M�������������� ���A��;��  �����H�L$@H�I��  H��H���  H�<��D��������H�T$@H���  H�������1�A����E�L�A��A9������M�WI)�I��E)�G�$
D��D��L��D�u�詸��A�   A���4H��  D��L��H�,�舸��H�Hc�A��H��H�H�� �  H��A�C�4D9w�I�WI�GH)�H��A9��|  D��H��D�(�@    A����E9��q���D��L��D)��{���H�D$�D$(    D�L$tD�`�PH�D$H�xH�H�����I�G����E��������|$? �����H�T$@���   ��������  �C���  �C����x���H�D$@�   H�x��������R������~�D��P��L$|��Hc�H�����   ��$�d  ����   ��t	������S��$�   P��$�   ��$�   D��$�   D��$�   ��$�   H��$�  �1���H�D$ D�`�PH�D$]A]H�xH�H�D$(    �D$t    �����E��������|$? �����H�\$@�   H�{�����������Hǃ�     �s���A���^����|$? �b���H��$�   1��
   HǄ$�      HǄ$�      H���H�D$hƄ$�   H��$�   ����A�������|$? tH�D$@���   ��������  ������t$|L���i�����$�d  �]���H�D$�D$(    �D$t   D�`�PH�D$H�xH�H�����H�D$@H��   ���  ����1��҉���1�����1��r���  �-���L���.���A���&���A������������E9�LƉ�����L��������������H�����  �����L�������Hc��۴�����z�������  �n���E���{���L��赴��H�\$@H�H�SHH�B衴��H�SHH�H�蓴����茴��H�S@�
�Hc�H�
�JƄ$�   �Hc�H�J�{[ �����H�L$�|$? �Q�e���D$|�$�d  ����E�������H�D$@L��L�t$L�@����A�������������D$����Hc�������|$p �D$����H�D$@�x[ ����H��`   ��  H�D$@H�@@HI���   H�xh �T  �������E�������H�D$@�xZ �{  H�H�   H��(  H�L$ H�H��H�T$�k��H�T$H�L$ ��A�������H���   HcD$H�L$(H�T$ �.H)�f�FH��H�F    D�f0f�F4 H�t$����H�t$Hc|$H���F8H�t$����H�T$ H�t$H��H�L$(�F<H�BXǁ�      H���   ǁ�   pmocǂ�      �����E�������E�������A���   �   IN��D$(L����   I��;t$(�$  L���u���A� ����L���ű������L�l$@��L��豞��D��L���褞��A������I���   H�xh �W���H�D$@H�@@H�e���L�l$@I�}�����I�}��L�l$@H��$X  蓻��A�Ņ�����H��$�   A�   L��E1�Uj H�T$`H�L$hH��$h  �
���L�l$PH��$p  H��$x  I�}H��$�   H)�H���   ��$   ^AXH�@hH��tH�xH� H��$�   �PI�}H�T$@D��H�B@H�RHH�H�L$0H�HH�L$(H�
H�RH�     H�@    H�T$ H��$X  H�L$踺��A�Ņ��@���U�D$A��A�   L��PH�L$hH�T$`D+L$ H��$h  �/���H�D$PH��$x  H�PH��$p  H��$�   H)�H���   ��$   ZH�@hYH��tH�xH� H��$�   �PH�T$@H�L$0E1�H�B@H�H�L$(H�HH�BHH�T$H�H�T$ H�P����H�D$�D$t    D�`�PH�D$H�xH�H����L���*���Hc��"���H�H��H�H�� �  H��� ���L�������������9�@��@���k�������L���ޯ������L���ѯ��1��������Hc�H���	~
��Hc��H��H��H���g���H�DH��H9�u������L��苯��=   �th�؉��r���L���s������l���)����Z���L��E��t�D$ uB�O���L��A���D���Ic�Hc���������)���L���*������#�������������	��������A��������D$  �L�������=   �tә1�)Љ������L���ۮ����蔮�������L���Ǯ���������A���x���D������L��訮��1���@�������>���L��莮����臮��	�@��@�����������L���k������d���������@��@��!��έ��������r��.���L���)���A���!����ƃ������H�D$M�_H�xH�HI�GL)�H��9���   D��E��xw���H�D$D�`����   ���A�   E1�E1�A���&)�Lc�A��O��A�(A�XE�E�PA��A��D9�tWA9�uA�ELc�A��O��E�E�P�9�~���y����ؙ�����I�GH��t�8 u� �   H�D$D�`�P�����H�D$��ff.�     f�AWI��AVAUI��ATUH��SH��   D�g\�D$4    E��tH��    ��  M��(  I�H���	  I�L���   L���   H���   H���   H�l$xH��$�   L�D�BpI�WH�D$p    D�H<H��$�   ��0   ��1  H�D$X    H�D$`    H�D$h    ��  �D$X   �D$d   E���
  �C D�c�C    ��tE��ty	E��u�K�P@���   ��  �PD��  �PH��  �PL��  �PP��  �PT��  �PX�@\���   ��  ��   ��tR�l$X����  D�d$dE����  ���  ��
  ���  �Hc��j���A9���
  9���
  L���   I�H�D$P    D���   E1��D$8    D���   H�D$H    M��   �D$<    H�D$@    �C    L;��   tL���   A�   �{ uI��  D���  E���y	  H���   �@��;C\t	�C\A�   �CH�{��   ��   H9|$X�f  �   ��  ������  H�L$`H�t$XH�       H�C$    H�CD   H�KH�K4H�L$hH�sH�s,H�K<H�{L9�t	����  D���   E���Q  �  ��A��H�H�$=�  I��A��I��   �{\   �   Mk\H���  ����$  ����
  H��  E��D�\$H��,  H�D$�  D��  ��$  ǃ,      E��tE��uH��E1���D���t$�/���XZI��   H�4$H���  ������~��9�$  ��
  �  n �I�����(  ��D��  E��ǃ0      ��E������u%E��u H��H��0  E����t$D��访��AZA[D��,  �   E��uD��0  E����H��@  ��  ��H���   H����  �Hǃ8      )�ƃ4   ���  1�Hǃ�      ���H��C8��8  H��   H���  �t���H��   ��D  ���  ����H  ���  ����L  ���  D��H  D��I  D��J  D��K  ��  E1�1�M��uI��   D  ��0  ƀ�   ���  򉐜  ���  ���  ����<  H��I9���   ��<  ���X  ���P  ��H��H��H����A�҉��  ���  A)�x�E9�EL�H���x������  ƀ�  ���  � L��8  A�s_A�� AI����t$XH��@  �V_�� I����T$dE���>  �C D�c�C   ����f.�     M��tsI��H���  I��I��N���  ���<  �H��H����H���F���  �����  )�x#A9�Ƃ�  DL����  �����  ��<  H��I9�u�Hc�8  �   ������<  H���  E1�H�<$��tz�    �~ ���  I��vS��0  A����A�   D�	B���  ����D�A��A)�)�AH�D9�E��DN�A9�~	���tA��I��M9�w�I��H��L;$u�Hc�D  E���%  Hc�8  9��D  ��   t
ǃP      D��<  M��tsLc�8  ��P  H���  1��!�    )�H��H�� �  f1��B�L9�t:HcI��H��H��?H��8 �  H���z uƍ� �  H��H��f1��B�L9�uƋ{���)  ƃ4   ��  L�d$8L���   H���   ǃ�       H�x�E���ATL��E1�j E1�H��H��$�   H�L$X�s����sZY����  @��t���   ����  H���   H�}(蓖��H�}�:����C�T$8����  H���   �y\ u�� �  H��0  ��H��H�H�Ę   []A\A]A^A_�D  ����M��tBE1� B��͈  A����A��A)�A)�EH�9�A��DN�E9�~
�>E��tXD��I��M9�w�I��������  ��A��A)�)�AH�9�N�9�������>I��H��L;$�l���������    1��@ 9��~���E���k����y���f.�     M�I�FP F H�T$4��  L��L�$�o9��D�L$4I��@   E�������I��(  L�$H�L�E��uI��  H��h  H���  H���   ��Hǃ�       Hǃ�       H���)����   1����H�H�CL���   H���   Hǃ�   �F Hǃ�   �AF Hǃ�   `3F � ��� E1�H�$   A�   A��  ����@ A��Hc�H�L$(Mc�H��H�T$ L��L�D$����Hct$L�D$H�T$ H�L$(H9�I����  ǃ,      ��$  A���  �����H����E1�E���t$D������Y^����H�s1�H9t$`���������f.�     ���  �C �C    �S�����fD  ���  �C �S����D  ƃ4  1�����f.�     Mc�   L������H9��G  ��D  Hc�8  9������ƃ@  Hcտ��  �������  )Ё��  ��  O�P  ����@ H���  D�$E1�1�H���  H�L$@H�t$<�PP�C���  I��   A��  H�L$@�T$<�UD�$��t I��  �T$<L��A�   H�L$@�UD�$I��(  �Ca I�H�ChA��  ���   �D$<���   H�D$@H���   �����@ ��   �'���fD  H��L��H�L$������$  H�L$ǃ,      ��A����������� L��   �S����ŉ�D  �a���fD  �   ����fD  M��tcE1�1�I���S�����P  ��=  ���?�����X  ��=  ���+�����`  ��=  p������h  ��=  p����@ Hc�8  ǃ�  ����ǃx  1   H��H�򉳐  H����p  H)�ƃA  ǃX  2   H��H)�H��H��?H�� �  H�� �  f1�- �  ���  ��0  ��  pHc�h  H��H�H�� �  H�� �  f1� �  ��l  �����fD  �   ����fD  H�4$�  K D�D$D�\$�����D�D$D�\$��$  ����� �  K �������(  �x���f�     �$   �/���fD  ���ωЁ����%���9�t�   w���    9��9Ѻ   G��f�     H�W �GH��H������H�rpH��H�<9�t^E1��,fD  H9�t;9�v.H�WH9�r.H��H)�H��H�<9�t-%���9�u�H9�tI��H�O�H9�s�1�M��u	��     L�ǋG�1��fD  S�_�����   ��L�_ D�@���M��A�
A9�txA��1�1��*�    v^�zD9�s0D��)���:M��H��A�
D9�tE�����A9�u�A��A�BD9�rЅ�u.E1�9�s'I��[D��BA�����D��D  A��� A�BD�[�1�E1�����   ��  w��H��?�wH H�yH Ð���  w��H��?�tH H�yH �fD  1��ff.�     f����G �6���fD  SD��4   E1�B����	H���G f����D����G L����G D����A9�tP~E�@  f�     A�	���H���G f����D����G L����G D����A9�tc��A9�|�1�[�H��H9�s/D��E�B�I�BE��A��E�ل�yID9�u�I��H��H9�u�1�E��x�A�z y�A�B[f�����@ ��D�JA9�����1��D  I��E��IH�H�PE���t���D�@fA��E��M����G E����G E��A��D9��z���E�C�N�L@�'�f����D����G L����G D����9��H���H��I9�u�1��������\���f��<utQ����   �WH����     ��.uH9�r�VH����u�H9�sv�0�����    �#���   ��D  �W��nt_L�GA�Ҿ   1�E��A�IЃ�	vA�I���w/A�IɃ�w&��I��E�ȃ�u�E��t�A��.�d����1�Ã��V����᐀iu�H�OL�O1�D�A�pЃ�	vA�p����w���A�pɃ��j�����H���L9�u��O��t��.�K����2����@ AW�B
AVAUM��ATA��1�USH��H��   �F    H�F     L�L$<H�t$�   H�L$H��L�D$E1�H�|$ H�D$@    H�D$H    H�D$P    H�D$X    H�D$`    H�D$(��N��H��H�C �D$<���  E����  1�f�     ��L��H�D$��I��H��tZE1�1��D  Jc<���G H�� �G L���Y�������   I��I��
u�L�������������   H�D$H��tL��L���Ѓ�A9�u�H�D$�L$@H�x 1��f�     �L@��u����G H���E��Dh�E�H��H��(u�H)�H������   A���A9���   �p�F �   H���J����D$<H�L$�iH�Ę   []A\A]A^A_�@ J��    H�D$@HЋ���'����    L���\h��������������1Ҿ�  ��    �4���G 9�tH��H��
u�E H���]������@ �E H���]��D�@   �����1�H��������    H��H�|$ �Ct��H�D$��   H�@     �D$<��D����� I��H�T$(H�|$ H��L�L$<�   �L���D$<    H��H�D$H�x ������     SH��H��S���H�C    H�C    H�    [�f.�     H��uH9wrEATUH��SH��L�gH9wu!L��H��H��[�   ]A\麂��f.�     1�L��������@ �   �f.�     H��騁���     H�������     H��H���%���D  H����   USH��H��H��H�s �0�H H�C    H�    H�C    H�C(    H�C0    �&���H�Ÿ   H��tB�   1�H���j���H���"���H�CH��t)1�1�H���M���H�k1�H�C(��F H�C0��F H��[]�H�������H���Q   []�@ �(   �f�H���    貀��H��tH�     H�@P�F H�@p�F H�@`�F H���f�     �����f.�     ��ff.�     @ 1��ff.�     f�1��ff.�     f��ff.�     @ �f.�     D  H��t'H�    H�G    H�G    H�G    H�G     � ��ff.�      AWAVAUATUSH���D$    H����  H����  H���  H9��6  �^�BA��A��A��A��A��A��H�~ ��   H�Չ�D�.I����L�EH�?1�)�Hc�L��M���V  ����1ȉE )�Hc�H��I9���   I�$H�E I�D$H�EI�D$H�EI�D$H�EI�D$ L�EH�E E9��  �E I��M�d$I�ݍx�H��H��I���u�$fD  ��L��L��H��I��~��I��M��u�D$H��[]A\A]A^A_��    H�H�H�FH�BH�FH�BH�FH�BH�F H�B E9�t�ۉZ1�H��[]A\A]A^A_��    L�L$L��   �G��H�E�D$��u�L�E������H���   []A\A]A^A_�@ H���!   []A\A]A^A_�@ H�T$L���G��H�E�D  I�t$L��L����}���D$�a���ff.�     @ AVAUATUSH���D$    H����  H���z  H���q  H���VH��D�mL�EH�Ѓ���vL�D$   �SL�c��y�����Hc�I)�E��y�M ��D��Mc�M)�<�  �$�8�H �    D��D��H�?�E���61�)C�U �u �ED�KA��E�ͅ�~D�ș������   ��D�Ҿ   A��L�L$�1F��I��H�E�D$����   D�ME���1  D�m�C�8���@ �;�   f�U��tq��C������  �r�1�L�N��     H��A�������A�@A�T@H�PH9�uދCK�K�H�t����HcCI�HcEI���u�@ �D$H��[]A\A]A^��    ��)�E�,E�������     D��   f�EE��t��    �C1�D�H���u�qf�     H��E�\�1�D��E��tEA��A�D�A�T�H��H��H��Hi�|  Hi��  Hi�m6  H�H�1�H��A��)ǉ�A�0H�FI9�u��SHc�I�HcEI�A���i�������@ D��   f�ME������ �C�����2  D�R�L��L��I��O���H��H���Ɖ�����@�r����������J����B�@�r�L9�uʋCM���s  HcCI�HcEI�A��u�����f�D�+�   D�sf�uE���g����    L��L��L���bz��I��HcCI�HcEI�A��u��6���fD  D��   f�}E������ �S�����:  D�P�L��L��I��O��     �H��H���ǉ�����@�z������J���@�z�������@�z�������@�z�������@�z������������B�@�z�L9�u��SK�Ѓ�u/HcCI�HcEI�A���O����b���f�A��������     ��A�	H�t@ ��H������P�H9�u�� ��A�I�L��I������A�A�I9�u��g���f�H���   []A\A]A^�fD  H���!   []A\A]A^�fD  L��M���A���D  M��M������D  L��L������D  1�H��t���   stibt�@ H��(  �Bu�SH���   H��H��0H�?H�D$    H�T$H�D$    H�D$    H�D$     H�D$(    �r�����uGH�T$H���   H�T$H���   H�T$H���   H�T$ H���   H�T$(H���   H��(  �JH��0[ÐH��tKH��t>SH��H�?H�v�i��H�    1�H�C    H�C    H�C    H�C     [� �   �f��!   �f.�     H���  H���  H�~ �  L�B �   I��I�����nL�A I��I�����]�� AW�� 1�AV��AUATUS������H��x	ʉ\$�L$��   ����  ����  �VH��H�����J  ���$�x�H �fD  A��D�A��H��A����_  D�t$H�t$(�L$�   HcSD�T$0L�D5 ��tEf.�     ����Hc�E��t&H��M��H)�I)��    �2
H��I9�u�HcS��D9�u�HՃ$��<$9���  T$�T$�D$C�D$�1�H��x[]A\A]A^A_ù   H�T$HH�D$H    H�D$P    H�D$X    H�D$`    H�D$h    �?�����u�H��H�������H�D$HH�H�D$PH�CH�D$XH�CH�D$`��H�CH�D$h��H�C �D$�sD�c�D$��H�E ��H�D$A�ϋA1�A��A)π���  ���$ո�H �   ø!   ø   �!����|$A�   F�t'A��D�L$E���a  E9��X  �|$B��    H�kB�'A��9��A  A��E����A� �  A��N�|5 A��I���  H�$D�ŉ��M�M�����  L���tE e I�}L9�s�L��1�H)���u���΋|$A�   F�t'A���N����|$�   D�f��NǉD$�D$�D$H�E H�D$��vA������A��A1�A)׋|$A�   F�t'A��������D$�@�D$�D$�sD�c�D$��H�E ��H�D$A�׋A1�A��A)׋|$A�   F�4'�����D$�@�D$�1������   �����|$L�L$HE1�1ҍD��H�|$H���)=��H�ŋD$H���p���D����{D��E��L�kL�H�$�D$A��A��A��D)�H�D$ ����  L;,$�3  Ic�I��H�D$(��H�D$0L�H�D$8L��L��L���=s��H�T$0K�<'1�Ll$(�8t��L|$8L;,$r�H�T$ 1�L���t��H�sH�|$�d���sH�k���:  D�s�E���  �T$A��Hc�HՅ������A�~��t$�$    A�   ��Hcǉ|$ ��H�zH�D$�D$�t$0H�|$(��H�|$�t$ H�A����������D�t$D�t$�   D�'E��uZ�|���D  D��)��l���Hc��D�[D�| ��E��D�A9��B���D���K�҃�9��2�����9��'����{u�D�����
�E��t�D�O�D��)�A��D	ʈ��H�$H�k��sA�������A�ލP�A��H������A�ދD�s����H��H��1��L$(�r��Ic�D�|$(H�D$ H�|$ K�<<H�H�|$(L;,$�b���H�\$0H��L��H��L���Zq��J�<#L��1�Ll$ �Wr��H\$(L;,$r�H�\$0�$���I������f.�     AWAVAUATUSH��   �D$d    H���>  M���5  H��H���)  M���   A�pH��@���  1��{ �  �{1�����   D�E����   H���A��H���H�@      �I��D��H�H9���   H����������I��H)�I)�I9���   A�@����   E�E����   I�QA��I�       �M�H���L9�|mI��������I��M�)M)�A��A��I���M)�M9�GM9�M��MN�M�L�L9�IL�M��L�\$ L)�M9�MN�H9�HM�L�T$(L)��dD  @��t"f��   H�Ę   []A\A]A^A_�f�     I�x t�1��{ t֋CA3@�������f�I��������L�t$(L�|$ M��H��H��H��H�T$���a  ���Y  H�U H�$���Y  A���t
L+l$ L+d$(@���H  9�u
;T$��  ��    H�L$H�t$Hc�L�L$0H��������H�щT$H�T$@H�H��Hc�H9������L$A�@L�D$HH�<$�D$PHc�H�L$dH�����H�D$8�D$d�������L�D$HL�L$0A�HM�P��H�L$��   �|$P�D$I��I��A�A��L)�A��H)�D1߉�H��H�T$@D)�H����N��L\$8Lc�M�M9�vYH�L$0Lc�L�L$PL�|$I��H�\$@L�� H��L��L��L���m��I��M�I9�w�L�D$HL�|$H�L$0H�\$@L�L$PM�PH�<$L��L�L$@L�D$0H�L$�l_��L�D$0H�L$�D$L�L$@A�PA�HA� ��y�\$�D$�D$H A�@H�D$8I�@�{�D$@ tp�   H�T$hH��H��L�$L�L$H�D$h    H�D$p    H�D$x    HǄ$�       HǄ$�       �t���L�$���D$d��  �D$@L�L$H�\$hA�@����  A�L+t$(�3I��L+|$ L)�I��H�{H���KH)�Hc�H��H�<$L�IPH�T$Hc�H�H�T$0H9��]  ��$�   H�l$PA�������$�   D��$�   H�\$L�D$8��D��$�   L�L$X��A��A��D��@ H�L$H�4$�iI��H�L$H�H9���   �     I��A�B�D�D���   �y�qH��A��D�I�I��H��')���D����I��M��I��H��'��I��'A��A�H��'D�A�E��I��D��I��H��'M��H��'I��'D�@�y�D�����I��H��'�@�q��A�L9��T���H�D$8�@H�L$HcQH$Hc�H�$HT$H9L$0� ���H�l$PL�D$8L�L$XH�D$ I��D$��HD$(I�A�D$d��t�|$H tL��H���'����    �|$@ tH�t$xH�} �\���D$d�7���f�1��.���f�     @��������   A�H��H��������fA�pH�Hc�H�|$H��L�L$A�8A�@A�HL�D$Hc�H9��������H�<$H�T$dHc����L�D$I�@�D$d��������D$HL�L$������|$H �����L��H���O����?����D$H ����H�A�" H���t3UH��S�`i H��D  ��H��H�H���u�H��[]�f.�     ��
l���                         r /initrd/close.bmp /initrd/shell.lef /dev/mouse0       Error initializing freetype r /initrd/montserrat.ttf    Error loading font /initrd/montserrat.ttf       Error loading font from memory /initrd/montserrat.ttf Error Setting Font Size Error loading custom font Error loading custom font from memory Freetype Error!        �o@      �?FREETYPE_PROPERTIES                             `�F     `�F     `�F      �F      �F     ��F     @�F     ��F     ��F     @G      )G     `eG     �eG     �gG     `gG     �fG     @�G      �G             properties font-format kerning glyph-dict postscript-font-name sfnt-table tt-cmaps type42 truetype truetype-engine darkening-parameters hinting-engine adobe no-stem-darkening random-seed .resource/ resource.frk/ .AppleDouble/ % ._ cff type1                        pt@     Pt@     �t@     �r@     �s@     (�@     k�@     k�@     k�@     �@     �@     k�@     k�@     �@     �@     Ȯ@     Ȯ@     ��@     ��@     ��@     ��@     ��@     ��@     ��@     ��@     ��@     ��@             ��     G	           ��     8�     *�      �r      L9      �      S      )      �      �      �       s       9                                                                 ��@             `�@             �@            ��@             �@            ж@            ��@            `�@            ��@            interpreter-version Weight OpticalSize Slant sfnt .notdef TrueType multi-masters metrics-variations tt-glyf     ��A     ��A     ��A     кA     �A     �A      �A     ��A     ĿA     ĿA     ĿA     ĿA     ĿA     ĿA     ��A     ��A     ��A     ��A     J�A     �A     ��A     ϾA     ��A     ��A     ��A     ��A     ��A     ��A     S�A     b�A     ��A     �A     ��A     ��A     ��A     �A     u�A     �A     R�A     !�A     ��A     ��A     ��A     {�A     b�A     e�A     ��A     ��A     �A     �A      �A     G�A     c�A     ��A     d�A     d�A     S�A     S�A     "�A     "�A     6�A     6�A     �A     �A     ��A     ��A     �A     �A     G�A     ,�A     U�A     U�A     ��A     %�A     �A     ��A     O�A     '�A     ��A     ��A     U�A     ��A     ��A     ��A     ��A     �A     e�A     S�A     0�A     �A     ��A     ��A     ��A     ��A     ��A     o�A     y�A     ��A     ��A     /�A     w�A     �A     f�A     T�A     �A     �A     4�A     ��A     ��A     r�A     ��A     ��A     ��A     ��A     ��A     ��A     @�A     @�A     @�A     @�A     \�A     �A     �A     ��A     ��A     ��A     ��A     ��A     ��A     j�A     ��A     �A     �A     ��A     ��A     ��A     �A     ��A     ��A     �A     �A     ��A     ��A     ��A     ��A     w�A     ��A     S�A     ��A     w�A     0�A     �A     �A     ��A     O�A                  
                                               "             
                                    X�    �      �;#(    ć      �D�    �      X�    �      �;#(    ć      �D�    �      ���    P      d    ��      c���    X      ���    P      �VY�    ��      �r�    E       F�W    P      `љ�    _q      h�"�    �      N�b    P      d]j�    @y      )�Px    �      
�-    P      �2=    ��      ;�?�    �      &�_    P      �ɬ�    �~      ����          ���    P      ;�0Z    c�      &�    ~       ���    P      ��    ��      &�    ~       ���    `      ����    n�      ���S    �       �C    P      0�
�    �t      	4��    {      F��          �|�@    *�      �t�`    z       8��          ����    og      ��    �      ����           �H��    ��      p           ����           �Z
    9|     p                           U%�@    �       �X��    |                      R�3    �       *��&    j                      e�m    �      Knl    �$                      U%�@    �       ��Q�    |                      dv�    �       1(Ʀ    �                      ��-    �      3F`�    �                      Lw�@    �      ��\�    �                      ��=    A      fw�    �"                      �&iJ    �      FC4    �                      �4�    f      F�l    �"                      S�]    �      _Zt@    �"                      H�U�    �      �� 9                `       n0��    �X      *HC�    5                       cpop                DFGirl-W6-WIN-BF    DFGothic-EB         DFGyoSho-Lt         DFHei-Md-HK-BF      DFHSGothic-W5       DFHSMincho-W3       DFHSMincho-W7       DFKaiSho-SB         DFKaiShu            DFKaiShu-Md-HK-BF   DFKai-SB            DFMing-Bd-HK-BF     DLC                 DLCHayMedium        DLCHayBold          DLCKaiMedium        DLCLiShu            DLCRoundBold        HuaTianKaiTi?       HuaTianSongTi?      Ming(for ISO10646)  MingLiU             MingMedium          PMingLiU            MingLi43                                    ��		             P    "                    !!  !!!!!! !!!!!!              3!!                                                                        @   @   @               @             D                       	                         �       ��F                            A     A      �A     �             0      ��A     �9A     �A     �A     �9A             ��A     P�@             �NA     ��A     PA     C�F     ��F     ��F     �F     ��F     ��F     ��F     ��F     ԥF     ��F     8�F     @�F                      A            �A                      �A                             �A                     0�A      �A     `�A     ��A     �A     �A                     �OA     � A     ��A     �MA     pshinter StandardEncoding ExpertEncoding ISOLatin1Encoding eexec closefile FontDirectory CharStrings dup put %!PS-AdobeFont %!FontType postscript-cmaps psaux Regular Black Notice FullName FamilyName ItalicAngle isFixedPitch UnderlinePosition UnderlineThickness UniqueID lenIV LanguageGroup password BlueScale BlueShift BlueFuzz BlueValues FamilyBlues FamilyOtherBlues StdHW StdVW MinFeature StemSnapH StemSnapV ExpansionFactor ForceBold PaintType StrokeWidth FontBBox NDV CDV DesignVector FontMatrix Subrs Private BlendDesignPositions BlendDesignMap BlendAxisTypes WeightVector postscript-info                               1%B     1%B     k%B     J%B     �%B     �%B     �%B     �%B     �$B     @:B     �:B     �9B     �9B     �9B     �9B     `9B     89B     �8B     �8B     `8B     88B     �7B     �7B     P7B     H=B     =B     �<B     �<B      ;B     �:B     h=B     �:B     �;B     �;B     �;B     `;B     8<B     <B     x<B     (7B     �6B     �6B      7B     p6B     @6B      6B      6B     �5B     �5B     h5B     @5B     5B     �4B     �4B     h:B             |�F                                         ��F                                        �F                                        �F                                        ��F                                         �F                   (                     #�F                   0                     0�F                   2                     B�F                   4                     ��F                                         U�F                                         ^�F                                        d�F                   �                     r�F                   �                     {�F                   p                     ��F                   x                     ��F                   |                     ��F        	                              ��F        	           (      
   	          ��F        	           <         
          ��F        	           X      
             ��F        	           �                    ƸF        	           �                    ̸F        	           �                    ׸F        	           �         �          �F        	           �         �          �F                   �                     ��F                   �                     ��F                                        �F                   �                    ηF                   �                    �F                                       �F                                         $�F                   X                    (�F                   \                    ,�F        	           �        �         9�F           @2B                            ��F           PB                            D�F           @.B                            ��F           �'B                            J�F           �B                            R�F            B                            g�F           �B                            v�F           p&B                            ��F            B                            ��F           `B                                                                                                  h       #�F                           @B     �B     �3B     x      X       P      �[B     0B     �GB     �GB     �B     0B     @B     P>B     �HB     �B     PGB             b�F     `�F     W�F     p�F     C�F     /�F     ��F     ��F     8�F     ��F     O�F     ��F     ��F      �F                     ��@     `�@     �3B             ��A      B       B     0 B     p4B                             P B     �DB     �FB      @B     �AB     PFB     �@B      GB     � B     �B             0B     ��A              >B     � B     /FSType cff-load CFF CID        ��B     ��B     p�B      �B     ��B     ��B       ( ) *                                                                                                  � �   � � � � � � � �    c � � � � � � � � � �   � � � �   � � �                	  
m n    !"#$%&'()*+,-./                                                                    012    34567  8    8    :;    <=>      � � � ?@ABCDE    F� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                                                                        	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _                                                                     ` a b c d e f g h i j k l m n   o p q r   s t u v w x y z   {   | } ~  � � � �   � �   � � � �                                 �   �         � � � �           �       �     � � � �            � � � � � �    c � � � � � � � � � �   � � � � � �  	
m n ,-.1:;� � � @ABCDEF� � � GHIJKLMNOPQRSTUVWXYZ                     � � � � � � � � � �    c � � � � � � � � � �   � � � � � � �  	
m n  !"#$%&'()*+,-./0123456789:;<=>� � � ?@ABCDEF� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                              	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _ ` a b c d e f g h i j k l m n o p q r s t u v w x y z { | } ~  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                                                                                        (                           0                           8                           <                                   ��B                  �                                   ��B                  �                           �                           �                           �                                   0�B                  �                           �                                   ��B                          `�B                  �                                                     !                          "                          #                          $                           %  (                        &  0                                                      x              
            �                       	   8             
         	!  �                        
!  �                        !  �                        
   �                           �                        !  �                �     !                   �     !  �                        !  �                        !  �                        !  �                        !  �                        !  �                           �                           �                           �                        1          ��B                0  �                         $1                           %1  (                        0  8                        0          0�B                @          0�B                A          ��B                P                          P  x              
         P  �                       	P  8             
         	Q  �                        
Q  �                        Q  �                        
P  �                        P  �                        Q  �                �     Q                   �     Q  �                        Q  �                        P          ��B                P          ��B                P  �                                                     ���������������G�z�G�S㥛�  e�c]�F ��#��S  �Z�{c  �Ք��   0�y   }�%                          
       d       �      '      ��     @B     ���      ��     ʚ;                          h       �F                           �dB     peB     �B     �      `       H      0�B     ��B     �}B     �{B     pfB     �dB      �B     �aB             `�B     0|B     �zB     C�F     ��F     ��F     `�F     ��F      �F     ��F      �F     b�F     ��F     W�F     0�F     ��F     ��F     ��F     ��F     8�F     ��F     ��F     ��F                                     �cB     0�B     �cB     �oB     �oB                             �bB                                                     �bB                     `bB     pbB     �bB     �bB     �bB     �bB     �bB     �bB     �dB     �dB     ��@     `�@     @wB     �aB     bB     �hB     PiB             �wB     0yB     �aB                             p�B     �mB     (       �`B     �eB     PaB     paB                                                                     ``B     �`B     �`B     �`B                                             CIDFontName StartData /sfnts (Hex) %ADOBeginFontDict t1cid CID Type 1 CIDFontVersion CIDFontType Registry Ordering Supplement UIDBase XUID CIDMapOffset FDBytes GDBytes CIDCount SubrMapOffset SDBytes SubrCount lenBuildCharArray ForceBoldThreshold FDArray   %!PS-Adobe-3.0 Resource-CIDFont                       h       %�F                           ��B     `�B     ��B     x      `       H       �B     `�B     ��B     ��B     @�B     ��B     ��B                             @�B             C�F     +�F     b�F     ��F     ��F     ��F     ��F     P�F     8�F     @�F                     ��@     `�@     ��B      �B     0�B                             ��B     ��B                             p�B                     ��F                                           6�F                                          E�F                                          Q�F                                          Z�F                                           c�F                    (                      n�F                    �                      v�F         	           �         �           {�F                                         ��F                                          ��F                    $                     ��F                    (                     |�F                                          ��F                                         �F                                         �F                                         ��F                                          �F                   (                      #�F                   0                      0�F                   2                      B�F                   4                      ��F                                          �F                                         ηF                                        ��F                   @                     ��F                   H                     ��F                   8                     ��F                   �                      ��F                   �                      �F                   �                      U�F                                          ^�F                                         d�F                   �                      r�F                   �                      {�F                   p                      ��F                   x                      ��F                   |                      ��F        	                               ��F        	           (      
   	           ��F        	           <         
           ��F        	           X      
              ��F        	           �                     ƸF        	           �                     ̸F        	           �                     ׸F        	           �         �           �F        	           �         �           ��F                   �                      �F                                          ��F           ��B                             9�F           P�B                             �F           p�B                             ��F           ��B                                                                                             sC     (
C     �C     �C     (
C     (
C     �C     �C     $C     C     C     C     CC     CC                            ��B            P�B            �B            ��B                                      :            $ ( , 0 4 8 < @ D H L P T X \ ` d h                       8       ��F                                           � C     �      X       h      �C     �C                      �B     ��B     �C      C                                     ��F     �F     C�F     ��F                     � C     ��B     ��B                             (       �B     p�B     ��B     ��B                                             pfr pfr-metrics PFR %!PS-TrueTypeFont known Type 42                             |�F                                          ��F                                         �F                                         �F                                         ��F                                          �F                   (                      #�F                   0                      0�F                   2                      B�F                   4                      ��F                                          ��F                                         �F                   �                     ηF                   �                     �F                                        �F                                          9�F            5C                             ��F           �;C                             ��F           �6C                             �F            0C                                                                                   @       ��F                           0/C     �+C     P6C     �      `       8      pCC     P-C     -C     0CC     �,C     �,C     p@C                              ,C     �+C     W�F     ��F     b�F     ��F     ��F     ��F     C�F     ��F                                      +C     P+C     `+C     p+C             �*C     `6C     `/C     Bold Italic winfonts Windows FNT                                      8       �F                                           PTC            X       0      �UC     @aC                                     `QC                             `TC     QC     C�F     �F     �F     0�F                     �PC                     �PC             �PC     �PC                                                              �    < L N P R T V X Z [ \ ^ ` b d f h j l m n o p x � � � � � � � � � �                                                                       (               �    
       n    h                   (   "                 @   :       Oblique SLANT WEIGHT_NAME SETWIDTH_NAME ADD_STYLE_NAME FAMILY_NAME RESOLUTION_X RESOLUTION_Y CHARSET_REGISTRY CHARSET_ENCODING 10646 8859 646.1991 IRV pcf bdf PCF                                                                         
                
                	                      	                                             
             
                                                       @       ��F                            cC     0cC     phC     8      X       0      ��C      jC                                     �dC                             �cC     @cC     ��F     ��F     C�F     ��F     8�F     ��F                      cC     cC     �bC     �jC             �aC     �aC     �aC      bC                                             COMMENT DEFAULT_CHAR FONT_ASCENT FONT_DESCENT SPACING ENDPROPERTIES %hd _XFREE86_GLYPH_RANGES  + STARTFONT STARTPROPERTIES FONTBOUNDINGBOX - CHARS ENDFONT ENDCHAR STARTCHAR SWIDTH DWIDTH BBX BITMAP BDF CHARSET_COLLECTIONS COPYRIGHT DESTINATION DEVICE_FONT_NAME FACE_NAME FONTNAME_REGISTRY FOUNDRY FULL_NAME ITALIC_ANGLE NOTICE RAW_ASCENT RAW_AVERAGE_WIDTH RAW_AVG_CAPITAL_WIDTH RAW_AVG_LOWERCASE_WIDTH RAW_CAP_HEIGHT RAW_DESCENT RAW_END_SPACE RAW_FIGURE_WIDTH RAW_MAX_SPACE RAW_MIN_SPACE RAW_NORM_SPACE RAW_PIXEL_SIZE RAW_POINT_SIZE RAW_PIXELSIZE RAW_POINTSIZE RAW_QUAD_WIDTH RAW_SMALL_CAP_SIZE RAW_STRIKEOUT_ASCENT RAW_STRIKEOUT_DESCENT RAW_SUBSCRIPT_SIZE RAW_SUBSCRIPT_X RAW_SUBSCRIPT_Y RAW_SUPERSCRIPT_SIZE RAW_SUPERSCRIPT_X RAW_SUPERSCRIPT_Y RAW_UNDERLINE_POSITION RAW_UNDERLINE_THICKNESS RAW_X_HEIGHT RELATIVE_SETWIDTH RELATIVE_WEIGHT RESOLUTION _MULE_BASELINE_OFFSET _MULE_RELATIVE_COMPOSE                       8       ��F                                           ��C            X       0       �C     ��C                                     ��C                             ��C     ��C     ��F     p�F     C�F     ��F                     p�C     0�C     (       ��C      �C      �C     ��C                                             ��������              �~   ~                         �                                                                         	       
                          
                                                         \�F                   F�F                   X�F                   n�F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   k�F                   ��F                   ��F                   ��F                   �F                   �F                   �F                   �F                   #�F                   ��F                   ��F                   ��F                   0�F                   ��F                   ��F                   %�F                   7�F                   B�F                   T�F                   j�F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   �F                   �F                   !�F                   0�F                   C�F                   X�F                   n�F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   	�F                   �F                   (�F                   8�F                   w�F                   ��F                   N�F                   <�F                   4�F                   �F                   G�F                   \�F                   r�F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   ��F                   1�F                   B�F                   �F                   C�F                   Y�F                                           �C      �C     0�C     H�C     P�C     ��C      �C     D     �D     D     �D     @D     ND     D     D     D     D     D     D     D     D     D     D     D     D     D     ND     �D     &D     �D     �D     �D     �D     &D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     zD     zD     zD     �D     �D     �D     mD     �D     �D     �D     ^D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     �D     D     �~D     '�D     .�D      �D     �~D     T�D     <�D     5�D     �~D     [�D     i�D     b�D     [~D     @~D     C�D     p�D              ,         ( * 0 8 @ H P                                    ����cinu    ����cinu       nmra       bmys   
   cinu      cinu      sijs        bg      5gib      snaw      ahoj                             $    
             " $ &                           
             "                    � �      
 x z | ~ �           h p                      N       
             ! " # $ % & ' ( ) 0 8 @ H P Q R S T V X Z \ ^ ` b                                ( 0 8                                                          6           , 4 	: 	; < =                                  6        " ( 0 8 @ H J L N P R T V X                                       
               �G     @G     �G     @G     �G     @G     �G     @G     �G                             (       0�C     �D     p�C     ��C                                             ����                                            H       ��C     PD     ��C     ��C      �C     ��C     � D     ��C     ��C            LD      �C                             P       ��C             p�C     0QD                                                    �JD     ��C                             P       �C             p�C     �PD                                                    `ID     ��C                             (       ��C              �C     @�C                                             
       �HD     ��C                             (       ��C             p�C     ��C                                                    �ED     ��C                             (       ��C              �C     p�C                                                     ED     @�C                             P       ��C             ��C     �PD                                                    �>D     ��C                             (       ��C             ��C     0�C                                                    p<D     ��C                             (       ��C             ��C     ��C                                                     �pD      �C                                            ��F                   �G                     `�C                             ��C     `_D      0D      D     `�C     �D     P^D     p,D     pQD     �+D     `^D     0+D     �'D     D     p�C     �D     �'D     @^D     pqD     �XD      D     ��C      ZD     ��C     �#D     ��C     p#D     @ D     �D     �D     �D     `D      �C     ��C     D     p�C     �D     ��C                     w�F     �G     b�F     XG     W�F     �G     ��F     @G     ��F     PG                     p�C     P�C     ��C     �wD     0123456789ABCDEF    �|���������W�YD     �XD     �D     ��C     0PD     glyph-to-script-map fallback-script default-script increase-x-height warping autofitter 田 囗 ꘓ ꖜ ꖴ า ๅ ๐ ⵔ ౦ ౧ ꪒ ꪫ ௦ ᮰ ට 𐑴 ꢝ ꣐ 𐒆 𐒠 𐓂 𐓪 𐰗 ᱛ ߋ ߀ ဝ င ဂ ᡂ ᠪ ഠ റ ꓳ ᵒ ᴼ ⁰ ₒ ₀ o O 0 ໐ ೦ ಬ ᧡ ᧪ ០ ꤍ ꤀ ם ਠ ਰ ੦ ટ ૦ ο Ο 𐌴 𐌾 𐍃 Ⱅ ⱅ Ⴖ Ⴑ ⴙ ი ე ა Ჿ ዐ 𐐄 𐐬 ठ व ट о О 𐠅 𐠣 Ⲟ ⲟ Ꭴ Ꮕ ꮕ 𐊫 𐋉 ᑌ ᓚ 𑄤 𑄉 𑄛 ᝋ ᝏ ০ ৪ ꛁ ꛯ 𐬚 ս Ս ل ح ـ 𞤌 𞤮                  #                      
                                                         ��������������������������������������������������������������������������������                                                          
                      *0  /0  �1  �1                     �  �.  �.   /  �/  �/  �/   0  ?0  @0  �0  �0  �0   1  /1  01  �1  �1  �1  �1  �1  �1  �1  �1  �1   3  �3   4  �M  �M  �M   N  ��  `�  �   �  ��  ��  ��   �  ��  �  �  0�  O�   �  ��   � ��  � /�  � _�    ߦ  � ?� @� �  � �� �� ��  � �                             5  5  7  7  9  9  >  ?  q  ~  �  �  �  �  �  �             �          �  �  �  �  �  �  %�  &�                   �  /�              <  <  ?  ?  A  D  M  V  b  c                                                  "  '  4  7  ;             O                           �  ?�                          0-  -                          1  1  4  :  G  N                                                 >  @  F  V  b  c                       ��  ��  ��  ��  ��  ��  ��  ��  ��  ��          ��  ߪ          �  �  �  �  �  �          �  �          �  �  �  �                  �  �  �  �                  �  �  �  �                  �  �                          P          ��  ��  ��  Ũ                  ��  ߨ                          � �                         � �                           O                         P                            �  �  �  �                  �  �                          -  0  2  7  :  :  =  >  X  Y  ^  `  q  t  �  �  �  �  �  �  �  �  |�  |�                                     �  �  ��  `�  �          �  �  �  �                     �  `                       ;  <  M  N  b  c                                               Ф  ��                                          �   �   �   �   �   �   �  �  �  �  ,  a  x  x  �  �  p      },  },  p�  p�  ��  ��  \�  _�                          b  j  �   �   |,  |,          ^   `   ~   ~   �   �   �   �   �   �   �   �   �   �   �  �  �  �     o  �  �  �  �        >   >   ��  ��  ��  ��                                         �   �   �   �   �   �   �   �        �  O  P  �  �  �  �  �     o  �  �     +  k  w  y    �  �  �  �     �      o   �   �   �   �   P!  �!  `,  {,  ~,  ,   .  .   �  o�  q�  ��  ��  ��  0�  [�  `�  o�   �  �   � ��                                 �  �  �  �  �  �          �  �                          �  �                          �  �  �  �  �  �  �  �                  �  �          �  �  �  �  �  �  �  �  �  �  �  �                  �  �          &�  -�           �  /�                          �  �  �  �  �  �  �  �  �  �          �  �  �  O�                                  
  
  <
  <
  A
  Q
  p
  q
  u
  u
           
  
          �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
  �
                  �
  �
                          z  z  �  �  �  �  �  �  �  �  �  �  �  �          p  �     �                  0 O          � /�          ,  _,   � /�                 �  �   -  --                  �  �  �  �                  ]  _                               �  �  �-  �-   �  /�                    O          	  	  :	  :	  A	  H	  M	  M	  S	  W	  b	  c	  �  �  ��  ��                                   	  ;	  =	  P	  S	  c	  f	  	  �   �   �  ��                  �  �  �-  �-  o�  �  ��  ��                                     �     /  �-  �-  @�  ��  �  �                            ?         �,  �,          �,  �,                          �  �  p�  ��                  � �                              �  �                     ' 4 F F           O         R  S          @  _                          �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	  �	                  �	  �	          �  �          ��  ��          9 ?           ?         Y  _          0  �  �  �                           K  _  p  p  �  �  �  �  �  �  �  �  �  �  �  �  ��  ��  p�  p�  r�  r�  t�  t�  v�  v�  x�  x�  z�  z�  |�  |�  ~�  ~�             �  P  �  �  �  P�  ��  p�  ��   � ��                 D� J�          � _�                H       �G                   `)G     ��D     @�D     ��D                                                     0�D     8�F     �)G                     ��D     �D                            ��      PE     ��D             P�D      �D     ��D            �r      �E      �D             @�D     0�D     ��D     �9G     p9G     P9G     09G     9G     �8G     �8G     �8G     �8G     p8G     P8G     08G     8G     �7G     �7G     �7G     �7G     p7G     P7G     07G     7G     �6G     �6G     �6G     �6G     p6G     P6G     06G     6G     �5G     �5G     �5G     �5G     p5G     P5G     05G     5G     �4G     �4G     �4G     �4G     p4G     P4G     04G     4G     �3G     �3G     �3G     �3G     p3G     P3G     03G     3G     �2G     �2G     �2G     �2G     p2G     P2G     02G     2G     �1G     �1G     �1G     �1G     p1G     P1G     01G     1G     �0G     �0G     �0G     �0G     p0G     P0G     00G     0G     �/G     �/G     �/G     �/G     p/G     P/G     0/G     /G                              HG     �GG     �GG     @GG      GG     �FG     �FG     @FG      FG     �EG     �EG     @EG      EG     �DG     �DG     @DG      DG     �CG     �CG     @CG      CG     �BG     �BG     @BG      BG     �AG     �AG     @AG      AG     �@G     �@G     @@G      @G     �?G     �?G     @?G      ?G     �>G     �>G     @>G      >G     �=G     �=G     @=G      =G     �<G     �<G     @<G      <G     �;G     �;G     @;G      ;G     �:G     �:G     @:G      :G     �9G                     @HG     �)G     �HG      *G                     T      9   �   
               S      8       
               R      7       
               Q      6       
               P      5       
               O      4   �   
               N      3   �   
               M      2   �   
               L      1   �   
               K      0   �   
               J      /   �   
               I      .   �   
               H      -   �   
               G      ,   �   
               F      +   �   
               E      *   �   
               D      )   �   
               C      (   �   
               B      '   �   
               A       &   �   
               @      %   �   
               ?      $   �   
               >      #   �   
               =      "   �   
               <      !   �   
               ;          �   
               :         �   
               9         �   
               8         �   	               7         �                  6         �                  5         �                  4         �                  3         �                  2         �                  1         �                  0         �                   /         �   
               .         �   
               -         �   
               ,         �   
               +         �   
               *         |   
               )         v   
               (         p   
               '         i   
               &         i   	               %         i                  $         i                  #         i                  "         i                  !         i                            i                           i                           i                            f   
                        a   
                        Z   
                        S   
                        P   
                        K   
                        E   
                        ?   
                        ?   	                        ?                           ?                           ?                           ?                           ?                           ?                           ?                           ?                            :   
                        5   
               
      
   .   
               	      	   +   
                        $   
                            
                           
                           
                           
                           
                        	   
                           
                              
                               9       �G     �G              G                             8       PG      G             ��F                             7       �G     `G             ��F                             6       �G     �G             ��F                             5        G      G             ��F                             4       @G     0G             G                             3       �G     �G             G                             2       `G     PG              G                             1       �G     �G             $G                             0       0G      G             ,G                             /       `G     @G             4G                             .       �G     pG             8G                             -       �G     �G             <G                             ,       �G     �G             @G                             +        G      G             EG                             *       @G     0G             MG                             )       `G     PG             WG                             (       �G     pG             aG                             '       �G     �G             fG                             &       �G     �G             �F                             %       �G     �G             jG                             $       �G      G             pG                             #       �G     �G            |G                             "       G     �G             �G                             !       0G      G             �G                                     `G     @G             �G                                    �G     �G             �G                                    � G       G             �G                                    �!G     �!G             �G                                    �"G     `"G             �G                                     "G     �!G             �G                                    P"G      "G             �G                                    �"G     �"G             �G                                    #G     �"G             �G                                    p#G     @#G            �G                                    �#G     �#G             �G                                     $G     �#G             �G                                    @$G     8$G            �G                                    `$G     P$G             �G                                    �$G     x$G             �G                                    �$G     �$G             
G                                    �$G     �$G             G                                    %G     %G             G                                    �%G      %G            (G                                     &G     �%G             4G                                    @&G     0&G             :G                                    `&G     P&G             DG                             
       �&G     p&G             LG                             	       �&G     �&G             XG                                    �&G     �&G             bG                                     'G     �&G             jG                                     'G     'G             yG                                    �'G     @'G            �G                                    �'G     �'G             �G                                    �'G     �'G             �G                                    �'G     �'G             �G                                    �(G      (G             �G                                     �(G     �(G             �G                                     H                                       ��D     ��D            �r      �E     ��D              �D     ��D     ��D                   (   	   A       �      i      {       �      �      �      �       �      �   	   �             �           .      �      8     X      �      �     �     x     x      �      �     �     �  	   �      �           4      M      �           4      T  	   t      �     �      �      �     �      �      �     �      �     �  	   �      �      �      �           >  	   ^      �      ~     �      �     �      �      �     �        	                �      �     �     �     �      �      �      )     B      [  	   t      �      �           �      5  	   U      u     �      u     �      �      �     �      �  	         5     U      �      �     �      �  	         �      5     ]      �      q     �      �     �  	   �      �      �      �  	   �      	     L	      m	     �      �	     �	     �	     �	      
     �      
     -
      ?
      �      �
  	   �
      �
     �
      �
      �      �
  	        /      O      q      �      �  	   �      �      N
     z
      �      �  	   �           (     4      �      L     \      l     z  	   �      �      �      �     �      �     �  	   �            �           7      T     n  	   n      �      �      �     �      �      �     �      �           J      �      N  	   n      �     �      �      �     �      �  	   �      �      �                 �           -      �      A     i      �      �  	   �      �     �      �           6      �      ^     ~      �      �     �      �      �  	   �      �      �           1      �      ]     u      �      �      �     �      �      �     �      �      �           �      �     �      �      5  	   M      i     u     �      �      �      �      �     �      �           �      �                              𞤌 𞤅 𞤈 𞤏 𞤔 𞤚 𞤂 𞤖 𞤬 𞤮 𞤻 𞤼 𞤾 𞤤 𞤨 𞤩 𞤭 𞤴 𞤸 𞤺 𞥀 ا إ ل ك ط ظ ت ث ط ظ ك ـ Ա Մ Ւ Ս Բ Գ Դ Օ Ւ Ո Դ Ճ Շ Ս Տ Օ ե է ի մ վ ֆ ճ ա յ ւ ս գ շ ր օ հ ո ճ ա ե ծ ս օ բ ը ի լ ղ պ փ ց 𐬀 𐬁 𐬐 𐬛 𐬀 𐬁 ꚧ ꚨ ꛛ ꛉ ꛁ ꛈ ꛫ ꛯ ꚭ ꚳ ꚶ ꛬ ꚢ ꚽ ꛯ ꛲ অ ড ত ন ব ভ ল ক ই ট ঠ ি ী ৈ ৗ ও এ ড ত ন ব ল ক ᝐ ᝈ ᝅ ᝊ ᝎ ᝂ ᝃ ᝉ ᝌ ᝀ ᝃ ᝆ ᝉ ᝋ ᝏ ᝑ ᗜ ᖴ ᐁ ᒣ ᑫ ᑎ ᔑ ᗰ ᗶ ᖵ ᒧ ᐃ ᑌ ᒍ ᔑ ᗢ ᓓ ᓕ ᓀ ᓂ ᓄ ᕄ ᕆ ᘣ ᕃ ᓂ ᓀ ᕂ ᓗ ᓚ ᕆ ᘣ ᐪ ᙆ ᣘ ᐢ ᒾ ᣗ ᔆ ᙆ ᗮ ᒻ ᐞ ᔆ ᒡ ᒢ ᓑ 𐊧 𐊫 𐊬 𐊭 𐊱 𐊺 𐊼 𐊿 𐊣 𐊧 𐊷 𐋀 𐊫 𐊸 𐋉 𑄃 𑄅 𑄉 𑄙 𑄗 𑄅 𑄛 𑄝 𑄗 𑄓 𑄖𑄳𑄢 𑄘𑄳𑄢 𑄙𑄳𑄢 𑄤𑄳𑄢 𑄥𑄳𑄢 Ꮖ Ꮋ Ꭼ Ꮓ Ꭴ Ꮳ Ꭶ Ꮥ ꮒ ꮤ ꮶ ꭴ ꭾ ꮗ ꮝ ꮿ ꮖ ꭼ ꮓ ꮠ ꮳ ꭶ ꮥ ꮻ ᏸ ꮐ ꭹ ꭻ Ⲍ Ⲏ Ⲡ Ⳟ Ⲟ Ⲑ Ⲥ Ⳋ Ⳑ Ⳙ Ⳟ Ⲏ Ⲟ Ⲑ Ⳝ Ⲱ ⲍ ⲏ ⲡ ⳟ ⲟ ⲑ ⲥ ⳋ ⳑ ⳙ ⳟ ⲏ ⲟ ⲑ ⳝ Ⳓ 𐠍 𐠙 𐠳 𐠱 𐠅 𐠓 𐠣 𐠦 𐠃 𐠊 𐠛 𐠣 𐠳 𐠵 𐠐 𐠈 𐠏 𐠖 Б В Е П З О С Э Б В Е Ш З О С Э х п н ш е з о с р у ф 𐐂 𐐄 𐐋 𐐗 𐐑 𐐀 𐐂 𐐄 𐐗 𐐛 𐐪 𐐬 𐐳 𐐿 𐐹 𐐨 𐐪 𐐬 𐐿 𐑃 क म अ आ थ ध भ श ई ऐ ओ औ ि ी ो ौ क म अ आ थ ध भ श ु ृ ሀ ሃ ዘ ፐ ማ በ ዋ ዐ ለ ሐ በ ዘ ሀ ሪ ዐ ጨ გ დ ე ვ თ ი ო ღ ა ზ მ ს შ ძ ხ პ ს ხ ქ ზ მ შ ჩ წ ე ვ ჟ ტ უ ფ ქ ყ Ⴑ Ⴇ Ⴙ Ⴜ Ⴄ Ⴅ Ⴓ Ⴚ Ⴄ Ⴅ Ⴇ Ⴈ Ⴆ Ⴑ Ⴊ Ⴋ ⴁ ⴗ ⴂ ⴄ ⴅ ⴇ ⴔ ⴖ ⴈ ⴌ ⴖ ⴎ ⴃ ⴆ ⴋ ⴢ ⴐ ⴑ ⴓ ⴕ ⴙ ⴛ ⴡ ⴣ ⴄ ⴅ ⴔ ⴕ ⴁ ⴂ ⴘ ⴝ Ნ Ჟ Ჳ Ჸ Გ Ე Ო Ჴ Ი Ჲ Ო Ჩ Მ Შ Ჯ Ჽ Ⰵ Ⱄ Ⱚ Ⰴ Ⰲ Ⰺ Ⱛ Ⰻ Ⰵ Ⰴ Ⰲ Ⱚ Ⱎ Ⱑ Ⰺ Ⱄ ⰵ ⱄ ⱚ ⰴ ⰲ ⰺ ⱛ ⰻ ⰵ ⰴ ⰲ ⱚ ⱎ ⱑ ⰺ ⱄ 𐌲 𐌶 𐍀 𐍄 𐌴 𐍃 𐍈 𐌾 𐌶 𐌴 𐍃 𐍈 Γ Β Ε Ζ Θ Ο Ω Β Δ Ζ Ξ Θ Ο β θ δ ζ λ ξ α ε ι ο π σ τ ω β γ η μ ρ φ χ ψ ત ન ઋ ઌ છ ટ ર ૦ ખ ગ ઘ ઞ ઇ ઈ ઠ જ ઈ ઊ િ ી લી શ્ચિ જિ સી ુ ૃ ૄ ખુ છૃ છૄ ૦ ૧ ૨ ૩ ૭ ਕ ਗ ਙ ਚ ਜ ਤ ਧ ਸ ਕ ਗ ਙ ਚ ਜ ਤ ਧ ਸ ਇ ਈ ਉ ਏ ਓ ੳ ਿ ੀ ਅ ਏ ਓ ਗ ਜ ਠ ਰ ਸ ੦ ੧ ੨ ੩ ੭ ב ד ה ח ך כ ם ס ב ט כ ם ס צ ק ך ן ף ץ ಇ ಊ ಐ ಣ ಸಾ ನಾ ದಾ ರಾ ಅ ಉ ಎ ಲ ೦ ೨ ೬ ೭ ꤅ ꤏ ꤁ ꤋ ꤀ ꤍ ꤈ ꤘ ꤀ ꤍ ꤢ ꤖ ꤡ ꤑ ꤜ ꤞ ꤑ꤬ ꤜ꤭ ꤔ꤬ ខ ទ ន ឧ ឩ ា ក្ក ក្ខ ក្គ ក្ថ ខ ឃ ច ឋ ប ម យ ឲ ត្រ រៀ ឲ្យ អឿ ន្ត្រៃ ង្ខ្យ ក្បៀ ច្រៀ ន្តឿ ល្បឿ ᧠ ᧡ ᧶ ᧹ າ ດ ອ ມ ລ ວ ຣ ງ າ ອ ບ ຍ ຣ ຮ ວ ຢ ປ ຢ ຟ ຝ ໂ ໄ ໃ ງ ຊ ຖ ຽ ໆ ຯ T H E Z O C Q S H E Z L O C U S f i j k d b h u v x z o e s c n r x z o e s c p q g j y ₀ ₃ ₅ ₇ ₈ ₀ ₁ ₂ ₃ ₈ ᵢ ⱼ ₕ ₖ ₗ ₐ ₑ ₒ ₓ ₙ ₛ ᵥ ᵤ ᵣ ᵦ ᵧ ᵨ ᵩ ₚ ⁰ ³ ⁵ ⁷ ᵀ ᴴ ᴱ ᴼ ⁰ ¹ ² ³ ᴱ ᴸ ᴼ ᵁ ᵇ ᵈ ᵏ ʰ ʲ ᶠ ⁱ ᵉ ᵒ ʳ ˢ ˣ ᶜ ᶻ ᵖ ʸ ᵍ ꓡ ꓧ ꓱ ꓶ ꓩ ꓚ ꓵ ꓳ ꓕ ꓜ ꓞ ꓡ ꓛ ꓢ ꓳ ꓴ ഒ ട ഠ റ ച പ ച്ച പ്പ ട ഠ ധ ശ ഘ ച ഥ ല ᠳ ᠴ ᠶ ᠽ ᡂ ᡊ ‍ᡡ‍ ‍ᡳ‍ ᡃ ခ ဂ င ဒ ဝ ၥ ၊ ။ င ဎ ဒ ပ ဗ ဝ ၊ ။ ဩ ြ ၍ ၏ ၆ ါ ိ ဉ ည ဥ ဩ ဨ ၂ ၅ ၉ ߐ ߉ ߒ ߟ ߖ ߜ ߠ ߥ ߀ ߘ ߡ ߠ ߥ ߏ ߛ ߋ ߎ ߏ ߛ ߋ ᱛ ᱜ ᱝ ᱡ ᱢ ᱥ 𐰗 𐰘 𐰧 𐰉 𐰗 𐰦 𐰧 𐒾 𐓍 𐓒 𐓓 𐒻 𐓂 𐒵 𐓆 𐒰 𐓍 𐓂 𐒿 𐓎 𐒹 𐒼 𐒽 𐒾 𐓵 𐓶 𐓺 𐓻 𐓝 𐓣 𐓪 𐓮 𐓘 𐓚 𐓣 𐓵 𐓡 𐓧 𐓪 𐓶 𐓤 𐓦 𐓸 𐓹 𐓛 𐓤 𐓥 𐓦 𐒆 𐒉 𐒐 𐒒 𐒘 𐒛 𐒠 𐒣 𐒀 𐒂 𐒆 𐒈 𐒊 𐒒 𐒠 𐒩 ꢜ ꢞ ꢳ ꢂ ꢖ ꢒ ꢝ ꢛ ꢂ ꢨ ꢺ ꢤ ꢎ 𐑕 𐑙 𐑔 𐑖 𐑗 𐑹 𐑻 𐑟 𐑣 𐑱 𐑲 𐑳 𐑴 𐑸 𐑺 𐑼 𐑴 𐑻 𐑹 ඉ ක ඝ ඳ ප ය ල ෆ එ ඔ ඝ ජ ට ථ ධ ර ද ඳ උ ල තූ තු බු දු ᮋ ᮞ ᮮ ᮽ ᮰ ᮈ ᮄ ᮔ ᮕ ᮗ ᮰ ᮆ ᮈ ᮉ ᮼ ᳄ ꪆ ꪔ ꪒ ꪖ ꪫ ꪉ ꪫ ꪮ உ ஒ ஓ ற ஈ க ங ச க ச ல ஶ உ ங ட ப ఇ ఌ ఙ ఞ ణ ఱ ౯ అ క చ ర ఽ ౨ ౬ บ เ แ อ ก า บ ป ษ ฯ อ ย ฮ ป ฝ ฟ โ ใ ไ ฎ ฏ ฤ ฦ ญ ฐ ๐ ๑ ๓ ⵔ ⵙ ⵛ ⵞ ⴵ ⴼ ⴹ ⵎ ꗍ ꘖ ꘙ ꘜ ꖜ ꖝ ꔅ ꕢ ꗍ ꘖ ꘙ ꗞ ꔅ ꕢ ꖜ ꔆ 他 们 你 來 們 到 和 地 对 對 就 席 我 时 時 會 来 為 能 舰 說 说 这 這 齊 | 军 同 已 愿 既 星 是 景 民 照 现 現 理 用 置 要 軍 那 配 里 開 雷 露 面 顾 个 为 人 他 以 们 你 來 個 們 到 和 大 对 對 就 我 时 時 有 来 為 要 說 说 | 主 些 因 它 想 意 理 生 當 看 着 置 者 自 著 裡 过 还 进 進 過 道 還 里 面                      P�F                   �eG     �E     pPE                      E     0E     @E     raster1                        �       �eG                           �cE                     ltuo    PzE     �|E     zE      dE     `fG             ltuo    �yE     �cE     �cE     �vE     @dE                     ~E     �~E     �~E     �~E     �~E     �~E     �~E     �~E            �       �hG                            }E                     ltuo    ��E     ��E     ЉE     p}E     `hG                    �       �hG                            }E                     ltuo    ��E     ��E     ЉE     p}E     `hG                    �       �hG                            }E                     ltuo    ��E     ��E     ЉE     p}E     `hG             ltuo    ��E     �|E     �|E     ��E     �}E                     @�E     �E     ��E     p�E                     smooth-lcdv smooth-lcd smooth unknown compression method invalid window size incorrect header check need dictionary invalid block type invalid stored block lengths invalid bit length repeat oversubscribed distance tree incomplete distance tree invalid literal/length code invalid distance code incorrect data check      too many length or distance symbols     oversubscribed dynamic bit lengths tree incomplete dynamic bit lengths tree     oversubscribed literal/length tree      incomplete literal/length tree  empty distance tree with lengths                ��E     �E     P�E     �E      �E     P�E     `�E     ��E     0�E     ��E      �E     0�E     x�E     ��E     w�E     �E     �E     A�E     ��E     ٫E     ֯E     رE     h�E     ��E     ̲E     ��E     ��E     ,�E     ��E     �E     5�E     =�E     �E     �E                                        	      
                                                                        ?      �   �  �  �  �  �  �?  �  ��                              P     W    S     [    Q     Y    U  A   ]  @  P     X    T  !   \     R  	   Z    V  �   �  `  P     W  �  S     [    Q     Y    U  a   ]  `  P     X    T  1   \  0  R     Z    V  �   �  `  `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �   `        P         T  s   R        p      0    	  �   P  
      `           	  �             �      @    	  �   P        X          	  �   S  ;      x      8    	  �   Q        h      (    	  �            �      H    	  �   P        T         U  �   S  +      t      4    	  �   Q        d      $    	  �            �      D    	  �   P        \          	  �   T  S      |      <    	  �   R        l      ,    	  �            �      L    	  �   P        R         U  �   S  #      r      2    	  �   Q        b      "    	  �            �      B    	  �   P        Z          	  �   T  C      z      :    	  �   R        j      *    	  �      
      �      J    	  �   P        V         �      S  3      v      6    	  �   Q        f      &    	  �            �      F    	  �   P  	      ^          	  �   T  c      ~      >    	  �   R        n      .    	  �            �      N    	  �   `        Q         U  �   R        q      1    	  �   P  
      a      !    	  �            �      A    	  �   P        Y          	  �   S  ;      y      9    	  �   Q        i      )    	  �      	      �      I    	  �   P        U         P    S  +      u      5    	  �   Q        e      %    	  �            �      E    	  �   P        ]          	  �   T  S      }      =    	  �   R        m      -    	  �            �      M    	  �   P        S         U  �   S  #      s      3    	  �   Q        c      #    	  �            �      C    	  �   P        [          	  �   T  C      {      ;    	  �   R        k      +    	  �            �      K    	  �   P        W         �      S  3      w      7    	  �   Q        g      '    	  �            �      G    	  �   P  	      _          	  �   T  c            ?    	  �   R        o      /    	  �            �      O    	  �                                                                   	   	   
   
                                               	            !   1   A   a   �   �     �                     0  @  `                                                                                                          p   p                         	   
                           #   +   3   ;   C   S   c   s   �   �   �   �                 ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     ��E     �E     �E     ��E     (�E     h�E     ��E     ��E     X�E     0�E     xF     xF     `F      F     �F     @F     P;F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F      ;F     [:F     [:F     [:F     [:F     [:F     ;F     [:F     [:F     [:F     [:F     [:F     �<F     [:F     [:F     [:F     `<F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     [:F     �<F     [:F     [:F     [:F     [:F     �;F     [:F     [:F     [:F     �;F     ;F     ;F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     8=F     8=F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �:F     �;F     pHF     0TF     pHF     �SF     0SF     �RF     (RF     (RF     (WF     �VF     �UF     �HF      XF     `HF     �PF     �PF     �OF     pHF     0TF     hNF     hNF     �MF     �MF     �SF     (WF     �LF     �KF     �JF     pJF     �UF     �TF     �TF     BNF     \]F     \]F     \]F     \]F     BNF     \]F     \]F     \]F     \]F     \]F     BNF     \]F     \]F     \]F     \]F     \]F     BNF     \]F     \]F     \]F     \]F     \]F     BNF     BNF     \]F     ]\F     2\F     '\F     �[F     bF     bF     bF     �pF     �pF     �pF     bF     bF     bF     RpF     pF     �oF     �oF     bF     �oF     GoF     3bF     3bF     joF     bF     ejF     FjF     jF     �iF     oF     bF     woF     mpF     �pF     `F     qF     bF     �bF     �bF     �pF     �pF     �pF     kF     �jF     bF     RpF     pF     �oF     �oF     bF     �oF     GoF     dF     �cF     joF     bF     ejF     FjF     jF     �iF     oF     bF     woF     mpF     �pF     `F     qF     bF     bF     �cF     kiF     �hF     �gF     iF     �lF     �lF     �lF     �lF     �lF     �lF     �lF     �lF     �gF     �gF     �fF     �fF     �fF     �fF     �fF     LfF     /fF     fF     �eF     �eF     3eF     �dF     �lF     �dF     CdF                                               (       @�E     ��E     ��E     ��E                                                             (       P�E     ��E     ��E     ��E                                                             8       �E     ��E      9F      9F                                                             8       ��E     ��E      9F      9F                                                             ������������������������������������������������ 	�������
 !"#������
 !"#�����               �F                   ��G                                                     ��G      �G     ��G     ��G     @�E     ��E     pF     �F     `�G     ��G      �G             `@F     �F     rF             p
F     p�E     �4F     ��E      5F     �F     p5F     �E     `�G      �G     ��G     @�G     ��E     ��E     �9F             `F     ��E     ��E     rF     @	F     @�E     @1F      �E     `1F     @F     �1F     ��E     p F     ��E                     ��E     0�E      �E     ��E      �E     P F      �E      �E      �E     0�E      �E     0�E     ��E                             ��E     ��E     � F     ��E     �G     /�G     9�G     B�G     v�F     g�F     R�F     S�G     R�G     D�G     G�G     Q�G     [�G     h�G     s�G     }�G     ��G     ��G     ��G     ��G     ��G     ͒G     ْG     �G     �G     �F     �F     ��F     �F     ��G     �G     �G     �G     �F     &�G     )�G     -�G     1�G     5�G     7�G     E�G     ��F     ��F     Q�G     U�G     _�G     p�G     ��G     �G     ��G     ��G     ��G     ��G     ̓G     ��F     ƸF     �G     0�F     B�F     ۓG     ޓG     =�F     ĸF     �G     �G     �G     �G     ��G     ��G     ��G     ��G     ��F     ��F     �G     Ascender true StartFontMetrics AxisLabel AxisType B CH CapHeight CharWidth CharacterSet Characters Descender EncodingScheme EndAxis EndCharMetrics EndComposites EndDirection EndFontMetrics EndKernData EndKernPairs EndTrackKern EscChar IsBaseFont IsCIDFont IsFixedPitch IsFixedV KP KPH KPX KPY L MappingScheme MetricsSets PCC StartAxis StartCharMetrics StartComposites StartDirection StartKernData StartKernPairs StartKernPairs0 StartKernPairs1 StartTrackKern VV VVector W0 W0X W0Y W1 W1X W1Y WX WY XHeight psnames                              
�G                   ��G                     @�F                             ׷F     ��G                     ��F      �F     ��F     @�F     ��F     �F     �rH     �pH                     #   &   5   ;   H                           Delta Omega fraction hyphen macron mu periodcentered space Tcommaaccent tcommaaccent            �  �  "  �   �  �  "  �                                4 j�?�}	�
���W��hXn GM�I� k �!7"�#�:
@zH�PmXh]=b�j[ros�z�������՞l�s�������̦���Q�A� A � � ����(9R[���E� � � � �����e�������n������l�������e� � �����l�������e� � � � � �����e���������c���������w������e����������e������e��c y����n����c(-�e�$������x� �BJU]iq����e���������w������e����������e������l�������e����e��������l���������c�d���������e� ������s� �����������c�������n������l����t������w�������n������e� ������l�����������e��i��������c�������������e����a��1����s��m?G����n� �������e��!�����k����g� �hpx����e������w� ����l�������l��a����e� ������l������������n�1B� B���
".6�����e�$���t�������t�����w�e����������c���������n�2�a�����k����������w���������e��"��������l�������l��b�����r��C� CU�������a]ho�������n�>���e���n���w����l���c������n������a� �������e�����l�����c���e�$������x���t�
������t�
����������l���h������������n�Ie#gs�����������������c���������c�'d)U�������r6J����������������c���������c����������������c����������n�C�����������������c�����������������������c��i����k���������������l�����������e��#��������n�Q����l��cD� D�
$`y���� 09Z������n��a�������n�4�����n��c.5>Y���n������a���cFK�e�$�����������w����t���thq�����t�
����w�e����������c�������c����a�"�����k�����k��i�������s����������e�������e�������l������������k�����������c���������w���������e��$������������l���s")���h����l��d�����r��z��CKp����n��eQe����������������c���������c����������c�E� E���Y����$^����	,	m	s����e� ������l�������e�c����O���n�����������e���������n�5��c���e�$������x� � +3?G����e������w��������w������e����������e������l�������e��������c�dak������e�������s� �w����l����t��������t�����w����������c�$����e� ������l���h���������n�7�������e��i����������n�!g�����������e���������������c�dl�������c���������n�!jm,HS����n�8@����e�����e��������c��������e��%nhs���������c�����������������c��g�J����������c�������������c��o������k���n�������n�������s��r���������c� ������d����������c�-s			!	%�������c�!����������������c��h�����l��et	4	N	\a��	<	F������n�8����s��h� �	T����l������e��	e����w���o� ��h��	|	�����n���������d��F� F	�	�	�	�	�	�

�����e�$���������t�e	�	���������n�V������c�����k��i	�	����������c�r������n�!d��������e��&�������n�!c����l��fG� G
3
=
k
s
�
�
�'4AZk������e�3�a
E
L
^���e����a��
T������n�����������c������e�c
}
�
�
����n�������a�"��c
�
��e�$������x����������t�"��t� 
������t� ��������c�h
�
�!���������n�Be
�
������������������c���������������c���������������c����k�����������n�3���������c�mGO����n� �������e��'���e���c����l��`sq����l��gz���k������e��H� H����(Mu������5����3�%ϴ3�%��1�%�����3�%�������e�3�a�� ����������������c������������������c���������������c�*b�r�&��������w�*c.7�����a�(��c?D�e�$������x�$dS]������s�&�tdm�����t�"����w�$��������e��(o���������n�@�������c������l��h����������t��������l���������e�3�I� I���%^�����0Vc�����������c�/J�2��������c�.����e� �����l�������e�,c-4T���n����c<A�e�$������x� �L����l���������c�dfp�������e�������s� ��������e�.�������c������l����t�0�������t�0����w��e��������������c���������c�������r�!����e� ������l�����������e��i �������c������������e�
������������c�m6K����n�*@�������c���������e��)���������n�;okv~�������c�����k�.�a�����������n���������s������s��s�����l��i����e������e�(�����w�,�����a���������c�t���������������c�vJ� J)5CO��������n�A���c �e�$������x�4��������c�����������n�K��������e��*����l��jK� Ks}�ALj�����������e�3�������e�3�a���������������������c��c����e�0������c�����������������c�������������c����a���������������c�����������������������c��c#,4���n�������a�6����e�$����������t�6�������w�2eR^��������n�T��������n�?hr~���������c�%�������c����k�����������c���������w�4��������e��+���a���������c������k��s����������c�n���l��kL� L	_�����J��L���a���e�9���a��c'.7R���n�=�����a�;��c?D�e�$�����������w�<���������t�;��t�?ir�����t�?����w�6|�����n�8����������n�<j�����������c�	��������w�:��������e��,s�����h�A�����l������l��lM� M��!:GS[d������e�3��c��n���
����l�����e�>�����e�$���t)2�����t�@����w�B���������n�D��������e��-����l��m�����d��u��N� N������!-:BTJ������e�Cc�������n�G�����a�E��c���e�$�����������w�J���������t�E��t�������t�D����w�F�������t���������n�!hj��	��������c�
��������w�H��������e��.���������n�F����l��n����e� �L����l���u��O� Ov���N��0E���5E�R|����l�������e� ������l���b������d���������c�����������������c�����e�Nc���D���n�������������e����c���e�$������x� � (4<����e���������w������e����������e������l�������e��������c�dVm��l]e����e�P����e�������s� �{��������c������l���������w��g����������l������e� ������l���h���"�������n�Um�!&o��������e���n��������e���������w������e����������e������e������������t�Pi��6�����������e�mOk������n�L[c����e�R����e�P��a�!&y����������c�`����k��������������c�zt�������������c�|���s������n�������s���������e��/������n�!`o������k��������n����n��s!(���h� �����e������l������l��o���������e��t;F�������c�~���e� �S[f����e�L�������s�N����l���P� P�����������e�T�����e�$���������t�Ve����������c���������n�J�����������������c��h��i����k��i������������n�S��������e��0si���������c�p���l��pQ� Q*3?�����e�$���������e��1����l��qR� R_w�����+aep�������n�L���e�Tc�������n�X�����a�V����e�$����������t�Vd��������e��t�������t�X����w�Z������n�\���������n�P������r�!�o���n������l�������������e���������w�^��������e��2����l��r5�������d��B�������r��S� Sg7���Tiu��Fu��Mw�0	��������ɱ���0�%����0�%����0�%����0�%����0�%<����0�%,����0�%4����0�%����0�%$1��鰰��0�% ����0�%����0�%a2	%-5=E����0�%b����0�%V����0�%U����0�%c����0�%Q����0�%W����0�%]����0�%\����0�%[3W_go����0�%^����0�%_����0�%Z����0�%T4
���������հ���0�%i����0�%f����0�%`����0�%P����0�%l����0�%g����0�%h����0�%d����0�%e����0�%Y5���	����0�%X����0�%R����0�%S����0�%k����0�%ja,���e�Z ��������t�d�������k��cCbk�����n�`NZ��������t�f����l��������a�^��a��u��������c�����������������c����c���e�$������x�\���������t���t�������t�`����w�b���������t�he����������n�M�������n�!fh"0;Ha�������n�G�������c�(����������c�)�������c�����������c����������c��iZ`��a�������n�!e��������e��3��������������c�,����l��s���������k��T� T��� `�����.�u����r�fc�������n�d�����a�b��c���e�$�����������w�p���������t�b��t�����t�j����w�le*5IR�������c�"����������������c�������n�!i����������c��hhn���a��oty�k���n� ������l����������n�!bi���������l������������n�O��������w�n��������e��4o���������n�9�e������e����x����o��������������k��s'��������c�&���������c����l��tw4@��������n�!k�����n�!aU� Ui{��EW����������e� �s����l�������e�lc������n����c���e�$������x� �������w�v����l���������c�#d��;�l������e�p����e�������s� ��"*3����e������w�rc���n��������c������e�������n������l���������w������e� �O����l���h]�ocm������e���n��|��������e���������w������e����������e������e������������t�p��������c��������������e���������c�xm�
����n�j���������c���������s�z�������e��5�����k�r�����n��15Zy�1��a;Q������������������k�������n���������s��g��������������k�����������l������s�����g�ns��������������c����l��u������t���������c���������������c������e�h������e�x����w�tV� V    < C O [ c�����e�$��������w�~e % 0�������c���������n�N���k����������e��6��������n�H����l��v����e�|W� W { � � � � �����e�����c � ��e�$������x�td � �������s���t � ������t������w������e����������e��7����l��wX� X � �!!!#!/�����e�$�d �!������s���������t�����������n�=i����������e��8����l��xY� Y!Q!t!�!�!�!�!�"("4"<"Da!W!h���e� �!`����l�����������c�b���c!}!��e�$������x�vd!�!�������s�x!�����l����t!�!������t������w���r!�!���������c�+����������������c������e�����k��!�����e��i"""�������n�E�������c����������n�R��������e��9����l��y����e���s"K"q��g"S"^�������c�j���������������c�l�����e"|"��������c�f���������������c�hZ� Z"�"�"�##Q#�#�#�a"�"��������n�6���e�yc"�"����n�}"�����l�����c"�"��e�$������x����t�{"�#�����t�{����w��e##!#L�������c�d#'#:���������������c����������������c���a���e#\#g#w#��������n�:������������c���������c�d#�#����������������c����������������c����������w����������e��:s#�#����l��z����e��a� a$&�''D'�'�((D(~(�)F)�*�*�+1�1�2 2�34`4�5{5�689929�9�1�'$2$r$�$�%%Z%�%�&&Z0�'!$J$N$R$V$Z$^$b$f$j$n0�'^1�'a2�'b3�'c4�'d5�'6�'e7�'f8�'g9�&`1�&$�$�$�$�$�$�0�&e1�&f2�&c7�'	8�'9�'2�&$�$�$�$�$�$�$�$�$�$�0�$`1�$a2�$b3�$c4�$d5�$e6�$f7�$g8�$h9�$i3�'$�$�$�$�%%%
%%%0�'v1�'w2�'x3�'y4�'z5�'{6�'|7�'}8�'~9�'4�'%2%6%:%>%B%F%J%N%R%V0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�5�'%r%v%z%~%�%�%�%�%�%�0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�6�'%�%�%�%�%�%�%�%�%�%�0�'�1�!�2�'�3�!�4�!�5�'�6�'�7�'�8�'�9�'�7�'%�%�%�%�&&&
&&&0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�8�'&2&6&:&>&B&F&J&N&R&V0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�9�'&r&v&z&~&�&�&�&�&�&�0�'�1�'�2�'�3�'�4�'�5�'�6�'�7�'�8�'�9�'�2�'&�&�&�&�&�&�&�&�&�' 0�'&�&�&�&�&�&�&�0�'�1�'�2�'3�'P4�'R5�'n6�'p1�'2�'3�'4�'5�'6�'7�'8�'9�'"3�''' '$'(','0'4'8'<'@0�'#1�'$2�'%3�'&4�''5�&6�')7�'*8�'+9�',4�&'\'`'d'h'l'p't'x'|'�0�'-1�'.2�'/3�'04�'15�'26�'37�'48�'59�'65�''�'�'�'�'�'�'�'�'�'�0�'71�'82�'93�':4�';5�'<6�'=7�'>8�'?9�'@6�''�'�'�'�'�'�'�'�'�( 0�'A1�'B2�'C3�'D4�'E5�'F6�'G7�'H8�'I9�'J7�'(( ($(((,(0(4(8(<(@0�'K1�%�2�'M3�%�4�'O5�'Q6�%�7�%�8�%�9�'V8�'(Z(^(b(f(j(n(r(v(z1�%�2�'X3�'Y4�'Z5�'o6�'q7�'r8�'s9�'h9�' (�(�(�(�(�(�(�(�(�(�0�'i1�'l2�'m3�'j4�'k5�'t6�'u7�'[8�'\9�']a(�(�(�(�(�))������i�	����e� ����a�	�u(�(������i�
������i�
������������i�
>�������e�3��������n)*)4);������i�	����a�	>�������i�
�b)P)y)�)����������n)_)n�����������n�_�������a�	p�����i�	�������o�1���e�)�)�)�)�)�)�����e���������c���������w������e����������e������e��c)�)�*9*���n����c)�)��e�$������x� �*
***%*1����e���������w������e����������e������e����e� �*I*T*e*l*u�������b�c*Z*_�b���b����a�	T�����d��������b�A������c�0d*�*�*�*�*�������e�����������i�
q��a�	������s� �*�*��������c�������n���t*�*�����w�������n��e� �*�*�+����e�������n�1P�����n����i+!+5-�-�.1o0+'+.���8� ���1� ��0+>-V-�0	+R+f+�+�, ,^,�,�-1+Z+^+b7�8�9�2
+|+�+�+�+�+�+�+�+�+�0�1�2�3�4�5�6�7�8�9�3
+�+�+�+�+�+�+�+�+�+�0�1�2�3�4� 5�!6�"7�#8�$9�%4
+�+�, ,,,,,,,0�&1�'2�(3�)4�*5�+6�,7�-8�.9�/5
,6,:,>,B,F,J,N,R,V,Z0��1�2�3�4�5�6�7�8�	9�
6
,t,x,|,�,�,�,�,�,�,�0�1�2�3���4���5�06�17�28�39�47
,�,�,�,�,�,�,�,�,�,�0�51�Q2�63�74�85�96�:7�;8�<9�=8
,�,�,�,�- -----0�>1�?2�@3�A4�B5�C6�D7�E8�F9�G9
-.-2-6-:->-B-F-J-N-R0�H1�I2�J3�K4�L5�M6�N7�O8��9�R1-`-�-�-�0
-v-z-~-�-�-�-�-�-�-�0�S1�T2�U3�V4�W5�X6�Y7�Z8�[9�\�0�^4-�-�-�-�5�6�b7�r8�t9-�-�-�-�-�2���3�_4�c5�s6�u8-�-�3-�-�1���2��ȴ6�ٲ�9� �0..0� 1� �7..b/�/�0�1"1i3.".08.(.,1�j8�9.B.F.J.N.R.V.Z.^2�`3�a4�b5�c6�d7�e8�f9�g4.r.�.�//./f/�0.~.�.�.�.�0�h1�i3�7�9�!1
.�.�.�.�.�.�.�.�.�.�0�"1�#2�$3�%4�&5�'6�(7�)8�*9�+2
.�.�.�.�.�.�.�///
0�,1�-2�.3�/4�05�16�27�38�49�53///"/&/*0�61�72�83�94�:4	/B/F/J/N/R/V/Z/^/b0�@1�A2�B3�C4�D5�E6�F8�H9�I5	/z/~/�/�/�/�/�/�/�0�J1�K2�L3�M4�N5�O6�P7�Q8�R�0�G5/�/�/�0/�/�/�/�/�5��6�~7��8��9��1/�/�/�/�/�1�y2��3��4��9�ҳ4��60 00
0050s0��6� ��5���8��600!0%0)0-014��5��6��7��8��9��7
0K0O0S0W0[0_0c0g0k0o0��1��2��3��4��5��6��7��8��9��8
0�0�0�0�0�0�0�0�0�0�0��1��2��3��4��5��6��7��8��9��90�0�0�0��4��*5��+70�0�0�0�00�0�0��K5��10�0�0�6��7��8��3��5911
111113��4��5��6��7��8��9��81*1V1[01:1>1B1F1J1N1R0��1��2��3��4��6��7���9��41a1e1��2����9��61w1�1�11�1�1�1�21�1��8�!�9�!��2�!�71�1�1�3� ,4� -5� .��4� ���7�m���7��g1�1����e� �u1�1������i�
������i�
h1�1�������a�0B�������e��i22)202<2U2e2�b22�����i�	�������o�1���a�	��������c���u2C2L�����i�
������i�
������������i�
Hn2q2z2�2�2������c�9����������c���������������c��������������c�������������e���������n2�2�2�������i�	����a�	H�������i�
�k2�2�������a�0�2���������h��q����n�1Ol34G4Pe34Bf��3)323A3O3�3�4%43�����c�'�����������w��0����������c���h3U3����a3^3����e3h3q�����c�#����������c�������w3�3������c�%����������c�������w������������w��O�a3�3��������e3�3������c�"����������c�������a3�3�44�����c�I����������c���������������c��������������c�������������w��.�����������w��/�h�!5�����l�"L��a��4X����s��m4j4r4}4�����n��������e��A������d� &4�4���������e������l��&�����e�3�n4�4�575A�������o�1"g4�4�4�5/�������o�1$����������i�Z�e�" 4�5 5'������t4�5���t�05 �������l��?����t�0	5�������l��@���t�#)����t�#*����m�!+������a��u5G5S��������a�	R����a5_5i5p������i�	����a�	�������i�
������k�p5�5�5�a5�5���������e�3 ��n�$��������e5�5��������n�Z��d��p5�5��e����o5�5�����s�"Px5�5�����l�"H5�������e�"R�����������l�"Er66*6.6[��a66!������n�1������n�1�c�#i646B����������g���g� �6K6S����e������w���w6o6v6�797k7�7�8���h�!�d6~6�6���h6�6�6�6����n�!����t�!�����t�!��p�!��l6�6�6�6�6����h�!����n�!����t�!�����t�!��p�!���n�!�6�6�6����t�!�����t�!�����e�!�h6�70��d7	777(������d��������d���������d������d�������x������t�!�7F7W7c��l�!�7N�����e�!���������t�!�����e�!�����t�!�7{7�7�7���������e�!�����y�'��������t�!�����e�!���b7�7����t�!�����t�!��p�!�7�7�7�7�d7�7�n�!�7���e�!�������e�!����t�!�7������n�!�����t�!�����e�!������x���s88e8�8�8�c88S�i8&8=�����m� ^81��������e��>����e� ~8G��������e��^���t�Q8\�����d�R���l8n8y�������a�0A�������a�0�8���������h��g����s8�8�k� *8�8�8�a8�8�����������c�m����c�mm8�8���h�"�������e��
����l��am� B������r�������������������l�"Ct� @999"9*���e� ���������e�� ����l��k����d�Pu9@9Y9`9y9�9�b9F9O�����i�	�������o�1 ���a�	�u9g9p�����i�
������i�
����������������i�	�������������i�
L��������n9�9�9�������i�	����a�	L�������i�
�����������a�	=y9�9���������n�a�n��9�:�����������w�� �����w��b� b:.:�:�:�:�<<I<�>H>T>>�>�@@'@0a:>:H:`:g:�:�:�������i�	�������h� \:T��������e��<���a�	,�u:n:w�����i�
������i�
,h:�:�������a�0p����i�?�������a�0�r� |:���������e��\�������o�1�����e�$���t:�:������t�����w�e:�;;;�;�;������������������s�&lc;;���e�"5������c�1h;(;1;?;];������c�(����������c���i;E;T�����������c��������a�0y�e;d;q���������c�����i;y;������������c���������������c����������������c��m�������a�0���������n�bt��;�;�;�;�a��;�����������k�������h��1;������w��1�����w�����������w��Lh<<Ca<<#<*������i�	����a�	-�u<1<:�����i�
������i�
-��k�Si<U<`<k<y<��������a�0s�������a�0�����������k������������i�
�������e�31l<�>7>Ba<�>2�k<�<�<�=r=�=������e�%�d<�<������d�%�������������������e�%�l<�=Je<�=���������g<�=������r�%��������e�%���������������t=!=5���t�0=*�������l��;����t�0=?�������l��<���r=S=b�����������e�%�������������e�%�r=x=��������e�%������������g=�=�������r�%��������e�%�s=�=�=�m=�=���������e�%���������e�&;����e�%���r�&��p=�>�r=�=������������e�%�������������e�%�������g>>'������������e�%��������e�%��k�$#�������w���k�%���������e��Bo>\>i>t���������i��������a�0|�������a�0�����n�$�������e�3�r>�?�?�@�c>�?8e>�>�>��x������t� {>�>�>�>�>��t���m>�>��d����������e��[����l��[�p����������l��7����t� }??
? ?(?-�t���m??�d����������e��]����l��\�p����������l��8��t?@?j���t� [?O?T?Y?e�t����x�����������e��;�p�������t� ]?z??�?��t����x�����������e��=�p�����e��?�?�?��������b�.��b��������d?�?�?��������b�/��b���������b�a���e?�?��������b�*���������������b�:������r� �s@@����e��������r��������r��u@8@C@N�������a�0v�������a�0��l@U@s�t� "@^@h������e�%��������r�"���e�%�c� c@�AiAtA�A�B0C�D�E+E\HTH\HfHrH�a	@�@�@�@�@�@�@�A*A3�������n�n������i�	����e����a�	�u@�@������i�
������i�
������e�3���������uAAAA������i�	���b����a�	�������i�
������k�!�rA;AAA[��f�!�n��AJAU�������b�,��b�����������n�!��������o�1cA~A�A�A����n������a� �A�����e�	��cA�A��e�$������x�	��l�UdA�A��t�A������t������e�3�eA�A�����a� �A���b�'�t� �A�BBB%iA�B����e�!������r�����������e����������e����������r���hB<B{B�C>C�aBFBQB[Bb�������n�y������i�	����a�	�uBiBr�����i�
������i�
�������o�1eB�B�B�CCC%����������������c��cB�B�����k�'������c�GdB�B��������rB�B�����������������c���������c����������������c����������n�s�����������������c�����������������������c��i��CD���hCQCtC�C�aCWCf�����������n�2w����������n�2�����������n�2i�����n�1J����������n�2	oC�C��hC�C�C��nC�C�����i�
���i�������i�	�����i��k��iC�DC��cC�DDD&D4aC�D �����������n�2v����������n�2�����������n�2h�����n�1H����������n�2�����������n�2�cDJD��e�%�DWDbDgD�������y�"��t�"�pDmDs��s�"���������k�06���hD�D�������������k�%��������������k�%������x��D�D��������b�-��b�lD�D�E��r�#'��kD�D�D�D��������r�������l��������l����������x���b�&cE���tEE#����k�&c����e�&gmE3EAEL����������e�3��������e��C������������e�3�oEnEyE�F�G�G�H=HF�������n����n� :E�E�E���nE�E�����y� ������e��sE�E���n� ����l��U���������rE�E�������d����d��mE�F��a� ,E�F'F2F>F\FsaE�F	F���eE�E���b��������b�����t���rFF���c������n�]�������r�����������e���������dFKFV�������b���d��sFbFi���l��P������r��������dF~F��������b���d�����s�&<nF�F������t�"EtF�F�����������l�".��l�#F�F�F�F�G+GXGfGkGpGuG{G�G�G���K� BF�F��L� S� CF�F��N� R� DGG!G&CGGGG1� 2� 3� 4� �L� �E� EG7G;G@GEGJM� �Q� �T� �C� TGPGTB� X� FG^GbF� S� �S� �T� 	�F� 
��K� �S� SG�G�G�G�G�I� O� G�T� �X� �B� �N� �S� �T� ������t� �G�sG�G���s������f���rG�H,���������tG�H	���t�0G�G���������h��b�������l��A����t�0HH!��������h��c�������l��B�������������e�3�����e�3�����������e�3�����n�$�������o� ���������d���rHyH��yH�H���d�"��r�"�����y� ��rH�H�H�H�����e������x�������e������x���d� dH�JnK�K�LrMDM�N;NHNQNkN�N�O�O�O�O�PaH�IIIYI�I�I�I�J1J7JU�������n�d������i�	�dII&I,I:IJ�����c�6��a�	&����������c���������������c��������������c���gIaIrI���h��Ii�����w����r�  Iz��l� !uI�I������i�
������i�
&�������a�0`�������a�0�lI�I�I������c�/�t��I�I������h��3I������w��3�����w������������c�����aI�JJ�����c�O��������c�O���aJJ)����������c�L����c�L��a�	d��aJ?JH�����w�����������w�����������������������b��bJvKsK}l	J�J�KKKK&K8KFKQ����e���aJ�J�����������tJ�J����t�0
J��������l��=����t�0J��������l��>rJ�J������������������b�+��wJ�J����t�!�����t�!�����a�	e����e���K��b��������l�",������e� K2��b�3����������b�?�������d���������lK^Kd��r� �����������b�������o�1	�����e�3�cK�K�K�K����n������a���cK�K��e�$�����������w����t�dK�LL'LZaK�K�K�L ������i�	����a�	!�uK�K������i�
������i�
!lLL�����c������������c���������a�	\�aL0L:LA������i�	����a�	"�uLHLQ�����i�
������i�
"�tLaLj�����t�����w�eL�L�L�L�L�L�MM?cL�L�������������rL�L������c�k������n�k������c�4���e� ��iL�L������w�������a�0g������c���������a�0�lL�M��eL�M���t�#+����t�#&�a��M�����d����������������������������������i�	��h��hMJM|aMRM\Mc������i�	����a�	'�uMjMs�����i�
������i�
'��k�WiM�M�M�NNNaM�M�����������s��M���b�D���d�&fM���������e�&b�����s� �M�M�M�M�M�����e����������b�$��b�����e�������s���������a�0b�������a�0�������k�0�iN$N/�e� �N+s�"#��������h�"���������c�R�����e�%�lNWNb�������w������e�3�mNqNy����n��������e��D�����k�%�o
N�N�N�N�N�OOO'O�O���������i�������i��������a�0i�������a�0����r� $N�N�N�O �������r�����������e���������e��$sOO���l��i������r����g� ��������e�3&tO5OFO\OgO�O������t��O@��b������cOQOV�b�#��b�#�������a�0����sOpOti�1j���Oz���������k�����h�"���������e�%������������h��O������w�������kO�O��������b���d������n�$��������r���tO�O���l�V����r��uO�P�������a�0e�������a�0�z��PP(P;P`�����e��cP.P5���n����l��ePAPU����������������c���������c�U���������c�_e� eP�P�P�Q�Q�RR%R<RqS�TT�T�U|U�U�V$VYWW�W�W�X8aP�P����e� ���h�&AbP�P�P������i�	�������o�1���e�cP�Q)Q7QWQ�aP�Q#���aP�P�Q���a�	�������i�
���������nQQ���a�	E�������i�
���n�����������e�hQ=QH�������n�e�����������n����cQ_Qd�e�$������x� �QyQ�Q�Q�Q�Q�����e������w��������w������e����������e������e��������c�TdQ�Q�Q�Q�������e���a�	������s� ��t�Q�Q������t�����w��eQ�R	�������i�
������������i�
G��������c�DgR+R2���e� �������i�
�hRFRQR\Rf�������n�g�������o�1������a�0H�������e��iR{R�S�S��������o�1��t� 8R�R�R�R�R�SSSLSnSzS�S�S�S������c�h������i�	������e�$gR����������������f�'����a�	n��nR�R������e�$qpR�R����n�$�����d�$��uSS�����i�
������i�
nhS%S?aS+S6�������c�h�����u�0(���������d�&kiSRSd��������������n�2'������r� ���������e���������e��8pS�S����n�${�rS�S���d�$����n������n�!w�������r� x���i�X�����������e���������������c�ekS�S�������a�0�S���������h��toTT�����������i�
t���n�1TlT#T.Tk�������c�;eT4T;���t�"��nTETNTc�����e�$jpTTT[���n�$~����d�$�����n�!z�����s� &Tv�������l�"�mT�T�T�T�T�����n�T�T�����e�����e��������c�<���h� T��������l��1�������e��EpT�T�����������������n�[����t�"nUUUUEUeUt�������o�1#�������c�=dUU2��h� U'�������l��2���������������c��g�KUMUX�������o�1%���������c�������������c������e� oU�U�U�����k������n�1S��n�[U�U������d���������d�\U�U������d�^���k�]pU�U����n�$�����n��U�����s���uU�V�l� =U�V��������e��sVV���l��f������r� |�������e�"arV,V7VB�������o�1&�������c�@������d�XVN�������c�MsVgVrV�V�WW�������c�A����������������c��h��V�V�V�V����l����tV�V����a�	������������a�	F�����������p��������������d�����lV�V��������a�0G�������a�0�V���������h��j������d�!.������r���tW$W>WBWSW�a��W,W6������n�h����s��h� ����e��WK����w�����aW_WW�����hWiWr�����w�����������w�������w�����������w������d��uW�W������n�1a�o� ���������nW�W�W�������i�	����a�	G�������i�
�xW�X,���m� !W�W�XX$�������n�\dXX�l� <��n� �X����l�����������e������l��!��������l�"�h��XCXVXacXIXP���n����l���������d�����l��f� fX�X�X�X�X�Y]Ym[u[�[�]!])aX�X�X�X����a�	^�������i�
^�������t�!	��aX�X�X������c�N��������c�N��������c�K�������o�1�����e�$���������t�eX�YLYVhYYY-Y=�rYY���c�A�����n������������c���������������c��������������c���������c�����e�&@f�� YeYii��l��i��Y�Y�Y�Y�ZDZUZ]Zj����nY�Y������e�$npY�Y����n�$�����d�$��������h� ���dY�Y���x�%����t�%���lY�Y�ZZ!Z1��f��Y�Y������h��:Y������w��:�����w����m��Z�����w����n��Z�����w���e��Z(�����w������i��Z;�����w���������������e������e�%����������c�s�e� 5Z�Z�Z�Z�Z�Z�Z�[[#[/[:[[[c[n�����c�e������i�	������e�$dZ����������������f�'����a�	k������s�!]�uZ�Z������i�
������i�
k�aZ�Z��������c�e�����u�0%i[[��������������n�2$������r� ���������e���������e��5p[@[G���n�$x�r[N[T��d�$����n������n�!t�������r� u���i�Ul��[{���n��m[�[��������e��F�����e�3�o[�[�[�[��a[�[�����i����i���������i�O���l�" �r� 4[�[�\\!\(\A\\\~\�\�\�\�\�\������c�d������i�	������e�$c\���������������f�'����a�	j�u\/\8�����i�
������i�
j�a\H\S�������c�d�����u�0$i\b\t��������������n�2#������r� ���������e�����������������i�	��������e��4p\�\����n�$w�r\�\���d�$����n������n�!s�������r� tt\�]��n\�\������e�$mp\�] ���n�$�����d�$�h]]�i�T����������e������n�$��a]0]8����n� D�c� �g� g]a^+^B^^�_A`:`�`�aa'aCaYb"b8b�a	]u]]�]�]�]�]�]�^������i�	����e�����a�	f]�]�]�]������c������������c���������������c��������������c����u]�]������i�
������i�
�������a�0L�������a�0���a��^^���������l�c�������r�����������c��b^1^;������o�1���e�c^L^S^\^r���n�������a�#��c^d^i�e�$������x����������t�#��t�!^������t�!e^�^�^�^�^�_8�������c�3�������a�0R�������a�0����������������l�"Qr^�__��h^�^�^������������w�������w�������������w��������s� ������m_ _/�����������w�������w�������k�0h_M_�``*`0a_W_a_x_�������i�	�d_g_r�������n�r��a�	�u__������i�
������i�
�n_�_�_�_������c�:����������c���������������c��������������c���e_�_�` �����������������c���������������c���������������c���a``���a�	Z�������i�
Z��k�`������e�3�i`B`M`X�������a�0N�������a�0�m`^`i�������n�c�l��`r`������h��2`}�����w��2�����w�����������c�S�����l`�`��������������e�����p��`�`�`�`��������d����d���������d��`�`���d���������r�������e��a�������d��maa����n�!�������e��Goa-a8�������a�0T�������a�0��aaJaP��n�$������e�3�ra_a�aaeam����t�"�e� `a~a�a�a�a�a��������b�ca�a��b� ��b� ���a�	S�����d����������e��@������b�@����r� >a�a�a�b����l�"ea������s�"���������e��oa�bra�b���������t�"s���s�"w�������l�"g����l��esb(b0����t�a����e��ubBbMb�b��������a�0P�lbTbm����tb^be���t� �����t� �����lbwb~���t� 9����t� :�������a�0����������e�3������e�3�h� hb�eZe}e�e�gZgnhKhWhci�i�i�i�jjab�ccc7cPc�c�c�c�c�c�d6d?ab�c���������������c������������c��������i�	��ec c2��������������c���a�	9�uc>cG�����i�
������i�
9hcZcccqc������c�-����������c���icwc������������c��������a�0o�����������c�����������e�3*�������a�0�c���������h��������������i�
M��ac�c������c�!��������c�!���������r�1drdd������������c�J���ndd(���������p�!�����������p�!������e�3���fdId�e ����h��d]dbdpdyd�d��6��2dhdl3��f�������w�������������w��������������w�����������w�������s��d�d�d�d�d�d�d�b���8���4�������w�������������w��������������w�����������w������l��eee e%e.e=eM�7���4���0�������w�������������w��������������w�����������w��bebegeq�r�'������o�1��������w�+ce�e������a�)��ce�e��e�$������x�%de�e�������s�'�te�e������t�#����w�%e��e�e�ff�gg5g>gK��t�&ee����te�e�����k�&e����e�&a�����h��4f
�����w��4hf!f=fEfwf�f�af'f5����������c������c�G����w�������afPfo�tfWfc��������c�����������c�������c������������ef�f�����������c����������������c���if�f�������af�f�����������c�������c��������a�0x������af�f�����������c�������c���������������e�3{kgg&������a�0�g��������h��������������e�36�����k�g���������e�39t��gQ�����w�����k�fgc�������r��igxg�g�g���hg�g�g�g�ag�g������������n�2{����������n�2�����������n�2m�����n�1N����������n�2�������a�0r�������a�0�g���������h�����q��hhhhh.h>�4��2hh1��d�������w�������������w��������������w�����������w����������w����������e��Ho	hwh�h�h�iiini�i��������n�p�ih�h�����i�+�����a�0{�������a�0�h���������h�����m��h�h�h�h�h�h�h��9���6���2�������w�������������w��������������w�����������w�����������i�.oiidki(i4i:iP��������b�	��b�	������������������b�!����������������b�"������e�3Briti�iizi������c����������r� ���b��������s�&h��e�#����n�$��������r�������d�eui�i�i�i��������a�0u���������e�33�������a�0�i���������h������������t��j��b�v������n� -j'j2j>jU�������r�����������e��sjDjK���l��c������r�����o� i� ij�j�j�j�n{n�oo3o�o�o�ppiqqYqaqnq�q�rrF�cj�j���e� �������c�Obj�j�j������i�	�������o�1'���e�-cj�j�j����n����cj�j��e�$������x� �������c�Vdj�knPnq������e�	eknK�����hk k.k;m�nn n,����������e�2����������e�2��ckZkjk�llElblrl�l�l�mmFm�m�������������n�2?cktkk�k��������n�2:����������e�2����e�0ok�k�k���a�0k����t��d����������������n�27����������e�2�ek�k�k���������n�2/�������������n�2=�������������e�2�fl	l�����������n�2@ill;������ll*l3�����e�2�����n�26������n�2+hlKlV�������n�22��������e�2�������������k�0llzl�l����rl�l������e�2�����n�28��������e�2��������e�2�ml�l�el�l������������e�2��������n�2.�������n�2*��������n�24pl�l�����d�0���������e�2�rm	m9emmm+�������n�2C�����������n�29����������n�2>���������e�2�smRmom}m�m�emXme���������e�2�������n�2B����������n�23pm�m���e�0 ���������n�25tm�m��������n�21�������n�2;um�m������n�20�����������n�2<wm�m���������n�2,�������n�2-���o�0mm�n���������e�2���������e�2����������e�2���������e�2�wn2n?���������e�2���������e�2��a�	������s� �n^nf����e�/�������c��������w��en�n�n�������������c���������c�5��gn�n�n�n�an�n������������n�2u����������n�2�����������n�2g�����n�1G����������n�2gn�o ���e� �uoo�����i�
������i�
hoo(������a�0D�������e��ioEoOoZoaozo�o�o�������i�	��������c�8���a�	�uohoq�����i�
������i�
������������i�
@�����������e�������������c�9��������no�o�o�������i�	����a�	@�������i�
�j�3ko�o�������a�0�o���������h��r����n�1clpp
�e���������w��mpp^ap#p7pP���n�+p,�������c�����������������������l�"S����������i�
?�������e��Inpupp�p�p�������t�"�����y�"��������n�ktp�p�ep�p����l�"+p�p�p�bp�p�����m�#!t�#!�x���tp�p��p�# p�# �������n�")������e�3vp�p�q�����t�%������e�%���������e�&;oqq!q)�������c�Q����k�/�a��q4qIqQ�������s��qA����s������n�i����s������n�$����������i�
rsqxq�q�q����lq�q��������a�0C�������a�0�q���������h��h����������i�	�����e�h������r���tq�q�������nq�q��������a�0��������a�0����e�)q�����w�-urr�������o�1)�������c�N��������nr*r4r;������i�	����a�	?�������i�
������arQr\�������c�u���������������c�wj� jr�r�r�sss�s�s�s�s�ar�r�r�r��������n�q������i�	����a�	�ur�r������i�
������i�
�������o�1cr�r�r����n����cr�r��e�$������x�5���������l��������������e�_ess&sg�������c�X�ms1s:sHsX�����c�,����������c���������������c��������������c���hsmsv�����c������������c���hs�s�as�s�s�������i�	����a�	�us�s������i�
������i�
���������n�{�s�0��������e��J����n�$��������r��k� ktvnvyv�v�ww*x�yZygy�y�z<zRz_zvz�z�at/tOtet�t�uu,uEu�u�v8vUbt5tF�������������c�������i�	�ctUt[��e�1������c�:�etlt~��������������c���a�	f��t�t�t�t�t�t�t������c�C�����h��;t������w��;����������c��������w��������������c��������������c������������w��M�ut�u�����i�
������i�
huu������a�0K����������c���������a�0�u9��������h��vpuKu`�a��uR����������k������nuluzu�����������n�1qpu�u������������n�1����������n�1x���������������n�1y����������e�3su�u�vvv(�������ou�u������c�@������������������c�@�����������a�0�����e�3��avv�����c�P��������c�M������������c���������������������������h��p���������������������c���������o�1cv�v�v�v�av�v�������e�3���n�������a�7����e�$����������t�7�������w�3ev�v�w whv�v��������n��������a�0Q�������a�0�v���������h��y��������n�o������������a�0�����������c�8hw8w�w�w�x4x�awDwNwYw`wy������i�	��������c�E���a�	�uwgwp�����i�
������i�
hw�w�w�w������c�.����������c���������������c��������������c����������c���aw�w����a�	Y�������i�
Y����hw�xxx&aw�x �����������n�2x����������n�2�����������n�2j�����n�1K����������n�2
ox>xoxyx~�hxIxRx[xe�����i������i�������i�������i�������i�[�k������������i�������e�3�ix�x�x�x��������a�0M�������a�0�x���������h��w�ox�x�x������������e�3������������e�3�����e�3���kyy'y6y?yMay
y�����������n�2n����������n�2�����������n�2`�����n�11����������n�2 ���������n�13���������c�\lymyx�������w�5�����e�3�my�y�y�����������e�3��������e��K������������e�3�oy�y�y�z
zhy�y�������a�0S������e�3��ay�y�����i������a�0�y���������h��z��������e�3����������c��rzz2����������������l�2������b�C�azCzI��n�$������e�3����������c�otzezn�����e�3�����d��uz|z��������a�0O�������a�0�z���������h��x������e�3�������e�3�l� lz�|�}}V}|~~~-~E~W~�~�}�����az�z�z�{{{-|�������i�	����e�:���a�	2�u{{�����i�
������i�
2������������i�Em
{C|||=|K|^|n|�|�|�a{I{���f{U{c{�{�����������c�������a{m{�����e{w{�����������c����������������c�������w{�{�����������c����������������c����������������c������������e{�{�����������c����������������c�������c�D��a��|�����e���d��| |4�����h��<|+�����w��<�����w������������c������������������c���������������c�������������������c�������������������c����������������������c����e|�|����������c����m|�|����������������c���������������c�����������e�%�b|�}}
�r����t�l������o�1c}}%}.}I���n�>�����a�<��c}6};�e�$�����������w�=���������t�<��t�@}`}i�����t�@����w�7}s�����n�9e}�}�~�t}�}�������������b������������b��s� <}�}�}�~����l�"d}���������r�"���������e��o}�}�r}�}����������t�"r������r�"v�������l�"f����l��d�h�n�����k�%�������������x�mi~3~8�a� ����������n�lj��~K��������c�Yl���~c~{~�~�a~i~p���a�	3�������i�
��������w�;�����a�	4������c~�~�~�������i�	����a�	a��������n~�~�������i�	����a�	cm~�~�~����������e�k�������e��L�����e�3�o:EKu��������i�,����l"5��d�"'��t� �*�������d�#�r�"(�������i�%��s�����eUlc[g��������e��N�b�2�����d��M����e�%�����n�$�s������h�B����e�!������r��������e�%�����i�&������c���������i�	����a�	��������n��������i�	����a�	b������e�3�m� m�#�����Ă݄�(�_�}����/�H�Q�l��a�=�G�������ׂ3�L�Q�_�k�p������i�	�c�M����n� ��[�f�l�u�������b�1��b������d����������e�����e�?���a�	.�u���������i�
������i�
.h��������h���������w�����������w��������a�0~i��(�g���'�������a�����w����������i�����������i������i�K������������i����k�1�P�W��w�9�D�������i�����������i������i�H������������i���������t�s�~�������i������i�1t����������u�����������i������i�G�o���с���w�����������i�����������i������i�I������������i����i�����w����������i�����������i������i�J������������i�����������i�F�������a�0ނ@��������h����e�&B����������e�3G��������w���s�&Bs�v����������������w������e�3�b����������o�1�����e�3�c��������e�$����������e�3���t�̂������t�A����w�Ce��l�w�����ă�e��_m�����$�����c�E����������c���������������c����e�+�8���������c�����i�@�O�����������c���������������c��H���������e�3M�������a�0������������e�3~�������a�0დ��������h���m�ރ��������h��>�������w��>�����w����������n�t���a�ۃ������w�������a��������w�����������w�����������w��h����k�q������e�3�i�6�[����A�d�=�V���������������������h��e�t� ���m�i��������a�o�~�����������n�2r����������n�2�����������n�2d�����n�1Ap����a��������������n�1p��������n�2���������n�1n���������n�1o�������a�0�������a�0߄���������h����u��<s�"��&�/�5�������b� �����e�"���d�����s�"�e� 2�i�H�V����������e�3J�����e�3Il�e�t�����������d�p�����e�3�m����������������e�3��������e��M������������e�3�o���ԅ��� h����������a�0�������e�3��������a�0����������h���������e�3������i�!���������e�3��������e�3��a� �&��n�$������e�3�s�5�>�����e�3�������r��������d�ou� ��o�s�}���������ن�����X�b1� �������e�3��h����������r�"k���s�"j������e�3�g�������k�������e�3��������a�0��������a�0�����������h���l�߆������e�3�����y� �������e�3���h�������w�����������w��s��O�c�'�8�C�����e�&j�2��l�&k�������n�&m��������n�&o�����e�3�������e�3�������e�3�v�r����������e�3������e�3�w�������������e�3������e�3�n� n�ԈZ�r���͉��T������̋��F�4�<�U�]�=�G�Qa������!�,�E�Qb��������i�	��a�"���e�D���a�	(�u�������i�
������i�
(�������a�0j�������a�0ʈ9��������h�����������e�I�����e�3�b�`�j������o�1����e� �c�|���������n�H�����a�F��c�����e�$�����������w�K���������t�F��t���������t�E����w�Ge�Ո����������a�0m�������a�0͈���������h�������������n� �������e�3�g��Ia��)�0������i�	����a�	�u�7�@�����i�
������i�
�������i�h�Z�d������a�0���k�l�s���t�r��������x�si���2�=�w��n�����މ����#a���������������n�2o����������n�2�i�ŉ���������n�15���������n�2a����������n�16�����n�14�a���
����������n�1h��������n�2���������n�1g�����������n�1f�������a�0kk�C�[������a�0ˊO��������h�������t�e�p�������i������i�M�e� 9�������ǊΊ��$�0�;�\�d�o�����c�i������i�	������e�$h�����������������f�'����a�	o�u�Պ������i�
������i�
o�a����������c�i�����u�0)i����������������n�2(������r� ���������e���������e��9p�A�H���n�$|�r�O�U��d�$����n������n�!x�������r� yt�u����n�}�������e�$rp�������n�$�����d�$���i�Yj�̋���������c�Z�������a�0����������h���l�ҋ�����������g���������w�Im����������e��N�����e�3�n��=a���$������i�	����a�	#�u�+�4�����i�
������i�
#�����a�	)o�T�_�x���q�(�������a�0n�������a�0Όl��������h���n������������������e� ������i�����i��n�����Ɍ���$�_�����c�F����������c��������a�Ԍ������c������������c���������������c�������i�������������c���������������c��K�e�+�8���������c�����i�@�O�����������c���������������c��N��������������c���t�������̍؍��������s�"e���������t�"	���f�"	���l�"`������r�"o����r��������l�"q���s�"y��������l�"b���s�"n���������l�"pp���������l�"&������s�"��u������t�"������s�"������t�"���������n�v����n�$�s�B�K�����e�3�������r� ����e� �u���i�t�ŏ�������a�0lk�z��������a�0̎���������h����a������������i�	����a�	<�u���������i�
������i�
<m�ˎ�������n� #�َ���������e������l��_�r�������n�������k�t���������k�uo�!n��� �4�����h��@�+�����w��@�����w��������e�3�������e�3��a�Z�d�k������i�	����a�	�u�r�{�����i�
������i�
o� o���Đ�����;���ˑ������H�i����G�Sa�������e� ������i�-b�Ώ�������d�u�ڏ��������c�����������������c�������i�	�������o�1���e�Oc��c��a� �]���a�+�2�=���a�	�������i�
���������n�K�R���a�	I�������i�
���n����c�k�p�e�$������x� ���������������e���������w������e����������e������e��������c�>d�Ɛݐ���l�͐�����e�Q����e���a�	������s� ����������c��������w��e�S�
�����n�1Zg��*�1���k�ۑ$��b�(���e� �������i�
�h�E�P�Z���������n��������a�0Jo�`�j������e���n���y������������e���������w������e����������e������e������������t�Qi���������������e�k�ё�������a�0�����������h��u����n�1W�������w��m�
�&�-����������n�M������e�S����e�Q���a�	P��a�ɒ=�A�L�Z�j1���������c�a����������d�w������������c�{t�p������������c�}���s���������i�
�����n��������s���������e��O�e� 1�Ւޒ���(�1�J�l���������ٓ��������c�a������i�	������e�$`�����������������f�'�d����a�	g���������r� $�����h�![�����d����u�8�A�����i�
������i�
g�a�S�^�c�������c�a�f� ������u�0!i�r����������������n�2 ������r� ���������e�����������������i�	��������e��1p�������n�$t�r�̓���d�$����n��������r� �����n�!p�������r� ��h����i�Q��d�!So��2�Bg��(���k�������n��������i�
������������i�
K��n�Tp�P�W�b���n�$��������t�%����n�#%r�o��d�u���������e� ���������e� ��������l�"s���Ôԕ����t�������a�	������������a�	J���h� �������e�����l�ݔ��������a�0I�������a�0�����������h��k���������e��������r���t��)�������c����e� ��4�<����e�M�������s�O��������o�1!v�Y���r�`�����e� >�m����c�s���������e��J�b�d��������d��I�����y��L���y��K����e� ��������n���Õ�������i�	����a�	K�������i�
�p� p���{�������P�Z�R�e���ٝ\�d��<�X�ba��9�C�J�Q���������Ԗ���oa��+��������e�3�����������e�3+������i�	����e�U���a�	*g�W�ie�]�d���n�!��p�!�u�o�x�����i�
������i�
*�������a�0q����������i�/�������a�0�l�������������������������b��������������c������������n�1r�����a�������h� ����l�"%�n��t���t� (��,�1�6�A�M�d�i�����������c��>�t����x����������r� ���������e��s�S�Z���l��Y������r� }�p����������l��5����t� )�������������ӗ������������c��?�t����x����������r� ���������e��	s�����l��Z������r� ~�p����������l��6�������f�"s�����������w����������w������e�3���h���'�5�:�C�R�b1�-�11��d���a�������w�������������w��������������w�����������w����������w���������o�1�����e�$���������t�We�䘱���Иܘ�V�a�v�I�������c�?�����h��D�������w��D��������e�3;����������������w��Ch�����)�G�r��
���c�~�����n�z����w������������c��Wi�/�>�����������c��X�����a�0z�����������c��Y�������a�0������������������c��r�������1�>��������w��N���t� %�����������c�j��������e������l��ji����d� .�ϙڙ�����������n���������d� ���������h��a�������r�����������e��s�����l��R������r�����������������b�B���������r�"��������d� 0���a� �������e�3�h�b���a�j�t�{������i�	����a�	+�u���������i�
������i�
+i�ƚ�������1�����h���֚��a���������������n�2z����������n�2�����������n�2l�����n�1M����������n�2����n�x�������i�:����������k��o�%�*�D�k���h�1�:�����i�������i�����������i� i���`�4�?�J�X��p�p�����ϛݜa�v�������������n�2s����������n�2�i������������n�1v���������n�2ek��������������n�1r����n�1B����������n�2���s��k�������������n�1t����n�1D�����������n�1ut��&�����������n�1w����������n�1s�������a�0t�������a�0�����������k�����������n����s� +�s�~�����������b������e�"�m�������s� �o����d��������e��s�������l��b������r� zm�Ŝ��������e��P�����e�3�o���3�>�H�������a�0}����������x����)��������e�&��������e�&���������e�&������e�&�������a�0�������i��������k�0�U���e�0 ����n�$�r�l����e�r�z����s�"z��������n�!��e������d���������d� 5o�����������t�"������e�#���������a�0�p�͝�e�ӝ����r�#��u������t�"������t�"������n�"7���l�"s��3i�Ȟ��������c�q��������������������b�������e�3�u�B�M�������a�0w�������a�0�������e�3�������e�3�q� q�������ş̟؟��a�����០d������a�	X�������w��f�����������c�B����������c���������������c��������������c������s��������$�-�<��1� ��0��a��c��2��7��9���3���e�������w�������������w��q�B�����n�O�X�g�w�����w�������������w��������������w�����������w�������������w�����������w���������������w���������o�1�����e�$����k����������e��Q�f���������h��G�������w��G�����w������n�$�u���u����������e�&i���s���1�6�;�@�I�X�h�8���5���1�������w�������������w��������������w�����������w�������n� ?�����������r�������c������n�^���n� �������l�������k�~��������e������l��?��e�ء�3�P��l� "���������e� ���t� ��������e������e�0��������d�0����t� ���t� �(�������d� r�9�C������d� ���t� �Ln�I����l�Z�a���e� e� '�g��������e��r� r�������ף
��3�����٦��#�ŧЧ�Wa�����ơ͢��7�B�[�r���������n�|������i�	����e�Ud�סݡ���a�	0���l�"���x�������������e�3���������e�3������e�3��e��������w���u�%�.�����i�
������i�
0�������a�0��������a�0�O��������h����������������������i�	�m�x���������������������i�	�����n�d��o�"6�������o�1c�����¢����n�Y�����a�W����e�$����������t�Wd�ݢ�������e��t��������t�Y����w�[������n�]e��E�h������f��+���������k� ;����u�5�<���t�"������t�"������r�P�U�d� �s�[�a��s������f���h�p�����r�w�~���c�1�����n������������c���������a�0��������a�0죬��������h����h����������������w��H�����w��v������������e�"=�a���������w��������������w�����������t�#�������k�~�(�������d�h�9�Pa�?�I������i�	����a�	]o���Z�w���k�}�a�����d�{�l�������r������������k�����������d��i���̥�������l	���٤���$�2������a���������������n�2q����������n�2�����������n�2c����������n�1@k�������k�������n�1:���������n�1i����n�19����������n�1;p�:�Z�ia�@�N����������n�1l��������n�2�����������n�1?���p�r�{�����n�1<���������n�1k���������n�1=t���������������n�1>����������n�1j����������������n�1m��t�ԥ�����e�"t�������������b�������e�"��������a�0��������a�0���������h���n�$��g�ڦ.�9�?�������b�%��b�
���f�H�v���t���U�`�k�������n�Y�������b��������d������t�������������b�9�������d������������e�����������e�3Ql�����������w�_�����g�|�������d�z��������e��Ro�����������a�0��������a�0���������h���������i�#����n�$�r�+�O�ma�3�=�D������i�	����a�	1�������i�
\�h�V�_�����c������������c���������c�}������������i�	����a�	`�������i�
���������n������������i�	����a�	D�������i�
��������r���t�֧�����k�%�����d�y���������r��u����!�P�������a�0��������a�0���������h���p�'�J�e�.�<����������i�	�����������i�	���h������i�$������c�g�q�x��������i�	����a�	�������i�
���������n������������i�	����a�	C�������i�
�s� s�٪��ƫD�k�1�<�˳U�����]�����˶��ηx��a	�����T�m�x������������i�	����e�[� ��������t�ed��!�'�5�E�����c�5��a�	8����������c���������������c��������������c����u�[�d�����i�
������i�
8�������a�0U�������a�0�����������h��{����������������������������c������h�᩼�������h��A�������w��A�����w���a��0�8�j�ra�����!�)����i�2����i�A����m���������i�D������i�C����i�3���i�0����i�@i�@�X�ci�F�Q�������i������i�5�������i������i�4����i�Bu�z����e������e�����������i������i�7�������i������i�6���i�8����i�9�������o�1c�Ҫ��!�7���n�a����������t�g�����a�_��a�Y�����������c�����������������c�����k�Z��c�)�.�e�$������x�]���������t���t�L�U�����t�a����w�c�_��������t�ie	�������Z�u���߬�������������b�<c������d� 3������������e�����n� ��n���ƫԫ������c�3����������c���������������c��������������c�����l������#�2�B�M1��3��f���c�������w�������������w��������������w���������w�����������w��h�`�k�������n�}������a�0[�������a�0�����������h��~�i��������n� ;�����������c���������e������l��T�������������a�0�����������h����t���������e�3"������e�3#��n� 7��%�/�M�T�^�w�������˭���������c�g������i�	������e�$f�:���������������f�'����a�	m������s�!^�u�e�n�����i�
������i�
m�a�~���������c�g�����u�0'i������������������n�2&������r� ���������e���������e��7p�ѭ����n�$z�r�߭���d�$����n������n�!v�������r� wt��+��n�������e�$pp��#���n�$�����d�$���i�W�������n� �h�L�2�=�K��!��a�Z�e�o�z�	�"�������n�w������i�	��������c�Hd�����a�������������c�Q����a���������c��a��������c��^����������c��`����a�ˮ������c��b��������c��_e�%���������k�%�����t�%������m�%��a�	6�u�������i�
������i�
6������������w���������o�1����������c�Ie�U�������n�`�i�w�������c�4����������c���������������c��������������c���������c����l� ��������w� ��a���¯ѯ߯���1�ȯͱ5��5��2�ׯ�2��e�������w�������������w��������������w�����������w�����������c��i�'�2�������c��n��<����d�B������h��I�N�W�����w��Is�]�q�����t��,�h�����w��,����t��-�{�����w��-�������w�������w��s���������t��*�������w��*����t��+�������w��+��k��i�ݱ	��-�K�S�`���a�ð���1������l������������������k���������a�0W�������a�0��!��������h��|��q�5�>�����w�����������w������r�"<���������w���s�o�����αܱ�a�u�������������n�2t����������n�2�i������������n�1~���������n�2fk��������������n�1z����n�1E����������n�1{p������������n�2���������n�1}�����������n�1|x� 6�)�2�<�Z�a�z�����òβ��������c�f������i�	������e�$e�G���������������f�'����a�	l�u�h�q�����i�
������i�
l�a�����������c�f�����u�0&i������������������n�2%������r� ���������e���������e��6p�Բ����n�$y�r�����d�$����n������n�!u�������r� vt��O��n��:c������e�$o������������������������i�	�p�@�G���n�$�����d�$���i�Vl�[�o��h� /�c��������e����g��w��������t��m����������e�&:�������e��So���޳��/�:f��������������w��t�Ƴ������n� ������������c�L�������a�0]�������a�0�����������h������s���������������b�8��������������b�7�������i�)s�B�L�T������i�(����i������i�*�a�f�z���e�  �m���������c�  �e�&`�����t��������k�&`����e�&d��n�$�����e���Ǵմ����(�I�d�����������b�;c�ʹ�c�3�m�3����������������������l�%��������������l�%�k��	g�3�m�3��������l�3�l��#n�3��g�3�m�2�6�;�?g�3��l�3�m�3�������d�3������������������������l�%�����r�n���������������������l�%��������������������l�%������������l�%�������������������k�%�������e�3�s�Ѷ{a�۵���������i�	����a�	7�������i�
��g�
��&�4�C�Q�_�l����������n�1I����������n�1�����������n�1������������n�12����������n�1e����������n�1C���������n�1F�����������n�18������r���t���������g� �����������e������e�����������������b�6��������������b�5u�޶����H�R�V���t�"�����������l�"�������l�"�c������s�"{����t�"�������a�0Yk�%�=������a�0��1��������h��}�������c�R������n�"n�&<�����t�"��c�n�������l�"�������l�"�������e�3��������������e�3|t� t�����չd�����F�����������9��å��a
�ͷ׷���Z�k������������i�	��k�޷����n�"����t�"����a�	$�u��������i�
������i�
$h���-�K�����c�7����������c���i�3�B�����������c��������a�0_�����������c����������������e�3}�������a�0��x��������h�������������c�@u��v�긞������s��J��h��J�������w��J�����w��b�Ƹ��r�g������o�1
c������<�W���n�e���l�������a�c��h����-�����c������������c��{������������c��|�����������c��}��c�D�I�e�$�����������w�q���������t�cd�j�t������s���t�{�������t�k����w�me	�������ɺ�"�e�j���������c�B����������������c��h�Ϲع��,�U�������c�*����������c������i��������������c���������������c��i��#�����������c��������a�0f����i�6�E�����������c���������������c��m�[�}�����a�f�o�����c�)����������c���e�������������c�����i���������������c���������������c����������������c��s�������a�0ƺ���������h���l��������e�!!������k�&���a�������������w�������������w��n�,�5�H�]�����e�$i���������������n�2)p�N�U���n�$}����d�$�����n�!y�h��t�ػt���������h��8������w��8�����w�����������c����r���������w�����������w��h�ʼb�ܽ`��<a�ֻ�� �������i�	����a�	%�u��������i�
������i�
%l�������c�0����������c����������t�,�K�R��w�4�?�������i�����������i������i�L������������i���e�j����h�t�}���������c�+����������c���������������c��������������c����e���������s�"���e�"4�a���ʼ�1������������k��i��8���h���!�*a��������������n�2y����������n�2�����������n�2k�����n�1L����������n�2����n�B�K�����e�$lp�Q�X���n�$�����d�$�o�n����������������������i��k������������i��n� ��h������a����������i�����i�������i�������i�����d�ֽ��������c�����������r��������c�l������n�l��e� 3�)�2�<�Z�a�k�������;���"�*�5�����c�c������i�	������e�$b�G���������������f�'����a�	i������s�!\�u�r�{�����i�
������i�
i�a�����������c�c�����u�0#i������������������n�2"������r� ���������e�����������������i�	��������e��3p������n�$v�r�����d�$����n���������s� �������h�������n�!r�������r� ����i�S������e�3�i�V�a���6�B�s���������a�0ak�g�������a�0��s��������h�����t��������a���������������n�2p����������n�2�����������n�2b�����n�17����������n�2��e�ܿ��� ��(�������b�0c�����b���b���������b�`o��������r�"<��������b�4����������b�>��������e�"�p�H�f��a�P�Y�����w�����������w�����������i�
p�������������b�����������n���������w�o��������e��To���������`�l���������n�i�������a�0h�������a�0�����������h���n���R�We���?�F�L��r��#�-�6����a��������d�������d��������d�������d�������d�����e����x����o���s�������e�3'��������i������������������t�������t�0��������l��]�������l��9����t�0��������l��^�������l��:������i��a������������k����n�$�r���
�������k�!"��s�����s������f��������������k����g�%�*�/�4�n�%��f�%��t�%��p�%�s���E�l������i���O�c�����h��F�Z�����w��F�����w��e�r�}�������c�F�e��¡ª¹��12��e���b�������w�������������w��������������w�����������w�����������c�[������r���t���)�jÝa���	�������i�	����a�	�u�� �����i�
������i�
�h�4�=�K�[�����c�y����������c��g������������c��h�����������c��i�a�s�}Ä������i�	����a�	 �uËÔ�����i�
������i�
 ����d��uíø���������a�0d�������a�0�����������h�������l�����������a�0c�������a�0�����������h��ow��ne��;��e���3�����e�$kp�$�+���n�$����d�$�����n�!{��y�E�N�Y�����e�$s�������u�SDp�_�f���n�$�����d�$�o� 2ĎėġĿ����'�I�U�h�sŔŜŴ�����c�b������i�	������e�$aĬ���������������f�'�d������a�	h�t�����������r� %�����r� %���������l��0�u��������i�
������i�
h�a���������c�b�����u�0"i�-�?��������������n�2!������r� ���������e�����������������i�	��������e��2p�yŀ���n�$u�rŇō��d�$����n������n�!qsŢŪ����e��������r� ��hŻ���i�R���s�!Tu� u������W���ǁǑ���
�[�d�����_�{������e� �b������r�������i�	�������o�1(���e�mc�&�-�M���n����c�5�:�e�$������x� ��E����w�w������c�Cd�c�nƅƋ���������a�	Q�l�u�}����e�q����e���a�		������s� �ƟƧƯ��������e������w�scƵƼ���n��������c������e�������n��������w��g�������e� �u���������i�
������i�
	h���f������a�0Fo��(������e���n���7�?�J�R�^����e���������w������e����������e������e������������t�q�v�������c��������������e�kǙǱǼ������a�0�ǥ��������h��s�������c�y����n�1\m����a�������n�k�����������c���������s�{����������i�
A�������e��Un��G�������e� _�#�)�5�@��l� ��������e��?�������l��3���y��Oi�M�R�n�"*�����l�" �����k�sp�p�w�Ȏ�����n�$�����k�%������������w������n��Ȝȱȹ�������s��ȩ����s������n������s�����k�����������b���d��r������������i�
s��g�os���
�7�����������c�^���l���������a�0E�������a�0��+��������h��i������t�C�N�������c���������������c������e�i�k�s����e�y����w�uuɇɑɘɱ��������i�	����a�	
�uɟɨ�����i�
������i�

������������i�
B��������n������������i�	����a�	B�������i�
���������n����������i�	����a�	A�������i�
�v� v�3������˔˛���	�m�ůa�=�D�]�h���a�	5�u�K�T�����i�
������i�
5�������a�0�v���tʏʯʻ�����h��5ʁʆ�5��5�����w��5hʕʝ����w�����m��Kʦ�����w��K��������w����������w�������e�$��������w�e�����4�?�Eˈ�������c�2h�����%�����c������������c��k������������c��l�����������c��m�������a�0���s�&@�����l�P�V��r� |���e�c�n�y˂�������b��������b�)�����d����d����������n�~���k��iˣˮ���������a�0����a˹����������i�	����a�	M�������i�
�����a������������i�	����a�	�������i�
���������e��Vo���b�������n�x���d�%�I��������n�3�>�������a�0��������a�0��������a�0��V��������h����������a�0�����n�$�t�{̂���e�}����d��u̛̐�������a�0��������a�0�w� w��ͱͻ�����=�E�(�Q�]Шаз����a����������<�H�l���e��������n�1Y�������a�0�k���������a�0����������h�������n�1X����l�&�1�������a�0��������a�0���������e�3Wv�N�V����h�0������������������l��4w�t�}͋�����c�H����������c������������e͚ͣ�����c�$����������c���������e�3����c�����e�$������x�ud����������s���t���������t������w��e����3�������a�0���������s�!k�!�+������a�0�����n�1^������n�1]����e�����e�Z�cη��eϒ���������t�%�c�i�}����e�%��s������e�%������������tΎ΢���t�0Η�������l��C����t�0ά�������l��Ddν�������d�%�����������������������������d�%�����������g���������������e�%��������e�%��e��B���������g�'�7������������e�%��������e�%���������������t�V�]���t�0����t�0������������g�wχ������������e�%��������e�%�sϚϸ��mϠϬ��������e�%���������e�&:����e�%���r�&t�����������e�&������������������t�������t�0����t�0���������g��������������e�%��������e�%�i�.�9�������a�0�k�?�I������a�0�����n�1_��������e��Wo�g�rЋН�������a�0��������a�0����������h��fn� �Б��������e����������i�'����n�$����g���������r�������d����n��x� x��������!�.�2�>�F�������b�=�������o�1�����e�$�d��������s���������t�����������n�mi����������e��X����n�$��������r��y� y�s�J�a҉�g�oԀ�������������aыїѡѨѯѹ�������>��������e�3N������i�	����e� ����a�	/������n�1R�u���������i�
������i�
/�������a�0�k����������a�0�����������h�������n�1Q���������i�N����l��%�������a�0��������a�0��2��������h��l��������c�c���c�S�X�e�$������x�wd�g�q������s� ��t�xҁ�����t������w��eҙӡӪӼ���(�[hҫҴ�����-�=�xӊ�����c�J�����eҿ�������c������������c�������������c������������e��� �������c�&����������c���������������c��������������c���������������c����e�D�Q���������c�����i�Y�h�����������c���������������c��X��������������c����������������������c�������n�1Vn� �Ӱ��������e���o���������n�1U�������������n�1�r������������o���������w�����������w����������c�K����������������c�������g�5�>�N�����n�1�������������n�1����������n�1���������w������e�����k���x����e��iԌԗԢԫԳ�������n�u�������c�W�����n�1b����g�&/���������n����������e��Yo���"�-�7�]ՋՔd������������h��9�������w��9�����w����d�������w������������w���������a�0�������n�1�k�=�U������a�0��I��������h�������n�1[����l�g�r�������a�0��������a�0����������h��n�����k��y՚տaՠժ������n�1�kհո����n�1����i�"������i�p�������n�$�����������i�z���������b�Er������g���������r��t�����e������d��u�)�4�>�d���������a�0�������n�1�k�D�\������a�0��P��������h�������n�1`s�lֻ֒��g�t��������c�k���������������c�m�����e֝֨�������c�g���������������c�i���l�����������a�0��������a�0�����������h��m�e���������n�1�������n�1��a�	�������i�	����a�	_z� z�:�B�M�xؓٶ�"�L�X�dڀڈژڡa
�P�[�b�i�t���������������n�f���e�z���a�	[�������i�
[h�~ׇו׳�����c�8����������c���iכת�����������c��������a�0V�����������c����n���������c�2����������c����������a�0���f�������������w������������w����������w����n���%�9�����h��6�0�����w��6�����w���������o�1c�U�\�r���n�~��c�d�i�e�$������x����l����t�|؂؋�����t�|����w��eءج������ٱ�������c�7dز�����������������c����������������c���������a�0\�������a�0��o� 0�
���$�=�J�U�a�l�vفو�����c�`������i�	����a�	f�u�+�4�����i�
������i�
f���������c�`�������r� ���������e���������e��0������n���������r� p���i�P����hٔٝ٩�����r�����������r� ����e� �a��hټ���������o�1e���������������n�j������������c���������c�6d������������������c����������������c��i�*�5�@�������a�0X�������a�0���������w����������w����������e��Zo�j�u�������a�0^�������a�0�����n�$�������������k�������e��uڧڲ�������a�0Z�������a�0�                                                                    � �   � � � � � � � �    c � � � � � � � � � �   � � � �   � � �                	  
m n    !"#$%&'()*+,-./                                                                    012    34567  8    9    :;    <=>      � � � ?@ABCDE    F� � � GHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz                                                                        	 
                        ! " # $ % & ' ( ) * + , - . / 0 1 2 3 4 5 6 7 8 9 : ; < = > ? @ A B C D E F G H I J K L M N O P Q R S T U V W X Y Z [ \ ] ^ _                                                                     ` a b c d e f g h i j k l m n   o p q r   s t u v w x y z   {   | } ~  � � � �   � �   � � � �                                 �   �         � � � �           �       �     � � � �         � &-5?JT_hmsz������������������������������ 
(2?KV`bdfhjlnprtvxz|~�����������������������+:=@GNXgqx�������������*17>AMT[^knw~����������������
!'+4BLS_ipv}�������������� $+2<CJV`gmt}���������������")3:FXgv��������� ,:HUcw������������				 	$	6	I	Y	h	s	z	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	�	



"
)
7
A
H
S
c
p
|
�
�
�
�
�
�
�
�
�
�
",9ER[er���������(6CP_n|����������
%1BQZfr~���������$,4<BGLRYag                  �    &-5�JT_hmsz������������������������������ 
(2?K�`bdfhjlnprtvxz|~��������������_p}���C`JVmgt}��������������G����qg�B�� >T  �) 3 ��@ L V ^ a A^j k~���p �x � ��� iv�[�@7�V?�� )2��+:=NXx��S�L��������� �$n�����*1Mw �<3��'+"��!+�
4���� � � � � � � � � � �                             .null nonmarkingreturn notequal infinity lessequal greaterequal partialdiff summation product pi integral Omega radical approxequal Delta nonbreakingspace lozenge apple franc Gbreve gbreve Idotaccent Scedilla scedilla Cacute cacute Ccaron ccaron dcroat .notdef space exclam quotedbl numbersign dollar percent ampersand quoteright parenleft parenright asterisk plus comma hyphen period slash zero one two three four five six seven eight nine colon semicolon less equal greater question at A B C D E F G H I J K L M N O P Q R S T U V W X Y Z bracketleft backslash bracketright asciicircum underscore quoteleft a b c d e f g h i j k l m n o p q r s t u v w x y z braceleft bar braceright asciitilde exclamdown cent sterling fraction yen florin section currency quotesingle quotedblleft guillemotleft guilsinglleft guilsinglright fi fl endash dagger daggerdbl periodcentered paragraph bullet quotesinglbase quotedblbase quotedblright guillemotright ellipsis perthousand questiondown grave acute circumflex tilde macron breve dotaccent dieresis ring cedilla hungarumlaut ogonek caron emdash AE ordfeminine Lslash Oslash OE ordmasculine ae dotlessi lslash oslash oe germandbls onesuperior logicalnot mu trademark Eth onehalf plusminus Thorn onequarter divide brokenbar degree thorn threequarters twosuperior registered minus eth multiply threesuperior copyright Aacute Acircumflex Adieresis Agrave Aring Atilde Ccedilla Eacute Ecircumflex Edieresis Egrave Iacute Icircumflex Idieresis Igrave Ntilde Oacute Ocircumflex Odieresis Ograve Otilde Scaron Uacute Ucircumflex Udieresis Ugrave Yacute Ydieresis Zcaron aacute acircumflex adieresis agrave aring atilde ccedilla eacute ecircumflex edieresis egrave iacute icircumflex idieresis igrave ntilde oacute ocircumflex odieresis ograve otilde scaron uacute ucircumflex udieresis ugrave yacute ydieresis zcaron exclamsmall Hungarumlautsmall dollaroldstyle dollarsuperior ampersandsmall Acutesmall parenleftsuperior parenrightsuperior twodotenleader onedotenleader zerooldstyle oneoldstyle twooldstyle threeoldstyle fouroldstyle fiveoldstyle sixoldstyle sevenoldstyle eightoldstyle nineoldstyle commasuperior threequartersemdash periodsuperior questionsmall asuperior bsuperior centsuperior dsuperior esuperior isuperior lsuperior msuperior nsuperior osuperior rsuperior ssuperior tsuperior ff ffi ffl parenleftinferior parenrightinferior Circumflexsmall hyphensuperior Gravesmall Asmall Bsmall Csmall Dsmall Esmall Fsmall Gsmall Hsmall Ismall Jsmall Ksmall Lsmall Msmall Nsmall Osmall Psmall Qsmall Rsmall Ssmall Tsmall Usmall Vsmall Wsmall Xsmall Ysmall Zsmall colonmonetary onefitted rupiah Tildesmall exclamdownsmall centoldstyle Lslashsmall Scaronsmall Zcaronsmall Dieresissmall Brevesmall Caronsmall Dotaccentsmall Macronsmall figuredash hypheninferior Ogoneksmall Ringsmall Cedillasmall questiondownsmall oneeighth threeeighths fiveeighths seveneighths onethird twothirds zerosuperior foursuperior fivesuperior sixsuperior sevensuperior eightsuperior ninesuperior zeroinferior oneinferior twoinferior threeinferior fourinferior fiveinferior sixinferior seveninferior eightinferior nineinferior centinferior dollarinferior periodinferior commainferior Agravesmall Aacutesmall Acircumflexsmall Atildesmall Adieresissmall Aringsmall AEsmall Ccedillasmall Egravesmall Eacutesmall Ecircumflexsmall Edieresissmall Igravesmall Iacutesmall Icircumflexsmall Idieresissmall Ethsmall Ntildesmall Ogravesmall Oacutesmall Ocircumflexsmall Otildesmall Odieresissmall OEsmall Oslashsmall Ugravesmall Uacutesmall Ucircumflexsmall Udieresissmall Yacutesmall Thornsmall Ydieresissmall 001.000 001.001 001.002 001.003 Black Bold Book Light Medium Regular Roman Semibold rb      ��F     ��F     `�F     ȎF     `�F     `�F     `�F     �F     A�F     Y�F     A�F     œF     œF     ��F     ��F     �F     �F     ��F     �F     A�F     ��F     �F     �F            zR x�  $      p���   FJw� ?;*3$"       D   ����I    A�CD     d   ����2    A�Cm       �   U���   A�CH��       �   5����   A�CH��     �   �����    A�C�      �   ����    A�CH��� (     ����J   A�CP�����5      <  ،��a   A�CJ��R   `  ���-    A�Ch      �  ���    A�CL      �  ���"    A�C]      �  ���-   A�C(    �  ����"    A�C]          �����    A�CE��      $  �����    A�C�     D  1���>    A�Cy      d  ���-    A�Ch      �  /���    A�CP      �  ՚��9    A�CA�s   �  ���3    A�CA�m   �  ���.    A�CA�h     ���5    A�CA�o   $  $���5    A�CA�o   D  9���4    A�CA�n   d  M���6    A�CA�p   �  c���1    A�CA�k   �  t���D    A�CA�~   �  ����)    A�Cd      �  ����)    A�Cd        ����    A�CV      $  ����    A�CZ      D  ����    A�CV      d  ����    A�CZ      �  ����8    A�Cs      �  �����    A�C�     �  >����    A�C�     �  ���u    A�Cp        X���[    A�CA�U      (  ����.    A�Ci      H  ����I    A�CD     h  Ɲ��   A�C    �  ����Q    A�CL     �  ���J   A�CE    �  ���j   A�Ce    �  c���W    A�CR       �����   A�C�    (  ����    A�C�     H  ����?   A�C:     h  ߥ��    A�C        �  ۦ��     A�C[       �  ۦ���   A�CE��      �  n����   A�CE��      �  ���k   A�CE�a        L����   A�CE��  $   <  ����3    A�I�I ]AA ,   d  �����   A�A�O�^
AAG   H   �  ����    B�B�D �A(�D0T
(D ABBFT(G DBB     �  l���&    F�SG�    �  ����1            ����H          $  ���       ,   8  ���k    B�A�D �D0X DAB(   h  $���X    B�D�D �IAB     �  X���z          �  Ķ��/    A�m      �  ض���          �  t���          �  ����#    TN $   	  �����    G�A��
DA   (   ,	  P����    G�A��
AAYA   X	  $���\       �   l	  p���7   j�E�F �E(�D0�A8�GPv8D�0D�(B� B�B�B�TP������P
8G�0A�(B� B�B�B�HI8A0A(B BBBE������PP������     
  ����          (
  ����   A��
D[   H
  �����       0   \
   ���   B�G�G �D@�
 AABA    �
  ����    H�y   (   �
  `���>    B�A�A �vAB      �
  t���<    A�\   D   �
  �����    B�B�E �B(�D0�A8�D@�8A0A(B BBB   <  ���(          P  ���-       D   d  (���m    B�E�B �B(�A0�A8�D@Q8A0A(B BBB   �  P���          �  \���          �  X���          �  T���\          �  ����V            ���           $  ����P       H   8  4���Q   [�B�B �B(�E0�E8��0f(I BFBL������      �  H����      L   �  ���!   T�I�E �B(�A0�A8�G`�8A0A(B BBBH������ ,   �  ����g   J�
HC
E��H�  <     $����    L�I�E �A(�A0�Y(A BBBD�����L   X  t����   F�B�A �A(�# AGBI����h(����} ADB   �  ���          �   ����          �  �����       @   �  h����    T�G�D �fABH���P ���ACBJ���    (  ����&          <  ����          P  ����#          d  ����          x  ����f       $   �  @���   A�A�G �AA$   �  (���#    A�A�G SDA    �  0���          �  <���w            ����Y       <     ����y    G�E�A �D(�D0W(A ABBF����      X  4���!    D\    p  L���#    D^    �  d���         �  `���          �  \���          �  X���f       4   �  ����[    F�D�D r
AAFDCAH��       ����          $  ����          8  ����    D8   L  ����A    G�A�C �b
�A�B�HAABD���   �  ���d    U�|G� ,   �  X���}    B�A�A �X
ABA   \   �  ����7   R�B�B �B(�A0�A8�D`�8A0C(B BBBG������P`������ $   4  ����    A�D�G PAA <   \  �����    J�A�D A
AAFbG�A�G ��   <   �  ����   B�B�E �A(�D0��
(A BBBF      �  �����          �  l���       D     x����    K�A�A �c
ABEI
CBJAFBG���  \   L  �����    K�B�A �A(�D0w
(A ABBHD
(F ABBIh����H0����    �  ����&          �  �����          �  ���^      D   �  T����   B�B�A �A(�q
 ABBD�
 ABBO     0  ����p    dK$   H  4����    e�G pAC�` �     p  �����    D0R
J    �  `���i    D0`
A @   �  �����   ~�G�D �
CBDCADH���h ���P   �  `����    _�J�D �C(�J0N
(L� A�B�B�GD(F ABBA����     @  �����          T  (���Q          h  t���3    R�UI� ,   �  ����i    B�D�A �D0V DAB$   �  ����u    A�D�D0iAA   �  0����       8   �  �����    b�D�G RG�A�Q ��_
CAE<   ,  p����    u�C�G0Q
F�A�ILFAE��h0�� (   l  0����    W�T
�E^
B`�H�4   �  ����c    _�H�J O
F�A�IDCAH��\   �  �����    `�E�E �D(�I0�`�(A� B�B�B�R0�����A(F BBBC�����L   0  �����    e�E�D �H(�J@^
(A ABBDD(F ABBI����  (   �  <���c    a�O [
ADDCI�  $   �  ����^    F�G |
AFI�  L   �  �����    K�B�A �A(�D0f
(A ABBAD(F ABBA���� 4   $  ���\    F�D�K r
AAGDCAA��  4   \  0���g    b�D�D �f
�G�B�GACB4   �  h���I    F�D�G b
C�A�BDFAA��    �  ����;    F�c
�GCE�  4   �  ����S    F�D�G g
C�A�DDCAH��4   (  ����S    F�D�G g
C�A�DDCAH��   `  ����6          t  ���a          �  t���6       H   �  ����p    B�B�A �A(�D0J
(D ABBCD(C DBB     �  ����'    DU
GF   @     �����    K�B�D �D(�F0b
(A ABBEP����  d   L  0����   J�E�B �B(�A0�A8�D@p
8C0A(B BBBK�������F@������      �  ����          �  ����          �  ����          �  ����            ����:       d     ����L   d�B�B �B(�D0�A8�D`�8C0A(B BBBI������A`������U������    �  ����+          �  ����C    Ii
FF      �  ����          �  ����;       �   �  ����   T�B�B �B(�A0�A8�G�U
8A0A(B BBBFP������F�������J������F�������      `  L���f       0   t  �����    [�D�G hCAF��X ��   0   �  $����    S�A�D }AAI��` ��     �  ����          �  ����/       4     �����    U�G�A �A(�� EBBA����    <  ����6          P  ����g    IpzMp     l  ���          �  ���       `   �  (����   B�B�B �B(�A0�A8�DXx
8A0A(B BBBAD8F0A(B BBB   T   �  t���/   Q�F�F �H(�G0�D8�D�U
8A0A(B BBBE�������     P  L���       X   d  H����   B�L�E �I(�A0�D`8
0C(A BBBES
0C(A BBBK     �  �����       D   �  X����    B�E�E �E(�D0�D8�FP�8A0A(B BBB     ����          0  ����(          D  ���       0   X  ���B    A�D�G \
CADJFA 4   �  0���^    F�D�D f
CAHJFAG��     �  X���       H   �  T���}    B�B�A �A(�D0w
(A ABBID
(F ABBA   $  ����       (   8  ����h    A�C�D s
DAH     d  ����+    A�i   X   �  ����1   a�B�A �D(�G0f
(A ABBEt(A ABBF����@0���� $   �  ����4    A�D�G eAA       ����6    A�t          ����          4   ���'          H   $���(          \   @���.          p   \���          �   h���       4   �   t���    A�D�G0u
CAKU
AAI  4   �   �����    A�D�D0U
AAHK
CAI l   !  ���$   B�E�E �D(�A0�G`�
0C(A BBBEN
0F(C BBBCS
0F(C BBBF  4   x!  �����    A�D�D0U
AAHK
CAI 4   �!  ,����    A�D�D0\
AAIK
CAA 4   �!  ����|    A�D�D0M
AAHK
CAA T    "  ����y   B�B�B �D(�C0�G@_
0C(A BBBC�
0F(C BBBF   x"  � ��&          �"  ��&       4   �"  ,��|    A�D�D0I
AADK
CAI L   �"  t���   T�E�D �D(�H@�
(A ABBH�����V@����    (#  ��    DS    @#  ��    DT    X#  ��~    Dy   p#  |��?    Tj    �#  ���       4   �#  ���Q   S�A�D(�
AAEcAAK��<   �#  ����    J�D f
DHC
CJG
ETlFN�      $  ���    DU <   ,$  ����    _�A�A �D0q AABF���H0���      l$  @��!          �$  \��/       4   �$  x��g    A�D�G i
DAFT
DAG  $   �$  ���3    A�I�G0]CA T   �$  ����    B�B�B �D(�D0�J@�
0D(A BBBJL0F(A BBB   0   L%  @��D    A�L�G ^
AADDFA 0   �%  \��D    A�L�G ^
AADDFA H   �%  x���    B�H�E �E(�D0�F8�DPm
8C0A(B BBBE  H    &  ����    B�H�E �E(�D0�F8�DPm
8C0A(B BBBE  (   L&   	��f    K�I�G0AAD��  l   x&  d	��Z   B�B�B �A(�A0�D@�
0D(A BBBB|
0G(D BBBCD
0G(D BBBK  <   �&  T
���    B�A�D �Dpf
 CABID HAB h   ('  �
���    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   h   �'  �
���    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   h    (  ���    B�M�E �A(�D0�D@|
0A(A BBBGH
0A(A BBBHD0F(A BBB   @   l(  @���    K�A�A �D@�
 AABHD FABK���    �(  ���6    IPa 0   �(  ��x    B�D�A �G0U
 AABI t   �(  P���   [�B�B �B(�A0�D8�G`u
8A0A(B BBBD�8A0A(B BBBE������``������  H   t)  ���   B�B�B �B(�A0�A8�Dpy
8D0A(B BBBA    �)  \��6       �   �)  ����   K�B�B �B(�D0�A8�D`"
8D�0A�(B� B�B�B�GT
8C0A(B BBBH������H`�������   X*  ����   K�B�B �B(�A0�D8�D@
8A0A(B BBBEJ
8C0A(B BBBB`������P@������T8J�0I�(B� B�B�B� h   �*  ����    ]�E�D �C(�G0z
(A ABBHO(Q� A�B�B�S0����J(M� F�B�B� (   \+  P��F    F�C�G dF�A�   H   �+  t��   B�E�B �E(�D0�A8�Dp\
8A0A(B BBBCT   �+  8��6   d�B�B �B(�D0�A8�GPD
8A0A(B BBBD�������   \   ,,   ���   g�B�B �B(�A0�D8�D`8A0A(B BBBJ������V`������    �,  ���1    A�Y
FP (   �,  ����    A�Z U
DDv
AA@   �,  ���x    B�E�B �D(�D0�G@o
0D(A BBBF     -  ����    A�Q |Ax   <-  0��9   B�B�B �B(�D0�A8�G`
8A0A(B BBBCL
8A0A(B BBBJD
8F0A(B BBBE0   �-  � ��    A�A�D0c
AAELAA   �-  @!��V    A�c pA X   .  �!��6   K�B�A �A(�D@C
(A ABBA�(A ABBB����H@���� `   h.  d"��;   B�B�B �B(�A0�A8�D`�
8A0A(B BBBID
8F0A(B BBBE h   �.  @#��F   K�B�B �B(�A0�A8�DP�
8A0A(B BBBID
8F0A(B BBBEx������H   8/  $$��>   B�B�E �H(�D0�A8�GPb
8C0A(B BBBE     �/  %��          �/  %��       H   �/  %��x   B�E�E �B(�A0�A8�Gp�
8C0A(B BBBD h   �/  D(���   B�B�B �B(�D0�D8�J�i
8D0A(B BBBHS�M�Q�B�J�N�V�A� l   d0  �/��C	   B�E�E �B(�A0�A8�G���L�\�A�V�L�U�B��
8A0A(B BBBJ    �0  �8��>    IPg |   �0  �8��F   K�B�E �E(�D0�I8�D��
8A0A(B BBBEh
8A0A(B BBBFT8A0A(B BBBJ������H   l1  �9��   B�E�B �E(�A0�A8�G�w
8C0A(B BBBF   �1  D=��F    IPu    �1  |=��       H   �1  x=��q   B�G�B �B(�A0�A8�DPy
8A0A(B BBBJ H   02  �>��c   B�G�B �B(�A0�A8�DPw
8A0A(B BBBA    |2  �?��V    A�c pA    �2  @��       8   �2  @��w    B�B�D �D(�D0e
(D ABBB  (   �2  `@��2    B�F�D �^AB      3  t@��O          ,3  �@��,          @3  �@��          T3  �@��.          h3  �@��          |3   A��F       d   �3  <A��   K�B�A �D(�D0�
(A ABBDD
(C ABBDD
(F ABBI`����  8   �3  �A��V    L�D�D �b
ABGACBJ���      44  B��              L4  B��3    \�QC�     h4  4B���    `�G0^AJ�     �4  �B���          �4  <C���          �4  D���         �4  �H��          �4  �H��          �4  �H��          5  �H��          5  �H��          ,5  �H��          @5  �H��G          T5  �H��M          h5  $I��          |5   I��          �5  I��(          �5  8I��\         �5  �J��8          �5  �J��8          �5  �J��          �5  �J��          6  �J���         6  �L���       H   06  M���   B�B�B �B(�A0�A8�GP6
8A0A(B BBBGL   |6  �O���   B�B�B �A(�D0��
(A BBBE
(A BBBB   �6  Q��!          �6  ,Q��
          �6  (Q��          7  $Q���       (   7   R��9   A�A�D #
AAE   H7  T��S    A�u
JR    h7  TT��    DT d   �7  \T���    L�O�E �E(�D0�C8�F@�
8A0A(B BBBE\8C0A(B BBBA������ \   �7  �T���    B�B�B �E(�D0�D8�G@^
8A0A(B BBBFg8A0A(B BBBH   H8  TU��+   B�B�B �B(�D0�D8�GP�
8A0A(B BBBH `   �8  8V���   B�B�B �B(�A0�D8�D`
8C0A(B BBBC�8F0A(B BBB  `   �8  �W��   B�B�B �B(�A0�A8�G`�
8A0A(B BBBJ�
8A0A(B BBBD$   \9  P[���    A�A�G �AA$   �9  �[���    A�A�D �AA$   �9  0\���    A�A�G �AA   �9  �\��    A�P   4   �9  �\���    B�B�A �A(�G0�(A ABBL   (:  �]��	   B�B�B �A(�A0��
(A BBBNA(A BBB   ,   x:  d_��W    R�G�H �P0a AAB 4   �:  �_��7   A�D�G0
AAHAA 8   �:  �d���   B�B�A �D(�F0�
(A ABBKd   ;  @g��i   B�B�B �E(�A0�A8�G@�
8A0A(B BBBK
8A0A(B BBBC  4   �;  Hk��R    B�G�D �Q
ABG_HB      �;  pk��	       H   �;  lk���   B�B�B �B(�D0�D8�G`�
8A0A(B BBBD H   <  �l��x   B�D�B �B(�A0�A8�D`�
8D0A(B BBBI    h<  $n���    Q�n  4   �<  �n��G    B�E�A �D(�G0m(A ABB (   �<  �n��0    B�D�D �bAB   $   �<  �n��9    A�D�G VAA    =  �n��&    A�P   H   ,=  �n���   B�B�B �B(�A0�D8�D`>
8A0A(B BBBG   x=  Ts��       <   �=  Ps��   K�B�A �A(�G0�(A ABBE����   `   �=  0t��   B�G�B �B(�A0�A8�D`z
8A0A(B BBBIE
8A0A(B BBBA H   0>  �u��y   B�B�B �B(�A0�A8�J��
8A0A(B BBBJ8   |>   }��   B�E�A �D(�G@x
(A ABBG  H   �>  �}��
   B�B�B �E(�D0�A8�Dpx
8A0A(B BBBJ  H   ?  ����7   B�B�B �E(�A0�A8�DPy
8D0A(B BBBI   P?  ����/          d?  ȅ��|       H   x?  4���   B�B�B �B(�D0�A8�FPj
8A0A(B BBBI    �?  ���f          �?  d���]          �?  �����           @  l���7          @  ����<          (@  Ĉ��:          <@  ����7          P@  ���7          d@  H���P          x@  ����U          �@  Љ���          �@  L����       H   �@  ����   B�B�B �E(�A0�A8�G@g
8A0A(B BBBKH    A  \����   B�H�K �K(�F0�H8�Dp
8A0A(B BBBDL   LA  �����   B�B�B �B(�A0�A8�G�&
8A0A(B BBBG   H   �A  �����   B�B�E �E(�D0�A8�J��
8A0A(B BBBCH   �A  ����   B�G�M �B(�D0�A8�Fp�
8A0A(B BBBE L   4B  X���   B�B�B �B(�A0�A8�D�3
8A0A(B BBBA   L   �B  (����    B�D�A �G0I
 CABC\
 CABFQ CCB H   �B  ȹ���   B�B�E �B(�A0�A8�DPE
8A0A(B BBBHL    C  L���?   B�B�B �E(�A0�A8�G��
8A0A(B BBBG   L   pC  <����   B�B�E �B(�D0�C8�I�Y
8A0A(B BBBB   H   �C  ����c   B�E�B �E(�A0�A8�FPi
8A0A(B BBBGT   D  ����    B�G�B �A(�C0�G@�
0A(A BBBGf
0A(A BBBB8   dD  ����   B�E�D �A(�F0�
(A ABBD 8   �D  ����   B�E�D �A(�F0�
(A ABBD `   �D  `����   B�D�F �B(�A0�A8�Dps
8A0A(G BEBGO8C0A(B BBB   h   @E  �����   O�B�B �B(�D0�A8�DP\
8A�0A�(B� B�B�B�LP������HP������  H   �E  ���u
   B�B�E �E(�D0�A8�J��
8C0A(B BBBK$   �E  D���7    A�H�G dAA H    F  \���l   B�B�E �B(�D0�A8�DpA
8D0A(B BBBF D   lF  ����   Q�B�A �A(�G0�(A ABBK����H0����   �F  X���
          �F  T���       4   �F  P���b    B�I�D �Q
ABEkGF   @   G  ����~    A�K�I X
CAG\
CAHG
CAE  $   XG  ����R    A�D�G0CAA   �G  �����    �RL   �G  ����	2   B�G�B �B(�A0�A8�G�D
8A0A(B BBBD   0   �G  T���    A�A�D0�
AAD^DAH   H   ��5   B�J�E �E(�A0�D8�G�W
8A0A(B BBBE\   hH  �#��,	   B�G�B �E(�A0�D8�I�A�h�L�B��
8D0A(B BBBE     �H  �,���          �H  �-��)          �H  �-��          I  �-��O          I  .��          ,I   .��          @I  �-��          TI  .��n           hI  d.���    Z��
FJF�    �I  @/���          �I  �/��    D�V      �I  �/��       \   �I  �/���    B�B�E �E(�D0�A8�G@Y
8A0A(B BBBCR8A0A(B BBB   0J  0��          DJ  0��x          XJ  t0��       $   lJ  p0��M    A�A�D BCAL   �J  �0��=   B�E�B �E(�A0�A8�J��
8A0A(B BBBG      �J  �2��Q    A�G@GAP   K  �2��!   B�F�B �D(�D0�G�h�B�B�K��0D(A BBB   L   XK  �3��T   B�B�D �A(�J�T�c�B�B�K��
(A ABBH`   �K  �4���   B�B�B �E(�D0�D8�DP{
8F0A(B BBBG�
8A0A(B BBBKH   L   7��   B�G�B �B(�A0�D8�J�N
8A0A(B BBBDL   XL  �7���   B�J�B �B(�A0�A8�J�g
8A0A(B BBBC   L   �L  49��   B�J�B �B(�A0�A8�J��
8A0A(B BBBF   $   �L  �:��P    A�D�G }AA H    M  ;��   B�B�B �B(�A0�A8�D@�
8A0A(B BBBE�   lM  �<���   B�E�B �B(�A0�D8�Dpd
8A0A(B BBBF�
8A0A(B BBBK|
8A0A(B BBBJ�
8A0A(B BBBJ  `   N  HA���   B�E�E �E(�A0�A8�J�m�Q�A�A�V��
8D0A(B BBBH (   hN  �F��Q   J�A�G 4AAH��L   �N  I��p    L�F�A �D(�F0s
(C ABBHD(C ABBA����  H   �N  (I���   B�E�B �B(�A0�A8�Hp
8A0A(B BBBF8   0O  �M��n    B�D�D �D(�G@t
(A ABBA  H   lO  N��&   B�G�B �E(�A0�A8�J��
8A0A(B BBBId   �O  �N���   B�B�E �B(�D0�A8�D��
8A0A(B BBBHu
8A0A(B BBBI  |    P  ,U��:   B�E�B �B(�A0�D8�D��
8A0A(B BBBDe
8A0A(B BBBAM
8A0A(B BBBA   (   �P  �W���    {�G�J POAA�� <   �P  �X��P   B�F�I �JP
 AABHK AAB   Q  �Y��
       \    Q  �Y���    B�B�B �B(�A0�A8�D@w
8C0A(B BBBGd8F0A(B BBB`   �Q  �Y���	   B�B�A �A(�I@t
(D ABBDi
(D ABBFl
(F DBBF     �Q  Hc��%    D`    �Q  `c���          R  �c��      0   $R  e���    A�A�D8~
CAHDFAT   XR  te���    B�B�B �A(�A0�DP�
0C(A BBBBD0F(A BBB   X   �R  �e���   B�B�B �A(�D0�G�g
0A(A BBBGA
0A(A BBBG  H   S  �g��   K�G�B �B(�A0�A8��0A(B BBBA������   H   XS  Th���   B�B�B �B(�A0�A8�G��
8A0A(B BBBA<   �S  �i��c    B�B�E �A(�F0�DPF0A(A BBB    �S  �i��1    A�C�kA      T  j��          T   j��<    A�r
EC (   <T   j��C    B�D�A �vCB      hT  Dj��H    A�G ~A    �T  tj��9    K�fG� H   �T  �j���    B�B�B �B(�D0�A8�DPx
8D0A(B BBBJ H   �T  �j��y   B�E�B �B(�A0�A8�G�Y
8A0A(B BBBI<   <U  0o���    B�F�D �G@M
 AABDi AAB L   |U  �o��~   B�K�G �B(�A0�A8�G��
8A0A(B BBBB   l   �U  �|���   B�B�B �A(�H0�G@0
0D(A BBBG�
0G(D BBBCL
0G(D BBBC   <V  0���          PV  <���	          dV  8���          xV  D���;          �V  p���V          �V  ����          �V  ȁ��          �V  ԁ��3    \�QC�    �V  ����
          �V  ���!          W  ���A           W  L���
          4W  H���
          HW  D���
          \W  @���
          pW  <���
          �W  8���
          �W  4���
          �W  0���
          �W  ,���	          �W  (���
          �W  $����          �W  ����          X  ̂���          $X  ����
          8X  ����          LX  ����          `X  ����x          tX  ���          �X  ���(    A�f   4   �X  ����    B�E�A �A(�G0�(A ABB$   �X  ����T    A�A�D ICA   Y  ؄���      (   Y  T���a    I�A�G LAAA�� 4   DY  ����~    U�I�G s
G�A�HDCAH��0   |Y  ����o    A�A�D b
AAFxDA H   �Y  ����   B�B�B �B(�A0�D8�DP�
8A0A(E BBBA H   �Y  ����
   B�B�A �D(�G0�
(D ABBHD(G ABB  0   HZ  t����    B�C�A �D0�
 AABE    |Z  0���;    _[ H   �Z  X����   B�B�B �B(�A0�A8�D�Z
8A0A(B BBBF H   �Z  ���   B�E�E �B(�A0�A8�G�v
8A0A(B BBBI    ,[  ����K          @[  ���       8   T[  �����    B�B�A �A(�D0b
(A ABBF 0   �[  l���6   B�C�A �D0_
 AABC 8   �[  x���    B�D�A �A(�D@o
(A ABBG      \  \���D    A�y
FC D    \  �����    B�B�B �B(�A0�D8�DP�8C0A(B BBBH   h\  D����    B�B�A �A(�D0[
(G ABBOD(A ABB  `   �\  ����D   B�B�B �B(�A0�D8�G` 
8C0A(B BBBHQ8A0A(B BBB   H   ]  t���>   B�B�B �B(�A0�D8�G�V
8D0A(B BBBI$   d]  h���Q    A�D�G0DA `   �]  �����   B�G�B �B(�A0�A8�D`�
8A0A(B BBBJj
8A0A(B BBBD @   �]  <����    A�A�G@c
DAGF
DAER
DAA x   4^  �����   B�B�E �E(�D0�A8�MPh
8A0A(B BBBFd
8A0A(B BBBJ�
8A0A(B BBBA0   �^  ���Z    A�D�G0p
AABWAA    �^  ���W    D l
H  l    _  \����
   B�B�B �B(�D0�C8�J�F
8D0A(B BBBDQ�E�Z�B���\�N�A�   p_  ����V       `   �_  ����   B�B�B �B(�D0�A8�F`�
8A0A(B BBBHZ
8A0A(B BBBD$   �_  4����    A�K�G qAA@   `  �����   K�B�B �A(�D0�x(A BBBE�����      T`  �����    I{
DhP(   t`  x����    B�F�A ��AB     �`  ���N    |M d   �`  $���T   B�E�B �E(�A0�A8�DP 
8A0A(B BBBB
8F0A(B BBBA  H    a  ����   B�B�B �B(�A0�C8�D�j
8C0A(B BBBJ    la  ����G    A�x
GF    �a  ����/    A�b
EF (   �a  ����^    B�F�A �QAB  $   �a  ����m    Y�A�G IAA@    b  <���j    B�F�A �O
ABEy
ABDAFB   l   Db  h���   O�B�B �B(�A0�A8�D`
8A0A(B BBBII
8A0A(B BBBE�������  L   �b  ���E   B�G�B �B(�A0�A8�D��
8A0A(B BBBB   4   c  ���Y    B�I�D �Q
ABEbGB   X   <c  @����    B�E�D �D(�F0@
(C ABBCm
(H ABBFL(L ABBL   �c  �����   B�B�E �B(�I0�D8�Q��
8D0A(B BBBC   p   �c  T���?&   B�B�E �E(�A0�A8�J��
8D0A(B BBBF��L�u�B���F�]�B�      \d   ���I    X�iG�    xd  T���          �d  P���          �d  L���x          �d  ����          �d  ����          �d  ����O          �d  ����          e  ����.          e  ���          ,e  ���
       $   @e  ���M    A�A�D BCAL   he  4���    B�B�B �B(�A0�D8�G��
8A0A(B BBBI   `   �e  �����   B�H�B �B(�A0�A8�G�_�A�G�A�R��
8D0A(B BBBF <   f  P����   K�B�A �A(�G0�(A ABBF����  @   \f   ����   B�B�B �A(�A0�D`c
0A(A BBBI8   �f  L���
   B�B�D �A(�D@V
(A ABBG    �f   ���
          �f  ���<    A�r
EC    g  <���4    A�r      ,g  `���Y    A�G OA   Lg  ����9    K�fG� H   hg  �����   B�B�B �E(�A0�A8�J�
8D0A(B BBBE    �g  h��V          �g  ���          �g  ���h          �g  ���          h  ���5       @   h  ���#   B�B�B �D(�A0�D@w
0A(A BBBB  8   \h  ����    B�D�A �A(�D@S
(A ABBK  `   �h  d���   B�B�F �B(�A0�A8�D`
8A0A(B BBBGI
8A0A(B BBBE$   �h  �
���    A�A�G tAA   $i  ��[    DVL   <i  P���   B�B�I �D(�G@;
(A ABBGL
(F ABBI  <   �i  ���u    B�C�A �D0S
 AABGH AAB L   �i  ���    B�E�D �D(�F@�
(A ABBIN
(A ABBD      j  ���
       <   0j  ����    B�B�E �D(�A0�i
(C BBBH       pj  ���    T�R
JhH�  4   �j  ���t    A�D�G k
CAEY
CAC  ,   �j  ����    K�D�G B
AAF`��H   �j  @���   B�E�I �H(�A0�A8�G�X
8D0A(B BBBJ L   Hk  ���'   B�B�B �B(�A0�C8�D��
8D0A(B BBBA   <   �k  d'���   K�B�A �A(�G0}(A ABBG����  H   �k  �(��J   B�B�B �B(�D0�D8�I�M
8A0A(B BBBH    $l  �5��          8l  �5��O          Ll  6��          `l  6��          tl  6��          �l  6��       (   �l  6��t    B�D�A �iAB  (   �l  d6��t    B�D�A �iAB     �l  �6��           m  �6��Q    V�J ZAE�   $   ,m  �6��6    A�A�G0hCA (   Tm  7���   J�A�G �AAH��   �m  �8��/    A�`
GF d   �m  �8���    P�E�M �E(�A0�A8�F@J
8A0A(B BBBED8C0A(B BBBA������ d   n  9��   B�B�B �B(�A0�G8�G��
8A0A(B BBBA7
8A0A(B BBBA <   pn  �=��0   B�C�I �JP
 AABCK AAB   �n  �>��
          �n  �>��%    D`    �n  �>��       H   �n  �>��
   B�B�E �B(�A0�A8�Dp
8A0A(B BBBD�   <o  �C���   B�B�E �B(�A0�D8�Dpd
8A0A(B BBBFt
8A0A(B BBBJ|
8A0A(B BBBJH
8A0A(B BBBF   H   �o  �G���   B�D�E �B(�D0�D8�D@�8A0A(B BBB       p  J��6    A�t   L   <p  @J��   B�B�B �B(�A0�A8�J�)
8D0A(B BBBF      �p  W��           �p  W��          �p  W��/          �p  4W��       $   �p  @W��L    A�C�G |CA X   q  hW��q   B�B�B �A(�A0�D@m
0A(A BBBGL
0F(A BBBG  (   `q  �Y��l    B�A�A �dAB     �q  �Y��
          �q  �Y���       <   �q  XZ���    A�D�G S
AAGn
KANMFAL   �q  �Z��k   B�G�E �B(�A0�C8�M�C
8A0A(B BBBB   ,   Dr  f��A    F�A�G kAAE��         tr  (f��          �r  $f��	          �r   f��c       ,   �r  |f���    f�A�A ��AEA���     �r  g��          �r  g��          s  g��          s  g��          0s  g��       $   Ds  g��N    A�A�G @CAL   ls  0g���    A�A�D f
AABD
FAEB
CAJYFA   `   �s  �g��-   B�B�B �A(�A0�
(A BBBFA
(F BBBCq
(F BBBC  (    t  �j���    J�M o
AIGAA�    Lt  0k��
       H   `t  ,k���   B�B�A �A(�G0d
(A ABBIW(A ABB    �t  �l��       P   �t  �l��h    F�E�E �D(�D0�e
(C BBBJH(A GBBA�����      u  �l��U    A�
HL (   4u  �l���    A�G b
AEXA   0   `u  Lm���   B�D�D �G@i
 AABB  H   �u  �n��?   B�B�B �B(�D0�D8�J�g
8D0A(B BBBB p   �u  ���E   B�B�E �G(�D0�GP�
0A(A BBBJe
0A(A BBBCh
0F(A BBBK         Tv  ȅ���          hv  �����          |v  @���          �v  L���          �v  H���           �v  T���          �v  `���{       $   �v  ̇���    A�y
fU
KF     w  t���       $   w  ����G    A�A�G yCA H   Dw  �����   B�G�B �B(�A0�A8�D@.
8A0A(B BBBE(   �w  �����    A�C�D0g
AAG    �w  `���6    A�t   4   �w  �����    B�J�A �D(�K@e(A ABB   x  ܊��
          $x  ؊��y          8x  D���g          Lx  �����       8   `x  ,���@   B�B�A �A(�G0,(A ABB   (   �x  0����    J�A�G �AAD�� d   �x  ���G   B�B�E �B(�D0�D8�D`�
8A0A(B BBBB	
8C0A(B BBBA     0y  ̑��4    A�f
IC 0   Py  ����    q�h
GQ
AF
HP
HPH� d   �y  x���   B�B�B �B(�D0�D8�G`[
8A0A(B BBBD�
8A0A(B BBBJ   H   �y   ����   B�B�E �B(�A0�A8�J�r
8A0A(B BBBE    8z  �����          Lz  0���I       H   `z  l���$   B�B�J �E(�I0�G8�G��
8C0A(B BBBBH   �z  P����   B�H�B �E(�D0�C8�G�~
8C0A(B BBBGH   �z  ����I   B�E�J �B(�A0�D8�O`�
8D0A(B BBBG   D{  �����          X{  $���"          l{  @���          �{  L����          �{  ����          �{  ����          �{  ����          �{  ����3          �{  (���$          �{  D���`          |  �����           |  ���]         4|  h���$          H|  ����(       H   \|  ����'   X�I�D �A(��
 AHBJA
 FBBAM���� l   �|  ����W   B�E�B �B(�A0�A8��
0E(B BBBHF
0A(F BBBEO
0E(B BBBDX   }  t����   B�E�B �B(�A0�A8��
0A(B BBBEA
0C(B BBBD L   t}  ����P   B�B�B �B(�A0�A8�D�p
8C0A(B BBBF      �}  ����:    Dd
HI      �}  ���$          �}  4���I          ~  p����           ~  ,���$          4~  H���e       D   H~  �����    q�F�A �I(�{
 ADBEV ADBK����     �~  \���          �~  h���3          �~  �����          �~  0���          �~  <���       L   �~  H���	   T�J�A �A(�� AFBE����H(����G AFB  4   D  ���!   B�D�A �A(��
 ABBK      |   ���    DT    �  ���          �  ���          �   ����       4   �  ����	   B�D�A �A(��
 ABBK      �  t���    DT     �  |���          4�  ����!          H�  ����          \�  ����	          p�  ����          ��  �����          ��  D����          ��  �����       X   ��  l����    B�B�F �C(�D0j
(C ABBE`
(A ABBBD(J ABB 4   �  ����x    B�A�E �q
CBBQ
ADJ   T�  ����6          h�  ���          |�  ���          ��  ���       D   ��  ���i   B�B�A �H(�s
 FBGAJ
 CBBG      �  @����       X    �  ����   B�I�B �B(�A0�H8�1
0D(B BBBK�0A(E BBB      \�  �����       p   p�  <���-   [�B�B �B(�A0�A8��
0A(B BBBFA
0F(B BBBI�������H8������ X   �  �����   B�B�B �B(�A0�A8��
0A(B BBBDy
0F(B BBBA    @�  ,���
       H   T�  (���E   B�E�B �B(�A0�I8�G`8D0A(B BBB      ��  ,���/    A�m      ��  @���V       H   Ѓ  ����   B�B�B �E(�D0�D8�Dp�
8D0A(B BBBA @   �  `���t    B�I�D �G@R
 AABDe
 FABB   8   `�  ����u    B�E�A �D(�D@G
(C ABBA H   ��  �����   B�H�B �E(�D0�A8�Np�
8A0A(B BBBK 4   �  D����    A�I�I0y
AABD
CAH @    �  �����    B�I�F �D0�
 AABHD
 CABF  (   d�  X���X    A�A�D0U
AAC  L   ��  �����    B�B�D �A(�D0�
(A ABBAD
(C ABBA   8   ��  ����    B�D�D �a
ABBA
CBJ   �   �  p���P   B�J�B �B(�A0�A8�D@�
8J0A(B BBBFD
8C0A(B BBBHJ
8D0A(B BBBI�
8A0A(B BBBA   H   ��  (���   B�E�H �B(�D0�A8�DP�
8D0A(B BBBF 8    �  �����    B�G�A �h
ABKA
CBJ   T   <�  P���B   B�G�B �A(�D0�G@[
0A(A BBBFR
0F(A BBBAH   ��  H����   B�B�B �B(�A0�D8�D`R
8A0A(B BBBC0   ��  ����G    A�A�D g
GAKDAA 0   �  ����G    A�A�D g
GAKDAA 8   H�  ����   B�B�A �A(�G0v
(A ABBG  4   ��  ����
   B�B�D �A(�D0�(A ABB4   ��  p����   K�A�A �R
ABF����      �  8���)    A�g      �  L���1    Z�TB�    ,�  p���(    A�f   `   H�  �����   B�B�B �B(�A0�A8�D`x
8A0A(B BBBH,8F0A(B BBB  H   ��   ���=   B�E�B �B(�A0�I8�Gpg
8A0A(B BBBC    ��  �����       x   �  ����(   T�B�E �E(�D0�D8�F�d
8A0A(B BBBDD8F0A(B BBBE������F�������   H   ��  D��K   B�K�B �B(�A0�A8�DP%
8A0A(B BBBAL   Ԋ  H��-   B�E�B �B(�A0�A8�G��
8A0A(B BBBA   H   $�  (��)   B�B�B �B(�A0�D8�G@�
8D0A(B BBBG    p�  ��
       H   ��  ���   B�E�B �B(�A0�I8�G`�
8A0A(B BBBB 0   Ћ  ���J    A�I�L N
AAJDPA H   �  ���Z   B�E�E �B(�A0�A8�G`g
8A0A(B BBBH  0   P�  ���J    A�I�L N
AAJDPA 8   ��  ���    B�G�I �A(�G0P
(C ABBF  (   ��  ���t    A�F�G H
AAH     �  ��   G��
GL
D L   �  ���g   B�E�B �B(�A0�D8�G�
8A0A(B BBBB   H   `�  &��v   B�F�E �E(�A0�A8�D`�
8C0A(B BBBAL   ��  P(��	   B�I�E �B(�A0�A8�D��
8A0A(B BBBF   <   ��  .���    B�B�B �D(�D0��
(C BBBD   H   <�  �.���   B�I�B �E(�A0�A8�GP�
8C0A(B BBBD<   ��  1���    B�B�E �D(�A0�^
(C BBBK   H   Ȏ  �1��j   B�B�E �B(�E0�D8�D`,
8C0A(B BBBHH   �  �2��2   B�E�B �F(�A0�D8�DP�
8C0A(B BBBF L   `�  �3��   B�F�B �B(�A0�A8�G�w
8C0A(B BBBH      ��  �7��V           ď  �7��U    y�D�VA       �  8��?    a�D�XA       �  08��?    a�D�XA   0   0�  L8��\    A�N�L N
AAEiAA H   d�  x8��n   B�G�B �B(�A0�A8�G�`
8D0A(B BBBE p   ��  �=��Q   B�B�A �A(�D0K
(C ABBCa
(C ABBGw
(C ABBA\
(F ABBI     $�  �>��&       8   8�  �>���    B�B�A �A(�D@c
(C ABBK    t�  �>��?    D n
FF   L   ��  ?��r    B�A�A �D0p
 DABAS
 DABFD JAB   H   �  H?���   B�B�B �H(�A0�A8�G�l
8A0A(B BBBC 0   0�  �B��B    A�I�J N
AADDPA    d�  �B��          x�  �B��       L   ��  �B���    B�G�I �A(�G0P
(C ABBF�
(L ABBI   L   ܒ  �C��K   B�E�B �E(�A0�A8�G��
8A0A(B BBBJ   ,   ,�  �T���    B�H�D �w
CBF   L   \�   U��   B�B�B �B(�A0�A8�D��
8C0A(B BBBK   H   ��  �X��   B�E�B �B(�D0�D8�G`�
8D0A(B BBBA H   ��  �Y��1   B�E�B �E(�A0�D8�G`�
8D0A(B BBBA L   D�  �Z��G
   B�B�B �B(�A0�A8�D�P
8D0A(B BBBE     D   ��  �d���   B�B�B �B(�A0�A8�x
0A(B BBBE     ܔ  0f��       @   �  <f���   D�I�B �I(�E0�A8�v0A(B BBB    4�  �g���          H�  4h��w          \�  �h��3          p�  �h��          ��  �h��          ��  �h��       @   ��  �h���   D�I�B �E(�D0�A8��0A(B BBB    �  <j���          �  �j��H          �  4k��       L   ,�  0k���   B�B�B �B(�A0�A8�G��
8A0A(B BBBA   L   |�  �l��m   B�B�E �B(�A0�A8�G�|
8A0A(B BBBA   L   ̖  �t���	   B�J�B �B(�A0�A8�G��
8A0A(B BBBJ   H   �  p~��x   B�B�E �E(�D0�C8�F`
8A0A(B BBBIH   h�  �����   D�I�B �B(�A0�D8�D`Y
8A0A(B BBBCH   ��  ����   B�B�B �B(�A0�A8�D@�
8A0A(B BBBE$    �  ����X    A�F�G xLA    (�  ���       L   <�  ����5   B�G�B �B(�A0�A8�D��
8A0A(B BBBG   H   ��  Љ��U   B�B�B �E(�A0�A8�D@<
8A0A(B BBBA$   ؘ  ���<    A�F�G \LA (    �  ����"   A�A�D AA   ,   ,�   ���}    G�A�D �b�G�B�      \�  P���
       ,   p�  L����   K�F
O��H�F
Z   d   ��  ���\   B�E�E �E(�A0�A8�I@}
8A0A(B BBBE[
8A0A(B BBBC      �  ���Q       (   �  0���   e�C��FN��H��$   H�  ���I    A�L�[ WHA 0   p�  <���K    A�D�M0M
AAG`AA L   ��  X����   B�G�B �B(�D0�D8�D�
8A0A(B BBBG   H   ��  ؝��   B�B�B �B(�D0�A8�GP�
8A0A(B BBBF H   @�  ����P   B�B�B �B(�A0�A8�Dp�
8A0A(B BBBA H   ��  �����   B�E�B �B(�D0�A8�D`Z
8A0A(B BBBHH   ؛  $���?   B�B�B �B(�D0�D8�Dpw
8A0A(B BBBK  L   $�  ���p   B�B�B �B(�A0�A8�G�h�
8D0A(B BBBB   ,   t�  8���f    F�D�G0[
AABp�� 4   ��  x����   A�W �
AJe
AJJ
AE   X   ܜ   ���4   B�E�B �K(�I0�D`x
0C(A BBBES
0C(A BBBK   \   8�  ����   B�B�B �B(�A0�A8�L�j�D�F�A��
8A0A(B BBBK  L   ��  d����   B�H�E �B(�A0�A8�G�{
8A0A(B BBBA      �  ����       \   ��  ����=   B�H�B �B(�A0�A8�L��b�X�A�
8A0A(B BBBE    \�  ����          p�  ����          ��  ����       8   ��  �����   B�D�D ��
IBJ�
IBD  D   Ԟ  ���    B�I�B �D(�A0�J���
0A(A BBBA  L   �  �����   B�B�B �B(�A0�A8�G��
8A0A(B BBBI   T   l�  P����    L�E�E �A(�D0�D`�
0A(A BBBAI0A(A BBB   (   ğ  ����`    B�A�D �q
CBC(   �  ���e    B�A�D �|
CBHD   �  P���    B�I�B �D(�A0�J���
0A(A BBBA  L   d�  (����   B�B�B �B(�A0�A8�G��
8A0A(B BBBG   H   ��  ����O   B�B�B �B(�D0�D8�G�v
8D0A(B BBBF (    �  ����:    A�A�G kDA     (   ,�  �����    f�A�QAG��H��   X�  4����       D   l�  �����   B�E�B �B(�A0�D8�
0A(B BBBF     ��  x���          ȡ  t���          ܡ  p���          �  l���9          �  ����9          �  �����       $   ,�  ����m    A�D�G ^AA4   T�  �����    B�E�A �D(�D0u(A ABB$   ��  @���C   @�F��AA��  \   ��  h����   P�I�G �E(�A0�A8��
0A(B BBBEP������H8������ `   �  ����#   B�G�H �E(�G0�H8�J`Z
8A0A(B BBBE�
8A0A(B BBBJ8   x�  d����    B�E�A �A(�G@t
(A ABBF  @   ��  �����    O�A�C �G0R
 AABH] AABG��� <   ��  $���t    B�D�D �D0]
 AABA AAB  (   8�  d���Q    B�A�D �`
ABF`   d�  �����   B�H�E �E(�D0�C8�Dpu
8A0A(B BBBBY
8A0A(B BBBEH   Ȥ  �����    B�G�D �D(�G0M
(A ABBEI(A ABB  ,   �  ���V    B�D�D �G0@ AABH   D�  8����    B�B�B �B(�A0�A8�G��8A0A(B BBB      ��  ����Q       T   ��  ����   Q�E�E �B(�E0�J8�Ip�
8A0A(B BBBE�������  8   ��  P���u    R�A�A �L
�A�B�MAAB   D   8�  ����f   B�B�B �B(�A0�C8��
0A(B BBBH   <   ��  �����   B�E�E �A(�A0��
(A BBBK  T   ��  \ ���   B�B�B �E(�A0�I8�G`�h]pUhE`/8A0A(B BBB |   �  ���z   M�E�B �B(�D0�A8�GpM
8A0A(B BBBG�������Hp������o
8A0A(B BBBG  H   ��  ���   B�J�B �B(�A0�A8�G��
8A0A(B BBBC   �  X��       \   ��  d��   M�B�B �B(�A0�A8�Gp�8A0A(B BBBJ������Hp������ $   X�  $���    A�A�K �AAt   ��  ���4   B�B�E �E(�D0�D8�FPs
8A0A(B BBBG�
8A0A(B BBBGa8A0A(B BBBX   ��  t ���    I�B�B �A(�A0�Q(A BBBI�����H0�����D(A BBB\   T�  � ���    I�B�B �A(�A0�Q(A BBBI�����H0�����E(A BBB       ��  � ���          ȩ  �!���          ܩ  @"���          �  #��d          �  h#���       d   �  $��   B�E�B �E(�E0�A8�G`,
8A0A(B BBBG�
8A0A(B BBBJ   (   ��  �%��[    B�D�D �MAB  H   ��  �%���   B�E�H �D(�G00
(A ABBH~(F ABBH   ��  �'��   B�B�D �H(�G0}
(A ABBFf(F ABB   D�  X)���          X�  �)��%          l�  *��	      4   ��  +���   B�B�A �A(�U
 ABBH      ��  �,��          ̫  �,��          �  �,��p       <   ��  �,���   F�B�E �H(�C0�V
(A BBBK      4�  �.��          H�  �.��          \�  �.��          p�  �.��!    GY    ��  �.��          ��  �.��       d   ��  �.���   B�E�E �B(�A0�A8�Dp�
8C0A(B BBBH�
8F0A(B BBBD   d   �  �0��   B�B�D �D(�G0m8c@F8A0h
(A ABBHt
(F ABBAP8C@W8A0   �   ��  �2��l   B�B�E �B(�A0�A8�D���E�G�B��
8C0A(B BBBDy
8A0A(B BBBE�
8F0A(B BBBEc�K�L�A�   $   $�  x?��:   ���l��I
G $   L�  �B��9    A�D�G0hCA    t�  �B��?       H   ��  �B��%   B�B�I �B(�A0�A8�J�O
8A0A(B BBBD,   Ԯ  �D��S    B�G�A �EAB         �  �D��          �  �D��          ,�  �D��g    Db   D�  8E��          X�  DE��          l�  @E��C   q�gH�   ��  tF���       (   ��  �F���    A�D Q
CG]C   L   ̯  PG���   B�B�B �B(�A0�A8�GЁ�
8A0A(B BBBA      �  �I���   |��V��  (   @�  �K��    A�G }
AJO
AH L   l�  �K���   B�B�E �B(�D0�A8�D��
8A0A(B BBBG      ��  `O��)    Dd (   ԰  xO��G    B�D�A �|AB   $    �  �O��9    A�D�G0hCA    (�  �O��?       H   <�  �O��j   B�B�I �B(�A0�D8�J�H
8A0A(B BBBH   ��  W��          ��  W��          ��  W��       @   ı  W���   B�J�J �I(�A0�G�t0A(A BBB     �  tY��*    DC b  @   $�  �Y���   B�U�D �K�t
 AABBt AAB      h�  $[��$    D_ (   ��  <[��S    B�G�A �EAB  L   ��  p[���   B�E�B �B(�A0�A8�G��
8A0A(B BBBB   $   ��  �`���    A�D�G qAA   $�  Ha��R    Ry (   <�  �a��~    X�A�G PCAD�� X   h�  �a��2   B�J�E �B(�A0�A8��
0A(B FBEGK0F(B BBB   4   ĳ  �c���    B�A�D �~
ABHMIB     ��  @d��          �  <d��          $�  8d��    H R    <�  @d��    H R (   T�  Hd��.   A�C�G0Q
AAB  H   ��  Le��A   B�B�B �B(�A0�D8�GP}
8A0A(B BBBE P   ̴  Pf���   K�B�B �A(�C0�
(A BBBD������F0������    �  �g��b   X�B�B �B(�A0�A8�D�

8A0A(B BBBHT
8F0A(B BBBE�
8A0A(B BBBHH�F�B�D�P���R�F�F�N�}������F���������Q�I�F�W�  L   ��  p����   B�M�H �A(�G0�
(A ABBKP
(C ABBH  `   L�  �����   B�B�E �D(�D0�e
(A BBBCo
(D BBBG[
(A EBBK      ��  ���	       \   Ķ  ���   T�B�B �B(�A0�D8�JPQ8A0A(B BBBD������HP������ T   $�  Ȇ���    `�A�G�s
DAHI
AAED
FAEX��P���       0   |�  p���c    A�I M
AHa
FIQA   (   ��  �����   A�A�G 
AAF0   ܷ  ����    R�D�S0]AAH��H0��     �  ����*          $�  ȉ���       P   8�  T���4   T�B�B �A(�D0�JP�0A(A BBBD�����HP����� $   ��  @����    A�H�G �AA(   ��  ����L    B�A�A �DAB  H   �  ܋���   B�B�B �B(�A0�C8�G`C
8D0A(B BBBE L   ,�  ����,   B�B�B �E(�D0�D8�D@�
8D0A(B BBBC        |�  p���)       D   ��  ����f   Z�B�A �A(�B����H(����\
 DBBD <   ع  ����p    B�I�A �D0i
 AABCi CAB     �  ���c          ,�  @����          @�  ���c    D^,   X�  t���$   A�G �
ACn
AA   4   ��  t���/   A�D�D(
AADP
AAF   ��  l���	       8   Ժ  h����   B�B�A �D(�G8�
(A ABBF `   �  �����    B�B�E �B(�D0�D8�Fp[
8A0A(B BBBB�
8A0A(B BBBA    t�  ����       L   ��  ����s   B�E�B �A(�D0�F
(C BBBC�
(F BBBB   ػ  Ԛ���          �  P���           �  L���D          �  �����          (�  T���D          <�  ����H          P�  ̜���          d�  ����D          x�  ԝ��P          ��  ���          ��  ���           ��  (���1          ȼ  T���1          ܼ  ����%          �  ����          �  ����          �  ����d          ,�  ���          @�  ���6          T�  8���          h�  4���          |�  0����         ��  ���      L   ��  ����   B�E�A �A(�D0�
(A ABBA�
(A ABBA 4   ��  Ȥ���   D��
Hi
GO
Ah
H{
E  $   ,�  `���f    Q�A�G JAA$   T�  �����    A�A�D |AA   |�  ���    A�X      ��  ���(    A�f   <   ��  (����    B�A�A �D0o
 AABE^ AAB 4   ��  ����g    B�E�D �I(�J@B(A ABBL   ,�  Ч���    B�E�I �G(�G@z
(A ABBBu
(A ABBE   <   |�  p����    L�C�A �G0o
 AABF` CAB (   ��  ���Y    A�D�G g
AAK  H   �  $����    B�B�B �A(�A0�Z
(A BBBGO(A BBBH   4�  h���   B�B�B �B(�A0�A8�Dph
8D0A(B BBBEH   ��  ,���]   B�B�B �B(�A0�A8�Dp�
8D0A(B BBBH    ��  @���)    D` H   ��  X���e   B�B�B �E(�A0�A8�J��
8A0A(B BBBJH   0�  |���_   B�E�B �B(�D0�D8�J��
8A0A(B BBBDH   |�  ����E   B�E�E �B(�D0�A8�D`�
8D0A(B BBBD    ��  ����     DW    ��  �����       0   ��  x����    B�A�D �G0_
 AABG     (�  4����   A��
Ge
[    L�  �����      (   `�  ����   A�C��
AK�A(   ��  ����    A�L
CG
IQ
GF   ��  ���x    A�G
Hg8   ��  t���$   B�B�A �A(�G0(A ABB   8   �  h���8   B�G�A �A(�G0(A ABB   L   P�  l����    U�E�A �A(�G0\
(C ABBID(F ABBA���� \   ��  ̿��   B�D�E �E(�D0�D8�NP�
8A0A(B BBBCD8F0A(B BBB8    �  �����    B�I�E �D(�A0�e(D BBB     <�  ����c          P�  <���x          d�  ����h       H   x�  ���{   B�B�E �E(�A0�C8�H`d
8C0A(B BBBF    ��  8����          ��  ���    A�R   ,   ��  ���	   B�A�D ��
ABG       $�  �����    D�T��E  l   H�  �����
   B�B�E �B(�A0�D8�J��L�}�B�y
8A0A(B BBBCo�L�I�A�   ��  ����          ��  ����          ��  ����2          ��  (���5          �  T���`          �  ����`          0�  ����>       (   D�  ���Q    F�A�G uAAK��  x   p�  L����   B�B�B �B(�D0�A8�Dpi
8A0A(B BBBD\
8F0A(B BBBEH8A0A(B BBB   H   ��  �����    B�H�E �B(�D0�A8�D`�
8A0A(B BBBC d   8�  4����   B�I�B �E(�H0�A8�G��
8A0A(B BBBB�
8A0A(B BBBH      ��  \���j    A�G E
AB    ��  ����i    A�|
C,   ��  �����    B�D�C ��
ABA   0   �  l����    B�D�D �Gpw
 AABD P   D�  �����   B�B�E �E(�D0�D8�D`AhE`a
8A0A(B BBBE \   ��  D���F   B�E�E �E(�F0�G8�G�R�U���B��
8A0A(B BBBF   T   ��  4����   B�B�B �B(�D0�D8�G���E�Y8A0A(B BBBD�     P�  ����'          d�  ����       <   x�  ����T    B�D�I �G0M
 AABI_ AAB  4   ��  ���J    R�D�D �W
ABDJ�A�B�   ��  ,���'          �  H���<       H   �  t����    B�B�A �A(�D@�
(A ABBJt(F ABB  8   d�  ���F   B�D�D �[
ABH�
ABA     ��  ���'          ��  8���       (   ��  D���d    B�D�I �QAB  4   ��  ����J    R�D�D �T
ABGJ�A�B�H   ,�  �����   B�E�B �B(�D0�A8�D`c
8A0A(B BBBG  H   x�  ���}    B�D�B �A(�A0�R
(C BBBKC(C BBB   ��  H���       4   ��  T���U    B�D�A �w
ABGIAB      �  |���b       L   $�  ����h   B�B�B �B(�A0�A8�G�
8D0A(B BBBD   (   t�  �����    B�J�K ��AB     ��  �����       H   ��  ���x    B�B�D �D(�D0H
(A ABBBD(J ABB      �  L���X       p  �  ����c/   B�B�E �B(�A0�A8�Q��_
8A0A(B BBBI��H��k��A�����R��_��B��	��Q��^��B����H��e��B����G��f��B��Y
��G��g���J��_��A��m��Q��a��A��\	��H��]��A��M��N��z��A��u
��A��Z���H��E��B�����B��J��B��y��Q��O��E��  �   ��  ���Z   B�E�B �E(�A0�D8�G�V�L�F�A�g�P�J�B���H�\�A�n
8A0A(B BBBF�L�I�A�    �  `(��7          0�  �(���           D�  )���    A��
VP
A    h�  �)��          |�  �)��#          ��  �)��
           ��  �)���   A��
AL
L   ��  $+��      L   ��  0,���   B�E�B �E(�F0�A8�J��
8A0A(B BBBE      ,�  �.��&    A�d   4   H�  �.��V    M�A�D �W
�F�B�OP���      ��  �.��          ��  �.��          ��  �.��       4   ��  �.���    J�A�J �
AAALFAE��    ��  X/��7    Dr    �  �/��              $�  x/��          8�  t/��          L�  p/��          `�  l/��          t�  h/��              ��  `/��-          ��  |/��       �   ��  x/��   B�B�B �B(�A0�A8�DP 
8A0A(B BBBHv
8A0A(B BBBHl
8F0A(B BBBED
8F0A(B BBBEl   H�  1���   B�B�B �A(�A0�D@�
0A(A BBBH�
0F(A BBBGD
0F(A BBBG   ��  �5���    f�N@�A   ��  46��V    K�yD� |   ��  x6��f   I�G�E �B(�A0�A8�K�}������G��������
8A0A(B BBBA�������L�������L   t�  h<���   B�B�B �B(�A0�A8�G�[
8A0A(B BBBJ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �"@     ��������        ��������                             p	@            �F             `i                          h@            p@            @@     
                                                  xai                                        p@                                                                                                     (`i                     �	@     �	@     �	@     �	@     �	@     �	@     �	@     
@     
@     &
@     6
@     F
@     V
@     f
@     v
@     �
@     �
@     �
@     �
@     �
@     �
@     �
@     �
@     @     @     &@     6@     F@     V@     f@     v@     �@                                                        �                                                           �   �                                                       �����   �                                                   ���������   �                                               �������������   �                                           �����������������   �                                       ���������������������   �                                   �������������������������   �                               �����������������������������   �                           ���������������������������������   �                       �������������������������������������   �                   �����������������������������������������   �               ���������������������������������������������   �           �������������������������������������������������   �       �����������������������������!!!�!!!�!!!�!!!�!!!�!!!�   �   �����������������!!!���������   �   �   �   �   �   �   �   �������������!!!�   �!!!�����   �                           ���������!!!�   �       �BBB�����   �                       �����!!!�   �           �!!!�����   �                       �!!!�   �                   �BBB�����   �                   �   �                       �!!!�����   �                   �                               �BBB�����   �                                               �!!!�����   �                                                   �   �                                      �bi                                            1   2   3   4   5   6   7   8   9   0   -   =      	   q   w   e   r   t   y   u   i   o   p   [   ]   
       a   s   d   f   g   h   j   k   l   ;   '   `       \   z   x   c   v   b   n   m   ,   .   /       *                                  	              
      -           +                                                                                                                                                                                                     d   d   @��                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `  GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o �             �@     �      �"@     I       #@     2       8#@     -       f#@            x#@     "       �#@     -      �$@     "       �$@     �       �%@     �       @&@     -                       ,     7       m&@     9                       ,    8       �&@     5                      ,    c;       �'@     u                       ,    =       P(@     �                       ,    �E       )@     E                      ,    wX       [6@     �                      ,    ws       �B@     �                           �s                       ,    at       �C@     �                      ,    ��       pF@     Ѹ                      ,    V      P�@     &                      ,    R�      ��A     �`                      ,    �w      ``B     o                      ,     �      p�B     �%                      ,    J4      �B     �5                      ,    �      �*C     �%                      ,    >H      �PC     �                      ,    }�      �aC     u#                      ,    ��      �C     �@                      ,    tY      ��C     W�                      ,    L�	      @�D     ��                      ,    "�
      �E     �=                      ,    �0      �SE     S)                      ,    �      �|E     #                      ,    �      �E     �0                      ,    B      ��E     �                      ,    �      ��E     ��                      ,    ��      p�F     H                      ,    R�      ��F     �                      ,    <�      ��F     A                       ,    �      ��F     �                                      7       �  S  �                  N  5   �  �  H   �  �  [   �  �
  n   �  V  	�   �  ;  �  �   int �   ,  C  �n   �  u   �  �   �  )   �  <   �  O   L  b   ;
  4�   �  P  5�  �    ��  �   bpp 	�   `�  �   
 K    i   �n   	std    
�  AAs  	�  	��  	�-  	�J  	�`  	��  	��  	��  	�  	�!  	�=  	�X  	�s  	��  	��  	��  	��  	�  	�  	�7  	�W  	�w  	��  	��  	�!  	�l  	��  	��  	�F  	��  	�  	�h  abs 
f/   �  �  �   abs 
TQ   �  �  �   abs 
N   �  �  �   abs 
J%   a  �  a   abs 
F   v    v   abs 
=~     !     abs 
89   �   ;  �    div 	��  �  Z  �   �    )�  *�  C  [  �  �  �   C  W  a  �  a   �  n�  �  �  �   �  j�  a  �  a   A  ��  �  �  �   A  }�  a    a     ��  �  '  �  �     �%  a  F  a  a   cos ��  �  `  �   cos ��  a  z  a   sin ��  �  �  �   sin ��  a  �  a   tan ��  �  �  �   tan ��  a  �  a     �   �     �     �  a    a   W
  ��  �  5  �   W
  ��  a  P  a   �  ��  �  k  �   �  ��  a  �  a   exp �  �  �  �   exp �  a  �  a     0A	  �  �  �  0     ,�  a  �  a  0   �  C@  �    �  �    �  ?!  a  :  a  �    log Vf  �  U  �   log Rp  a  p  a   0  i�   �  �  �   0  e�   a  �  a   _  |�  �  �  �     _  x�	  a  �  a     pow �y  �    �  �   pow �   a  &  a  a   �   �c  �  A  �   �   �n  a  \  a   M  �'  �  v  �   M  �2  a  �  a   o	  ��  �  �  �   o	  ��  a  �  a   �  �  �  �  �   �  �  a  �  a   "     �    �  �   "  �   a  :  a  a   v  #  �   U  �   v  �  �   p  v   v  !  �   �  a   d  :�  [  �  �   d  6�  [  �  v   d  2�  [  �  a   @  U�  [  �  �   @  P�  [  	  v   @  H�  [  -	  a   �  p�
  [  H	  �   �  k�
  [  c	  v   �  c�
  [  ~	  a     �  [  �	  �     ��  [  �	  v     ~  [  �	  a   U  �\  [  �	  �   U  �[   [  
  v   U  �p   [   
  a     ��	  [  @
  �  �     ��  [  `
  v  v     �E
  [  �
  a  a   �  ��  [  �
  �  �   �  �  [  �
  v  v   �  ��  [  �
  a  a   2  �t  [     �  �   2  ��  [     v  v   2  �  [  @  a  a   �  }  [  `  �  �   �  ��  [  �  v  v   �  �y  [  �  a  a   �  ,  [  �  �  �   �  B  [  �  v  v   �  +	  [     a  a     5  [     �  �     1~  [  @  v  v     -i  [  `  a  a     �!  �  {  �     �-  a  �  a   V
  ��  �  �  �   V
  ��  a  �  a   �  ��  �  �  �   �  ��  a    a   W  ��	  �    �   W  ��	  a  8  a   �  
{  �  X  �  �   �  d  a  x  a  a   erf U  �  �  �   erf 8  a  �  a   6
  0�  �  �  �   6
  ,�  a  �  a   �  B  �  �  �   �  >  a    a   H  Tt  �  5  �   H  P�  a  P  a       f]  �  p  �  �       bF  a  �  a  a   fma z�  �  �  �  �  �   fma v�  a  �  a  a  a   �  �c  �  �  �  �   �  �  a    a  a   �   ��  �  :  �  �   �   ��   a  Z  a  a   �H  �  �  z  �  �   �H  ��	  a  �  a  a   S  ��  �   �  �   S  �m  �   �  a   +  �  �  �  �   +  �  a    a   �  ��    !  �   �  ��    <  a   �  c    W  �   �  �q    r  a   +  �  �  �  �   +  �  a  �  a   �  &F  �  �  �   �  "Q  a  �  a   T  8�  �  �  �   T  4 	  a    a   �  J#  �   /  �   �  F/  �   J  a   �  \  �   e  �   �  X#  �   �  a   �  n&  �  �  �   �  j6  a  �  a   N  ��   �  �  �  �   N  |�  a  �  a  a   �  ��  �    �  �   �  �q  a  6  a  �   �  ��  �  V  �  �   �  ��  a  v  a  a   d  ��  �  �  �  �  0   d  ��  a  �  a  a  0   �  ��  �  �  �   �  ��  a  �  a   �  �	
  �    �   �  �
  a  ,  a   �  ��  �  L  �  �    �  ��  a  l  a  �    E  �  �  �  �  �    E   C   a  �  a  �    -  \
  �  �  �   -  i
  a  �  a   �  (  �  �  �   �  $  a  a    j  �  
�  AA"  	�!  	��  	��  	��  	�  	�F  	�h  div 	��  !        >  �    �    rem �    ?  �  �	  �    �    rem �    �	  �  3         rem    '  4  �  m  I�   C  C   I  �  J�   `  C   �  'v  v  }   �  �  �  �  �  (�   �  }   E@ )�   �  }   R  V�  �  �  �  \  \  �   �  �  �     �  �   div a�  !  �   �    �	  M7  7  }   �  �   b�  X  �   �    	  g�   s  }  \   �  m\  �  �  }  \   �  �  �  \  h�   �  �  }  \   �  X�  �  \  \  �   �  N#�  �       5�     7  [      +v  1  }  1   7  $  .�   W  }  1  �    �  0n   w  }  1  �    2� O�   �  }   J  n\  �  7  �  \   �    i�   �  7  �   �   c	!  �       j  *  �  }   W  /    }  1  �    �  1?  ?  }  1  �    �    ,a  a  }  1   \   -�  �  }  1   �  '-  +J  .�  3�  4�  abs ]�   �  �    6�  v
  6�  4  6�  6�  6�  6�  6  6!  7`  8�  9�  :�  <l  <  <;  >!  @=  CX  Ds  E�  G�  H�  J  K  L7  MW  Nw  P�  Q�  	  v  �  a  &�  &�  &�  &�  &�  &�  &  &!  C  uv  ,  v   '  'l  '�  �  yv  Z  v   (D  (�  (�  A  }v  �  v   )r  )�  )�    �v  �  v  v   *�  *  *'  cos �v  �  v   +�  +F  +`  sin �v    v   ,  ,z  ,�  tan �v  E  v   -/  -�  -�    �v  s  v   .]  .�  .   W
  �v  �  v   /�  /  /5  �  �v  �  v   0�  0P  0k  exp �v  �  v   1�  1�  1�    �v  0  v  0   �   2  2�  2�  �  �v  i  v  �    3N  3�  3  log �v  �  v   4�  4:  4U  0  �v  �  v   5�  5p  5�  _  �v  �  v  �   v  6�  �  6�  a  6�  pow �v  =  v  v   7"  7�  7  �   �v  k  v   8U  8&  8A  !M  v  �  v   9�  9\  9v  o	  �v  �  v   :�  :�  :�  !�  v  �  v   ;�  ;�  ;�  !"  9v  +  v  v   <  <�  <  ?:  ?U  ?p  ��  @�  @�  @�  A�  A�  A	  B-	  BH	  Bc	  C~	  C�	  C�	  D�	  D�	  D
  E 
  E@
  E`
  F�
  F�
  F�
  G�
  G   G   H@  H`  H�  I�  I�  I�  J   J   J@    �v  �  v   Nj  N`  N{  V
  �v  �  v   O�  O�  O�  �  �v  �  v   P�  P�  P�  W  �v  
   v   Q�  Q  Q  !�  Gv  >   v  v   R"   R8  RX  erf �v  l   v   SV   Sx  S�  !6
  v  �   v   T�   T�  T�  �  �v  �   v   U�   U�  U�  H  �v  �   v   V�   V  V5  !    Yv  +!  v  v   W!  WP  Wp  "fma gv  d!  v  v  v   XC!  X�  X�  !�  ]v  �!  v  v   Y|!  Y�  Y�  !�   av  �!  v  v   Z�!  Z  Z:  �H  �v  �!  v  v   [�!  [Z  [z  S  ��   -"  v   \"  \�  \�  !+  v  \"  v   ]E"  ]�  ]�  !�  #  �"  v   ^t"  ^  ^!  !�  /  �"  v   _�"  _<  _W  +  �v  �"  v   `�"  `r  `�  �  �v  #  v   a #  a�  a�  T  �v  D#  v   b.#  b�  b�  !�  �   s#  v   c\#  c  c/  !�  +�   �#  v   d�#  dJ  de  !�  v  �#  v   e�#  e�  e�  !N  Ov  $  v  v   f�#  f�  f�  !�  Sv  9$  v  �   g$  g�  g  !�  =v  m$  v  v   hQ$  h6  hV  !d  Av  �$  v  v  0   i�$  iv  i�  !�  v  �$  v   j�$  j�  j�  !�  'v  %  v   k�$  k�  k  �  �v  7%  v  �    l%  l,  lL  E  �v  j%  v  �    mO%  ml  m�  !-  	v  �%  v   n�%  n�  n�  !�  3v  �%  v   o�%  o�  o�  1  (R&  x �    y 	�   5�  �   ��  �   `�  �   �V 
�   _| 	R&  '  

�     �   �  �%  3  �&  x 	�    y �    ^  	d&  �&  �  �&  r �    g �   b �   a �    �  �&  (.  |'  6  /�    5�  0
�   ��  1
�   �  2�   bpp 3�   \  4�   ֳ  5�   �  6
�   =  7
�   �
  8�    9  9�   $ 
  :�&  #i  2  �  X&  |�  $(  x �    y �   5�  �   ��  �   �1  �     $(  �  �   l�  �'  t$�  �  (  %q6    &�  4(  'n   _ �  �'  �   @�(  �  7   p   	\  �  #	\  X  &	\  �  )	\   �  ,	\  (�  -	\  0/  2�   8�  5�   < �  8"@(  (+  K�(  �(  (%  L�(  (�  M�(  (]  H)  �  �    �  �   msg �   Kl  �     �     _  �(  (�  �1  (9  �7  (�	  ��   (�  ��   (Z  ��   )�  [   *S  [   �b*  +Y   ,�  bmys,�  cinu,�
  sijs,    bg,�  5gib,F  snaw,  ahoj,�    bg,�  sijs,=    bg,�  5gib,�
  snaw,k  ahoj,�  BODA,t  EBDA,�  CBDA,  1tal,�  2tal,�   nmra &�&  s*  -n   g .  !b*  	�bi     .�  <X&  	`hi     &�   �*  'n    .  D�*  	�hi     8  �l+  �  m�'   �  n4(  pos o�&  �&
  p[  � /fb s
R&  	 ui     .�  tP  	(ui     .�  uX&  	@ui     &�   X+  'n    .�  wH+  	hui     .�  x�&  	�ji     .�  y[  	kui     .a  z[  	lui     .  {�&  	pui     .�  }[  	�ji     .�  �  	xui     .�  ��&  	�ji     .v  �X&  	�ui     .s  ��   	�ui     0�
  �-  1�j  �  V,  \,  %�-   1'    q,  |,  %�-  %�    1O�  !z  �,  �,  %�-   1�	  *o  �,  �,  %�-  .   1<  ;*  �,  �,  %�-  .   2�	  L5  .  �,  �,  %�-  [    2Z  P�  .  -  -  %�-  [    1}  ZP  4-  D-  %�-  [   .   2�  d   �   ]-  c-  %�-   2�  hX  .  |-  �-  %�-  [    2  }B  .  �-  �-  %�-   2=  �R  .  �-  �-  %�-   3@  �_.   3�	  �_.  4num �[   5T .   4,  �-  �*  0B  _.  3�W 	_.   3�� 
_.  4obj .  6�"  �  Q.  W.  %_.   5T .   .  _.  .;  �4,  	�ui     .&
  �.  	�ui     7�  �  8   �"@            �9\,  �.  �.  :!
  �-  :.  �    ;�.  E  �.  @&@     -       �/  <�.  �h =�  i"@     >       �?/  >�
  ��   �l>�	  ��   �h ?�,  ^/  �%@     �       ��/  @!
  �-  �XApos P[   �TB�  S_.  �hC�%@     8       Di U[   �d  E�,  �/  �$@     �       ��/  @!
  �-  �HAobj *.  �@B�K  +_.  �X F?.  0  0  :!
  e.   G�/  �  00  �$@     "       �90  <0  �h Ec-  X0  �#@     -      ��0  @!
  �-  �HApos h[   �DB�  n_.  �hDobj r.  �XH�#@     	       �0  B�S  j.  �P C�#@     8       Di p[   �d  E�,  �0  x#@     "       �1  @!
  �-  �hApos L[   �d ?D-  01  f#@            �=1  @!
  �-  �h 9A,  K1  U1  :!
  �-   G=1  �  x1  8#@     -       ��1  <K1  �h IF  �   @     a      ��3  JM  �'  ��J�  �(  ��J]	  �   ��~J_  R&  ��J�  �3  ��J�	  !�   ��C�@     �      Kmsg �H)  ��~H�@     7       s2  Ki /�   �\C�@            Kwin 0.  ��  Ha@     d      $3  Ki K�   �XC{@     A      Kwin L.  ��Hc@     >       �2  J�  SH)  ��~ C�@     �       Jy  [H)  ��~Jh  ]�   �TJo  ^�   �P   Hh@     �       k3  Jy  yH)  ��~Jh  {�   �LJo  |�   �H H�@     �       �3  Jy  �H)  ��~Jh  ��   �DJo  ��   �@ C� @     �       J  �H)  ��~Kkey ��   ��   |'  L8  �(  �@     J      �14  Awin �.  ��~BF  ��&  �� M�  ��  [  �@     �       ��4  Awin �$.  �HNc �4�&  �@B�  ��   �\ MO	  �2  [  b@     �       ��4  Awin �.  �XNc �.�&  �PB3  ��   �l L�  ��  �@     �      ��5  Br  ��   ��C@     H      Dj �
�   �\C@     )      B1  �[  �[B  �4(  ��~B`  ��'  �HH\@     �       �5  Di ��   �T C\@     �       Dwin �.  �@    L�  �a  �@           �q6  Br  ��   �DC@     �       Di �
�   �\C#@     �       B1  �	[  �[C'@     u       Dj ��   �TC9@     ]       B  �4(  ��~B`  ��'  �H     4(  q6  F(  �6  �6  :!
  w6   G|6  	  �6  #@     2       ��6  <�6  �h O�  t	  �&  �"@     I       �7  Al 07  �hAr E7  �` P�&  !  -
  �   �      9  �  �  m&@     9         N  9   �  �  �  �  �  ;  int ,  C  �N   �  -   ;
  4q   �  
�  �   m&@     9       ��   �  &�   �Pptr �   �` }   	�  �    S   �  9  �  �  �&@     5      �  �  �  �  G   �  �
  Z   �  �  ;  int ,  C  �Z   �  ;   L  N   ;
  4}   i   �Z   '  �  i  n  v   9  �  �  �    }W   b �   � 	    
Z    �    �  �     !#  o   �'@     6       ��  fd !o   �T/� !$�   �H?  !;�  �@ret "�   �` +  �  �  �   q'@     4       �  fd o   �T�   �   �H�  ,o   �Pret �   �` �  t  o   <'@     5       �c  fd o   �T_| %c  �H/� 4�   �@ret 	o   �d i  �  [  o   '@     5       ��  fd o   �T_| �   �H/� -�   �@ret 	o   �d O  �  �&@     .       ��  fd o   �d �    o   �&@     3       �P  F  P  �P�1  *o   �Lfd 	o   �d &   �   �  9  ;  �  �'@     u       �  �  �  �  �
  N   �  �  ;  int ,  C  �N   L  B   ;
  4q   (]  �   �  }    �  }   msg }   Kl  }     }     _  �   $  
�  (@     D       �\  	pid 
}   �@	msg 
.�   � 
m }   �`Kl  }   �X  }   �P   
J  }   �'@     1       ��  	msg (�  �P0  }   �` �    �   �  9  �  �  P(@     �       �  ,  i   �@   �  '  �  i  std    �  AAe   �  ��  �-  �J  �`  ��  ��  ��  �  �!  �=  �X  �s  ��  ��  ��  ��  �  �  �>  �^  �~  ��  ��  �!  �l  ��  ��  �M  �  �&  �o  	abs N   N   �  
N    	abs J%   h  �  
h   	abs F   v  �  
v   	abs =~   G   �  
G    	abs 89   -   �  
-    div ��  �  
-   
-     j  �  �  AA"  �!  ��  ��  �  �&  �M  �o  div ��  !  
G   
G     >  �    �   rem �   int ?  �  �	  �    -    rem -    �	  �  3  !    G    rem G    4  �  m  I�  C  
C   I  �  J�  `  
C   �  'v  v  
}   �  �  �  �  �  (�  �  
}   E@ )-   �  
}   R  V�  �  
�  
�  
4   
4   
�   �  �  �    
�  
�   div a�  !  
�  
�   �	  M7  7  
}   �  �   b�  X  
-   
-    	  g�  s  
}  
4    �  m4   �  
�  
}  
4    �  �  �  \  h�  �  
�  
}  
4    �  X�  
�  
4   
4   
�   �  N#�  
�     5�    7  
   �    +v  8  
}  
8   7  $  .-   ^  
}  
8  
�   �  0@   ~  
}  
8  
�   2� O�  �  
}   J  n4   �  
7  
�  
4    �    i�  �  
7  
�   �   c	!  �  
G   
G    j  *G     
}   W  /G   &  
}  
8  
�   �  1F  F  
}  
8  
�   �    ,h  h  
}  
8   \   -N   �  
}  
8   '-  +J  .�  3�  4�  abs ]�  �  
�   6�  6w  6�  6�  6�  6�  7`  8�  9�  :�  <l  <  <�  >!  @=  CX  Ds  E�  G�  H�  J  K  L>  M^  N~  P�  Q�  s  )�  �(@            ��  p )�  �h@   �` s  #�  �(@            �  p #�  �h �  �  �(@            �@  p �  �h@   �` �  �  �(@            �p  p �  �h �  �  �  y(@     )       ��   ֳ  (@   �h !�  m  �  P(@     )       � ֳ  &@   �h  �   �	  9  �  �  )@     E      �  N  9   �  �  L   �  �  _   �  �
  r   �  �  ;  int ,  �  -   �  @   �  S   L  f   1  (7  x �    y 	�   5�  �   ��  �   `�  �   �V 
�   _| 	7  '  

�     �   �  �   �  �  5�  �    ��  �   bpp 	�   `�  �   
 K  I  3  �  x 	�    y �    ^  	�  �  �  pos �   ֳ  �   �  �  �  5  r �    g �   b �   a �    �  �  	'u  �  �  (�   ֳ  )�   Y  *�   �  +�   
 
�  �  r    �  �  w  ,A  i   �r   std  r  �  
A
A�    �C  ��  ��  ��  ��  ��  �  �W  �r  ��  ��  ��  ��  �  �7  �I  �U  �g  ��  ��  ��  ��  �  �~  ��  �  �:  ��  �P  �p  ��  abs 	N   �  �  �   abs 	J%   �    �   abs 	F   �  "  �   abs 	=~   w  <  w   abs 	89   �   V  �    div ��  C  �   �     j  
�  �  
A
A  �~  �  �:  �P  �p  ��  ��  div ��  ~  w  w    	>      �    rem �    ?  �  	�	  C    �    rem �    �	    	3  w    w   rem w   '  4  O  m  I�   �  �   �  �  J�   �  �   �  '�  �  �   �  �  �  (�   �  �   E@ )�     �   R  V�  6  6  6  �  �  =   <  C  �   W  6  6   div a  r  �   �    �	  M�  �  �   �  �   bC  �  �   �    	  g�   �  �  �   �  m�  �  �  �  �   �  �  �  \  h�     �  �  �   �  X7  �  �  �  =   �  N#I  �      5�     7g  _      +�  �  �  �   �  $  .�   �  �  �  �    �  0r   �  �  �  �    2� O�   �  �   J  n�  �  �  �  �   �    i�     �  �   �   c	~  :  w  w   j  *w  P  �   W  /w  p  �  �  �    �  1�  �  �  �  �    �    ,�  �  �  �   \   -�  �  �  �   �  '�  +�  .7  3  4C  abs ]�   	  �    6	  6�  6�  6  6"  6<  7�  8�  9�  :  <�  <W  <V  >r  @�  C�  D�  E�  G  HI  JU  Kg  L�  M�  N�  P�  Q  �  �  ;5@            ��
  F  �'�
  �H src �8�
  �@�  �H�  ��!b  ��
  �`!z  ��
  �X"c5@     �       #i �
�   �l"�5@     �       #j ��   �h   =  �   $�  ��  �3@     ?      �V  F  ��
  �X src �-�
  �P�  �=�  �H�  �L�  ��!�  �	�   �h!<  �	�   �d!_  �	�   �`"�4@     �       #i �
�   �l  $�  �  #3@     �       ��  F  ��
  �X src �-�
  �P�  �=�  �H"73@     �       #i �
�   �l"e3@     �       !_  ��   �h   $�  ��  �1@     �      ��   x ��   �\ y �&�   �X5�  �-�   �T��  �8�   �P c1 �N5  �L c2 �`5  �H�  �o�
  � "�1@     #      #j ��   �l  $�  �  ?1@     W       ��  �  �"�  �` c1 �65  �\ c2 �H5  �X�  �W�
  �P $K  ��  �/@     j      ��   x ��   �\ y ��   �X5�  �%�   �T��  �0�   �P c1 �F5  �L c2 �X5  �H�  �g�
  � "0@     %      #j ��   �l  $�  �K  �-@     J      ��   x ��   �� y �!�   �� w �(�   �� h �/�   ��Kl  �;7  ���  �L�
  ��!�  ��  �B!X  �
�   �_!_  ��   �X!�  ��   �l!n  ��   �h!�  ��   �T".@     �      #i ��   �d";.@     ~      #j ��   �`"e.@     K      !�  ��   �P    $l  �&  :-@     Q       �:   x ��   �l y ��   �h5�  �!�   �d��  �,�   �`�  �B5  �\�  �U�
  �P $l  �^  ",@           �;   x ��   �L y ��   �H5�  �!�   �D��  �,�   �@ r �<�   �� g �G�   �� b �R�   ���  �`�
  �!�  ��   �h!_| ��
  �`"�,@     �       #i ��   �l"�,@     l       !�  ��   �\!4�  ��   �X   $l  �g  �+@     I       ��  �  ��  �`�  �*5  �\�  �=�
  �P %�  �T  �   �+@     .       ��   num ��  �X#x ��   �l %�  ~;    P+@     [       �  �  ~�  �Pc ~*�  �H ��  &�  p�  �
  �*@     u       �n  �  p/�  � �& p=�  �X!�  q�
  �h $�  ]�  �)@     �       ��  F  ]�  �X src ])�  �P/� ]5�  �H!��  c	�  �h!�  d	�  �` $�  I9  N)@     �       �H  F  I�  �X c I.�   �P/� I8�  �H!��  R	�  �h!�  S	�  �` '(  5�  )@     8       �F  5�  �h c 5.�   �d/� 58�  �X  �   �  9  K"  �  [6@     �      �  N  9   �  �  �  S   �  �  �  ;  int ,  C  �Z   �  -   �  G   ;
  4}   1  (  x o    y 	o   5�  o   ��  o   `�  o   �V 
�   _| 	  '  

�     �   �  �   �  	1  i   �Z   '  �  
i  �   @�  �  �   p   	=  �  #	=  X  &	=  �  )	=   �  ,	=  (�  -	=  0/  2o   8�  5o   < 1  �  8"^  +  K�  �  %  L�  �  M�  std  �  �  	A	A(  s  ��  ��  �  �  �=  �S  �i  ��  ��  ��  �   �  �M  �m  ��  ��  ��  ��  ��  ��  �  �5  �[  ��  �/  �v  ��  ��  ��  ��  �  abs N   P  T  P   abs J%   	  n  	   abs F   0  �  0   abs =~   I  �  I   abs 89   v   �  v    div ��  �  v   v     j  	K  �  	A	A�  ��  �v  ��  ��  ��  ��  �  div ��  �  I  I    
>  s    
o    rem 
o    ?  
K  
�	  �    
v    rem 
v    �	  
  
3  �    
I   rem 
I   4  
�  m  
Io   �  �     �  
Jo     �   �  
'0  0  7   �  8  �  
(o   S  7   E@ 
)v   i  7   R  
V\  �  �  �  =  =  �   �  �  o   �  �  �   div 
as  �  o   o    �	  
M�  �  7   �   
b�     v   v    	  
go     7  =   �  
m=  ;  ;  7  =   A  �  	A  \  
ho   m  ;  7  =   �  
X�  \  =  =  �   �  
N#�  o      
5o     
7�  S      
+0  �  7  �   �  $  
.v   �  7  �  o    �  
0Z     7  �  o    2� 
Oo   5  7   J  
n=  U  �  U  =   H    
io   v  �  A   �   
c	�  �  I  I   j  
*I  �  7   W  
/I  �  7  �  o    �  
1�  �  7  �  o    �    
,	  	  7  �   \   
-P  +  7  �   '�  +  .�  3s  4�  abs 
]o   i  o    6S  6:  6T  6n  6�  6�  7  8=  9S  :i  </  <�  <�  >�  @�  C   D  EM  Gm  H�  J�  K�  L�  M�  N  P5  Q[  �  S   )  A"Z	  `	  �   ��	  �  �\   ��  ��	  <h ��	  �I  ��	   �  X�	  �	  \  �	  N	  v    �   m�	  �	  �	  N	  \   f  ��	  �	  \  
  N	  v   v   \   J   �"&
  ,
   �  PH�
  !Ǟ  J)   !ֳ  KZ   "pos LZ   !  N�
  !/[  O�
   !�K P�
  (!�R Q/  0!ڰ  SN	  8!O�  T)  @!��  U)  H #�  ��
  $<v �v   $��  �\   �  ��
  ""  �    Z   )  
  Z   )  Z    9   �   <  B  M  
   v  :v   �  L}  x NM   y OM   �  QY  ~   w�  
  yM   �!  yM  �   zM  H  zM   "  |�   �  (V  !M} S    !5�  S   !`�  	o   !_| 
)  !
!  @   !?   9   !2   9   !B  \    �  �   �  (Q�  !   Sh    !0�  Th   !N5  V�  !�   W�  !H� X�  !�1  Zo     }  h   �  \c  %�  S   �  &�!   '�   pmoc'�  stib'u!  ltuo'�  tolp :  ��    �1  {"  �h   !  �@   \   �o   �  �S   }  �v   �   v   c   ��  �  �  \    �  ��  !Kl  �\   !�  �   s  ��  �"  $�  �   �   +!  !�� -�   !�W .�  !Kl  /\    %  DL  !uR F�   !�
 G�   }  I!   �  @<�  !5�  >M   !��  ?M  !�"  AM  !�"  BM  !i!  CM   !%!  EM  (!2!  FM  0!�  GM  8   IY   �"   s:  !��  u6   !5�  v6  !ֳ  xM  !!  zM  !m  {M   v  }�  J  �#T  Z  (�!  U  �"l  r  (�  T   � �  �   _  �K  !�!  f   !�  f  !�  f  !  f  !�  f   !�U F  (!�  F  0!3"  N  8!�  L  @!`  !N  H!d  "R  P!�@  $�  X!�;  )�  h!�   +B  �!�  ,6  �!
  -6  �!��  .6  �!?!  06  �!�  16  �!�  36  �!�  46  �!ȩ  6�  �!ֳ  7K  �!�� 8  �!K <_  �!ڰ  =N	  �!^�  >
  �!U  @L  �!t  B�  �!k  C\  �!�L  E.  � "   X  ^   1  Xm�  !��  ow   !�@  p�  !�e q�  !�L  rX  P @  $%�  �  )  0\  !�-  ^G   !��  _w  !�W `�  !x aZ  !�@  b�   !�e d�  0!�"  er  p!i"  fr  x!� g}  �!��  i  �!.a kV  �!�  lN  �!J  mN  �!Mj  o�  �!�  qZ  �!�  r�  �*M  t\   *Z  uv   *_"  wM  *(   xM  *Ud z\   *�L  |  ( �!  F#     Z!  A\  !��  Cw   !T D!  !�!  EB  !"  FB   %S  S   �!  &Y   '�  bmys'�  cinu'�
  sijs'    bg'�  5gib'F  snaw'  ahoj'�    bg'�  sijs'=    bg'�  5gib'�
  snaw'k  ahoj'�  BODA't  EBDA'�  CBDA'  1tal'�  2tal'�   nmra �  \  0  `);  A  (�"  *  :    �  �)e  k  (�!   b  8H�  !!  JB   !m  KB  !A� Mr  !�� Nr  !�  PM  !
  QM   !��  RM  (!�  SM  0 �  Up  x   �$	    (�!    �)!  '  (�"  +�   7  , 3  	,  +�   Y  -Z   -Z    .�  	C  	�ji     /�  �o   	�ui     /�-  �G  	�ui     /�  �w  	�ui     0=  �  X>@     �      ��  1str �  ��1x )S   ��1y 9S   ��1r D�   ��~1g O�   ��~1b Z�   ��~2�  h�  � 3�  �   �L3_| �  �@3C"  !	o   �X4�   �  3C"  o   �\ 5�?@     ]       �  6err *o   �� 7�?@     �      6i 0o   �T79@@     u      3�  1�   ��7i@@     E      6j 3o   �P7@A@     e      6val 80  ��3�!  9�   ��3  :o   ��3(  ;o   ��3�  <o   ��3   =�   ��     %  �   8A  ��   o   �9@     k      ��  9�  �1  ��:x �"o   ��:y �)o   ��:r �4�   ��:g �?�   ��~:b �J�   ��~9�  �X�  � /�  ��   �H/_| ��  �@5S:@     �       �  ;i �o   �\7d:@     w       /� ��   �[7�:@     Y       ;j �o   �T   5;@     \       �  ;err �o   �� 7v;@     �      ;i �o   �P7�;@     �      /�  ��   ��7�;@     O      6j  o   �L7�<@     _      6val 0  ��3�!  �   ��3  o   ��3(  o   ��3�  	o   ��3   
�   ��     <�  �   28@     �      �K  9Rl ��  ��/Q!  ��  �X/�  �	=  �P/�  �  �H5D9@     Q       )  ;err �	o   �D 7�9@     G       ;err �	o   �@  <�  �M  {6@     �      ��  /Q!  ��  �X/�  �	=  �P/�  �  �H5�7@     Q       �  ;err �	o   �D 7�7@     G       ;err �	o   �@  =-  ��"  [6@             � Q    �  �B@     �C@     g'  ../src/gfx/sse2.asm NASM 2.13.02 ��B@              �    �  9  #  �  �'  N  )   �  �  �  �  �  ;  int ,  �     a   ~   >   � 3  	m   	�ni      <&     &  �$  �:  �C@     �      �(  ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  s&  G   �  N   )  A"]  c  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  Q  -    �   m�  �  �  Q  U    f  ��  �  U     Q  -   -   U    J   �")  /  �  PH�  Ǟ  J,   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q9  0ڰ  SQ  8O�  T,  @��  U,  H �  ��  <v �-   ��  �U    �  ��  ""  �    @   ,    @   ,  @    2  �  �   F  L  W     v  :-   �  L�  x NW   y OW   �  Qc  	�  ~   w�  
  yW   �!  yW  �   zW  H  zW   "  |�  �  (e  M} N    5�  N   `�  	G   _| 
,  
!  0  ?   2  2   2  B  U     �  �  	e  �  (Q�     S)   0�  T)  N5  V�  �   W�   H� X�  �1  ZG     �  )  �  \w  �  �  N   �7  �!   �   pmoc�  stibu!  ltuo�  tolp :  ��  �8  5"Q  W  �$  �4  S�  x U)   len V0  e� W2   �#  Y\  	�  �%  {�  �  �  G   G   �  U    �  �#  ��  �  G     G   G   U    �.  �    ,  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(  �  (�/    0�  U   8*  �  @ r  �  u(  
,  	�  �2  (�  �  G   �  U   �   D  �3  ;    #  D   v)  ]0  6  K  D  ,  @    �3  yX  ^  G   w  D  @   U    H7  ��  �  G   �  D  �   �  51  0�  y2  �7   � ��   �#  *
 �K  / �w   $ �  ( 2$  ��  -4  l2  +  �,  �  $8  �2  	3  ?    ��   	J  {"  �)  !  �0  \   �G   �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U    :   �	  xx ��   xy ��  yx ��  yy ��   5  ��  		  8  �J	  ��  �D   ��  �s   $  �	  c   �d	  j	  u	  U    �  ��	  Kl  �U    �  �W	   s  �u	  �"  $�	  �	  �   +�	  �� -�	   �W .�	  Kl  /U    %  D$
  uR F�	   �
 G�	   }  I�	  N   �t  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<�  5�  >W   ��  ?W  �"  AW  �"  BW  i!  CW   %!  EW  (2!  FW  0�  GW  8   It  �"   sU  ��  u[   5�  v[  ֳ  xW  !  zW  m  {W   v  }   J  �#o  u  �!  �	}3  ڰ  	Q   {3  	�s  S0  	�s  �/  	�s  �1  	�  �1  	�z!  Y/  	�$
  �*  	��  (�)  	�3  0+:  	��!  8<8  	��!  X�*  	�s  � �3  �"@  F  �(  	�  Oe 	�a!   �-  	�b  ڰ  	�Q   U  �"�  �  �  8	�  ah 	!g!   Oe 	"b  U1  	#$
   ;+  	$�  0 i(  �$�  �  l;  �	�]  ah 	�g!   Oe 	�t!  y2  	�7   {:  	��  (�� 	�D  h/ 	�w  p�� 	��  x T   � j  p  _  �1  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"  s  8�  �  @`  !s  Hd  "�  P�@  $�	  X�;  )�  h�   +g  ��  ,[  �
  -[  ���  .[  �?!  0[  ��  1[  ��  3[  ��  4[  �ȩ  6�  �ֳ  71  ��� 8�  �K <  �ڰ  =Q  �^�  >  �U  @$
  �t  B�	  �k  CU   ��L  E  � "   >  D  1  Xm�  ��  o]   �@  p�	  �e q�  �L  r�  P @  $%�  �    0\�  �-  ^b   ��  _]  �W `�  x a  �@  b�	   �e d�  0�"  e�  pi"  f�  x� g�  ���  i7  �.a ke  ��  ls  �J  ms  �Mj  o�  ��  q  ��  r�  �M  tU    Z  u-   _"  wW  (   xW  Ud zU    �L  |�  ( �!  F#�  �  Z!  AB  ��  C]   T D  �!  Eg  "  Fg   S  N   �  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  B  0  `)!  '  �"  �	e�  �1  	g	   H+  	h�   x+  	is  0��  	k�  8�)  	n#[!  h�'  	q   p��  	r7  t�*  	ys  x J  U  �  �  �)�  �  �!  H	�  $  	�U    7:  	��  s4  	��   b  8H�  !  Jg   m  Kg  A� M�  �� N�  �  PW  
  QW   ��  RW  (�  SW  0 �  U  x   �$�  �  �!  0
'�  ad  
)s   �1  
*g  &D  
+s  2B  
,s  x� 
-	     �)�    �"  P	�v  ��  	��   �1  	�  �&  	�  �3  	�	  ]7  	��  0�7  	�U   @�1  	�7  H P6  �  tag �   Kl  �   �6  	v  �  �5  N   
�  i7   �&  9  F9  8%  �*   �,  
�  ./   6
N  b 8
�   5�  9
�  ��  :
�  5  ;
  Q(  <
    -  I
([  �  �8  N   ��  �:   4,  �6  $  �/  l9   �2  �a  �#  ��  �'  ��  �  �  �  3   �2  ��  �  �  3   l/  ��    �    3     �   ;)  H��  �#  ��   :  ��  �5  ��  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  ��  8��  ��  @ V  �-  �  	�  d)  s�  �  �  �  U    9  F#�  	�  �$  @J_  �#  L�   y2  M7  W� O�  �� P�  �,  QQ   M4  R�  (�;  S)  0�*  Tw  8 c/  X!k  q  �-  (q�  �-  sb   Oe t�  ��  u7  � v�   �  �/  )�  �  �  �  _  �   g%  .�  �  �  _   �.  1    #  _  #  �   	  73  65  ;  K  _  K   �  �8  :]  c  �  w  _  _   "3  >�  $)  Y�  �  �  �  �  �  �  �   �6  _�  �  �  �  �  �  #  �   �3  f�  �  
  �  �  K   ;0  l    �  5  �  �  �   �&  x��  ah � �   y2  � 7  H�8  � �  P�8  � �  X�'  � �  `� � 
  h�9  � �  p   �.  �5  	�  "9  H
2  Mj  
4�   H5  
5�  (�)  
6�  0�  
7  8�  
8�  @ �0  
:�  T%  �
=�  ڰ  
?Q   �0  
@  q5  
A  L)  
B  )  
C  Ǟ  
E  �  
F  `Ud 
HU   � X+  
J�    1  �  �  �  �    ]  s  s  �   �&  &�  �  �  ]   �1  *�  �  �    1   �6  -    (  1   w-  14  :  �  I  �   �;  4U  [  f  �   =;  8r  x  �  �  1  N   B$  <�  �  �  �  1  �   2  @�  �  �  �  �  1    7   7  G�  �  �    ]      �   q8  N  $  �  8  ]     )2  SD  J  �  m  ]      7  m   �  k.  ��Q  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q ��  hZ)  ��  p�#  �  x'0  �(  �.  �I  ���  ��  �� ��  �`9  �  ���  �8  �5  �f  �U#  ��  � �/  �s  	Q  �2  �n  s  �&  0��  y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  �t  *  V'�  �  �0  �*   u=   |#  w�   �#  x�  � y�  C4  z�   �&  |�  �'  �U   [   �  t   �    t    J	  �9  ��   �   �   �  t    A2  ��   �   �  �   �      �    =   8(  !  ��  )I    $�  )z   �-  )�    )  �   	!  3  <H!  �� >%H!   ��  ?%�   !  #  A!  N!  �  �(  	�F  �  3  �!  @    �  �!  @    �  �!  @    H'  	�%  
�7  ]  
k3  ]  
�1  ]  
�)  ]  
�8  ]  
�4  ]  
!1  ]  
2  	]  
g+  
]  
�7  �  
�-  �  
]4  �  
!+  �  
�$  �  
�#  �  
�.  �  
�(  �  
�/  �  �"  �"  @    	�"  �  	�"   y6  F!�"  	��F     !;  ��  @F@     &       �=#  "�-  �!b        #ڰ  �Q  d   b   $NF@     �%  (#  %U�U &VF@     �%  %Us   !�4  ��  �E@     �       �S$  "�-  �"S$  �   �   #�U ��      #ڰ  �Q  r  j  '^%  �E@      �E@     $       �$  (k%  �  �  )�E@     $       *w%  +�%  �  �  &�E@     �%  %Uv    ,�E@     &  $�E@     &  1$  %Us %T|  ,�E@     Y$  &F@     �%  %Us   b  -4  p D@     �      �N%  "�-  p*b  j  b  .env r  �  �  .p s     �  .q t  �  �   �5  vN%  ��| �1  wN%  ��} �,  xN%  ��~.i z
G   5    $D@     &&  $%  %U	p�F      &RE@     2&  %Us %T��|%Q��}%R��~  �   ^%  @   � /�3  P�%  0�-  P'b  1�U R$�  2cur S$�%   �"  3^%  �C@     3       ��%  (k%      *w%  +�%  r  j  &�C@     �%  %Uv   4�+  �+  Q4b8  b8  	�4�1  �1  4�:  �:  	�4|&  |&  85�	  �	  M4B/  B/  	> �|    y&  Nr  �:  pF@     Ѹ      �-  R�  (\  �@   R,  i   �-   zint R�  {!�   @�   	�  �    	p   	G   	�  #	G   	X  &	G   	�  )	G    	�  ,	G   (	�  -	G   0	/  2S   8	�  5S   < �   R�  +�   �  8"c   c+  K  �   c%  L  c�  M  R'  �M  A  /@   Q  0-    R;  �s  �d  R�  s&  S   +k  �  Z   \i  g@   �<  h-   )  A"�  �  !�   ��  	�  �a    	��  ��  	<h �  	�I  �@   �  X  
  a     �  @    �   m*  0  2@  �  a    f  �L  R  a   p  �  @   @   a    J   �"|  �  �  PH  Ǟ  J   ֳ  K-   Epos L-     NC  /[  OC   �K PO  (�R Q�  0ڰ  S�  8O�  T  @��  U  H i�  �C  j<v �@   j��  �a    �  �  ""  �[  a  -     p  -     -    �  R�  �   �  �  2�  p   v  :@   !�  L�  Xx N�   Xy O�   �  Q�  +�  !~   w-  	
  y�   	�!  y�  	�   z�  	H  z�   "  |�  ]N`  Z   ��  
�T   
jt  
�C  
�H  
�H  
�K  
RR  
Zs  
WO   �o  �9  �  (  M} Z    5�  Z   `�  	S   _| 
  
!  d  ?   �  2   �  B  a     �  �  +  �  (Q�     SQ   0�  TQ  N5  V�  �   W�   H� X�  �1  ZS     �  Q  �  \  +�  �P  ��  �  S   �  �  a    �  m\  �  �N  4�  �  S     �  �  a    �s  X    S   7  �  �  �  a    K[  0��   ��   - ��  �
 ��  Q �  m�  �S    �� ��  ( �l  �7  +�  S�  Z   ��  
�!   3�   pmoc3�  stib3u!  ltuo3�  tolp :  ��  �8  5"  
  Y�$  �4  SF  Ex UQ   Elen Vd  e� W�   �#  Y  +F  �%  {e  k  2�  S   S   �  a    S  �#  ��  �  S   �  S   S   a    �.  ��  �  2�  S   S   a    �8  `�l  .   l   �; r  �1  S   �5  X  �+  X   `(  �  (�/  �  0�  a   8*  -  @   x  |u(  
�  +y  �2  (�  �  S   �  a   �   �  �3  ;�  �  2�  �   v)  ]�  �  2�  �    -    �3  y	  	  S   *	  �  -   a    H7  �7	  =	  S   Q	  �  Q	   �  51  0��	  y2  ��   � ��   ��  *
 ��  / �*	   $ ��  ( 2$  �W	  -4  l�  +  ��	  R�  $8  ��  +�	  �	  Ab  �}    ��   +	
  {"  �Q  !  �d  +&
  \   �S   �  �Z   }  �@   )$  �-   _]  @   �   @   c,  +S   C*  6a   +D  CG   �]  P4    :   ��
  Exx �t
   Exy �t
  Eyx �t
  Eyy �t
   5  ��
  +�
  8  �5  ��  ��	   ��  �7
   $  �
  c   �O  U  2`  a    �  ��  Kl  �a    �  �B   s  �`  �"  $�  �  �   +�  �� -�   �W .�  Kl  /a    �j   �  �  %  D"  uR F�   �
 G�   }  I�  }Z   ;�r  
10   
�(  
Q;  
�4  
�(  
�0  
*  
/  
d2  
�+  	
a0  

~5  
�0  
k*  
�,  
U5  
l1  
�.  
�)  
�/  
l,  
a-   
.  !
�5  "
-5  #
�%  $
�*  %
�-  &
_:  '
N*  (
�8  0
a#  1
(  @
�$  A
I,  Q
.  R
6  S
^6  T
�9  U
L3  V
�(  W
�:  X
�7  `
Z'  a
�,  b
�7  c
�%  p
U.  �
I8  �
�,  �
�5  �
+  �
r'  �
�9  �
U$  �
-  �
�4  �
�4  �
�1  �
i$  �
@-  �
#(  �
�0  �
/7  �
�+  �
�+  �
E:  �
x0  �
+'  �
'  �
�'  �
�)  �
�%  �
,  �

8  �
9.  �
0  �
|;  �
�:  �
54  �
�5  �
+-  �
�2  �
�-  �
�2  �
+6  �
�3  �
�9  �
�6  �
�%  �
39  �
�$  �
8#  �
�:  � �  @<�  5�  >�   ��  ?�  �"  A�  �"  B�  i!  C�   %!  E�  (2!  F�  0�  G�  8   Ir  �"   sS  ��  u
   5�  v
  ֳ  x�  !  z�  m  {�   v  }�  J  �#m  s  ^�!  �}1  ڰ  �   {3  �7
  S0  �7
  �/  �7
  �1  �C
  �1  ��(  Y/  �"  �*  ��  (�)  �1  0+:  ��(  8<8  ��(  X�*  �7
  � �3  �">  D  �(  �}  Oe ��(   �-  �`  ڰ  ��   U  �"�  �  �  8�  ah !�(   Oe "�"  U1  #"   ;+  $/   0 i(  �$�  �  l;  ��[  ah ��(   Oe ��(  y2  ��   {:  �1  (�� ��  h/ �*	  p�� ��  x T   � h  n  _  �/  �!  O
   �  O
  �  O
    O
  �  O
   �U �  (�  �  03"  7
  8�  �  @`  !7
  Hd  "�  P�@  $�  X�;  )-  h�   +&
  ��  ,
  �
  -
  ���  .
  �?!  0
  ��  1
  ��  3
  ��  4
  �ȩ  6�  �ֳ  7/  ��� 8�  �K <}  �ڰ  =�  �^�  >p  �U  @"  �t  B�  �k  Ca   ��L  E  � "   <  B  1  Xm�  ��  o[   �@  p�  �e q�  �L  r�  P @  $%�  �  ^  0\�  �-  ^`   ��  _[  �W `�  x aC
  �@  b�   �e d�  0�"  et
  pi"  ft
  x� g�  ���  i�  �.a k  ��  l7
  �J  m7
  �Mj  o�  ��  qC
  ��  r�  �M  ta    Z  u@   _"  w�  (   x�  Ud za    �L  |
  ( �!  F#�  �  Z!  A@  ��  C[   T D  �!  E&
  "  F&
   SS  Z   �  
Y   3�  bmys3�  cinu3�
  sijs3    bg3�  5gib3F  snaw3  ahoj3�    bg3�  sijs3=    bg3�  5gib3�
  snaw3k  ahoj3�  BODA3t  EBDA3�  CBDA3  1tal3�  2tal3�   nmra �  @  �C  H�  0  `),  2  �"  �e�  �1  g�
   H+  h�   x+  i7
  0��  k�$  8�)  n#g&  h�'  q�	  p��  rk  t�*  y7
  x 	
  S  �  �S  In  �  �)�  �  �!  H�  $  �a    7:  �O  s4  ��   b  8H�  !  J&
   m  K&
  A� Mt
  �� Nt
  �  P�  
  Q�   ��  R�  (�  S�  0 �  U  x   �$�  �  !�!  0'
  	ad  )7
   	�1  *&
  	&D  +7
  	2B  ,7
  	x� -�
     �)    �"  P��  ��  �/    �1  �C
  �&  ��	  �3  ��
  ]7  ��  0�7  �a   @�1  �k  H P6  �  Etag [
   Kl  �
   �6  	�  c  @KE  �1  MC
   %_  N�	  c  OO
  /[  P�  ^�  Qp   K R1  (�[  S7
  0\  TE  8 �  �e  V�  +K  S�5  Z   
�  
i7   
�&  
9  
F9  
8%  
�*   �,  
]  ./   6
�  b 8
�   5�  9
O
  ��  :
O
  5  ;
C
  Q(  <
C
   'b  >
�   -  I
(  �  S�8  Z   �O  
�:   
4,  
�6  
$  
�/  
l9   �2  �  S�u  Z   Z�  
�R   
�l  
�]   �\  ��  b<  �C
   1S �C
  Ep ��   �	  p  ��  �#  ��
  �'  ��  �  �
  �  1   �2  �    2  1   l/  �"  (  �  <  1  <   �   !;)  H��  	�#  �[
   	:  �O
  	�5  ��  	F1  �t
  	,8  �t
   	2*  �r  (	�*  ��  0	`1  ��  8	��  �  @ 
  �-  �B  +�  d)  s�  �  �
  �  a    S�j  Z   �$  
jb   
�U  
�P   �B  ��  9  F#B  +1  !�$  @J�  	�#  LO
   	y2  M�  	W� O  	�� P8  	�,  Q�   	M4  RU  (	�;  S�  0	�*  T�  8 c/  X!�  �  !�-  (q  	�-  s`   	Oe t  	��  u�  	� v�   =  �/  )  $  �
  8  �  �   g%  .D  J  2U  �   �.  1a  g  2|  �  |  �     73  6�  �  2�  �  �   -  �8  :�  �  �
  �  �  �   "3  >  $)  Y�  �  �
    �  �  O  �   �6  _    �
  <  �  �  |  �   �3  fH  N  2c  �  �  �   ;0  lo  u  �
  �  �  [
  �
   !�&  x��  	ah � �   	y2  � �  H	�8  � �  P	�8  �   X	�'  � <  `	� � c  h	�9  � �  p �	  �.  ��  ]�@  Z   �@  
e   
,J  
f  
�f  
i  
.F   �C  �	  !"9  H2�  	Mj  4�   	H5  5�  (	�)  6�  0	�  7C
  8	�  8�  @ �0  :L  7<  :�  L  !T%  �=/   	ڰ  ?�   	�0  @C
  	q5  AC
  	L)  BC
  	)  C�	  	Ǟ  E�  	�  F�  `	Ud Ha   � X+  J;   �  1   M   S   �
  v   p  [  7
  7
  E   �&   &�   �   2�   [   �1   *�   �   �
  �   /   �6   -�   �   2�   /   w-   1�   �   �
  �   �   �;   4�   !  2!  �   =;   8!  !!  �
  5!  /     B$   <A!  G!  �
  [!  /  [
   2   @g!  m!  �
  �!  �  /  C
  k   7   G�!  �!  �
  �!  [  C
  C
  �   q8   N�!  �!  �
  �!  [  p   )2   S�!  �!  �
  "  [  C
  C
  k  "   t
  !k.  � ��"  	ah  ��   	#,   �O
  H	�4   �O
  P	,;   �O
  X	EY  �A   `	/q  �v   h	Z)   ��   p	�#   ��   x	'0   ��   �	.   ��   �	��   �[!  �	�  ��!  �	`9   ��!  �	��   ��!  �	5   �!  �	U#   �5!  � �2   �#  "  0t  !P&#  #  Y�h  �V  !m/#  5#  2O#  #  [  O#  U#   a   @   EU  !�g#  m#  2}#  #  a    j]  !��#  �#  2�#  #  [   �l  !��#  �#  �
  �#  #  �  /  C
  k   !t>   !�$  	�=  !�$}#   	[I  !�$##  	�d  !�$[#  	��  !�$�#   H  !�""$  �#  !8S  "�P$  	�d  "�<   	�W  "�r   C  "�($  +P$  �F  "�%m$  \$  �&  0"��$  y%  "��
   �/  "��
  �'  "��
  �6  "��
  �+  "��
   �6  "��
  ( �7  "�s$  *  #V'�$  �$  Y�0  !�*   #u<%  	|#  #wO
   	�#  #xO
  	� #yO
  	C4  #zO
   �&  #|�$  �'  #�T%  Z%  �
  s%  �$  C
  s%   5  �9  #��%  �%  2�%  �$  s%   A2  #��%  �%  �
  �%  �$  C
  �	  �%   <%  8(  #
&  ��  #)H%   $�  #)y%  �-  #)�%   )  #�%  +
&  3  #<G&  �� #>%G&   ��  #?%�$   &  #  #A&  �o  #M*g&  M&  �U  �,y&  &  !�B  ��&  	�� �   	Oe ��&   fP  �,�&  I'  !4I  P�I'  	ֳ  �[
   	�� �N'  	�q �t'  	R` ��'  	�W ��'   	P �#�'  (	�U  �#(  0	�v  �#>(  8	�v  �#d(  @	�J  �#�(  H +�&  wq  �Z'  `'  �
  t'  m&  �
   �J  ��'  �'  2�'  m&   �\  ��'  �'  C
  �'  m&  }   \  ��'  �'  C
  �'  m&  �'   }  U  ��'  �'  C
  (  m&  m&  }  }   �O  �(  %(  7
  >(  m&  }  }   �n  �J(  P(  �'  d(  m&  �   ;O  �p(  v(  �'  �(  m&  �  }   -k  �p(  �  �(  �D  �  �D  &�  /1  �(  0-    /�  �(  0-    /�  �(  0-    �(  <  )  [   )  �
  *)  [  C
  �
  C
   0)  C
  D)  [  �   ~H'  �%�	  nq  $4t
  +Q)  !�I  `%UM*  	Q  %Wt
   	�g  %Xt
  	�;  %ZO
  	�U  %[O
  	�B %]&
   	�o  %^&
  "	Y  %`M*  (	+I  %aM*  8	
  %c
  H	�!  %d
  J	�   %e
  L	H  %f
  N	�`  %h&
  P	�X  %i&
  R	O  %k
  T	,G  %l
  V	�t  %m
  X /[
  ]*  0-    I  %ob)  !�g  8%�G+  	��  %�t
   	)r  %�
  	dS  %�
  
	�B  %�
  	�P  %�&
  	�p  %�
  	�K  %�
  	=  %�
  	me  %�
  	+^  %�
  	�]  %�
  	�u  %�G+  	
h  %�
  $	^K  %�&
  &	tR  %�a   (	%?  %�a   0 /
  W+  0-    �]  %�i*  �S  8%?R,  ��  %At
   )r  %B
  dS  %C
  
�B  %D
  �A  %F&
  �n  %H
  �n  %I
  �W  %J
  me  %K
  +^  %L
  �]  %M
  �u  %OG+  
h  %Q
  $�V  %R&
  &tR  %Xa   (%?  %Ya   0 �u  %[c+  JW  �%x�.  ��  %z&
   =  %{
  �<  %|&
  tB  %}&
  �k  %~&
  �m  %
  
�D  %�
  gJ  %�
  !X  %�
  �S  %�
  5f  %�
  ?X  %�
  �a  %�
  �_  %�
  �a  %�
  Gf  %�
  �=  %��.   �E  %�[
  0F  %�[
  8�A  %�[
  @F  %�[
  H�E  %��.  P5D  %�&
  TH  %�&
  V#l  %�&
  X$r  %�
  Z_S  %�
  \'N  %�
  ^?_  %�&
  `L  %�&
  b�O  %�[
  h�O  %�[
  p~e  %�
  x [  %�
  z0m  %�&
  |�M  %�&
  ~rM  %�&
  �]  %�&
  ��g  %�&
  � /�	  �.  0-   	 /�	  �.  0-    �X  %�_,  kE  @%�J/  �^  %�t
   zp  %�t
  dv  %�
  �i  %�
  �<  %�[
  �F  %�[
   �D  %�[
  (�p  %�[
  03X  %�[
  8 �b  %��.  K_  @%�80  ��  %�t
   �J  %�[
  �<  %�&
  e  %�&
  $� %�&
  dk  %�&
  ![  %�&
  L^  %�&
  �`  %�80  yN  %�H0  ,ma  %�X0  4�Z  %��	  :�q  %��	  ;r  %��	  <�u  %��	  = /�	  H0  0-    /�	  X0  0-    /�	  h0  0-    	l  %�W/  �M  (%8V1  ��  %:t
   �T  %;&
  �P  %<&
  
�K  %=&
  B  %>&
  ^  %?&
  �g  %@&
  /o  %A&
  %B  %B&
  �O  %C&
  �<  %D&
  �]  %E&
  *w  %F&
  dW  %G&
   �F  %H&
  " e=  %Ju0  Sm<  Z   %m�1  
nA   
ZY  
TE  
�U  
�R  
{H  
b  
�c   �`  %yc1  !|[  &O�1  	�� &Q�	   	�\  &R�	  Xred &S�	  	q  &T�	   �[  &V�1  !�?  (&�Q2  	`a  &�&
   	�L  &�Q2  	r  &�Q2  	&W  &�&
  	�F  &�Q2    2
  Ik  &�2  +W2  O
  !>i   'J�2  Xtag 'L[
   	��  'Mt
  	/� 'NO
  	�f  'O�2   [
  2\  'Qn2  !G   '�3  XTag '�[
   	g  '�[
  	�=  '�[
  	Ja  '�[
   mn  '�3  �2  !�v   '�3  	�T  '�&
   	�Y  '�&
  	D  '�&
  	S  '�&
  	E]  '�&
  	;C  '�[
  	�: '��   �[  '�3  M  '��3  3  DQ  '�3  E]  '&
   ;C  '[
  �: '�   �i  '�3  hh  '�3  �3  >M  0'.g4  ��  '0&
   �Z  '1C
  vv  '2C
  �r '3g4  =P  '4C
  �Q  '5m4   ^�  '6p  ( 3  �3  �p  '8�3  CE  'Y�4  �B  '[&
   b  '\&
   Pq  '^�4  �4  �m  'x�4  ��  'z&
   �R  '{&
  Up  '|�4   �=  '~�4  �i  '��5  ��  '�&
   5�  '�&
  �"  '�
  �"  '�
  i!  '�&
  %!  '�
  
2!  '�
  �  '�&
   W  '�5  �U  '96  �  '�	   
  ' �	  Sd  '!�	  �Q  '"�	  �G  '#�	  �v  '$�	  �=  '%�	  sD  '&�	  �\  ''�	  �X  '(�	  	`N  ')96  
 /�	  I6  0-    �T  '+�5  &
  >t  '��6  �>  '�I6   � '�I6  !  '��	  m  '��	  �[  '��	  SX  '��	   �<  '��6  \6  x@  '"7  �  '$&
   �`  '%&
  TL  '&V6  �o ''7   7  �	  �h  ')�6  �Z  '<]7  �  '>&
   �f  '?7   fR  'A27  'Z�7  kj '\%7  k�Y ']]7   ms   'V�7  �  'X�	   �r '_j7   J  'a�7  �t  'r!�7  �7  YU<  �c  ('�B8  �B '��   �c  '��  �y '��  �Y  '�[
  cC  '�C
   �  '��	  $ 	\  '��7   L  '� \8  b8  ^�i  �'�=  ah '��   �u  '��2  ��v  '�[
  �R  '�&
   o  '�3  (�& '�]*  0�Q  '�W+  �@  '�V1  �5�  '��	  �<  '�R,  ��`  '�&
  0�a  '�s4  8Uos2 '��.  hF�  '�J/  �j  '��  0 M  '�[
  8w_ '��>  @�>  '�!?  H�A  '�t?  P^Z  '�R?  X�f  '�R?  `KT  '�R?  h�i  '�a   pQ  '�a   xUmm '�a   �Uvar '�a   �g  '�a   ��Y '��4  �Fq '�h0  �jQ  '�[
  �nQ  '��6  �m  '�7  ��P  'W2  @  '&
  @B  '�?  H�u  '�	  P�u  '�1  Q�;  '[
  XzQ  '�  `FN  '[
  hT  '�  p!u  '[
  xUcvt '�?  �2i  '=  �)  ')�  ��  '+<  ��j  '-[
  �:>  '.[
  ��_  '0�	  �S?  '3�	  �E�  '4�7  ��W  '6}  �XA  '8<  �	K  '9C
  ��c  '?[
  �][  '@[
  ��J  'B[
  �'<  'C�  �	Z  'E�   �q  'F[
  �G  'GC
  �T  'H[
  �a  'I�   �\  'K�  (�u  'L[
  0o  'M�?  8^C  'NC
  <:W  'O�?  @_  'Q�  H�@  'R[
  P>  'SC
  X}?  'T}  \m?  'U}  `Ubdf 'XB8  h�k  '\[
  ��Z  '][
  �Pl  'h[
  �(a  'i[
  �i 'ma   ��d 'na   � �Q  '��  �g  '�"9=  ?=  ^�t  x'��>  ��  '�O8   ֳ  '��@  ȩ  '��  �m  '�/   �1  '�[
   x '�C
  (^�  '�p  0��  '�7
  8   '�
  <�;  '�-  @�C  '�7
  `� '�7
  d"f '�7
  h�I  '��	  lEpp1 '��  pEpp2 '��  �Ǟ  '��@  ��y  '��@  �BJ  '��@  �<  '��  bL  '�[
   Ud '�a   (�W  '�7
  0r�  '�7
  4Upp3 '��  8Upp4 '��  HO�  '��  X��  '��  `�k  '�"  h �^  '�>  ?  �
  !?  O8  [
  p  �2   �D  '*.?  4?  �
  R?  ,=  C
  [
  C
   �b  'A_?  e?  �
  t?  ,=   SQ  'Q�?  �?  2�?  ,=   S�=  Z   'T�?  
�G   
�v  
k_  
<L  
ok   �`  '_�?  �1  k  C
  �j  @'��@  ڰ  '��   �0  '�&
  q5  '�
  
0�  '�&
     '�
  Eorg '��  Ecur '��  " '��   �   '��  (H� '�V6  0�>  '�&
  8 ,L  '��?  @\  '�'�@  �@  Y�r  �d  '� �@  �@  Y�a  <e  (I�@  �@  �
  �@  p  O8  7
  7
  E   l  (s�@  Z  (�A  A  2'A  O8   -H  (�3A  9A  �
  \A  O8  [
  O
  �  �2   �e  (2iA  oA  �
  �A  O8  [
  C
  C
  p  �A  �A     �5  �h  (S�A  �A  �
  �A  O8    �2   �^  (p�A  �A  �
   B  O8  [
   B   �  eN  (�B  B  �
  2B  O8  C
  2B   �  Ub  (�EB  KB  �
  dB  O8  p  �	   #K  (�qB  wB  2�B  O8  �	  C
  �B  V6   
  3l  (��B  �B  �
  �B  O8  C
   �d  (	�B  �B  �	  �B  O8  C
  �?  �?  �B   �  �J  (0C  C  �
  0C  O8  C
  �  �   CZ  (N=C  CC  �
  \C  O8  &
  2B   :=  (piC  oC  �	  �C  O8  &
  �C  �C   7
  �Z  (��C  �C  �
  �C  O8  p   �^  (�A  GK  (��C  �C  7
  �C  O8  C
  C
   ^N=  0(�F  w_ (�"�>   EY (�"�@  �e (�"�@  /q (�"
A  ��  (�"   ob (�"'A  (pR (�"�C  0�^ (�"8B  8D_ (�"�C  @x` (�"�C  HPr (�"�C  P1s (�"�C  X�k (�"�C  `�S (�"�C  h�O (�"�C  p�Y (�"�C  xAq (�"�C  ��b (�"�C  �ar (�"\A  ��[  (�"B  � Q  (�"�C  �� (�"�C  �X (�"�C  ��U (�"8B  �`H  (�"�C  ��W  (�"�C  ��n (�"�A  ��T (�"�A  �zi ( "�C  ��d ("�C  ��Q ("�C  ��] ("�C  �B  ("�B   UU ("�B  �p  ("�B  �[ ("dB  ]o (
"0C   4P ("\C  ( sh  (�C  AD  (7F  F  l�P  
c2  (                                        ihG  )5�F  mnum )77
  mstr )8<   *f  ):rF  !�_  )=�F  Xkey )?�F   	Kl  )@G    �K  )D$�F  �F  �d  )H�F  �F  [
  �F  �F   �F  �r  )KG  G  �	  +G  �F  �F   !Uj  ()O�G  	��  )QC
   	ֳ  )RC
  	[M )SC
  	�V  )U�F  	�F  )VG  	�B )X�G    �F  �@  )\ �G  +G  ]<  Z   *9H  
�?   
Mm  
2a  
�=  	
2r  
�u  
0@  
�>  
gd  
�e  
Lo  
s  
�Y  
�^  
�f  
�l  
E  
�M   !_c  *VSH  	<v *X�	   	ֳ  *Y�	  	�  *Z&
   yK  *\H  +SH  �p  +�pH  vH  �
  �H  �  a    `  +��H  �H  2�H  �  a   a    S�[  Z   ,�H  
 Y   
zS  
�e   
ti  
�M   �m  ,%�H  �u  -*.�H  QI  !�R  X-XQI  	�Y  -Z5   	Ǟ  -\�	  @	��  -]�	  H	gY  -^|I  P	�U -_�
  T �I  ]�G  Z   -F|I  
X   
�t  
*u   �k  -LWI  !�h  .,�I  	�s  ..
   	�  ./O
   a  .1�I  �i  .6�I  �I  �
  �I  `  p  �   �I  h2   �   ]�B  S   .<LJ  n	m  ~n�c  
�\   
�h  
TB  
#j  
�F  
 W  
�?  
}T  
Ch   *S  .H�I  !�m  .N�J  	3 .O�I   	b .PLJ   �X  .QXJ  +�J  �  �  !xX  h/*�J  	ah /,�(   	�q  /.C
  8	�'  //�	  <	iO  /0�J  @	��  /1k  ` /7
  �J  0-    Y  /3K  �J  �<  0K   K  �
  >K  1  <  r  �	   s=  0$JK  PK  �
  iK  1  <  a    !#P  0)�K  	R  0+K   	bD 0,>K   +iK  8`  0)�K  �K  �g  1(�K  �K  �
  �K  [  [
  O
  �  �2   3?  12�K  �K  a   L  [  �1   �K  1:L  L  �
  8L  [  C
  �2  �2  �2   !6q  1AmL  	�s  1C�K   	I  1D�K  	Y 1EL   +8L  �Q  1A~L  mL  �d  2)�(  !`p  2,�L  	g 2.�L    +�L  �e  2,�L  �L  �A  3&)  �V  3,*)  !tG  30M  	]o 32!�L   	�  33!�L   +�L  T  30M  M  !V^  49AM  	�L  4;[
   	��  4<O
   �`  4>M  {V  4BYM  _M  �
  sM  �  sM   AM  !�N  4F�M  	�  4HMM    +yM  ]g  4F�M  �M  'd  5 �M  �M  �
  �M  [  t
  7
  "   !T_  5%�M  	F  5'�M    +�M  �L  5%N  �M  !�p  6'(N  	�B  6)$    +N   >  6'9N  (N  lHj  	&�  (                                        /�J  �N  0-    +tN  \m  ��N  	�F     !OP  7l�N  	�!  7n&
   	"  7o&
  	�q  7p&
  	8P 7q&
  	�: 7s�  	��  7tC
   �i  7v�N  !v  7�0O  	�: 7��   	��  7�C
   �_  7�O  /])  LO  0-    +<O  F]`  1LO  	 �F     I�M  ��O  �q  �)�  �� �)�H  ڰ  �)�  �  �)a   'cur ��  >�W ��  Kl  �a     �J  }�
  ��@     V       ��P  �q  }&�  �  �  ��  ~&dH  7  +  �  &a   �  �  cur ��  [  S  �U ��
  �  �  %��@            �W ��      �@     T|    I�i  \�P  �q  \�  �K  ]�  �j  _�  R  _�   I�g  AQ  �q  A �  �K  B �  �j  D�  R  D�   6�T  ' �@     .       �pQ  �q  ' �  U�K  ( �  TR  *�  F  B   I
^  �Q  �q  �  �K  �  �j  �   J\u  ��  �Q  "�q  ��  "Kl  �a   *cur ��   )u  �7
  ��@     O       �;R  Bdst � �   �  |  Bsrc � <  �  �  ֳ  � [
  	  	   )=T  ��
  @�@     2       ��R  ڰ  ��  L	  D	  Bstr �<  �	  �	  >H  ��R  
  
  #len �[
  {
  y
  \�@     | �R  Us  .r�@     �R  U�UT�TR�Q  �
  )!G  ��
  ��@     w       �T  ڰ  ��  �
  �
  �& �r      ֳ  �[
  �  �  >H  ��R  6  *  (�U ��
  *p ��
  7�V  ��@      pU  ��S  �V  �  �  �V  �  �  �V  ~  v  pU  K�V   �V  �  �  ��@     U�UTv    �@     $| T} Qv   _�s  �(T  "ڰ  ��  AP �r   )Cs  r�
  `�@     �       ��U  ڰ  r�  m  [  Kp  sO
  D  4  q  tO
  
  �  �F  uO
  �  �  *�  va   |  h  >H  w�R  c  Q  �U y�
  3  %  ?�@     5       ;U  ^=  ��
  �  �  (wO  �O
  (v  �O
  '�@     U�UT�T�QRw   7T  ��@      �D  ��U  T  �  �  T  3  /  ��@     U�UT�X  ��@     U�UT�R�T  )�I  \�
  P�@     x       ��V  ڰ  \�  p  l  Kp  ]O
  �  �  q  ^O
  0  (  �F  _O
  �  �  *�  `a       >H  a�R  �  �  F�U c�
  �Lz�@     (T  �V  U�UTv Q~ Rs X�XY�L ��@     /| U} v "T0Qs �T  J�U  B�
  �V  "ڰ  B�  "ֳ  CO
  ">H  D�R  (�U F�
  (*�  G�
   )�`  2�
   �@     g       ��W  ڰ  2�      ֳ  3O
  |  p  >H  4�R      (�U 6�
  (*�  7�
  7�V   �@      @:  7�W  �V    }  �V  �  �  �V  @  8  @:  K�V   �V  �  �  �@     U�UTs    )�@     /| T0Qs   G  �Q)  д@     /       �TX  �D  �Q)  U�D  �Q)  T�� �Q)       6tP  ���@     !       ��X  ;vec �%�  H  B  ��  �%t
  �  �  �  �%Q)    �  .��@     �Z  U�UT�Q  6UG  ���@     �       ��Y  ;vec �#�  V  N  ��  �#"  �  �  �  �#�Y  >  4  m�  �7
  �  �  Lv ��  �P`  "�@       :  ��Y  +`    �  :  7`  �  �    �@     �T �Y  Uu Tt 1�_  u  �@     T Uu 1_  u   Q)  @a  �t
  ��@     �       ��Z  ;vec �!�  9  /  m�  �7
  �  �  Lv ��  �``  ��@       �9  �lZ  +`  =  -  �9  7`     
     �@     �T �Z  Uu Tt 1�_  u  ��@     T Uu 1_  u   6zL  z@�@     Q      �\  ;vec z!�  i   ]   �  {!Q)  �   �   m�  }7
  `!  X!  Lv ~�  �X?�@     3       F[  �� �k  �!  �!   `  ��@       `9  ��[  +`  �!  �!  `9  7`  �"  �"    `  ��@      �9  ��[  +`  %#  #  �9  7`  �#  �#    ��@     �T �[  Uu Tt 1�_  u  ��@     �S Uu Q�T1�_  u   IdD  i1\  `vec i�  �  jQ)   "I  TQ)  �@     ?       ��\  ;dx Tt
  K$  E$  ;dy Ut
  �$  �$  Lv W�  �h�@     �T �\  Uu Tt 1�_  u  �@     T Uu 1_  u   Hb  Ft
  `�@     ~       ��]  �  FQ)  �$  �$  Lv H�  �hN ��@       ��@     K       M�]  /N C%  =%   $N %��@     K       :N �%  �%  EN &  &  PN 9&  1&  [N �&  �&  fN �&  �&    ��@     �S Uu Tt Q�U1�_  u   :b  8t
  @�@            �j^  �  8Q)  �&  �&  Lv :�  �h<\  G�@       G�@            =#\  O'  I'  \  �'  �'  O�@     D] Uw T�U   GJ  *t
   �@            �
_  �  *Q)  �'  �'  Lv ,�  �h<\  '�@       '�@            /#\  (  (  \  f(  d(  /�@     D] Uw T�U   a�p  �p_  Avec �(�  (I  �Q)  *i �7
  *x �t
  *y �t
  (�S  �t
  *b �#t
  (V  �p_   ])  a-s  ��_  Avec �&�  "I  �&Q)  *i �7
  *x �t
  *y �t
  (�S  �t
  *b �#t
  (V  �p_   Z$c  �7
  `  Avec � �  *x ��  *y ��  (m�  �7
   Zt  =t
  B`  Aval = t
  *s ?7
   dd  ��
  @�@     �      ��a  ^�  �0p  �(  �(  �k �0�a  &)  )  HC  �0a   �)  �)  �U ��
  M*  =*  �N  ��	  +  �*  O�  ��  �+  �+  ,�  [��@     &�8  na  <v �[
  �-  �-  "s  �7
  j.  Z.  p ��  #/  /  &�8  Ya  len �C
  �/  �/   4�@     nh  Uv   <Ch  ��@      ��@     :       ^Qh  Q0  O0  9�m ��@     #       _h  v0  t0  4T  ��@       09  VT  �0  �0  T  �0  �0      _H  �f  �[
  ��@     |       ��b  ^�  �%p  �0  �0  �U �%�R  X1  L1  Mi  ��b  �\p ��  �1  �1  �Y  �[
  ~2  x2  ,WD  ��@     ��@     Us Q�\R4  /�	  �b  0-    �[  x[
  `�@     |       �oc  ^�  x#p  �2  �2  �U y#�R  <3  03  Mi  {�b  �\p |�  �3  �3  �Y  }[
  b4  \4  ,WD  ���@     ��@     Us Q�\R4  �=  K[
  Щ@     �       �!d  ^�  K%p  �4  �4  �U L%�R   5  5  Mi  N!d  �]p O�  �5  �5  �Y  P[
  F6  @6  ,WD  m@�@     �@     Us Q�]R3  /�	  1d  0-    �G  &
  @�@     �       ��d  ^�  &p  �6  �6  �U &�R  7  �6  Mi  !�d  �^p "�  �7  �7  �Y  #&
  *8  $8  ,WD  @��@     u�@     Us Q�^R2  /�	  �d  0-    Hg  �&
  ��@     �       ��e  ^�  �$p  }8  u8  �U �$�R  �8  �8  Mi  ��d  �^p ��  |9  p9  �Y  �&
  :  :  ,WD  �@     ��@     Us Q�^R2  �k  ��	   �@            �4f  ^�  �"p  e:  Y:  �U �"�R  �:  �:  �Y  ��	  �;  �;  ,WD  �6�@     0�@     Us Q�_R1  �s  �[
  �@            ��f  ^�  �$p  Up ��  �;  �;  �Y  �[
  �;  �;   �]  �[
  ��@            ��f  ^�  �"p  Up ��  8<  2<  �Y  �[
  �<  �<   FI  �[
  ��@     .       �Eg  ^�  �$p  Up ��  �<  �<  �Y  �[
  =  =   �c  �&
  `�@     (       ��g  ^�  �%p  Up ��  P=  J=  �Y  �&
  �=  �=   KS  p&
  0�@     '       ��g  ^�  p#p  Up r�  �=  �=  �Y  s&
  +>  '>   �X  `�	  �@            �Ch  ^�  `!p  U�Y  b�	  d>  b>   I�a  >nh  ^�  >#p  >ڰ  O�    )@G  ��
  P�@     1      ��i  ^�  �$p  �>  �>  /� �$[
  E?  1?  �U ��
  (@  @  Qu  �[
  �@  �@  ,�  8>�@      5  ڰ  ��  A  A  �V  {�@      p5  {i  �V  ?A  9A  �V  �A  �A   �V  p5  �V  B  �A  �V  nB  dB  ��@     U| Tv    T  ��@      ��@            	�i  T  �B  �B   T  Ģ@     U|   8��@     �i  Us Rv  	�@     Us Q0R0   �!`  � �@     +       ��j  ^�  �&p  	C  C  �^  �&�J  HC  BC  %0�@            ڰ  ��  �C  �C  $T  3�@       �4  �T  �C  �C  T  �C  �C     )]>  ��
  ��@     4       �(k  ^�  �&p  5D  /D  /� �&[
  �D  �D  �^  �&�J  �D  �D  �U ��
  E  E  ��@     nh  Us T�T  )�h  �[
  ��@     h       ��k  ^�  �!p  =E  5E  _| �!�  �E  �E  /� �![
  <F  0F  Qu  �[
  �F  �F  e�  ���@     8�@     �k  Us Q�TR�Q �@     $| U�TQv   )�^  w�
   �@     }       ��l  ^�  w p  �G  �G  Bpos x [
  H  H  _| y �  vH  nH  /� z [
  �H  �H  �U |�
  ZI  TI  Qu  }[
  �I  �I  8K�@     �l  Uv Ts Q�QR}  ��@     $| U�QQ|   J�D  n�
  �l  "^�  np  "_| o�  "/� p[
   J�Z  g[
  m  "^�  gp   Jw  \�
  Cm  "^�  \p  "d�  ]O
   JM  9�
  ym  "^�  9p  Apos :[
  (�U <�
   _~l  1�m  "^�  1p   _)p  #�m  "^�  #)p  "Ǟ  $)�	  "ֳ  %)[
   )pg  `�
  ��@     c      ��o  ��  `)[  �I  �I  CB  a)C
  OJ  KJ  eX  b)�o  �J  �J  (�U d�
  T  �H  iO8  �J  �J  PT  �, r�3  ]K  YK  �T  ڰ  y�  �K  �K  ^�  zp  �K  �K  7Cm  ��@       �T  ~�n  `m  �K  �K  Tm  2L  ,L  �T  lm  �L  {L  ��@     U} T Q0R0   7�l  ��@        U  Ro  �l  �L  �L  �l  �L  �L  �l  #M  M  ��@     �k  U} T   NT  ��@      ��@            ��o  T  [M  YM  T  �M  M  ��@     U|   ��@     �U  U| T1Q0X0Y��     0O  );^  -�
  P�@     q      ��q  ��  -#[  �M  �M  Bidx .#C
  N  N  Y  /#�q  SN  KN  �U 1�
  �N  �N  �R  �H  6O8  �N  �N  0S  �, ;�3  FO  BO  `S  ڰ  A�  ~O  |O  ^�  Bp  �O  �O  7Cm  ,�@       �S  Fq  `m  �O  �O  Tm  P  P  �S  lm  jP  dP  >�@     U} T Q0R0   7�l  `�@       �S  Glq  �l  �P  �P  �l  �P  �P  �l  Q  Q  e�@     �k  U} T   NT  ��@      ��@            I�q  T  =Q  ;Q  T  cQ  aQ  ��@     U|   �@     �U  U| T1Q0X0Y��     �N  )�C  $C
  �@            �"r  C��  $$[  U D,h  f�   ��@     �       ��s  ڰ  f(�  �Q  �Q  �B  g(<  R  R  �e  h(<  �R  �R  �^  j�   $S  S  tmp k<  �S  �S  �d  l<  �S  �S  Yk  mG   2T  0T  �U n�
  �Lյ@     |  s  Uv  �@     | s  U|  �@     �V  6s  Us Q�L 
�@     :| Ts  Uv T/ +�@     F| ys  Us T�TQ~ <�@     R| �s  Us T|  G�@     R| Us Tv   DQV  L�
  0�@     �       �v  �-  L:`  ^T  ZT  9h  M:�   �T  �T  �=  N:h2  �T  �T  �@  PK  ��qK  Qp  ��i@  R�   lU  jU  �U S�
  �U  �U  �  b�@       �:  \�t  V�  V  	V  I�  wV  sV  <�  �V  �V  /�  �V  �V  "�  5W  1W  �:  c�  uW  qW  t�@     �m T Qv 1'v  �U1Av  �T   P" {�@      {�@     "       _�u  k" �W  �W  ^" �W  �W  9�c ��@            y" X   X  ym  ��@      ;  
�u  �m  'X  %X  ��@     Uv   <T  ��@      ��@            	T  LX  JX  T  qX  oX  ��@     U| Tv     W�@     �" U�UT��Q��  =�@  
�
  �v  �-  
,`  ^�  ,p  Qa  ,�   �  ,k  �=  ,h2  4N  k  �U �
  �;  k  �s  &
  'i S   �d  k  R]  k  �D  (k  �d  x   DjU  ��
  ��@     �       �Lx  �-  �-`  �X  �X  ^�  �-p  DY  @Y  Qa  �-�   �Y  }Y  ?  �-�I  �Y  �Y  �=  �-h2  �Z  {Z  �b  ��   5[  '[  �U ��
  �[  �[  ڰ  ��  $\  \  T  �@      �@            �w  T  o\  m\  T  �\  �\  �@     U| Ts   �@     "r  +x  U| T�QQ	�F      ��@     �s  Uv Ts Q~   D C  ��
  `�@     �       ��y  �-  �+`  �\  �\  ^�  �+p  g]  c]  Qa  �+�   �]  �]  ?  �+�I   ^  �]  �=  �+h2  �^  �^  �b  ��   X_  J_  �U ��
  �_  �_  ڰ  ��  G`  A`  T  ��@      ��@            �oy  T  �`  �`  T  �`  �`  ��@     U| Ts   ��@     "r  �y  U| T�QQ	�F      ��@     �s  Uv Ts Q~   D�E  ��
  ��@     D       ��z  �-  �(`  �`  �`  ^�  �(p  a  a  Qa  �(�   Za  Ta  ?  �(�I  �a  �a  �=  �(h2  /b  %b  �b  ��   �b  �b  ڰ  ��  c  c  ��@     "r  T�QQ	�F       D�[  ��
  ж@     D       �n{  �-  �#`  5c  1c  ^�  �#p  rc  nc  Qa  �#�   �c  �c  ?  �#�I  d  �c  �=  �#h2  �d  |d  �b  ��   e  �d  ڰ  ��  de  be  �@     "r  T�QQ	��F       D�q  r�
  ��@     �       ��|  �-  r,`  �e  �e  ^�  s,p  �e  �e  Qa  t,�   4f  ,f  ?  u,�I  �f  �f  �=  v,h2  g  �f  �U {�
  ���b  |�   gg  ag  ڰ  }�  �g  �g  (e  ~O
  �g  �g  ׷@     | b|  U|  �@     �V  �|  TsQ�� �@     $| T| Qs   D&Z  N�
   �@     �       ��}  �-  N-`  .h  &h  ^�  O-p  �h  �h  Qa  P-�   �h  �h  ?  Q-�I  9i  1i  �=  R-h2  �i  �i  �U W�
  ���b  X�   j  �i  ڰ  Y�  Qj  Oj  (e  ZO
  {j  uj  G�@     | �}  U|  c�@     �V  �}  TsQ�� ��@     $| T| Qs   D�Y  0�
   �@     �       �:  �-  00`  �j  �j  ^�  10p  tk  pk  Qa  20�   �k  �k  ?  30�I  l  �k  �=  40h2  �l  �l  �b  6�   em  Wm  �U 7�
  n  �m  ڰ  8�  Tn  Nn  T  F�@      F�@            G�~  T  �n  �n  T  �n  �n  Q�@     U| Ts   (�@     "r    U| T�QQ	�F      >�@     �s  Uv Ts Q~   D�I  �
  `�@     &       ��  �-  +`  �n  �n  ^�  +p  ,o  $o  Qa  +�   �o  �o  ?  +�I  �o  �o  �=  +h2  5p  /p  ��   k    .|�@     �m U�TT  Q�X1'v  �U1Av  �Q  ="T  �
  q�  �-  +`  ^�  +p  Qa  +�   ?  +�I  �=  +h2  �  
k   =�L  ��	  ��  �-  �.`  �n  �.C
   =vn  �LJ  ˀ  �-  �6`  �n  �6C
   6�H  � �@     �       ��  �-  �!`  �p  �p  ^�  �!p  �p  �p  p  �!�   )q  %q  �b  �!�I  eq  aq  �f  �!h2  �q  �q  �>  �!�R  �q  �q  i �7
  Lr  Br  Cm  P�@      P4  ��  `m  �r  �r  Tm   s  �r  P4  lm  :s  6s  d�@     U~ T0Q0R0   ��@     U T~ Q��RvxXs 3$} "  )�X  ��
  ��@     x      �P�  �-  �+`  zs  rs  ^�  �+p  �s  �s  �  �+O
  Qt  Ct  Zv  �+O
  �t  �t  Btag �+O
  gu  Wu  �s  �+�	   v  v  C�f  �+P�  � C/� �+h2  �F�U ��
  ��#i �S   �v  �v  #j �S   �v  �v  #cnt �S   �w  �w  �^  �S   +x  %x  [  �O
  �x  �x  �O  �!O
  y  y  ڰ  ��  �y  y  �S  �O
  z  �y  �m  �h2  lz  bz  #ref �V�  �z  �z  ,�  BX�@     7Cm  ��@      �F  ��  `m  �{  �{  Tm  �{  �{  �F  lm  =|  9|  ��@     Us T Q0R0   Cm  �@      0G   ��  `m  y|  u|  Tm  �|  �|  0G  lm  �|  �|   �@     Us T Q0R0   m  1�@      pG  �  6m  )}  %}  *m  e}  a}  $Cm  9�@       �G  b`m  �}  �}  Tm  �}  �}  �G  lm  A~  9~  ��@     Us T~ Q0R0    m  ��@      �G  ��  6m  �~  �~  *m  �~  �~  $Cm  ��@        H  b`m      Tm  l  f   H  lm  �  �  ��@     Us T~ Q0R0    T  X�@      X�@            C	�  T  	�  �  T  .�  ,�  k�@     U��T}   �@     �d  .�  Us T�� M�@     �d  M�  Us T�� g�@     �d  l�  Us T�� ��@     �b  ��  Us T�� R�@     �U  ��  U��T@Q0X0Y�� ��@     �b  چ  Us T�� %�@     �d  ��  Us T�� ��@     �U  )�  U��T8Q0X0Y�� #�@     ^| U} Q@R	@I@       h2  �I  V�;  �S   @I@            ���  Oa �-V�  UOb �-V�  T )�V  3�
  �@     $      ���  �-  3*`  [�  S�  ^�  4*p  ̀  ��  �I  5*O
  ��  ~�  �  6*h2  <�  *�  Zv  7*h2  �   �  �U 9�
  ؃  փ  FuR :��  ��F(F  :��  �@�`  ;O
  �  ��  �@  ;O
  y�  u�  z<  ;&O
  ��  ��  OM  <S   �  �  <v  <S   �  �  #i <(S   L�  H�  �q  =O
  ��  ��  7Cm  �@      06  BB�  `m  ��  ��  Tm  �   �  06  lm  S�  O�  A�@     Us T| Q0R0   7�l  f�@      p6  F��  �l  ��  ��  �l  ��  ��  �l  �  �  k�@     �k  Us T| Q��R@  7Cm  ��@      �6  ��  `m  ,�  (�  Tm  f�  b�  �6  lm  ��  ��  ��@     Us T| Q0R0   7�l  �@      �6  �y�  �l  ڇ  ؇  �l  �  ��  �l  >�  :�  �@     �k  Us T| Q�@R@  7m  3�@       7  ��  6m  x�  t�  *m  ��  ��  $Cm  ;�@       P7  b`m  �  �  Tm  (�  $�  P7  lm  b�  ^�  T�@     Us Tv Q0R0    7Cm  ��@       �7  �z�  `m  ��  ��  Tm  ؉  ԉ  �7  lm  �  �  ��@     Us T| Q0R0   t�@     �d  Us T��  /�  ��  0-    )�Q  ��
  `�@     �       �ڌ  ϖ �!1  N�  J�  �1  �!<  ��  ��  C<v �!a   Qo�U ��
   K ��J  ��  ��  ?О@     @       ]�  iO  ��C  �  �  #val ��C  �  �   ?��@            ��  �q  C
  2�  0�  val �?  W�  U�   %��@            �'  �	  |�  z�  val ڌ  ��  ��    �	  )�T  '�
  ��@     �      ��  ϖ '!1  Ћ  ċ  �1  (!<  Z�  X�  <v )!r  ��  }�  �h  *!�	  *�  &�  o�U ,�
   K -�J  o�  c�  ?ԛ@     !      Ŏ  iO  6�C  ��  ��  #x1 77
  J�  H�  #y1 77
  q�  m�  #x2 77
  ��  ��  #y2 77
  ю  ͎  #x3 7 7
  �  �  #y3 7$7
  G�  C�  #x4 7(7
  ��  ~�  #y4 7,7
  ��  ��  [dp :�J  ��%�@     m       #s ?<  �  ߏ  [ep @�   ��*i AS   �@     j| ��  U~ T��Q: ,�@     j| U~ T��Q:   ?,�@     &       �  #s ~<  �  �   & 4  �  �q  ��?  E�  A�   ? �@             e�  #s �<  }�  {�  #nsd �@   ��  ��  /�@     j| U~ T0Q:  ?ԝ@            ��  �'  �ڌ  ǐ  Ő   �3  ��  �k  �  �  %@�@            #s �<  M�  K�  O�@     j| U~ T0Q:    �_  	�H  ��@     �      ���  Mj  	,�J  v�  p�  �'  	-  ��<B  	7
  Ƒ    {A  	7
  �  �  N5  	�  B�  @�  �D  	�  o�  e�  _  	�  ��  ��  c 	7
  :�  8�  n 	7
  `�  ^�  ��  	7
  ��  ��  �r  	�  ٓ  ӓ  ?��@     �       �  ��  	47
  %�  #�   4?�  ��@      �.  	"Z�  J�  H�  M�  q�  m�  �.  g�  t�  ��  ��   �@     �W U{ Tt     %O  	��
  `�@     /      ���  Mj  	�'�J  ��  ��  �t  	�'�  +�  %�  M  	�'�  ��  w�  N5  	��  �  	�  c 	�7
  ��  ��  ��  	�7
  �  ֖  ��  	�7
  g�  e�  �l  	��H  ��  ��  & /  l�  in 	��  ��  �  Lout 	��  ���`  	��  G�  ;�  m�  	�#�  �  ��  L 	�t
  J�  @�  � 	�t
    ��  �`  	�t
  $�   �  l 	�-t
  a�  ]�  q 	�0t
  ��  ��  d 	�3t
  X�  J�  i 	�7
  ��  �  j 	�7
  [�  Y�  k 	�7
  ��  ~�  sN �@      �/  	�ɓ  �N ՝  ӝ   �N $ES �@       0  �`S ��  ��   VS  0  jS #�  �  vS f�  d�     sN &�@      p0  	�*@�  �N ��  ��   �N $ES &�@      �0  �`S ��  ��   VS �0  jS ݞ  ٞ  vS  �  �     sN �@       1  	�ǔ  �N ]�  [�  �N ��  ��  $ES �@      �1  �`S ��  ��  VS П  Ο  �1  jS ��  ��  vS <�  8�     sN �@      @2  	�/>�  �N y�  w�  �N ��  ��  $ES �@      �2  �`S à  ��  VS �  �   3  jS vS    sN L�@      `3  	�ŕ  �N �  �  �N 3�  1�  $ES L�@      �3  �`S Z�  X�  VS ��  ~�  �3  jS ��  ��  vS �  �     ��@     b> ݕ  Uu  B�@     dO ��  T��Q�� ��@     dO )�  U��~T��Q�� >�@     dO P�  U��~T} Qw  a�@     dO T} Qw   @     �  U��  �a  	�
  ��@            ���  Mj  	%�J  +�  '�  �t  	�%�  h�  d�  .��@     ��  U�UT�TQ�T  ICA  	�7�  Mj  	�,7�  �3  	�,|  'vec 	��  ��  	��   �  I�C  	�~�  ��  	�*�  �3  	�*|  'xz 	��  'yz 	��    q  	��
   �@     g       �m�  �-  	�,`  ��  ��  Mj  	�,�J  ��  �  Ue  	�,l  O�  E�  \  	�y  ��4m�  -�@      �.  	���  ɣ  ã  ��  �  �  �  m�  g�  �.  ��  ��  ��  ͘  ?�@     �X U�UT�TQw     W?u  	R�
  ۘ  �-  	R)`  Mj  	S)�J  \  	T)ۘ  �U 	V�
  eo  	W�  �K  	X�  �'  	Y-   y  6�S  	��@     �       ��  Mj  	$�J  Un 	&
  ��  ��  ��  	7
  '�  �  ��  	7
  ��  ��  &�.  ��  p 	&�  ��  ��  q 	'�  �  ��  uL  	(�  P�  L�   %\�@     .       p 	7�   ��  ��  q 	8�   �  �  %p�@            uL  	=�   3�  1�     I�a  	�?�  Mj  	�,7�  C"  	�,�  �  	�,�  'n 	 &
  'vec 	�   I@  	�К  Mj  	�+7�  N  	�+�  
  	��  �!  	��  �   	��  H  	��  >'vec 	��  ��  	��  >'x 	��  'y 	��     s  	��
  ��@     �       �%�  �-  	�!`  \�  V�  Mj  	�!�J  ��  ��  ڰ  	��  �  �  T  �@       �@            	���  T  K�  I�  T  p�  n�  ��@     Uv   T  �@      �@            	�֛  T  ��  ��  T  ��  ��  �@     Uv   <T  �@      �@            	�T  ߨ  ݨ  T  �  �  *�@     Uv    �v  	��
  �@     �       ���  �; 	�'7�  1�  '�  .  	�'�J  ��  ��  �H  	�7
  M�  I�  G��@     $| G��@     $| G��@     $|  �v  	V�
  ��@     f       �g�  Mj  	V"�J  ��  ��  �Bad 	{�@     P.  0�  	Z7
  ʪ  ƪ     	[7
  �  �  �J  	\7
  C�  =�  end 	\7
  ��  ��  n 	]7
  ߫  ۫    �Y  	&�
   �@     F      �Ҟ  �-  	& `  #�  �  �E  	' C
  ��  ��  �n  	( 7
  Z�  N�  JB  	) �J  �  ߭  �U 	+�
  ��ڰ  	,�  x�  p�  ,WD  	K��@     ��@     �U  I�  U} T@Q0R X0Y�� ��@     �U  }�  U} T1Q0R X0Y�� ��@     К  ��  Uv Ts  "�@     �U  U} T2Q0R|  $ &X0Y��  )�c  	,�
  ��@           ��  Mj  	,2�J  �  ծ  ei  	-2�  ܯ  ȯ  �  	.2a   ˰  ��  w  	3�  ��  ��  FnX  	4�  ��~FJ  	5�  ��c 	7�  ²  ��  ��  	8�  ٳ  ͳ  �   	9�   }�  ]�  �U 	;�
  �  ͵  #n 	=7
  ��  ��  ��  	>C
  �  y�  #tag 	?7
  ݷ  ɷ  m�  	A7
  �  ��  �� 	B�  u�  _�  @M�  	@�  	e?j  	�	�@     ,�l  	��@     �,  ��  	Q7
  b�  V�  &p-  ��  [vec 	��  ���@     U��T��~  &.  �  [vec 	��  ��F�R  	��  ��8z�@     �  U~ T��Q��~ >�@     U��~T��Q��~  &�-  ��  F<  	��  ��F"<  	��  ��&�-  l�  [vec 	��  ��4�@     U��T��Q��R��~  ��@     U��T��Q��R��~  8��@     ��  U��T��~ 8��@     Ρ  U��T��~ ��@     U~ T��Q��~   �  W�g  ��	  c�  ��  �0[  Oq �0C
  �j  �0�?  �e  �0�?  ��  �0�B  �H  �O8  �i  �*F   �f  i�
  ��@     �       �?�  ȩ  i'�  U]d  j'C
  &�   �  =  k'�C  x�  r�  o  l'�?  ʻ  Ļ  $D  m'�C  X0B  n'�C  Y�c  o'?�  � �U q�
  �  �  %��@     P       7B  y�  l�  h�    �
  �X  J$  `�@     C       ��  �-  J,`  ��  ��  �Y  L$  
�  �  �,  ϖ Q1  W�  U�  ?x�@            ��  �b  V$-N  |�  z�  ��@     �  T	��F     Q0  s�@     ��  U�UT	��F        6RW  <0�@     +       �h�  �-  <)`  UjL  =)C
  T�=  >)�  Q �+  ��
  ��@     L      �ܥ  �-  � `  ��  ��  ڰ  ��  4�  .�  @�  4&p,  m�  m �C
  ��  ��  n �C
  ��  ��  �?  �ܥ  ��%d�@     G       ϖ �1  *�  &�  �5  �<  b�  `�  �!   �  }�@     v| ^�  T}  G��@     f�    T  �@      �@            2ǥ  T  ��  ��  T  ��  ��  ��@     U��T|   ��@      �  U|   /<  �  0-    6pZ  ���@     :       ���  �-  �$`  USs  �$�C  T�E  �$�C  Qa  �$�C  R�3  �7
  ؿ  ҿ  [0  �7
  )�  #�  �/  �7
  z�  t�   |&  ��
  `�@     f       ��  ڰ  � �  ��  ��  �-  � �  4�  ,�  �-  �`  ��  ��  �U ��
  �\��@     �V  Us T
�Q�\  `  n  ��
  ��@            �T�  �-  �%`  U B/  c�
  `�@            � �  �-  c-`  ��  ��  �5  d-�  :�  6�  �1  e-�  w�  s�  <v f-�  ��  ��  .q�@     X�  U�UT�TQ�QR�RX1Y1  �;  O�
  P�@            ���  �-  O&`  ��  ��  �5  P&�  .�  *�  �1  Q&�  k�  g�  <v R&a   ��  ��  .[�@     X�  U�UT�TQ�QR�RX0Y0  E  >�
  @�@            �X�  �-  >&`  ��  ��  �5  ?&�  "�  �  �1  @&�  _�  [�  <v A&r  ��  ��  .N�@     X�  U�UT�TQ�QR�RX1Y0  =h  ��
  ��  �-  �%`  �5  �%�  �1  �%�  <v �%a   `set �%�	  �h  �%�	  'cur ���  ��  ���  ��  ��  �b  ��K  �R  ��	   1  d�N  ��
  p�@     �      ��  �-  �!`  ��  ��  ϖ �!1  K�  ?�  0*  cur ���  ��  ��  ��  ���  D�  6�  4��  ��@      �*  ���  ��  ��  �*  ��  F�  @�  ĳ  ��  ��  ѳ  ��  ��  T  +�@      +�@     
       �$�  T  /�  -�  T  T�  R�  5�@     U} Ts   � P�@      P�@             �׫  � y�  w�  4gO  T�@        +  ��O  ��  ��  �O  ��  ��  �O  ��  ��  uO  �  �   +  �O  j�@     �_ Us T	pl@     Rs     ��  0+  ��  �  k�  g�  0+  &�  ��  ��  3�  ��  ��  @�  �  �  �Q  p�@      p�@            T��  �Q  �  }�  �Q  ��  ��  %p�@            �Q  ��  ��    HM�  `+  N�  ��  ��  �P  ��@      �+  `��  �P  +�  )�  �P  P�  N�  �+  Q  Q  ��@     ^_ Uu Tv    T  ��@      ��@            a;�   T   T  ��@     U   4ߺ  ��@      �+  c�  z�  v�  �+  ��  4O�  ��@      ,  {�  ��  ��  n�  ��  ��  a�  4�  0�  ,  ��  n�  j�  ��  ��  ��  M��  �@     H�g @,  ��  ��  ��          +�@     Us      W�b  ��
  u�  ϖ �'1  �E  �'<  V� �'�	  �Y  ��
  >�-  �`  'cur ���  ��  ���    �?  �r  ��@     '       ���  �-  �)`  �  �  �j  �)<  [�  W�  ϖ �1  ��  ��  ��@     ��  U�UT�T  $i  d1  0�@     p       ���  �-  d`  ��  ��  �5  e<  �  �  P�Y  g1   cur h��  _�  ]�  ��  i��  ��  ��  |�@     v| T|   d�1  ��
  @�@     �      ���  �-  �*`  ��  ��  Oe �*��  [�  M�  �U ��
  ��ڰ  ��  ��  ��  ϖ �1  Z�  D�  nn �C
  C�  ?�  ,�  M��@     ,WD  P��@     ?D�@            w�  K =}  }�  {�   ?��@     "       ��  eo  S�  ��  ��   ]�  ��@      C  1ز  o�  ��  ��  C  |�  �  �  ��  i�  c�  5��  ����  ��  ��  M��  ��@     M��  u�@     pº  PC  j�  ú  o�  k�  к  ��  ��  pQ  *�@      �C  8��  �Q  ��  ��  ~Q  !�  �  �C  �Q  9�@     '_ Uu T    ߺ  9�@      �C  :R�  �  ^�  Z�  �C  ��  4O�  9�@       D  {�  ��  ��  n�  ��  ��  a�  �  �   D  ��  R�  N�  ��  ��  ��  M��  j�@     H�g 0D  ��  ��  ��       �@     U| Ts�   T  u�@      `D  ?��  T  �  ��  T  h�  b�  �@     U| T   ��@     �V  U| THQ��   T  ��@      ��@     
       \0�  T  ��  ��  T  ��  ��  ��@     U} Ts   ��@     v| H�  T|  ��@      �  f�  Uv T  �@     �V  ��  U} Q�� ^�@     Us   �  T�R  �߳  ϖ �1  ڰ  ��  Oe ��(  �-  �`   ]e  ��
  �@     6       �^�  �  �$�  �  ��  �L  �$O  �  w�  �-  �`  ��  ��  .6�@     ^�  T�UQ�T  �t  ��
  �@           ��  �-  �-`  �  �  �  �-�  ��  ��  �L  �-O  ��  ��  �U ��
  h�  R�  ��  �[  O�  M�  eo  ��  {�  s�  &`<  x�  ��  ��  ��Oq �C
  ��  ��  �]  ��	  �  �  x �C
  ���e  �C
  ��&�<  +�  �H  �O8  �i  �*F  R�  L�  &�<  ݵ  �1  �k  ��  ��  8��@     ȵ  U} Qs  <�@     � U}   �@     ��  �  U} T~ Q��R��X�� GL�@     � G�@     �  ��@     ��  ^�  U} T~ Q��R��X�� ��@     � U} T0  �;  �K  	�  ��  ��  O�  ,�@      ,�@     D       5�  {�  p�  n�  n�  ��  ��  a�  ��  ��  %,�@     D       ��  ��  ��  ��  	�  �  \��  9�g =�@     %       ��  3�  -�     O�  ��@       ��@     ?       #̷  {�  �  }�  n�  ��  ��  a�  ��  ��  %��@     ?       ��  ��  ��  ��  �  �  \��  H�g 0<  ��  B�  <�     �@     Ts Q| R0   U  w�
  ��@           �"�  �-  w#`  ��  ��  eo  x#�  �  �  �[  y#C
  ��  ��  �Y  z#E  _�  W�  �K  |�  ��  ��  �U }�
  �  ��  � c  ��  ��  ,�  ���@     �Q  �@       �U  ���  �Q  ��  ��  �Q  �  �  �U  �Q  8�  6�    $�@     �P  �  Tt  f�@     Uv   �U  k�  ��@     6       ��  �-  k%`  U��  l%�  T<O�  ��@      ��@     4       p{�  _�  [�  n�  ��  ��  a�  ��  ��  %��@     4       ��  �  �  ��  I�  E�  M��  $�@     9�g �@            ��  ��  ��      Tj  G]�  ϖ G"1  �-  I`  ڰ  J�  �K  K�  >�� W�    =^o  �
  ߺ  ϖ 1  �-  `  ڰ  �  �U �
  �K  �  @�  A@WD  =>�� #�  Oe $�(    T�q  �  �-  (`  eo  �   =4c  ��  O�  �  �+�  ��  �[  �-   `  �Y  �   Ww  ��  û  �-  �(`  ��  �(�  �K  �(û  'cur ��  �Y  ��  ,�  �م@     >eo  ��    �  no  ��
  @�@     6       ��  ֳ  �/  U��  �[  ��  ��   �M  �O
   �@     ^       ��  �� �#�  V�  L�  �b  ��M  ��  ��  ��  �[  ��  ��  �  �AM  �`?5�@            ڼ  ϖ �1  *�  (�  6e  ��
  Q�  M�  O�@     T	��F       \�@     Us Tw   `T  �[
  ��@     c       �Ž  �� �(�  ��  ��  �b  ��M  �  �  ��  �[  E�  A�  �  �AM  �`&0'  ��  ϖ �1  ~�  |�  6e  ��
  ��  ��  �@     T	��F       �@     Us Tw   �l  h�
   �@     �       �վ  ��  h"[  ��  ��  �f  i"C
  |�  p�  ;tag j"�2  �  �  ��  k"�2  ��  ��  �b  mrL  0�  ,�  �  n[
  �H&�&  ��  ϖ v1  j�  f�  6e  v�
  ��  ��  b�@     T	w�F       z�@     Us Tv Q| R�HX}   �O  Q�
  ��@     �       ��  ��  Q"[  �  �  ;tag R"[
  ��  ��  �  S"O
  ��  ��  _| T"�  P�  @�  ��  U"�2  �  ��  �b  WrL  ��  ��  &�&  ��  ϖ ]1  ��  ��  6e  ]�
  8�  0�  π@     T	w�F       :��@     U�UT�TQ�QR�RX�X  [?  <a    �@     c       ���  ��  <#[  ��  ��  ;tag =#�1  M�  ?�  P�B ?a    �b  @rL  ��  ��  &P&  ��  ϖ E1  $�  "�  6e  E�
  M�  G�  S�@     T	w�F       :i�@     U�UT�T  oC  <  �@     �       ���  ��  $[  ��  ��  P�Y  !<   ,�  4�@     `%  �b  )�L  p�  j�  &�%  ��  svc ,�
  ��  ��   &  ϖ ,1  8�  4�  6e  ,�
  v�  n�  �@     T	b�F        :�@     U�U   �]  ��
  �~@     �       ���  ��  �"[  ��  ��  x �"C
  ��  ��  _| �"�
  q�  e�  �H  �"C
  �  ��  �U ��
  P�b   M  ��  ��  &�$  ��  svc �
  ��  ��  %0@     "       ϖ 1  H�  D�  6e  �
  ��  ~�  R@     T	W�F        :�~@     U�UT�T  S  �C
  �}@     �       ���  ��  �([  ��  ��  { �(�  ��  ��  P�Y  �C
   �#  �b  �M  f�  `�  &P$  ��  svc ��
  ��  ��  �$  ϖ �1  �  �  6e  ��
  U�  O�  W~@     T	W�F        :~@     U�UT�T   �m  ��'  ��@     S       ���  ��  �([  ��  ��  �I  �([
  @�  4�  P�Y  ��'   p)  �� ��  ��  ��  &�)  ��  =E  �m&  �  �  ڰ  ��  +�  '�  :�@     Q�T  ��@     �f 1Q s    Pt  ��'  ��@     S       �l�  ��  �([  o�  c�  �_ �([
  �  ��  P�Y  ��'   �(  �� ��  ��  ��  &0)  T�  =E  �m&  ��  ��  ڰ  ��  ��  ��  :��@     Q�T  ��@     �f 1Q s    q�A  ~�'  @�@     ;       ��  ��  ~)[  2�  &�  P�Y  ��'   �(  �� ��  ��  ��  &�(   �  =E  �m&  ��  ��  ڰ  ��  �  �   U�@     �f 1Q s    �b  S7
  ��@     I       ���  ��  S.[  [�  U�  �_ T.[
  ��  ��  �I  U.[
  G�  ;�  ��Y  W7
  �'  �� \�  ��  ��  &@(  ��  =E  am&    	  :)�@     T�TQ�Q  �@     �f 1Q �U   qlI  %C
  ��@     g       ���  ��  %*[  8  .  �_ &*[
  �  �  �I  '*[
  6 , P�Y  )C
   p'  �� 0�  � � �n  1m&  � � &�'  ��  =E  6m&  T R  ��@     �f 1Q s    8[  ��
   }@     �       �L�  ��  �&[  U�b  �&C
  y w �  �&E  � � �U ��
  � � ,�  �}@      �n  �[
  |@     i       �&�  ��  �[    �_ �[
  � y \D  ��?  � � �Y  �[
  c _ J�  �C
  � � %6|@     *       �* �}  �\I_ �m&     O|@     Us T�\   PF  �[
  �|@     u       �3�  ��  � [  + % \D  � �?  } w �Y  �[
  � � J�  �C
  �\3�  �|@      �#  ��  R�  3 / E�  o k �#  _�  � � 9�f �|@            m�    �|@     T0    �|@     L�  Us T0Q�\  W�Q  C
  |�  ��   [  �_ � [
  �Y  �C
  >I_ �m&    2n  I�
  ��@     ;      �m�  Oe I�&  < 0 �h  J�
  � � �� K�  6 , �D  Lm�  � � �U N�
  ����  O[  (	 $	 ڰ  P�  b	 ^	 I_ Qm&  �	 �	 ,WD  u��@     ,�  o��@     �  ��@       F  v�  &�  W
 S
  F  3�  �
 �
 @�  �
 �
 M�  �
 �
 T  ��@      PF  ��  T   �
 T  : 8 ��@     Us   ��@     U~    �@     �V  0�  U Q�� 8J�@     L�  U~ T�� r�@     �U  U T8Y��  m&  6o[  ��@     6      ��  I_ m&  k ] �E  ��  [    ڰ   �  Y U �U !�
  �Li "7
  � � j "7
  ) % �E  bF  )�  c _ �  n�@      n�@     &       ?��  &�  � � %n�@     &       3�  � � @�  � � M�  "   T  ��@      ��@     	       ��  T  G E T  l j ��@     Us Tv   ��@     Uv    
�@     �U  T8Y�L    T'E  [�  I_ #m&  Oe �&  ��  [  ڰ  �   �I  �7
  p{@     Q       ���  �� �%�  Ui �7
  � �  �E  ��
  ��@     �       �-�  ��  �[    �� ��  { s cur ��  � � ��  ��  - + ւ@     �  Uv   @R  ��
  �z@     �       ���  ��  �#[  UT �#  V P cur ��  � � ��  ��    fe{@     �  �M  ��
  @z@     �       ���  ��  �$[  P B �' �$t
  � � N  �$7
  � � 6_  �$"  K = �b  ��M  � � P�U ��
   &P#  ��  ϖ �1  $   6e  ��
  b Z |z@     T	O�F       :�z@     U�UT�TQ�QR�R  �A  ?�
  Px@     �      ���  ��  ?[  � � sl  @C
  y i �J  AC
  5 - c  BC
  � � 6_  C�  N @ �U E�
  � � K F}  j d &�"  ��  �j  c�  � � �j  d�  %  dO y@      �"  k0�  �O � � �O � � uO + # �"  �O � � �O �O � � �O E A �O � } �O < 6   4dO Ty@       #  n�O � � �O � � uO P H  #  �O � � �O �O    �O i e �O � � �O _ Y    sN �x@       �!  ^C�  �N � � �N � � $ES �x@      "  �`S     VS =  ;  "  jS g  a  vS �  �     sN �x@      @"  _��  �N A! ?! �N g! e! $ES �x@      �"  �`S �! �! VS �! �! �"  jS �! �! vS 3" /"    �x@     Us T�TQ�QRv   yJ  �
  �w@     i       �v�  ��   [  t" n" �@   C
  �" �" p   C
  1# '# Lreq �  �P@x@     '�  Tw   D<  ��
  Pw@     �       �'�  ��  �![  �# �# N  �!g
  �# �# �I  �!g
  V$ J$ oF  �!C
  % �$ @F  �!C
  �% �% Lreq ��  �P�w@     '�  Tw   �q  ��
  pv@     �       ���  ��  �%[  & & ;req �%  �& �& �U ��
  $' ' Oe ��"  �' �' m �[
  �h��   w@       w@            �L�  ��  �' �' ��  K( G( ��  �( �( ��  �( �( % w@            �  �  �  w@     SW Us T�TRr    8�v@     a�  T�T *w@     ��  y�  Us  Hw@     ��  Us   W6U  n�
  ��  ��  n[  m o7
  �U q�
  Oe r�"   6R   0r@     �      �Z�  ��   ([  ) ) ;req (  �) �) �e  B  �* �* ,	S  U�s@       w 
O
  8+ + h 
O
  g, G, Si  
O
  �- �- j  
,O
  �. �. N Ps@      P  ;�  /N 0 0 $N ?0 ;0 P  :N {0 u0 EN �0 �0 PN 1 1 [N Z1 T1 fN �1 �1   N �s@      �  ?��  /N B2 <2 $N �2 �2 �  :N �2 �2 EN K3 C3 PN �3 �3 [N �3 �3 fN s4 m4   sN �s@       �  Y�  �N �4 �4 �N 5 5 $ES �s@      0  �`S L5 J5 VS q5 o5 �  jS �5 �5 vS �5 �5    sN t@         Z��  �N 66 46  �N $ES t@      �   � `S VS \6 Z6 �   jS �6 �6 vS �6 �6    N �t@      `!  Q/�  /N �6 �6 $N %7 !7 `!  :N a7 [7 EN �7 �7 PN 8  8 [N >8 :8 fN �8 �8   gFt@     �  ,�  Uu Tt  �t@     dO D�  Uz  �t@     dO U{    6f  ��p@     ^      ��  ��  � [  Um � [
  �8 �8 �e � B  A9 59 �d  ��  �9 �9 N q@      �  �D�  /N �: : $N �: �: �  :N 7; 1; EN �; �; PN �; �; [N =< 3< fN = =   N 6q@      �  ���  /N �= �= $N .>  > �  :N �> �> EN h? X? PN 6@ ,@ [N �@ �@ fN �A �A   g^q@     �  ��  Tt  g�q@     �  ��  Tt  ..r@     �  Tt   h�W  ��H@     �       �\�  ��  �2[  U�e �2 B  TsN �H@      `  ���  �N �B �B �N �B �B $ES �H@      �  �`S C C VS =C ;C �  jS oC kC vS �C �C    sN �H@         �Q�  �N �C �C �N D D $ES �H@      `  �`S ED CD VS kD iD `  jS �D �D vS �D �D    sN �H@      �  ���  �N E E �N GE AE $ES �H@      �  �`S �E �E VS �E �E �  jS  F �E vS CF ?F    4sN I@      �  ��N �F ~F �N �F �F $ES I@         �`S G 	G VS 1G /G `  jS cG _G vS �G �G     6mY  �Pp@     �       ���  �e �6��  U� �6�  �G �G ��  ��  9H 3H  �  Wva  g�
  2�  ��  g#[  `req h#  >p  i#�	  �H  j#�2  'i l7
  'w mO
  'h mO
  >�d  ��    �t  7�
   o@     �       ���  ֳ  7/  �H �H �U 9�
  I I K :}  ZI PI ڰ  ;�  �I �I ��  <[  1J 'J �K  =�  �J �J �Q  Oo@      Oo@             N4�  �Q  �J �J �Q  2K ,K %Oo@             �Q  �K �K   �P  to@      P  Q��  �P  �K �K �P  �K �K P  Q  Q  �o@     ^_ Uu Tr    T  �o@      �o@            R��   T   T  �o@     U}   �o@     ] U} Ts Q|   �B  �
�
   �@     6      �`�  ��  �
[  L L �p  �
`�  �L �L �U �
�
  ��ڰ  �
�  
M M K �
}  BM @M Oe �
�"  iM eM ֳ  �
/  �M �M �K  �
�  AN /N �L  �  O  O @�  )T  d�@      d�@            -4�  T  �O �O T  �O �O r�@     Uv T}   T  ��@      ��@            ,��  T  �O �O T  P P ��@     Uv T   pQ  �@      �B  &��  �Q  *P (P ~Q  OP MP �B  �Q  �@     '_ Uu Tt    Y�@     �V  �  Uv Q�� ��@     �V  *�  Uv THQ�� ��@     �V  O�  Uv THQ�� ��@     U}   /  �Z  �
�
  pn@     �       ��  ��  �
[  zP rP �U �
�
  �P �P K �
}  /Q -Q ڰ  �
�  TQ RQ �K  �
�  |Q xQ �Q  �n@      �n@            �
S�  �Q  �Q �Q �Q  �Q �Q %�n@            �Q  R �Q   �P  �n@         �
��  �P  &R $R �P  KR IR    Q  Q  �n@     ^_ Uu Tr    T  �n@      �n@            �
��   T   T  �n@     U|   �n@     � U| Ts Qv   �`  �
�
  Pn@            �I�  ��  �
[  U �N  �
�
  ��@     �       ��  ��  �
$[  xR pR �Y  �
$�  �R �R ^�  �
p  �X�U �
�
  FS >S K �
}  �S �S Oe �
�"  �S �S @�  �
P" �@       �@     6       �
��  k" 2T 0T ^" cT _T 9�c �@     1       y" �T �T ym  !�@      @;  
��  �m  �T �T /�@     U|   <T  ;�@      ;�@     	       	 T  T  �T �T D�@     Us T|     ּ@     �" ��  Ts Q�X ��@     Uv T|   K  �u  }
�
  ��@     6       ���  ��  }
 [  U U +[  ~
 <  eU ]U ��  �
K  ����@     I�  U�UTw   ��L  C	�
   �@     C	      ���  �-  C	/`  �U �U E�  D	/��  NX &X �  E	/O
  �Y �Y �]  F	/��  �Z �Z �@  G	/�	  =[ [ �U I	�
  ��|K J	}  �\ �\ ڰ  K	�  �^ �^ ^�  L	p  ��|��  M	[  ��}�K  N	�  /` ` 7K  O	�	   a �` cur P	��  �a �a ��  Q	��  Db <b ,Ob  �	�@     ,�n  �	�@     ,WD  `
I�@     ,Z  �	��@     ,�  f
��@     & L  �  �[  }	7
  �b �b \  ~	E  �b �b ��@     � U��|T��|Q} R��|  &�L  b�  �[  �	7
  Hc Bc \  �	E  �c �c Cm  �@       M  �	�  `m  �c �c Tm  d d M  lm  wd sd .�@     U��|T0Q0R0   P" �@       �@     1       �	�  k" �d �d ^" �d �d 9�c �@     (       y" e e ym  �@      @M  
��  �m  6e 4e (�@     Us   <T  1�@      1�@     	       	T  [e Ye T  �e ~e :�@     Uv Ts     g�@     � ;�  U T��|Q} R��| a�@     et U��|Q��|R��|  ?e�@     2       ��  ֳ  

/  ��~w�@     ��  T��~  ?��@     �       ��  i $
7
  �e �e `L  �d  )
�  �e �e   &PO  �  �L  D
  f f  pQ  4�@      0L  �	\�  �Q  Af =f ~Q  yf wf 0L  �Q  B�@     '_ Uu Tt    P" ��@      ��@     4       �	6�   k" ^" �f �f 9�c ��@     /       y" �f �f ym  ��@      �L  
��   �m  ��@     Us   <T  ��@      ��@     	       	 T  T  g g ��@     Uv Ts     ��  ��@      pM  �	�  ��  =g )g ��  h h ��  �h �h ��  i i ��  Ei ;i pM  ��  �i �i ��  ��@      ��@     �       	=�  #�  Sj Qj �  zj xj 	�  �j �j ��  �j �j %��@     �       50�  ��~=�  �j �j J�  0k (k W�  �k �k \d�  Cm  ��@      �M  ���  `m  |l zl Tm  �l �l �M  lm  �l �l ��@     Us T0Q0R0   �l  ��@      N  ��  �l  �l �l �l  m m  �l  ��@     �k  Us T0Q��|R�  ��@     ~�  U��|Ts R��|X��|   ��  c�@      @N  -	��  ,�  tm hm �  n �m �  mn en  �  ��  �n �n @N  9�  io _o F�  �o �o S�  �p �p 5^�  ��}5k�  ��~5x�  ��}��  uq mq ��  �q �q 5��  ��}5��  ��}P" (�@       (�@     A       ���  k" Nr Lr ^" vr rr 9�c -�@     <       y" �r �r ym  5�@      �N  
��  �m  �r �r M�@     U��|  <T  _�@      _�@     
       	T  (s &s T  Ms Ks    q�  ��@      �N  ��  ��  zs ps ��  �s �s  T  ��@      ��@            �	j�  T  t t T  5t 3t ��@     U~   ��@     ˀ  ��  Us R��}X��|Y��} ��@     �" ��  U~ T��}Q��} #�@     ~�  U~ R��|X��|   ��@     ~�  U��|Ts Q0R��|X��|   P" ��@      ��@     -       �	��   k" ^" Zt Xt 9�c ��@     $       y" �t t ym  ��@       O  
��  �m  �t �t ��@     Us   <T  ��@      ��@     	       	 T  T  �t �t ��@     Uv Ts     P" �@       �@            �	;�  k" �t �t ^" u u  ��@     �" `�  Us Tv Q��| �@     �V  ��  U��|THQ��| Y�@     � ��  T0 ��@     � ��  U��| G��@     f�  G��@     f�   X  [  �S  9	�
  @�@            ���  �-  9	&`  Cu ?u E�  :	&��  �u |u �  ;	&O
  �u �u �]  <	&��  �u �u .K�@     ��  U�UT�TQ�QR�RX1  =�j  
	�
  ��  �-  
	'`  ^�  	'p  �  	'O
  �]  	'��  E�  	'��  �U 	�
   = v  ��
  ��  �-  �5`  ^�  �5p  �  �5O
  �]  �5��  E�  �5��  ڰ  ��  �U ��
  'i �C
  �L  ���  �f  ���  �>  ���  a  ��	  �R  ��	  �@  �K  qK  �p   /�   ��  0-    /O
  ��  0-    /�
  ��  0-    =nS  t�
  n�  �-  t`  ^�  up  �  vO
  �]  w��  �& yn�  �U z�
  �_  {O
  �  {O
  @�  � /�  ~�  0-    D>n  8�
  0�@     �      �;�  �-  8`  Wv 3v ^�  9p  �w �w �k  :O
  y y �  ;O
  Xy Hy �]  <��  z z ڰ  >�  Wz Gz �U ?�
  '{ 	{ �  @O
  ��Zv  @O
  ���f  Ah2  ��/� BO
  ��&0H  ��  ?d  bO
  d| \| ;�  �@      �H  e��  ��  �| �| ��  �} |} t�  '~ ~ g�  �~ �~ Z�  �~ �~ M�  � � �H  ��  @� 0� ��  � �� 5��  ����  ց ȁ ��  � q� ��  ��   � � M��  ��@     Cm  %�@      0I  ��  `m  �� �� Tm  � � 0I  lm   � � C�@     Us T} Q0R0   Cm  ��@       pI  2�  `m  \� X� Tm  �� �� pI  lm  Є ̄ ��@     Us T} Q0R0   �l  <�@      �I  ��  �l  
� � �l  1� -� �l  k� g� A�@     �k  Us Q| R   T  ��@      ��@     <       !��  T  �� �� T  ȅ ƅ ��@     U��~T|   o�@     �b  �  Us T�� ��@     et H�  Uv Ts Q| R��~1F 01S 0 �@     �V  o�  U��~T Q�� ��@     t Uv T| Q R0Y��~   4T  ��@       J  gT  �� � T  \� T� ��@     Uw       ��@       `J  Qf�  S  Ȇ ��  F  9  \� V� ,  �� ��   �� |�   g� U� `J  5`  ��m  G� 7� z  � �� �   � � �  6� &� �  � � �  &� � �  � � �  � �� �  �� w� �  j� \� �  S� O� M�  ��@     M ��@     Cm  ��@       �J  ,c�  `m  �� �� Tm  Ǔ Ó �J  lm  � �� ,�@     Us Tv Q0R0   Cm  �@       `K  f��  `m  ?� 9� Tm  �� �� `K  lm  Ȕ Ĕ ��@     Us T��~Q0R0   �l  ��@      �K  �P�  �l  �  � �l  e� a� �l  �� �� ��@     �k  Us R'��~20��~#������������������+(   T  <�@      <�@            ���  T  Ǖ ŕ T  � � J�@     U��~T   J�@     �b  ��  Us T�� U�@     �V  ��  U��~T��~Q�� ��@     �b  �  Us T�� �@     �d  0�  Us T�� ��@     t Uv T R0X	#�F     Y��~   T  ��@      �K  S��  T  � � T  Q� M� ��@     Uw T~   e�@     ��  ��  Uv Ts Q�QR��X�� ��@     �  �  Uv Ts XTSOPY1 ��@     �  Uv Ts XtnfsY0  =�>  ��
     �-  �'`  ^�  �'p  �f  �'h2  �O  �'O
  �  �'O
  �]  �'��  ڰ  ��  �H  ��  �U ��
  !k  �[
  Pe  �O
  FH  �S   A  �O
  @�  - =L  �
   �-  '`  ^�  'p  �f  'h2  �O  'O
  �  'O
  �]  '��  �U �
  ڰ  �  Gl  �  'i S   b S   �1  S   'len [
  �C  [
  �c  [
  `E  "[
  Pe  [
  �S  [
  @�  �@*t  � =aj  ��
  � �-  �1`  ^�  �1p  �  �1O
  �[  �17
  \  �1E  �]  �1��  �U ��
  ڰ  ��  �  �[
  ��  �[
  'pos �[
  RC  ��	  �^  ��  @�  �>P  ��
    =�W  t�
  t ^�  t+p  �  u+O
  �  v+�2  ��  w+�2  RC  x+ڌ  �U z�
  yd  {&
  �f  |O
  'tag }[
  'i ~S    D2g  .�
  ��@     F      �{ �-  .'`  �� �� Ǟ  /'�  Z� J� ֳ  0'[
  � � �  1'O
  ܘ ̘ �?  2'<  �� �� �]  3'��  � �� E�  5K  ���U 6�
  �� �� ^�  7p  =� 5� ڰ  8�  �� �� { ��@      �O  ;L � ۛ כ � '� #� � m� g� � �� �� � � � �O  5� ��� � \� T� \� �m  ��@      �O   ) �m  �� �� �m  �� ޝ �m  � �  ��@     �V  U TPQ��   ym  p�@      p�@            a� �m  *� (� ��@     Us   T  ��@      ��@            b� T  O� M�  T  ��@     U Ts   T  ��@      P  B- T  x� r� T  Ǟ Ş ��@     U Tv   1�@     ��  M U} T��~ M�@     ��  U} T��Qw R| X0  =3]  
�
  � �-  
+`  Ǟ  +�  ֳ  +[
  �R +�  C  +� �U �
  ڰ  �  ^�  p  @�  & p  r*M  �`H@     /       �y ^�  �#p  � � ڰ  ��  ?� =� 4T  dH@          �T  e� c�  T    n  ��
  ��@     F       �E �-  �'`  �� �� �   �'�	  � ڟ �>  �'O
  K� C� �  �'O
  �� �� �]  �'��  � � E�  �K  ��*�@     ��  U�UTw Q�RR�XX1  �=  ��
  P�@     >       �� �-  �`  � y� /[  �<  ӡ ˡ �  �O
  9� 3� �]  ���  �� �� E�  �K  ��|�@     ��  U�UTw Q�QR�RX1  DTZ  F�
  ��@           �? K F}  � ע C  G� s� k� 7K  H�	  ֣ ң �  IO
  � � �[  J7
  S� K� \  KE  �� �� �]  L��  � ڰ  N�  � � Oe O�"  ,� (� ��  P[  v� b� �L  Q  T� F� �U S�
  ��P  S�
  � � @WD  �?��@     I       Y	 i lS   � �   p�@      `B  ��	 5 >� 8� ( �� �� `B  B %�@     �] �	 U~ Ts  ��@     �] �	 U~ Ts  ��@     �] U~ Ts    T  3�@      �B  �<
 T  �  � T  ?� ;� A�@     Us T   T  A�@      A�@            ��
 T  w� u� T  �� �� O�@     Us T~   1�@     �V  �
 Us Q�� z�@     �V  �
 Us T�Q�� 8�@      T~ Q���R} X�� 83�@      U~  ��@     � / Uu  ��@     U0  =c^   �  � ��   +[  ��  "�  'end #�  'cur $�   D�k  ��
  �G@     z       �� ��  �"[  U��  ��  �� �� cur ��  � �  T�v  �� K �}   rJ  }pl@           � ڰ  }�  R� H� ��  ~[  Ω ĩ K }  F� @� Oe ��"  �� �� gO  �l@        �� �O  �� �� �O  ު ܪ �O  � � uO  5� /�   �O  �l@     �_ Us�T	�G@     Qv R}     �l@      �l@            �n 5 �� �� ( �� �� %�l@            B �l@     �] Us Tv    P" m@       @  �H k" ԫ Ϋ ^" E� ?� H�c �  y" �� �� ym  m@      �  
� �m  ˬ ɬ $m@     U|   <T  pm@      pm@     
       	T  � � T  � � zm@     U~ T|     T  Hm@      Hm@            �� T  :� 8� T  _� ]� Mm@     Uv   T  \m@      �  �� T  �� �� T  ڭ ԭ :lm@     U�UT�T  G�l@     � 8�l@     	 Us   m@     Us   T]q  c] ��  c [  ڰ  d �  'n f7
  >I_ nm&    h�_  M�G@     X       �� ڰ  M�  .� &� ֳ  N/  �� �� K O}  �� �� T  �G@       �G@            Y T  H� F� T  m� k� �G@     Uv   T  �G@      �   Z[ T  �� �� T  � � :�G@     U�UT�T  8�G@     o Us  �G@     Us   �_  9�
  ��@     F       �� ��  9[  >� 4� ��  :[
  �� �� �1  ;k  � � x =C
  �� ~� 3�  ��@      ��@            E� R�  Ա б E�  � � %��@            _�  8� 2� 9�f ��@            m�  �� �� ��@     T�T    .��@     � U�UQ�Q  �J  �
  P�@     �      �� ��  [  �� �� x C
  �� �� �1  k  �� �� �U !�
  � �� K "}  a� W� �  #�  ۷ ѷ �-  $`  R� J� Pt  %�	   �)  &1  �� �� �H  'O8  A� +� ,NJ  ��@     @�  1&�?  ~ t nO  3� +� �O  o�	  �� �� 9; J�@       @  ub J; Ӻ Ϻ  @  V; � 	� Hjb P@  c; `� Z� o; �� �� f�@     Uw T	C�F         ��@     �| T	/�F       &�@  	 n�  � $  � � & A  � �L  �  � � x+  �7
  M� K� ��@     U Ts R~ Xv   ,�@     Us Q~   &p=  R �e � B  y� q� dO ]�@       �=  �!� �O � � �O '� #� uO e� ]� �=  �O ͽ Ž �O 8� .� �O �� �� �O � � �O I� A� �O �� ��   4dO ��@       �=  �!�O � �� �O @� <� uO ~� v� �=  �O �� �� �O h� ^� �O �� �� �O O� K� �O �� �� �O �� ��    & >  � �L  �  L� F� @>  eo  ��  �� �� �  ��@       �>  �!� �  �� �� �  �� �� �>  '�  ;� 5� 4�  �� �� A�  �� �� <O�  ��@      ��@     '       {�  Q� K� n�  �� �� a�  �� �� %��@     '       ��  l� h� ��  �� �� \��  H�g �>  ��  �� ��      =�  7�@      �>  	� X�  1� /� K�  V� T� �>  e�  q�  <�@     6Z Uu T|    �  0�@        ?  C �  {� y� �  �� �� ��  �� ��  ?  &�  �� �� 1�  =� ;�   ��  ��@      P?  �� �  b� `� �  �� �� P?  �  )�  ��@     �\ U} T|    (�@     Ts Q| R|    &�?   t O  �� �� f��@     ߳  ��@     � Us Q0  C ��@      �<  1C Q D� B� ��@     �! Us   � %�@      �@  �� � k� g� � �� �� �@   �� ��  3� '�  �� ��   8��@     � Us Q~ Rv   �@     ��  U}   Tr`  �+ �  �0�  <  �0�	  �e ���  c� ��  v� ��   6jH  ��m@     �       �� ��  �![  P� J� �3  �!?�  �� �� �� �!�  � � �L  �  A� =�  6Mc  ��k@     �       �� �  �$�  �� w� p  K �}  �� �� ڰ  ��  o� e� �� ��  �� �� cur ��  m� a� T  Bl@      �  �s T  �� �� T  H� D� :Tl@     T�U  8:l@     � Us  Bl@      Us    IY  T�
  @�@     �      � ��  T$[  �� ~� �B  U$ 5� '� �U W�
  ��K X}  �� �� Oe Y�"  �� �� ڰ  Z�  !� � �  [�  |� j� ,�  ��@     �! ��@      p;  m� �! B� <� p;  " �� �� " �� �� " G� A� 5," ��9" �� �� MF" %�@     �: ��@      �;  ;J �: '� #� �: g� a� �;  �: �� �� 5�: ����@     �V  U~ T�Q��   �@     �V  o U~ TPQ�� %�@     U|    T  ��@      ��@     
       q	� T  �  � T  '� %� ��@     U} T|   ��@     �V  � U} Q�� ��@      U|   �  h�B  5�g@     }       �C �  5$�  R� J� K 7}  �� �� Oe 8�"  �� �� ڰ  9�  � � T  8h@      8h@            L� T  M� K� T  t� r� @h@     U|   38 Sh@       Sh@            H	 @8 �� �� G]h@     �b  8h@     . Us   h@     �! Us   T]  _ �  %�   �<  �
  ��@     x       �D �  ,�  �� �� ֳ  ,[
  +� #� ڰ  �  �� �� �U �
  �\T  �@       �@            # T  �� �� T  �� �� ��@     Uv   �@     �V  Uv T| Q�\  6[l  ��k@            �� �  �*�  � � _| �*�  f� `� �k@     �! Us   �_  \�	  ph@     7      ��! �  \1�  �� �� t ]1O  "� � �t  ^1�  �� �� Mj  `�J  � �� .a a�A  v� n� ?   c�  �� �� �'  e-  ��1_  e-  �� p� yW  f�  � � �b  g�  �� �� R  h�  � � O� h�  s� k� 5�  i�  �� �� ��  i�  E� =� `�  i�  �� �� ,�;  �ai@     ?�  �h@      @  wx! Z�  �� �� M�  2� .� @  g�  t�  ��  ��  �h@     �W U{�Tt    �j@     �& �! Uu T{ Q3 "k@     �& Uu T{ Q4  I�o  F�! �  F+�  >ڰ  J�    =P  *�
  P" �  *$�  K ,}  Oe -�"  ڰ  .�  �U /�
  �L  0
  @�  @ IO  �" ^�  p  Er  7
  >ڰ  �    )�E  ��
  и@     Z      �P$ �-  �'`  v� n� E�  �'��  �� �� C  �'� u� i� F�U ��
  �Lڰ  ��   � �� ^�  �p  [� I� e�  �_�@     N�m  +�@       +�@     ,       �{# �m  � � �m  @� >� �m  f� d�  NT  ��@      ��@            ��# T  �� �� T  �� �� ��@     U~ Tv   7T  ��@      �:  �$ T  �� �� T  &� "� ڹ@     U~   �@     �V  ;$ U~ TPQ�L ��@     �| Uv   b�r  �g@            ��$ ��  �%�H  `� \� �U �%�
  �� �� �Y  ��$ �� �� !g@     �| U�UT1  A  )�K  �7
   g@            ��$ C��  �#�H  U b�k  ��f@            �S% C��  �*�H  UCǞ  �*�	  TC��  �*�	  QCgY  �*|I  R )F>  n�
  �f@     [       ��% �r  n+a$  2� *� �E  o+<  �� �� �Y  q�
  +� %� I  ra$  |� v� �f@     v| Tv   Sn  ��
  f@     f       �& �-  �*`  Ussub �*�  T �r  ��
   f@            �^& �-  �*`  Uo  �*@  T �Z  ��
  �e@            ��& �-  �3`  U�� �3  T 6�o  u�d@           �' �'  u#�  U�  v#�  �� �� t w#O  7� /� sub y�  �� ��  �o  G�' �d@     #       ��' ;num G 7
  � � ��  H �G  R� N� hk J�F  �� �� <�( �d@       �d@            O�( �� ��  �( %�d@            �( � � �d@     �/ U	�U����T�T    G   t  :�' �d@     !       ��( ;key :$<  6� 2� ��  ;$�G  s� o� hk =�F  �� �� 4�( �d@      P  B�( �� ��  �( P  �( ,� *� �d@     �/ U�UT�T    =�V  .�' �( `key .�F  ��  /�G  'np 1�G   MH  �
  ��@            ��) ;num "7
  S� O� Kl   "G   �� �� ��  !"�G  �� �� ڰ  ""�  
� � 'hk $�F  .��@     C* U	�U����T�TQ�QR�R  V@  �
  ��@            �C* ;key $<  G� C� Kl  $G   �� �� ��  $�G  �� �� ڰ  $�  �� �� 'hk �F  .��@     C* U�UT�TQ�QR�R  V�>  ��
  P�@     >      �m, Bkey ��F  =� 7� Kl  �G   �� �� ��  ��G  O� G� ڰ  ��  �� �� #nn ��F  � � #bp ��G  �� �� �U ��
  �� �� ,�  
{�@     }/ ��@      �F   ., �/ � � �/ W� S� �F  �/ �� �� �/ �� �� �/ � � �/ ?� ;� �/ {� w� 5�/ ��M�/ k�@     7T  \�@      �F  ��+ T  �� �� T  �� �� k�@     U~ T   �@     �U  , U~ T8Q0R
| 1$����X0Y�� L�@     �/ Ts    r�@     �/ L, U| Ts  ��@     �V  U~ T@Q��  bTf  � d@     y       ��- ��  � �G  -� %� ڰ  � �  �� ��    #sz �C
  �� �� #bp ��G  0� .� #i �C
  U� S� NT  3d@       3d@            �	A- T  {� y� T  �� �� >d@     Uv   tT  Rd@      Rd@            �T  �� �� T  �� �� `d@     Uv Ts     )
A  ��
   �@     V       �c. ��  � �G  � � ڰ  � �  f� `� $0/ *�@       `E  �Y/ �� �� M/ � � A/ .� *� `E  Ke/ �5p/ �lh�@     �U  U�TT8Q0R�X0Y�l    )2A  ��
  @�@     V       �0/ ��  � �G  j� d� ڰ  � �  �� �� $0/ J�@       0U  �Y/ � � M/ \� Z� A/ �� �� 0U  Ke/ �5p/ �l��@     �U  U�TT8Q0R�X0Y�l    Z�G  ��
  }/ "��  ��G  "�Z  ��	  "ڰ  ��  *sz �C
  (�U ��
   Z�f  ��
  �/ "��  ��G  "ڰ  ��  *obp ��G  *bp ��G  *nbp ��G  *i �C
  *sz �C
  (�U ��
  ��  � V�D  j�G  G@     k       ��0 Okey j�F  �X��  k�G  �� �� #res m[
  � � #bp n�G  I� G� #ndp o�G  p� l� 8,G@     �0 U�X PG@     T�X  V�F  _�	   G@            ��0 Oa _"�F  UOb `"�F  T V)=  S�	  `I@     #       �(1 Ba S"�F  �� �� Bb T"�F  �� �� GyI@     v|  V�o  B[
  �F@     H       ��1 Okey B!�F  U#num D[
  &�  � #res E[
  �� y�  Vt  3[
  pF@     1       ��1 Okey 3!�F  U#kp 5<  `� ^� #res 6[
  �� ��  6�>  H�c@     Y       �|2 ��  H'/   UǞ  J�  �� �� �  K�  �� �� sm  M7
  '� #� �Q  N7
  r� p� n O7
  �� �� f�c@     |2  6:V  8 c@     w       �f3 ��  8+/   U�  :�  �� �� 8 :c@      �  A3 8 �� �� �  8 � � &8 9� 7�   <
7 �c@      �c@            B7 a� _� %�c@            #7 �� �� /7 �� ��    O\  �
  ��@            ��4 ��  2/   �� �� Ln  2C
  V� R� ڰ  �  �� �� �U �
  �\�N  C
  �� �� -Q  C
  K� G� Ǟ   �  �� �� �  !�  � 
� ,�  1��@     
7 �@      0E  .�4 7 �� �� 0E  #7 �� �� /7       ��@     �U  T0Rs ����Y�\  )�?  ��
  `�@     9      �
7 ��  �//   f  V  0�  �/C
       �/C
  ` T ڰ  ��  � � F�U ��
  ��Ǟ  ��J  \ L �  ��J  -  t�  ��	  � � �N  �C
  � � -Q  �C
  b V ,�  ��@     8 ��@      ��@     F       
6 8 � � %��@     F       8  	 &8 2 0   ��@     �U  76 U} T@Q��R~ Y�� '�@     �U  i6 U} T1Q��R~ Y�� ��@     �U  �6 U} T2R| ����Y�� �@     [8 �6 Us  f�@     �U  �6 U} T@Q
 1$����R
v 1$����Y�� ��@     �| Q��4$  aef  �<7 "��  �4/   (Ǟ  ��  (�  ��   )�S  ��
  ��@     �       �8 ��  �//   ^ X F�U ��
  �lڰ  ��  � � 78 A�@      �D  ��7 8 � � �D  8 � � &8     ��@     �U  T@Q0X0Y�l  aV  �38 "��  �1/   (Ǟ  ��J  (�  ��J   _�C  �[8 "��  �(/   >(ڰ  ��    bEv  i�a@           �{: ��  i)/   J D ڰ  k�  � � NT  �a@      �a@            n�8 T  � � T  � � �a@     Uv   NT  �a@      �a@            oC9 T    T  , * �a@     Uv   NT  �a@      �a@            p�9 T  Q O T  v t 	b@     Uv   NT  b@      b@            q�9 T  � � T  � �  b@     Uv   NT  ,b@      ,b@            r6: T  � � T  
	 	 7b@     Uv   ${: �b@         z�: /	 -	    �: V	 R	 �: �	 �	    _�W  X�: "��  X*/   (Ǟ  Z�  (�  [�   J�N  F�
  �: "ڰ  F(�  "`h  G(�: (��  I/   (�U J�
   /   �iu  +<  9; "��  +$[  (�Y  -<  >(ϖ 11  (6e  1�
    JC@  <  }; "��   [  (�Y  <  >(ϖ "1  (6e  "�
    )�K  <   a@            ��; CH?  �
  U )k  
_�
  �`@     &       �< C��  
_.[  UC�u  
`.�1  T�H  
bO8  �	 �	  )�P  
7�
  @`@     �       ��< ��  
7"[  
 �	 @  
8"&
  �
 �
 ND  
9"�< 0 " �U 
;�
  � � �H  
=O8    �i  
>*F  � � h`@     Us T�T
��  �?  )�\  
#�
  �_@     �       ��< C��  
#*[  UC�m  
$*�< T W2  Q  7
  �^@     �       ��= �j  �  � � C  �  l ^ �o  �  3 ' �o  �  � � ax �  � } ay �  � � xT  �  D > �T  �  � � �H  �  � �  �l  �7
  �^@            �b> �j  �"�  UC  �"�  � � �o  �"�  Q�o  �"�    �� ��  U Q  �E  N}  �\@     �      �? ��  N"�  Ux_ Pk  � � y_ Qk  � � b Rk  4 2 z Rk  [ W x S}  � � y S}  � � u S}  [ Y v S}  � ~ l S}  � � sx T7
  � � sy T7
  � � m�  T 7
  B <  6�t  50\@     �       ��@ ��  51�  � � �3  61|  � � �  71O
  G A xz 9�  � � yz 9�  � � val ;O
  I A ]\@     dO 8@ Uv Qz  s\@     dO V@ U} Qz  �\@     dO t@ Uv Qz  �\@     dO U} Qz   �[  ��	  �Y@     g      �gD �3  �&|  � � m ��
  !  Lval �gD �P�\  �t
  � � �d  � t
  2 , g  �t
  ~ | M  �t
  � � 'i �C
  �  1� t
  � � N �Z@      �Z@     %       �A /N   $N D B %�Z@     %       :N i g EN � � PN � � [N � � fN     N [@        uB /N = 9 $N w s   :N � � EN    PN V R [N � � fN � �   N ([@      @  �B /N & " $N d \ @  :N � � EN !  PN � � [N � � fN M G   N A[@      p   oC /N � � $N � � p  :N f  `  EN �  �  PN >! :! [N z! t! fN �! �!   N Z[@      �  !�C /N b" ^" $N �" �" �  :N 
# # EN a# W# PN �# �# [N $ $ fN �$ �$   4N o[@      �  "/N % % $N D% <% �  :N �% �% EN & �% PN �& �& [N �& �& fN �' '     /t
  wD 0-    6XM  ��X@     !      �WF ;a �0|  �' �' ;b �0?�  a( [( �  �0O
  �( �( xx �t
  �( �( xy �t
  +) )) yx �t
  W) U) yy �t
  �) �) val �O
  �) �) �X@     dO \E Uv T��Qz  �X@     dO �E U~ T| Qz  Y@     dO �E Uv T Qz  Y@     dO �E U~ T} Qz  5Y@     dO �E U~ T��Qz  LY@     dO F Us T| Qz  _Y@     dO 6F U~ T Qz  pY@     dO Us T} Qz   zE  ��
  �U@     �      ��I �3  �!?�  U�� ��  G* C* xx ��  �* �* yy ��  &+ + sN �U@       �  �MG �N , , �N 4, 2, $ES �U@      @  �`S Y, W, VS ~, |, @  jS �, �, vS �, �,    sN �U@      �  ��G �N %- #- �N J- H- $ES �U@         �`S o- m- VS �- �-    jS �- �- vS �- �-    N &V@      �  �QH /N A. 9. $N �. �. �  :N =/ // EN �/ �/ PN �0 �0 [N X1 J1 fN 72 /2   N UV@      �  ��H /N �2 �2 $N $3 3 �  :N �3 �3 EN �4 �4 PN �5 �5 [N fN �5 �5   N ~V@         �3I /N 66 ,6 $N �6 �6    :N �7 �7 EN 8 e8 PN [N fN �9 �9   4N �V@      �  �/N �9 �9 $N Z: P: �  :N �: �: EN �; �; PN [N 5fN P   6�r  �`T@     Q      �N ;a �)|  S< M< sb �)?�  Txx �t
  �< �< 'xy �t
  yx �t
  H= B= 'yy �t
  sN rT@      �  �
�J �N �= �= �N > > $ES rT@      p	  �`S 5> 1> VS n> l>  
  jS �> �> vS �> �>    sN �T@      �
  �
$K �N ? ? �N <? :? $ES �T@         �`S b? `? VS �? �? �  jS �? �? vS �? �?    sN �T@      @  �
�K �N 0@ .@  �N $ES �T@      �  �`S V@ T@  VS @  jS vS    sN �T@      �  �
L �N |@ z@ �N �@ �@ $ES �T@      `  �`S �@ �@ VS �@ �@    jS A A vS WA UA    sN �T@      �  �
�L  �N �N |A zA $ES �T@      @  �`S �A �A VS �A �A �  jS �A �A vS 2B 0B    sN OU@      �  �
M �N \B ZB �N �B �B $ES OU@         �`S �B �B VS �B �B    jS vS    sN �T@      p  �
�M �N �B �B �N "C C $ES �T@     ! �  �`S _C ]C VS �C �C p  jS �C �C vS 	D D    4sN OU@      �  �
�N FD DD �N lD jD $ES OU@      `  �`S �D �D VS �D �D `  jS �D �D vS )E %E     J\P  �O
  sN Aa_ �O
  Ab_ �O
  's  7
  'a �  'b �  'q �  'q_ O
   J�A  �O
  �N Aa_ �O
  Ab_ �O
   )-R  �O
  �S@     V       �dO Ba_ � O
  jE dE Bb_ � O
  �E �E Bc_ � O
  +F #F #s �7
  �F �F #a ��  ;G 9G #b ��  dG ^G #c ��  �G �G #d ��  H H #d_ �O
  RH NH  Je  �O
  �O Aa_ �O
  Ab_ �O
  Ac_ �O
  *s �7
  *a ��  *b ��  *c ��  *d ��  *d_ �O
   )WN  �t
  ��@            �<P Bx �t
  �H �H By �t
  �H �H [v ��  �h��@     �Y  Uw   )&g  jt
   S@            �kP Oa jt
  U )Ao  at
  S@            ��P Oa at
  U )�s  Xt
  �R@            ��P Oa Xt
  U Joc  q�
  ^Q "��  q[  "�k rC
  "/� sC
  "�1  tk  "�H  u"  (�U w�
  (3 y�!  *num {C
  *end {C
  *nn {C
  (��  |7
   )>m  K�
  ��@     �       ��R ��  K[  /I I J�  LC
  J J �1  Mk  K K o@  N"  3L L 3 P�!  4M 0M & B  �R �U _�
  nM jM 7�R P�@      B  d�R �R �M �M !S �M �M S MN KN 	S wN qN B  -S 9S .v�@     _V U�U#�T�RQ1R�Q1�R �U   ��@     Us T} Q1Rv X|   .B�@     �P U�UT�TQ1R�QX�R  Z�@  �
  ES "��  '[  "�@  '"  "/� 'C
  "�1  'k  (1�  t
  *nn !C
   ZVJ  �k  �S Aa �k  Ab �k  *ret �.  *tmp �.   v_  �I@     �       �T �_  �N �N  �_   �_  �_  JO FO �_  �O �O �_  �P �P �_  �Q �Q �_  \R XR �_  �R �R  
_  pJ@     �       ��T  _   _  #_  �S tS /_  NT JT 9_  �T �T C_  �U �U M_  �V �V Y_  �V �V c_  DW 8W  �_  pK@     \       ��T  �_   �_  �_  "X X `  �X �X `  �X �X  X�  �K@     7      �_V j�  uY iY w�  Z  Z ��  [ �Z ��  \  \ ��  !] ] ��  �] �] ��  ũ  ҩ  ߩ  �  HX�  �  ��  E^ C^ ��  r^ j^ ��  �^ �^ ��  �_ �_ w�  �` �` j�  ma ea �  ��  �a �a ũ  >b 6b ҩ  �b �b ߩ  �b �b �  KL@     v| V Ts  8nL@     V T	8�F      u�L@     DV T�QQ�RR���� :�L@     T�QQ�R    �R M@     �       �SW 	S c c S fc `c !S �c �c  �R -S d d 9S +d )d $dO aM@       @  3�O Ud Od �O �d �d uO �d �d @  �O �e �e �O 'f f �O �f �f �O 7g 1g �O �g �g �O %h h    ��  �M@           ��W ��  vh nh ��  �h �h ��  i i -��  R�  Yi Oi �  �i �i �  )j !j H"�  �  #�  �j �j   ?�  �N@     �       ��X M�  �j �j -Z�  Tg�  ak ]k t�  �k �k ��  �k �k ��  &l  l 9��  �N@     Q       ��  ql ol ��  �l �l 9��  �N@     #       ��  �l �l   m 
m    m�  PO@           �6Z �  7m /m ��  �m �m ��  n n ��  �n yn ��  �n �n ��  wo oo 5͘  �@?�  dO@       �  	ezY Z�  �o �o M�  �o �o �  g�  t�  ��  ��  lO@     �W U{ Tw    O�  P@      P@     0       	�Z {�  Ip Gp n�  sp qp a�  �p �p %P@     0       ��  �p �p ��  �p �p \��  H��  �  ��  &q  q    8P@     %Z Tv  SP@     Tv   =�  pP@     �       ��\ -K�  UX�  tq pq e�  q�  �q �q sN pP@         	�
�Z �N �r �r �N �r �r $ES pP@      �  �`S s s VS =s 9s �  jS xs ts vS �s �s    sN �P@        	�
�[ �N �s �s �N t t $ES �P@      �  �`S Dt Bt VS jt ht �  jS �t �t vS �t �t    sN �P@      @  	�
�[ �N u u  �N $ES �P@      �  �`S 8u 6u  VS �  jS `u \u vS �u �u    4sN �P@         	�
�N �u �u �N v v $ES �P@      p  �`S Gv Cv VS �v �v p  jS �v �v vS �v �v     ��   Q@     >       �D] �  .w *w �  mw gw �  �w �w )�  �w �w <=�   Q@       Q@            	�X�  x x K�  *x (x % Q@            e�  q�  0Q@     6Z Us T|     \  @Q@     <       ��] -\  U#\  Sx Mx \Q@     �S Uu Tt Q�T1�_  u    �Q@     �       �'_ ( �x �x 5 �x �x B Gy Cy vM �Q@     D       �^ N �y ~y <�  �Q@      �Q@     3       q&�  �y �y %�Q@     3       3�  �y �y @�  �y �y M�  z z T  �Q@      �Q@            �^ T  ;z 9z T  `z ^z �Q@     U Tv   �Q@     Uv     <T  �Q@      �Q@            vT  �z �z T  �z �z �Q@     U~    pQ   R@     (       �^_ -~Q  U-�Q  T�Q  �z �z  �P  PR@     -       ��_ -�P  U-�P  TQ  �z �z Q  { {  gO  �R@     m       ��` uO  D{ >{ �O  �{ �{ �O  �{ �{ �O  :| 4| �O  �| �| 9�O  �R@     "       �O  �| �| �O  } } T  �R@      �R@            �` T  :} 6} T  r} p} �R@     Uv   ��R@     } Uv Q~    dO 0S@     \       �,a uO �} �} �O �} �} �O \~ T~ �O �~ �~ �O l j �O � � �O � � �O [� W� �O �� ��  sN �S@             ��a �N Հ р �N � � tES �S@      �S@            �`S O� K� VS �� �� %�S@            jS �� �� vS � ��    N T@     P       �<b $N 5� /� -/N T:N �� �� EN � � PN ,� (� [N f� b� fN �� ��  9; a@     #       ��b J; �� ܃ KV;  %a@            c; � � o; @� >� :/a@     T	C�F        {: Pa@     f       ��b -�: U�: f� d� �: �� ��  38 �b@     #       ��c @8 �� �� HL8 `  M8 � � 7T  �b@      �  �oc T  Z� T� T  �� �� :�b@     T�U  �b@     [8 Us    38  c@            ��c @8 � �� .c@     �b U�U  P" 0g@     A       ��d ^" @� 2� k" � ۆ �  y" u� o� ym  Fg@      �  
Cd �m   �� Mg@     Us   4T  Qg@      �  	T  �� �� T  N� J� :bg@     T�U    w�! �g@     d       �De �! �� �� ?�g@     *       e �! � � 4T  �g@        MT  1� /� T  X� T�   9�! �g@            �! �� �� 9�d �g@            �!    ��   p@     &       ��e ��  ۉ Չ ��  -� '� ��  � y� -��  R�  �  �  .4p@     SW U�UT�TQ�Q�Rr   ��   v@     p       �pf ��  ъ ˊ ��  %� � K��   ��  H��  �!  ��  �� �� ��  �� � �!  5��  P��  I� C� u7v@     `f T	�T $ & Giv@     Z�     3�  �{@     3       ��f E�  �� �� R�  � � _�  c� ]� %�{@            m�  �� �� �{@     T�T   ?  �@     \       �=g  Q  Q ^ ׍ Ӎ k � � x M� G� GZ�@     �   O�  ��@     a       ��g -a�  U-n�  T-{�  Q��  �� �� K��    *  ��  ؎ Ў   �  І@     �       ��h �  =� 5� $�  �� �� 1�  � � >�  �� �� v�  �@     @       �h 1�  Ր Ӑ $�  �� �� �  "�  � %�@     @       >�  K� E� 9K�  �@     @       L�  �� �� Y�  ӑ ё f�  �� �� 9�@     T|     ��@     Uv T|   ��  @�@     ;       ��i �  !� � �  s� m� !�  Œ �� .�  � � ;�  i� c� H�  U�  9��  _�@            ;�  �� �� .�  �� � !�  3� /� �  p� l� �  �� �� %_�@            H�  � � U�  %� #� :t�@     U�UT�TQ�QR�RX�X    ?�  ��@            �j M�  P� J� -Z�  Tg�  t�  ��  ��  .��@     �W U�UTt   �  ��@     /       �nj ��  �� �� -�  T-�  Q&�  ߕ ٕ 1�  +� )�  m�  ��@     6       ��j �  T� N� ��  �� �� ��  �� � ��  ��  ��  ͘  .Ԕ@     �X U�UT�TQ�Q  =�  p�@            �=k -K�  UX�  J� D� e�  q�  .�@     6Z Uu T�T  ��  ��@            ��k �  �� �� �  � � �  )�  .��@     �\ U�UT�T  �m  �@     (       ��k -�m  U-�m  T-�m  Q ym  @�@            �l �m  @� :� :P�@     U�U  Cm  `�@     B       �`l Tm  �� �� `m  � � Klm   {�@     Us Tv Q0R0  m  ��@     ^       ��l *m  �� �� 6m  S� I� $Cm  ɠ@       �4  b`m  К Ț Tm  =� 1� �4  lm  Ǜ ś נ@     Uv Ts Q0R0    �l  �@            �m -m  U �l  ��@            ��m �l  � � �l  .� (� �l  �� z� .��@     �k  U�UQ�TR�Q  wCh  У@     6       ��m Qh  Ҝ ̜ %ۣ@            _h  "� � 4T  ޣ@        6  VT  [� Y� T  �� ~�    v  �@     y      ��p 4v  ŝ �� Nv  W� M� [v  ؞ ̞ Av  b� `� 'v  �� �� hv  �� �� 5uv  �L�v  � � �v  0� *� �v  � y� �v  ͠ ɠ �v  � � �v  .� (� K�v  m  5�@      �7  )Uo 6m  ~� z� *m  �� �� $Cm  =�@       �7  b`m  �� � Tm  0� *� �7  Klm   V�@     Us Tv Q0R0    m  ث@      08  A�o 6m  �� |� *m  �� �� $Cm  �@       `8  b`m  �� � Tm  0� ,� `8  lm  j� f� ��@     Us Tv Q0R0    ��@     �b  p Us T�L -�@     �b  +p Us T�L x�@     �d  Ip Us T�L ǫ@     �b  gp Us T�L %�@     �b  �p Us T�L A�@     �b  Us T�L  �  ��@     &       �>q "�  �� �� /�  � ߣ <�  L� F� I�  �� �� V�  � � �c�   .��@     �m U�TT Q�X1'v  �U1Av  �Q  \   �@            ��q -\  U#\  B� <� .*�@     D] Uu T�T  �: p�@     3       ��q �: �� �� �: � � �: 6� 2� 5�: �\��@     �V  Us T�Q�\  �P ��@     �      ��s �P �� m� �P q� [� �P v� ^� �P �� v� 
Q �� �� KQ  "Q .Q �� �� :Q 3� #� FQ QQ H�P @A  
Q � �� �P �� �� �P R� D� �P �� � �P �� �� @A  Q K� ?� "Q Ӱ ϰ .Q :Q FQ � 	� QQ ]� [� 7�R �@      �A  ��s �R �� �� !S � � S Y� Q� 	S �� �� �A  -S 9S .��@     _V U�U#�T�XQ�QR�R1�R �U   8r�@     �s U| Ts Q R} Xv  ��@     � U| Ts Q}     �V   �@     1       �et �V  %� � �V  w� q� �V  ˳ ó �V  2� *� �V  �� �� ,�@     U�UT�T   ��@           ��y  
� �� , � � 9 k� c� ` ߶ ۶ S � � F C� A� 5m ��z q� k� � ׷ �� � � � � A� 9� � �� �� � ]� K� M� ��@     � �@      @P  ��w ' *� �  ּ ʼ  �� v�   .� "� � �� �� @P  54 ��A a� S� N 
� �� [ �� �� h P� F� m  ��@      �P  �
jv 6m  �� �� *m   � �� $Cm  ��@        Q  b`m  <� 6� Tm  �� ��  Q  lm  �� �� ��@     U Tv Q0R0    m  ^�@       pQ  �(w 6m   � �� *m  <� 8� $Cm  f�@       �Q  b`m  v� r� Tm  �� �� �Q  lm  � � �@     U T~ Q0R0    #�@     �b  #w U T�� ��@     �d  Bw U T�� O�@     �b  aw U T�� ��@     �b  �w U T�� ��@     �b  U T��   �l  �@      �Q  ��w m  |� x�  p�  R  Gx � �� �� 4Cm  ;�@      PR  �`m  �� �� Tm  � � PR  lm  R� N� U�@     U Tw Q0R0    Cm  ��@       �R  ��x `m  �� �� Tm  �� �� �R  lm  � �� ��@     U T~ Q0R0   �l  !�@      �R  �y  �l  �l  <� :� �l  a� _� 3�@     �k  U Qv R��  T  ��@      ��@     '       �gy T  �� �� T  �� �� ��@     U��Tv   
�@     �V  �y U��T��Q�� u�@     t U} Tv Q��Rs 0s 0,( X'�F     #�F     ���0.( Y��  T  ��@            �;z T  �� �� T  (� "� :��@     U�UT�T  �Q  ��@     ,       �rz -�Q  U-�Q  T�Q  x� t�  pQ   �@            ��z -~Q  U-�Q  T�Q  .�@     '_ Uu Tt   �P  P�@            �	{ -�P  U-�P  TQ  Q  ._�@     ^_ Uu Tt   �P  p�@     F       ��{ -�P  U-�P  T�P  �� �� �P  �� �� 9�P  ��@            �P  :� 8� �P  _� ]� %��@            �P  �P     gO  0�@            �| uO  �� �� �O  �� �� �O  ,� &� �O  ~� x� �O  .?�@     �_ U�UT�TQ�QR�R  QNe  Ne  92xBY  8Y  8 xD  D  8 Q}t  }t  9&QN  N  9Q j   j  9Q�  �  :XQ$  $  :.Q�  �  9Q?  ?  9(�5Q  5Q  *cQbU  bU  #Qn  n  9 ��  �  &  ��  �:  P�@     &      �  (\  �9   ,  i   �L   �  int �  �   @	�   �  	�    p  	 	@   �  	#	@   X  	&	@   �  	)	@    �  	,	@   (�  	-	@   0/  	2S   8�  	5S   < �   �  	�   �  	8"c   
+  	K  �   
%  	L  
�  	M  '  ��  
�A  ;  �s  
�T  �  s&  
S   �  
Z   )  A"�  �  �   ��  �  �a    ��  ��  <h ��  �I  �   �  X�  �  a   �  u  9    �   m�      u  a    f  �  #  a   A  u  9   9   a    J   �"M  S  �  PH�  Ǟ  JP   ֳ  KL   pos LL     N  /[  O   �K P   (�R Q]  0ڰ  Su  8O�  TP  @��  UP  H �  �  <v �9   ��  �a    �  ��  ""  �,  2  L   P  A  L   P  L    V  �  �   j  p  {  A   X�  WS  v  :9   �  L�  x N�   y O�   �  Q�  	�  ~   w  
  y�   �!  y�  �   z�  H  z�   "  |�  N`  Z   �`  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} Z    5�  Z   `�  	S   _| 
P  
!  T  ?   V  2   V  B  a     �  `  	�  �  (QT     SA   0�  TA  N5  VT  �   W�   H� XZ  �1  ZS     �  A  �  \�  �  �  Z   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  �s  �8  5"�  �  �$  �4  S  x UA   len VT  e� WV   �#  Y�  	  �%  {,  2  L  S   S   L  a      �#  �_  e  S   ~  S   S   a    �.  ��  �  �  S   S   a    �8  `�3  .   3   �; 9  �1  S   �5    �+     `(  R  (�/  ~  0�  a   8*    @ �  ?  u(  
�  	@  �2  (_  e  S   y  a   y   �  �3  ;�  �  �  �   v)  ]�  �  �  �  P  L    �3  y�  �  S   �  �  L   a    H7  ��    S     �     M  51  0��  y2  ��   � �R   ��  *
 ��  / ��   $ �  ( 2$  �  -4  lV  +  ��  	�  �  $8  �V  	�  �  Ab  �h    ��   	�  {"  �A  !  �T  	�  \   �S   �  �Z   }  �9   )$  �L   �z  A  _]  9   �   9   c,  +S   C*  6a   +D  C@   �]  P-   {�  c�	  x e3	   y f3	   ��  h�	   :   �
  xx �M	   xy �M	  yx �M	  yy �M	   5  ��	  	
  8  �B
  ��  ��   ��  �	   $  �
  c   �\
  b
  m
  a    �  ��
  Kl  �a    �  �O
   s  �m
  �"  $�
  �
  �   +�
  �� -�
   �W .�
  Kl  /a    �j   �
    %  D/  uR F�
   �
 G�
   }  I  Z   &�  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<�  5�  >�   ��  ?�  �"  A�  �"  B�  i!  C�   %!  E�  (2!  F�  0�  G�  8   I  �"   s`  ��  u�   5�  v�  ֳ  x�  !  z�  m  {�   v  }  J  �#z  �  �!  �}>  ڰ  u   {3  �	  S0  �	  �/  �	  �1  �	  �1  �p#  Y/  �/  �*  ��  (�)  �>  0+:  ��#  8<8  ��#  X�*  �	  � �3  �"K  Q  �(  ��  Oe �J#   �-  �m  ڰ  �u   U  �"�  �  �  8�  ah !P#   Oe "!  U1  #/   ;+  $0  0 i(  �$�  �  l;  ��h  ah �P#   Oe �]#  y2  ��   {:  �u  (�� ��  h/ ��  p�� �   x T   � u  {  _  �<  �!  	   �  	  �  	    	  �  	   �U �  (�  �  03"  	  8�  �  @`  !	  Hd  "�  P�@  $�
  X�;  )  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7<  ��� 8�  �K <�  �ڰ  =u  �^�  >A  �U  @/  �t  B�
  �k  Ca   ��L  E  � "   I  O  1  Xm�  ��  oh   �@  p�
  �e q�  �L  r�  P @  $%�  �    0\�  �-  ^m   ��  _h  �W `�  x a	  �@  b�
   �e d�  0�"  eM	  pi"  fM	  x� g�  ���  i�  �.a k�  ��  l	  �J  m	  �Mj  o`  ��  q	  ��  r�  �M  ta    Z  u9   _"  w�  (   x�  Ud za    �L  |  ( �!  F#     Z!  AM  ��  Ch   T D  �!  E�  "  F�   S  Z   �  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  M  0  `),  2  �"  �e�  �1  g
   H+  h�   x+  i	  0��  k�!  8�)  n#D#  h�'  q�  p��  r[  t�*  y	  x �  `  �  �S  I{  �  �)�  �  �!  H�  $  �a    7:  ��  s4  ��   b  8H�  !  J�   m  K�  A� MM	  �� NM	  �  P�  
  Q�   ��  R�  (�  S�  0 �  U   x  tO  x   �$�  �  �!  0'  ad  )	   �1  *�  &D  +	  2B  ,	  x� -
     �)$  *  �"  P��  ��  �0   �1  �	  �&  ��  �3  �
  ]7  ��  0�7  �a   @�1  �[  H P6  �  tag '	   Kl  g	   �6  	�  �  �5  Z   
  i7   �&  9  F9  8%  �*   �,  
�  ./   6
s  b 8
   5�  9
	  ��  :
	  5  ;
	  Q(  <
	    -  I
(�    �8  Z   ��  �:   4,  �6  $  �/  l9   �2  ��  �\  �  b<  �	   1S �	  p �   �  p  ��  �#  �g	  �'  �-  3  Z	  B  >   �2  �N  T  _  >   l/  �k  q    �  >  �   �   ;)  H�  �#  �'	   :  �	  �5  �  F1  �M	  ,8  �M	   2*  �9  (�*  �!  0`1  �B  8��  �_  @ �  �-  ��  d)  s-  3  Z	  B  a    �j  Z   �h  jb   �U  �P   �B  �B  9  F#�  	u  �$  @J�  �#  L	   y2  M�  W� OV  �� P|  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!    �-  (qP  �-  sm   Oe tP  ��  u�  � v�   �  �/  )b  h  Z	  |  �  �   g%  .�  �  �  �   �.  1�  �  �  �  �  m   
  73  6�  �  �  �  �     �8  :�     Z	    �  �   "3  >b  $)  Y,  2  Z	  P  �  �  �  m   �6  _\  b  Z	  �  �  �  �  m   �3  f�  �  �  �  �  �   ;0  l�  �  Z	  �  �  '	  g	   �&  x�;  ah �    y2  � �  H�8  �    P�8  � P  X�'  � �  `� � �  h�9  � ;  p �  �.  ��  "9  H2�  Mj  4`   H5  5T  (�)  6T  0�  7	  8�  8�  @ �0  :M  7<  :�  M  T%  �=0  ڰ  ?u   �0  @	  q5  A	  L)  B	  )  C�  Ǟ  E�  �  F�  `Ud Ha   � X+  J<  �  1  N  T  Z	  w  A  h  	  	  �   �&  &�  �  �  h   �1  *�  �  Z	  �  <   �6  -�  �  �  <   w-  1�  �  Z	  �  �   �;  4�      �   =;  8  "  Z	  6  <  s   B$  <B  H  Z	  \  <  '	   2  @h  n  Z	  �  �  <  	  [   7  G�  �  Z	  �  h  	  	  T   q8  N�  �  Z	  �  h  A   )2  S�  �  Z	     h  	  	  [      M	  k.  ���   ah �   #,  �	  H�4  �	  P,;  �	  XEY �B  `/q �w  hZ)  ��  p�#  ��  x'0  ��  �.  ��  ���  �\  �� ��  �`9  ��  ���  ��  �5  �  �U#  �6  � �/  �   	�   �2  �!     a   8S  �L!  �d  ��   �W  �9   C  �$!  	L!  �&  0��!  y%  �g	   �/  �g	  �'  �g	  �6  �g	  �+  �g	   �6  �g	  ( �7  �]!  *  V'�!  �!  �0  �*   u&"  |#  w	   �#  x	  � y	  C4  z	   �&  |�!  �'  �>"  D"  Z	  ]"  �!  	  ]"   B
  �9  �o"  u"  �"  �!  ]"   A2  ��"  �"  Z	  �"  �!  	  �  �"   &"  8(  �"  ��  )2"   $�  )c"  �-  )�"   )  �"  	�"  3  <1#  �� >%1#   ��  ?%�!   #  #  A#  7#    �(  �Q  A  �D  &�  >  �#  L       �#  L    �  �#  L     H'  �%�  <  Z   9,$  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  Va$  <v X�   ֳ  Y�  �  Z�   yK  \,$  	a$  �I  `U]%  Q  WM	   �g  XM	  �;  Z	  �U  [	  �B ]�   �o  ^�  "Y  `]%  (+I  a]%  8
  c�  H�!  d�  J�   e�  LH  f�  N�`  h�  P�X  i�  RO  k�  T,G  l�  V�t  m�  X '	  m%  L    I  or$  �g  8�W&  ��  �M	   )r  ��  dS  ��  
�B  ��  �P  ��  �p  ��  �K  ��  =  ��  me  ��  +^  ��  �]  ��  �u  �W&  
h  ��  $^K  ��  &tR  �a   (%?  �a   0 �  g&  L    �]  �y%  �S  8?b'  ��  AM	   )r  B�  dS  C�  
�B  D�  �A  F�  �n  H�  �n  I�  �W  J�  me  K�  +^  L�  �]  M�  �u  OW&  
h  Q�  $�V  R�  &tR  Xa   (%?  Ya   0 �u  [s&  JW  �x�)  ��  z�   =  {�  �<  |�  tB  }�  �k  ~�  �m  �  
�D  ��  gJ  ��  !X  ��  �S  ��  5f  ��  ?X  ��  �a  ��  �_  ��  �a  ��  Gf  ��  �=  ��)   �E  �'	  0F  �'	  8�A  �'	  @F  �'	  H�E  ��)  P5D  ��  TH  ��  V#l  ��  X$r  ��  Z_S  ��  \'N  ��  ^?_  ��  `L  ��  b�O  �'	  h�O  �'	  p~e  ��  x [  ��  z0m  ��  |�M  ��  ~rM  ��  �]  ��  ��g  ��  � �  �)  L   	 �  �)  L    �X  �o'  kE  @�Z*  �^  �M	   zp  �M	  dv  ��  �i  ��  �<  �'	  �F  �'	   �D  �'	  (�p  �'	  03X  �'	  8 �b  ��)  K_  @�H+  ��  �M	   �J  �'	  �<  ��  e  ��  $� ��  dk  ��  ![  ��  L^  ��  �`  �H+  yN  �X+  ,ma  �h+  4�Z  ��  :�q  ��  ;r  ��  <�u  ��  = �  X+  L    �  h+  L    �  x+  L    	l  �g*  �M  (8f,  ��  :M	   �T  ;�  �P  <�  
�K  =�  B  >�  ^  ?�  �g  @�  /o  A�  %B  B�  �O  C�  �<  D�  �]  E�  *w  F�  dW  G�   �F  H�  " e=  J�+  |[  O�,  �� Q�   �\  R�  red S�  q  T�   �[  Vs,  �?  (�-  `a  ��   �L  �-  r  �-  &W  ��  �F  �-    �  Ik  ��,  	  ��  L]-  }W N�   ��  O	  ��  P	   ��  R(-  8y  hl�-  �~  n	   ��  o	  �~  p�-   ]-  �-  L    `�  ri-  ,�  0�.  }W ��   ��  �M	  def �M	  ��  �M	  tag �'	   cy  �	  ( ˣ  ��-  ��  �W.  Ԛ  �    cy  �	  �}  �	   	�  �".  U�   ��.  �~  �	   ��  �	  ˧  �	  �~  ��.  i{  ��.   .  W.  �  �c.  >i   J/  tag L'	   ��  MM	  /� N	  �f  O/   '	  2\  Q�.  G   �`/  Tag �'	   g  �'	  �=  �'	  Ja  �'	   mn  �l/  /  �v   ��/  �T  ��   �Y  ��  D  ��  S  ��  E]  ��  ;C  �'	  �: �   �[  �r/  DQ   0  E]  �   ;C  '	  �:    �i  �/  >M  0.�0  ��  0�   �Z  1	  vv  2	  �r 3�0  =P  4	  �Q  5�0   ^�  6A  ( �/   0  �p  8-0  CE  Y�0  �B  [�   b  \�   Pq  ^�0  �0  �m  x.1  ��  z�   �R  {�  Up  |�0   �=  ~�0  �i  ��1  ��  ��   5�  ��  �"  ��  �"  ��  i!  ��  %!  ��  
2!  ��  �  ��   W  �;1  �U  p2  �  �   
   �  Sd  !�  �Q  "�  �G  #�  �v  $�  �=  %�  sD  &�  �\  '�  �X  (�  	`N  )p2  
 �  �2  L    �T  +�1  �  >t  ��2  �>  ��2   � ��2  !  ��  m  ��  �[  ��  SX  ��   �<  �3  �2  x@  "P3  �  $�   �`  %�  TL  &�2  �o 'P3   V3  �  �h  )	3  �Z  <�3  �  >�   �f  ?V3   fR  Ai3  !Z�3  "j \\3  "�Y ]�3   ms   V�3  �  X�   �r _�3   J  a�3  �t  r!4  4  U<  �-T5  �~  /	   Ԛ  0   ��  1   ;�  3�I  ��  4t	   ��  6   (z�  9�  0��  :�R  8��  <�  @*�  =�  A��  >Z	  D��  ?eT  H�  A�  P|�  B�  Q��  CZ	  T��  DeT  X�  F U  `_�  H	  hˊ  I   p�{  K	  x��  L/  ���  N'	  � �c  (��5  �B �   �c  �  �y �  �Y  �'	  cC  �	   �  ��  $ 	\  �T5   L  � �5  �5  �i  ���:  ah ��   �u  �/  ��v  �'	  �R  ��   o  �`/  (�& �m%  0�Q  �g&  �@  �f,  �5�  ��  �<  �b'  ��`  ��  0�a  ��0  8#os2 ��)  hF�  �Z*  �j  �  0 M  �'	  8w_ �e<  @�>  ��<  H�A  ��<  P^Z  ��<  X�f  ��<  `KT  ��<  h�i  �a   pQ  �a   x#mm �a   �#var �a   �g  �a   ��Y �.1  �Fq �x+  �jQ  �'	  �nQ  ��2  �m  �3  ��P  -  @  �  @B  F=  H�u  �  P�u  �,  Q�;  '	  XzQ    `FN  '	  hT    p!u  '	  x#cvt L=  �2i  �:  �)  )�
  ��  +�  ��j  -'	  �:>  .'	  ��_  0�  �S?  3�  �E�  4�3  ��W  6h  �XA  8�  �	K  9	  ��c  ?'	  �][  @'	  ��J  B'	  �'<  C  �	Z  E   �q  F'	  �G  G	  �T  H'	  �a  I   �\  K  (�u  L'	  0o  M9=  8^C  N	  <:W  OR=  @_  Q  H�@  R'	  P>  S	  X}?  Th  \m?  Uh  `#bdf X�5  h�k  \'	  ��Z  ]'	  �Pl  h'	  �(a  i'	  �i ma   ��d na   � �Q  �-  �g  �"�:  �:  �t  x�e<  ��  ��5   ֳ  �KB  ȩ  ��  �m  �0  �1  �'	   x �	  (^�  �A  0��  �	  8   ��  <�;  �  @�C  �	  `� �	  d"f �	  h�I  ��  lpp1 ��  ppp2 ��  �Ǟ  �>  ��y  �>  �BJ  �!>  �<  �  bL  �'	   Ud �a   (�W  �	  0r�  �	  4#pp3 ��  8#pp4 ��  HO�  �  X��  �  `�k  �/  h �^  r<  x<  Z	  �<  �5  '	  A  /   �D  *�<  �<  Z	  �<  �:  	  '	  	   �b  A�<  �<  Z	  �<  �:   SQ  Q�<  �<  =  �:   �=  Z   T9=  �G   �v  k_  <L  ok   �`  _=  �,  [  	  �j  @�>  ڰ  �u   �0  ��  q5  ��  
0�  ��     ��  org �T  cur �T  " �T   �   �  (H� ��2  0�>  ��  8 ,L  �X=  ��  �>  X=  @\  �'.>  4>  $�r  P�KB  ��  ��5   ֳ  �KB  ڰ  �u  �U �Z	  top �	   �  �	  (�� �"-  0E�  �	  8/�  �	  @zp0 �>  Hzp1 �>  �zp2 �>  �%pts �>  & �  �>  H&ٙ  �	  �&�e ��  �&��  ��P  �%GS �$O  &�  �	  x&�* �  �%IP �	  �&�z  �	  �&�|  ��  �&��  �	  �&��  ��  �&�  �'	  �%cvt �"-  �&*�  �	  �&	�  �  �&��  �	  �&Ӣ  �	  �&č  �%P  �&��  �	  �&��  �	  �&��  �%P  �&��  �	  �&�  �	  �&̞  �	  �&}�  �	  �&և  �"R  �&�P  ��   &�K  ��  &Ex  ��O  &@�  ��  8&�y  �"-  @&C�  �@	  H&^�  �@	  P&�  �@	  X&�  ��  `&��  �$O  h&�w  ��  �&e�  ��  �&�|  �	  �&߅  ��P  �&��  �5Q  �&!�  �5Q  �&(�  �5Q  �&��  �	Q  �&W�  �	Q   &8�  �`Q  &��  ��Q  &�}  ��Q  &�  ��Q   &}~  ��  ()�  q�  )��  v�  *�  {�  +|  �  ,#}  ��  -��  ��  .�  �'	  0T�  �'	  8��  �'	  @��  �'	  H �d  � XB  ^B  �a   �C  ah �   �e E  X�  �  `q�  �P  �m '	  ��' "	  �%�  $	  ��  %	  �)�  &%P   ��  (	  ��  )	  ��  *%P  7�  ,	  %�  -	  Ex  /�O   #GS 1$O  P!u  3'	  �#cvt 4"-  �9z  6�  ��y  7"-  � �  9>  �B�  ;!>  �  ?Z	  Fz  @Z	   /�  ��:  <e  I�C  �C  Z	  D  A  �5  	  	  �   l  s�C  Z  �'D  -D  8D  �5   -H  �DD  JD  Z	  mD  �5  '	  	    /   �e  2zD  �D  Z	  �D  �5  '	  	  	  A  �D  �D   �  �1  �h  S�D  �D  Z	  �D  �5  s  /   �^  p�D  �D  Z	  E  �5  '	  E   �  eN  �$E  *E  Z	  CE  �5  	  CE   �  Ub  �VE  \E  Z	  uE  �5  A  �   #K  ��E  �E  �E  �5  �  	  �E  �2   �  3l  ��E  �E  Z	  �E  �5  	   �d  	�E  �E  �  
F  �5  	  R=  R=  
F     �J  0F  #F  Z	  AF  �5  	  �  �   CZ  NNF  TF  Z	  mF  �5  �  CE   :=  pzF  �F  �  �F  �5  �  �F  �F   	  �Z  ��F  �F  Z	  �F  �5  A   �^  �'D  GK  ��F  �F  	  G  �5  	  	   N=  0�.I  w_ �"e<   EY �"�C  �e �"D  /q �"D  ��  �"_   ob �"8D  (pR �"�F  0�^ �"IE  8D_ �"�F  @x` �"�F  HPr �"�F  P1s �"�F  X�k �"�F  `�S �"�F  h�O �"�F  p�Y �"�F  xAq �"�F  ��b �"�F  �ar �"mD  ��[  �"E  � Q  �"�F  �� �"�F  �X �"�F  ��U �"IE  �`H  �"�F  ��W  �"�F  ��n �"�D  ��T �"�D  �zi  "�F  ��d "�F  ��Q "�F  ��] "�F  �B  "�E   UU "�E  �p  "F  �[ "uE  ]o 
"AF   4P "mF  ( sh  G  AD  HI  .I  ��   'ZI  `I  Z	  tI  h  tI   �-  �z   +�I  �I  Z	  �I  h  �I   �I  �.  9~   /�I  �I  Z	  �I  h  	  "-   "�   6�I  �I  Z	  J  h  	      ��   =�I  �   B�I  ��   G&J  ,J  Z	  @J  h  	   Ӏ   K�I  ݓ   PXJ  ^J  Z	  �J  h  R=  �J  �J  �I      `�   W�  ��   Z�I  3�   _�J  �J  Z	  �J  h  R=      >�   d�J  	�J  y  ` d�K  �~   f"NI   -�   g"�I  g�   h"J  ��   i"@J  7�   j"zI   Y�   k"�I  (�   l"J  0&�   m"J  8U�   n"�J  @A�   o"�J  HY�   rLJ  P��   s�J  X �  !'�K  �K  Z	  �K  h  	  �F   ¦  !,�K  ۧ  !1�K  r�  !8�K  ��  !=�K  ��  !B�K  ʍ  !G�K  �  !N�  ֈ  !QL  	L  ��  @!Q�L  H�  !S�K   ��  !T�K  -�  !U�K  ��  !W�K  ݖ  !X�K   p�  !Y�K  (#�  !Z�K  0��  !\�K  8 ͂  "'�L  	�L  �p  "'�L  �B  ")h    ��  # �L  �L  '	  �L  h  	  /   s�  #$�L  	�L  ��  #$M  ��  #&�L    �<  $M   M  Z	  >M  >  �  9  �   s=  $$JM  PM  Z	  iM  >  �  a    �  $)zM  	iM  #P  $)�M  R  $+M   bD $,>M   
�7  %!  ��  '"�M  �M  \�  �K�M  ah Mc#   �y  O>  8��  Q	  x ��  6�  �  `A$O  rp0 C�   rp1 D�  rp2 E�  �w  G�	  �y  H�	  
��  I�	  Ǥ  K	  \�  L@	   ��  M	  (��  O�  ,�}  P@	  0c�  Q@	  8��  R@	  @��  S�  Hg�  T�  J�~  V�  L��  [�  Mף  \	  P
�  ^�  T�  _�  V>�  `�  X �  bN  	$O  W�  Z   �`O  ��   �x  ۡ  D�   �{  ��O  Ǟ  �   ֳ  �	   3�  �`O  ��  ��O  �O  �O  L    ��  (�P  x  �	   �k �	  end �	  opc �	  &
  ��  �w  ��  ��  �'	    �  ��O  '�  �1P  �O  ��  P��P  U�  �	   a{  �	  � �  � 	  1� M	   �y  �P  (��  �  H�|  	�  I�  
�  J @	  �P  L    �  7P  -�  5�P  �P  @	  	Q  !>  @	  @	   �  ;Q  Q  5Q  !>  >  �  @	   z  BAQ  GQ  @	  `Q  !>  �  �   o�  HlQ  rQ  	  �Q  !>   \�  L�Q  �Q  @	  �Q  !>  '	   C�  R�Q  �Q  �Q  !>  '	  @	   �z   [R  Q�  ]	   J{  ^	  ��  _	  Def aR   P  �y  c�Q  V�  c.R  �Q   .�  �"0O  �{  )iR  �  +M	   {�  ,M	   ��  .!uR  AR  ��  :�R  �  <�   �  =iR   �  ?�R  {R  ݗ  B�R  ɢ  D	   ��  E	  ��  FR=  �  H�E   F�  KS  �R  &�  O>S  z  QM	   �  RM	  �  SM	   j�  UJS  	S  �~  XkS  ّ  Z>S    !�  \wS  PS  �{   `�S  ��  b	   ��  c�R  �  e�  ��  f	  ��  gkS   �  i}S  ,�  i�S  }S  Ń  lT  ��  n	   "�  oR=  �y  pR=   x�  r�S  S|  r7T  �S  �w  8}eT  �  �S   ��  �T    М  �qT  =T  b�  ��T  tag �'	   "�  ��  �y  ��  
p�  ��   *�  ��T  wT  ��  0� U  9�  ��   �  ��S  
Q ��T  ( +�  �U  �T  ��  Z   [;U  'S�   �'y   p'�  � ̐  Z   mrU  '��   �'�~   @'��    'Iy   'k�  � Z   &��W  �   ��  ��  ��  �  3�  &�  >�  @w    	��  
(�  s�  ��  j�  X�  �  Y�  8�  P�  �}  l�   �  !��  "<}  #��  $��  %׊  &C�  'j�  (�  0��  19�  @d�  AV�  Q��  R>�  Sn}  TTx  U�  V��  Wc�  Xy�  `�  a�x  b��  c��  pڌ  �̤  ��  ���  �.�  �%�  ��w  ���  �ۋ  �֠  �}�  ���  ��x  ���  �u�  ��x  �O~  ��y  �&�  ��|  �,�  �{  �Uw  �ř  �/�  �(�  ��  �d�  �?�  ���  �{w  �n�  �vz  �զ  �az  ���  �+x  ���  �~  �l�  ��  �2�  ���  �p�  �a�  ��  ��  � (#z  �uM  	@�F     )4�  ��J  	�F     )��  L  	��F     )�  .�L  	��F     )�  $�L  	��F     X!  7X  L    	'X  )G�  ,7X  	 �F     *�M  o	`�F     ;�  (��X  ��  �	   �  ��  �  ��  
�  �'	  x�  ��  �1  ��  �  �'	    t�  �eX  ͛  �FY  ��  �	   �  ��  �  ��  
�x  ��  ��  ��  a}  ��   ��  ��X  ��  (��Y  f�  �'	   �  �M	  b�  �M	  ��  �M	  �1  ��   S  ��  " �  �SY  +4R  H	 �F     �  �Y  L   � 	�Y  )ɟ  ��Y  	 �F     �  Z  L   � 	Z  )��  �Z  	 �F     ڝ   �uZ  K�  �T   t�  �T  "  T  �0  	   ��  .Z  i�  �Z  .Z  R�  �Z  g  '	   Ja  '	   �  �Z  	�Z  ,I�  u  ?[  -��  u(�5  -� v(	  -J�  w(	  .nn y	  /�Y  z  /U  {'	  /w� |   0y�  du[  -��  d�5  /^�  fA  /ڰ  gu   ,�  Z	  \  -��  !�5  -^�  !A  /�U Z	  /ڰ  u  .nn 	  /��  	  /�@  '	  /U  '	  .p   /��    1�  Y1WD  \ ,�{  �Z	  i\  -��  �!�5  -^�  �!A  /�U �Z	  /ց  �'	  1�  � ,τ  �Z	  �\  -��  �!�5  -^�  �!A  /�U �Z	  /ց  �'	  1�  � 2W�  BZ	  �DA           �F^  3��  B �5  �� �� 3^�  C A  ;� 1� 4�U GZ	  �� �� 4ڰ  Hu  �� �� )ց  I'	  �H5�  s�EA     68EA     1       �]  7cur cL=  (� "� 4��  dL=  u� s� 8\EA     �� 9Uv   :�DA     �]  9Us 9T tvc9Qv 9R�H ;EA     �� �]  9U| 9T49Q09X09Y�D ;0EA     Ă ^  9Uv  ;qEA     т +^  9Uv  8�EA     ��  9Us 9Tv   0�  #o^  -��  #�5  /^�  %A   <��  �'	   A     �       �_  =��  �#�5  U>J�  �#	  �� �� =�p  �#R=  Q?r� �'	  2� &� ?{� �'	  �� �� @p �  �� �� ?��  �  h� ^�  A�w  @Z	  �_  B��  @!�5  B^�  A!A  C�U CZ	  Cց  D'	  Cm�  E	  D�  �ECޜ  �'	  C�, �`/  C��  �`/  Fpos �	  C�  �	  C�  ��  EC  �	     26�  �Z	  �9A            �`  3�  ��  �� �� G�9A     ނ  H�|  �A            �3`  I��  �>  U 2[�  �Z	   A     
       �{`  I��  �>  U4K ��M  &� $�  2�w  Z	  A     9      ��b  3ֳ  KB  O� I� 3n�  �  �� �� 4��  �5  6� 2� 4I�  E  p� l� Jk �A      �A     "       5 `a  K k �� �� Kk �� �� L�A     "       M*k � � M6k J� F�   Jk �A      �A            8!�a  K k �� �� Kk �� �� L�A            M*k �� �� M6k #� �   Nk �A      @V  ;$b  K k `� ^� Kk �� �� O@V  M*k �� �� M6k � �   Nk A      pV  R#zb  K k V� T� Kk }� {� OpV  M*k �� �� M6k �� ��   PqA     � P�A     � P�A     � PA     �  H7�  ��A            �c  3��  �<  3� -� 4ֳ  �KB  �� � 8�A     ed  9Us   2T{  �Z	  �A     !       �cc  I��  �<  U4ֳ  �KB  �� �� Q�U �Z	    ,b�  �Z	  �c  -ֳ  �$KB  -ؘ  �$�  /�U �Z	  1�  �E.i �	    ,Ά  )Z	  Yd  -�  )#<  -ؘ  *#�  /�U ,Z	  /ֳ  -KB  /��  .�5  /ڰ  /u  /��  1�  /}` 2Yd  1�  �RId  /��  R_d   E/�-  |m    f,  �P  H@�   �A     �       �[e  3�   #<  �� �� 4ֳ  KB  N� H� 4��  �5  �� �� 4ڰ  u  �� �� P�A     ��  ;A     �� �d  9Uv  ;3A     �� e  9Uv  ;SA     `v  .e  9Us� ;bA     �� Fe  9Uv  8|A     �� 9Uv   2�  �Z	  p(A     �      ��g  3ֳ  �KB  �� �� 3ؘ  ��  P� L� 4��  ��5  �� �� 4BJ  �!>  �� �� 4�U �Z	  � �� 7i �	  =� 7� 41� �M	  �� �� Jk �(A      �(A            �uf  S k Kk �� �� L�(A            M*k �� �� M6k 9� 5�   JX�  1)A      1)A            ��f  K��  v� t� K}�  �� �� Kq�  �� �� Ke�  �� ��  J2�  A)A      A)A            �g  KK�  � 	� K?�  1� /�  JO�  i*A      i*A     �       �tg  Kj�  V� T� K]�  {� y� Li*A     �       Mw�  �� ��   N��  +A      `Y  ��g  K��  �� �� K��  � � K��  >� <� O`Y  M��  c� a�   ;�(A     ��  �g  9U| 9T} 9Qv  TB+A     9U|   ,Pz  HZ	  oh  -ֳ  HKB  -ؘ  I�  /��  K�5  /BJ  L!>  /�U MZ	  E/I�  cE  /��  d_d    U�  �9A           �8j  3�H  h  �� �� 4��  �5  �� �� 4ڰ  u  Y� W� 4^�  A  ~� |� 4�i  ;I  �� �� NF^  :A      P[  Hi  KT^  �� �� OP[  Ma^  �� �� 80:A     � 9Ts�	   N?[  B:A      �[  �i  KM[  � � O�[  MZ[  9� 7� Mg[  ^� \� PS:A     �� 8m:A     � 9U| 9Ts�
   ::A     �i  9Us  ;|:A     �� �i  9U}  ;�:A     � j  9Uv 9Ts� ;�:A     � #j  9Uv 9Ts� 8�:A     ��  9Us   2K�  ^Z	  ��A     u
      ��s  3^�  ^ A  �� �� 3�H  _ h  � �� 3�  ` 	  �� �� 3�[  a 	  &� � 3\  b �  �� �� 4�U dZ	  �� �� 4�-  em  � � 4�i  f;I  O� A� 4��  g�5  �� �� 1�  �1��  �VPr  uk  4�' �	  �� �� ;_�A     ��  `k  9Us  8q�A     � 9Us   N`t  ��A      �o  �
�m  Krt  ;� /� W�u  ԥA     ,       
�k  S�u  LԥA     ,       X�u  8�A     � 9U| 9T~    Y�t  �A      0p  
K�t  �� �� O�p  M�t  T� H� Z�t  ��~M�t  �� �� M�t  �� �� M�t  .�  � M�t  �� �� Mu  ~� |� Mu  �� �� YDu  �A      �p  �Kau  �� �� KUu  � � Nlu  +�A        q  tm  K�u  b� V� K}u  �� �� O q  M�u  &� "� M�u  d� \� M�u  �� �� ;;�A     Ă .m  9U} 9T|  ;\�A     � Fm  9U}  ;��A     )� ^m  9U}  8��A     т 9U}    T�A     9Us 9R0     Nu[  ��A      @q  �o  S�[  K�[  1� )� O@q  Z�[  ��~M�[  �� �� M�[  �� �� M�[  `� V� Z�[  ��~M�[  �� �� M�[  "� � M�[   � �� [\  �A     [\  @�A     :̧A     dn  9Us 9Txmdh9Q 9R��~ ;
�A     6� �n  9U 9Q}  ;��A     �� �n  9U| 9T19Q09R	��~�
��9X09Y��~ ;M�A     � �n  9U��~9T}  8ìA     �� 9U| 9T19Q09R09X09Y��~   Ni\  �A      �q  ��o  S�\  K{\  � {� O�q  M�\  �� �� Z�\  ��~[�\  ��A     :4�A     �o  9Us 9Tmgpf9Q��~9R��~ 8��A     6� 9U��~9Qs�   N\  R�A     	 �q  �Pp  S8\  K+\  � � O�q  ME\  \� T� ZR\  ��~[_\  ��A     :j�A     1p  9Us 9Tperp9Q��~9R��~ 8��A     6� 9U��~9Qs�   \�s  r  �Mq  S�s  Or  M�s  �� �� X�s  Zt  ��~Mt  �� �� Mt  7� /� M&t  �� �� ]3t  �A     D       +q  M4t  )� '� ZAt  ��~;��A     C� q  9Us 9T} 9Q��~9R8 8�A     P� 9U��~9T	��F       8��A     o^  9Uu 9T~ 9Qq    J[] ��A      ��A     <       ��q  Ki] N� L�  N_  `�A      �r  �s  S-_  K!_  y� q� O�r  M9_  �� �� ZE_  ��~MQ_  o� c� []_  3�A     ^e_  �r  }r  Mf_  �� �� Mr_  H� D� M~_  �� ~� M�_  �� �� M�_  �� �� M�_  _� [� ]�_  L�A     "       fr  M�_  �� ��  8@�A     [� 9U��~  :z�A     �r  9Us 9Tfylg9Q��~9Rs�	 :��A     �r  9Us 9Tacol9Q��~9R��~ ;)�A     6� �r  9U��~9Qs�	 8��A     [� 9U��~   ;�A     h� .s  9T	��F      ;��A     u� Ks  9U~ 9T0 :�A     zs  9U~ 9Ts 9Q��~�9R| 9X}  :��A     �s  9U��~9Ts 9Q��~�9R| 9X}  8�A     �\  9Us 9T��~  ,�  �  Pt  -�H  $h  /�Y  �  /��  �5  /�p  	  .i '	  /x '	  //� 	  E/�U /Z	  .buf 0Pt    �   `t  L    ,Ŕ  ��  �t  -��  �!h   ,�}  �  u  -��  *�5  )x  !/u  	`�F     /�  �'	  /��  �4u  /�  ��  /�  ��  /��  �#�  .i ��  .j �S   .k �S    �Z  /u  L   L    	u  S   Du  L    A�  �'	  lu  B��  �$�5  _i �$�   A
�  �h  �u  B^�  �&A  B��  �&'	  C�U �Z	  C�  �h  Fi �	   A��  ��  �u  B}W �1  (�  �v  	�F     Fnn �
S    �   v  L   L    	�u  A7�  uZ	  `v  Bڰ  u#u  B�P  v#�  B�K  w#�  B�y  x#>  C�U zZ	   `��  G@A     �       �w  >�y  G$>  �� �� ?ڰ  Iu  � � ;]A     �� �v  9Uv  ;qA     �� �v  9Uv  ;�A     �� �v  9Uv  ;�A     �� w  9Uv  8�A     �� 9Uv   aN�  iZ	   �A     	2      ��  bexc i!>  f� 2� 4ʠ  k'	  u� g� 4�  l'	  � � 7i m�  8� 2� 5@�  �!?�A     5�  �!?�A     5J�  �!��A     5O�  �!.�A     V u  �  4E�  X"-  �� �� 4�|  Y�  �� �� N��  ��A      �v  � �x  K��    K��  L B O�v  MǪ  � � MԪ  < 4 Mߪ  � � M�  � � M��  d X M �  � � [�  O�A     :��A     �x  9U  T��A     9U    N��  e�A       w  �y  K��  "
 
 K��  \
 X
 O w  M	�  �
 �
   Nܿ  ��A      0w  W 3{  K��  �
 �
 K�  N F O0w  M�  � � M�    M�  � � ^E�  �w  �z  MF�  � � MS�  � � ]`�  C�A     Z       ^z  Xa�  Nk C�A      �w  z  K k U S Kk � x O�w  M*k � � M6k A =   Nk l�A      px  �Mz  S k Sk Opx  M*k � | M6k � �   T��A     9U   Jk ��A      ��A            x�z  K k   � Kk ' % L��A            M*k N J M6k � �   T��A     9U   ]%�  ��A     .       !{  M*�  � � M7�  � � T�A     9U   TW�A     9U    J��  �A       �A     	       �u{  K��    K��  = ;  N�  ��A      �x  T!�{  K+�  d ` K�  � � O�x  M8�  � � ME�    MR�  h ^   N^�  �A       y   �|  Ky�  � � Kl�  2 , O y  Z��  ��Z��  ��~Z��  ��~Z��  ��~M��   { Mĺ  � � ;��A     �  �|  9U 9T��~9Q��~9R��9X��~ 8��A     ̻  9Uu 9Ty 9Qq 9Rr 9Xx    JF�  j�A      j�A            � }  Ka�    KT�  C A 8��A     ��  9Uu 9Tt   N��  ��A      `y  _ T}  K��  h f K��  � � T��A     9U   N�  ��A      �y  ��  K�  � � K�  � � O�y  M,�    M9�  7 5 ME�  ] [ MQ�  � � M]�  � � Mi�  � � Mv�  ; 1 M��  � � M��  � � M��  b \ M��  � � M��  � � Mµ   � Mϵ  a _ Xܵ  ;��A     �� q~  9U��~9T��~9Q@ ;��A     �� �~  9U��~9T��}9Q@ ;νA     �� �~  9U��~9T��}9Q@ ;�A     �� �~  9U��~9T��~| 9Q@ ;G�A     ��   9U	��~��~9T��~9Q@ ;c�A     �� D  9U| ��~9T��}9Q@ ;{�A     �� j  9U| 9T��~9Qv  8��A     �� 9U| 9T��~9Qv    J��  ��A      ��A            ��  K��  � � 8ƾA     h�  9Uu   J��  ׾A       ׾A     !       ~&�  K��  � � K��  � � K��  � �  J��   �A        �A     !       zu�  K��  � � K��  � � K��     J}�  !�A      !�A     1       �.�  K��  ? = K��  ? = K��  d b ck !�A      !�A     "       3"K k � � Kk � � L!�A     "       M*k � � M6k      J��  V�A       V�A            �p�  K��  X V K��  } {  JC�  f�A       f�A            ���  KQ�  � � K^�  � �  Jl�  {�A      {�A     !       ��  Kz�  � � L{�A     !       M��      J��  ��A      ��A            �;�  K��  L J  J��  ��A      ��A            �p�  K��  q o  J��  ĿA      ĿA     S       dނ  K��  � � LĿA     S       M�  � � M�  � � M#�      J��  �A      �A     3       vՃ  K	�  , * K��  Q O L�A     3       M�  x t M!�  � � M,�  � � Y'�  �A      �y  �KQ�  8 2 KQ�  8 2 KE�  � � K9�  � � O�y  X\�  8E�A     �� 9Q�9R�dQ�  �     J8�  J�A      J�A     =       r̄  KS�    KF�  2 0 LJ�A     =       M`�  Y U Mk�  � � Mv�  � � Y'�  R�A       z  �KQ�    KQ�    KE�  l h K9�  � � O z  X\�  8t�A     �� 9Q�9R�dQ�  �     J��  ��A      ��A     $       n)�  K��  � � K��      8��A     1�  9U 9R�  J��  ��A      ��A     >       i��  K��  8  6  K��  ]  [  ;��A     1�  ��  9U 9R� 8��A     h�  9U   J��  ��A      ��A     5       A ��  K��  �  �  K��  �  �  L��A     5       M��  �  �    J��  �A      �A     5       = `�  K��  ! ! K��  ,! *! L�A     5       M��  Q! O!   Jg�  h�A       h�A     u        *�  K��  x! t! Ku�  �! �! Lh�A     u       M��  �! �! M��  " " M��  C" A" :��A     �  9U  :��A     �  9U 9Ts  T��A     9U 9T� 9Qv 
��   N��  ��A      0z  ��  K��  l" f" O0z  M��  �" �" c��  ��A       ��A     !       _K��  e# a# K��  �# �# K��  �# �# L��A     !       X��  8��A     �n 9U 9Tt 9Qq      N��  @�A      pz  � p�  K��  �# �# K��  $$  $ Yf�  Q�A       �z  �K��  b$ Z$ K��  �$ �$ Kx�  H% D% O�z  M��  �% ~%    N��  ��A      �z  6!ƈ  K��  �% �% O�z  M��  & & M��  8& 6& M��  ]& [&   J��  ��A      ��A     (       � �  K��  �& �& K��  �& �& T��A     9U   J$�  ��A      ��A            � M�  K2�  �& �&  J�  ��A      ��A     !       � ��  K�  �& �&  J]�  ��A      ��A            !ĉ  Kk�  ' ' Kk�  ' '  Jy�  �A      �A            !�  K��  <' :' K��  <' :'  JF�  0�A      0�A     x       F!��  Ka�  a' _' KT�  �' �' L0�A     x       Mn�  �' �' My�  �' �' M��  �' �'   JA�  ��A      ��A            � Ê  KO�  �( �( KO�  �( �(  Jo�  ��A      ��A            � �  K��  �( �( K}�  �( �(  J��  ��A      ��A     0       � b�  K
�  ) ) K��  )) ') 8��A     ��  9U 9T
A-  J{�  �A       �A     %       ���  K��  N) L) K��  N) L) K��  s) q)  J��  ,�A      ,�A            , �  K��  �) �) K��  �) �)  N�  G�A       {  ( u�  K��  �) �) O {  M�  �) �) M�  * * e�  :��A     S�  9U  T�A     9U 9Ts 9Qv 
��   N��  �A      0{  $ �  Kҹ  [* W* KŹ  �* �* O0{  M߹  �* �* M�  + + :��A     ݌  9U  :��A     ��  9U 9T�9Q|  T��A     9U 9T�9Q|    N��  ��A      `{   �  K�  D+ @+ K�  ~+ z+ O`{  M"�  �+ �+ M.�  �+ �+ M:�  ., (, MG�  {, w, eT�  ;H�A     ��  ��  9Uy  ;[�A     ��  ��  9Uy  ;-�A     ̻  �  9Uu 9Qq 9Rr 9Xx  8��A     ̻  9Uu 9Qq 9Rr 9Xx    Nк  C�A       �{   �  K�  �, �, K޺  �, �, O�{  Z��  ��Z�  ��~Z�  ��~Z�  ��~M)�  7- 3- X6�  MC�  q- m- MP�  �- �- M]�  �- �- ;��A     �  ݎ  9U 9T��~9Q��~9R��9X��~ 8��A     ̻  9Uu 9Ty 9Qq 9Rr 9Xx    Ni�  "�A      �{   ҏ  Kw�  I. G. O�{  Z��  ��Z��  ��~Z��  ��~Z��  ��~M��  p. l. [»  ^�A     ;X�A     �  ��  9U 9T��~9Q��~9R��9X��~ 8��A     ̻  9Uu 9Qq 9Rr 9Xx    N��  ��A       |  5 (�  K��  �. �. K��  �. �. O |  M��   / / M��  v/ n/   N�  U�A      0|  1 ]�  K �  �/ �/ K�  B0 :0 O0|  M�  �0 �0 M�  �0 �0 M'�  �1 ~1 M4�  �1 �1 MA�  ;2 12 [N�  �A     ]W�  ��A     -       �  MX�  �2 �2 T��A     9U 9T|   :��A     �  9U  :��A     �  9U  :�A     :�  9U 9T� 9Qs 
�� P��A     ��  8�A     ��  9U|    JB�  %�A      %�A     �       9 	�  K]�  3 3 KP�  43 23 L%�A     �       Mj�  ]3 W3 Mu�  �3 �3 c��  {�A      {�A            �K��  �3 �3 K��  �3 �3    J�  ��A      ��A     0       � f�  K3�  4 4 K&�  74 54 8��A     ��  9U 9T
 @  N��  ��A       �|  ���  K��  ^4 Z4 K��  �4 �4  Jx�  ��A      ��A            � �  K��  �4 �4 8��A     �� 9Q@  N�   �A      �|  �ړ  K�  �4 �4 K�  _5 W5 O�|  M+�  �5 �5 M6�  &6  6 MC�  �6 �6 [P�  G�A     ^Y�   }  n�  MZ�  ^7 Z7  Y��  ��A      0}  K��  �7 �7 K��  �7 �7 K��  #8 8 O0}  X��  8��A     �n 9U 9Tt 9Qq      J#�  �A       �A     9       �H�  K>�  [8 Y8 K1�  �8 ~8 L�A     9       MK�  �8 �8 MX�  �8 �8   Jq�  U�A      U�A     �       R �  K��  9 9 K�  +9 )9 LU�A     �       M��  P9 N9 M��  u9 s9 :��A     Ȕ  9U  T��A     9U 9T�9Qs 
��   N��  ��A      `}  N e�  K��  �9 �9 K��  �9 �9 O`}  M��  : : M��  c: ]: :�A     S�  9U  T!�A     9U    N�  '�A      �}  I ��  K�  �: �: K�  �: �: O�}  M,�  �: �: TB�A     9U    Jl�  O�A      O�A     (       E /�  K��  ; ; Kz�  B; @; LO�A     (       M��  g; e; Tn�A     9U    N��  w�A      �}  2!��  K��  �; �; K��  �; �; O�}  M��  C< =< M��  �< �< 84�A     7�  9Uu    N��  c�A      ~  ��  K�  �< �< K�  = = O~  M �  }= y= M+�  �= �= M8�  > > 8�A     7�  9Uu    J^�  ��A      ��A     �       .!~�  Ky�  >> <> Kl�  c> a> L��A     �       M��  �> �> M��  �> �>   N5�  ��A      `~  *!l�  KP�  �> �> KC�  j? d? O`~  M]�  �? �? Mh�  �@ �@ Ms�  �A �A M~�  7B /B M��  �B �B M��  FC >C ^��  �~  .�  M��  �C �C M��  )D !D  N'�  8�A      �~  ���  KQ�  �D �D KQ�  �D �D KE�  rE jE K9�  �E �E O�~  X\�  8��A     �� 9Q�9R�dQ�  �   ^��     ֘  M¿  8F 2F Mο  �F �F  N'�  ��A      `  �V�  KQ�  �F �F KQ�  �F �F KE�  HG @G K9�  �G �G O`  X\�  8��A     �� 9Q�9R�dQ�  �   8��A     h�  9Uu    J��  ��A       ��A            ���  K�  
H H K�  /H -H  J��  ��A      ��A            ��  K��  TH RH K��  TH RH  Ni�  G�A      �  ��  K��  }H wH Kw�  �H �H O�  M��  I I M��  kI eI M��  �I �I [��  G�A     ]��  w�A     3       ��  M��  �J �J  Y��  �A      �  �K��  �J �J K��  K  K K��  >K :K O�  X��  8�A     �n 9U 9Tt 9Qq      J�  /�A      /�A            � &�  K�  vK tK  N-�  ��A      �  � O�  K;�  �K �K  J��  `�A      `�A            ^!��  K�  �K �K  N��  y�A      @�  � �  K�  �K �K K�  #L L O@�  M�  tL lL M)�  �L �L 8��A     7�  9Uu    J��  ��A      ��A     #       { #�  K��  M M  J��  ��A      ��A     #       w X�  K��  5M 3M  J�  �A      �A     #       s ��  K�  ZM XM  J'�  0�A      0�A     #       o   K5�  M }M  N��  S�A      p�  k �  K��  �M �M  JE�  e�A      e�A            g  �  KS�  �M �M  J@�  r�A      r�A            � U�  KN�  �M �M  J\�  ��A      ��A     %       � ��  Kj�  N N  J��  ��A      ��A            � ��  K��  8N 6N  J��  ��A      ��A             ��  K��  ]N [N  N��  w�A      ��  � �  K�  �N �N  J!�  ��A      ��A            �_�  K/�  �N �N K<�  �N �N  JJ�  ��A      ��A            ���  KX�  �N �N Ke�  O O  Js�  ��A      ��A            ��  K��  ;O 9O K��  `O ^O  W��  �A     D       �9�  S��  L�A     D       M��  �O �O 89�A     7�  9Uu    N�  W�A       Ѐ  �o�  K��  �O �O K�  P P  N�  ��A        �  ���  K'�  OP KP K�  �P �P  N��  f�A       0�  �۟  Kվ  �P �P KȾ  �P �P  J��  ��A      ��A            ��  K��  5Q 3Q K��  5Q 3Q  Ja�  �A      �A            c R�  Ko�  ZQ XQ  N��  �A      `�  !��  KŽ  �Q }Q O`�  Mҽ  �Q �Q e߽    JT�  ��A      ��A     #       >!Ƞ  Kb�  #R !R  J��  ��A      ��A     �       ���  KѴ  LR FR KĴ  �R �R L��A     �       M޴  �R �R M�  �R �R M��  US OS :�A     U�  9U  :?�A     ��  9U 9T�9Q| 
��9Rs  TS�A     9U 9T� 9Qv 
��9Rs    J8�  \�A      \�A     Q       � ]�  KS�  �S �S KF�  �S �S L\�A     Q       M`�  �S �S Yk m�A      ��  kK k T T Kk 9T 7T O��  M*k aT ]T M6k �T �T     N�  ��A      Ё  %!��  K-�  �T �T K �  U U OЁ  M:�  WU SU   J�  {�A       {�A            B!�  K��  �U �U K�  �U �U  N#�  ��A       �  !K�  K>�  �U �U K1�  V V O �  MK�  MV KV MV�  rV pV Ma�  �V �V   Nm�  ��A      0�  !��  K��  �V �V K{�  W 	W O0�  M��  EW CW M��  jW hW M��  �W �W   J��  X�A       X�A            � ��  K��  �W �W K��  �W �W K�  �W �W  JI�  o�A      o�A     !       � T�  Kd�  X X KW�  8X 6X T�A     9U 9Q0  Jr�  ��A      ��A     *       � ��  K��  ]X [X K��  �X �X T��A     9U 9Q0  N�  ��A       `�  ��  K0�  �X �X K#�  �X �X O`�  M=�  Y Y MH�  UY SY P��A     ��   J��  �A      �A            � C�  K��  zY xY  J��  �A      �A            � x�  K��  �Y �Y  N��  4�A      ��  � ¥  K��  �Y �Y K��   Z �Y 8��A     �� 9T@  Jp�  S�A      S�A            :!��  K~�  8Z 6Z  J�  f�A      f�A            � 9�  K �  ]Z [Z K-�  �Z �Z  J�  ��A      ��A     C       l!��  K�  �Z �Z K�  �Z �Z L��A     C       M+�  �Z �Z M6�  [ [   J��  -�A      -�A     t       j!S�  K��  R[ P[ K��  w[ u[ L-�A     t       M��  �[ �[ M��  �[ �[ c��  j�A      j�A            �K��  \ �[ K��  \ �[    ;�A     �  k�  9Uu  ;��A     �  ��  9U 9Tv  ;[�A     �  ��  9U  ;��A     f�  ��  9U  ;��A     �  ѧ  9Uu  ;2�A     '�  �  9U 9Tv  8��A     bt 9U dO�  v   VЂ  Ũ  7def y!R  =\ 9\ 4��  z!R  �\ �\ O �  4�  �!�  �\ �\ Y��  ��A      p�  �!K��  $]  ] K��  ]] [] K��  �] �] Op�  X��  8ջA     �n 9U 9Tt 9Qq      NL�  o�A      �t  ���  Kg�  �] �] KZ�  (^ �]  8o�A     h�  9Uu   R  HY�  #�PA     �       ���  fexc # !>  U7def %R  �_ �_ 4��  &R  2` *` O^  4��  -�  �` �` Y��  QA      @^  =	K��  �` �` K��  0a ,a K��  la fa O@^  X��  80QA     �n 9Uu 9Tt 9Qq      0ٔ  �  -E�  "-   0��  �^�  gexc �%!>  -E�  �%"-  /�  �	  /Ԛ  �   .i �	   0�y  ��  gexc  !>  -E�   "-  .K 	  /K �M   0�  ��  gexc �!>  -E�  �"-  /��  �'	  .k �'	  .A �'	  .C �'	  .P �'	  .B �	  1WD  � HN�  A     �      ��  bexc !>  �a �a 3E�  	"-  Qb Ib 4��  '	  �b �b 7k '	  c �b 7A �  �c �c 7C '	  d d 7P '	  �d �d 7B 	  e e 5WD  ��A     :$A     ��  9Us  TA     9Us 9Ts�   H��  ���A           ���  bexc �!>  \f Nf hV �uZ  ��4�� ��  �f �f 4�>  �	  ^g Zg 4t�  �	  �g �g 4��  �	  �g �g 4��  �	  �g �g 4c �	  ch Wh 42 ��  �h �h N��  ��A       �k  ���  K�  Pi Ji K�  �i �i Kٯ  j �i Kͯ  Tj Pj K��  �j �j O�k  X��  X
�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  8L�A     �x 9U��9X|    J��  ��A       ��A     7       �i�  K�  �j �j K�  k k Kٯ  Ck Ak Kͯ  jk fk K��  �k �k L��A     7       X��  X
�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  8ʃA     �x 9U��9T
��9Qv 9R 9Xs    J��  ۃA       ۃA     *       �8�  K�  �k �k K�  "l  l Kٯ  Il El Kͯ  �l �l K��  �l �l LۃA     *       X��  X
�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  8�A     �x 9U��9Qs9R 9Xs    YͰ  �A        l  �K۰  �l �l K۰  �l �l K �  ?m ;m K��  ym um K�  �m �m O l  M�  n n M�  �n n    0��  Ͱ  -�  (�Z  gp1 (	  gp2 (	  -~�   (	  -�|  !(	  .i #	  /��  $@	  /��  $@	  /��  $@	  /��  $%@	  /ɀ  $+@	  /΀  $1@	  /��  $7@	  /P�  $?@	  R��  /V�  3@	  /�  4	   R��  .x M@	   E/1� ^M	  /��  _�  E.x e@	     0$�  #�  -�  "�Z  gp1 "	  gp2 	"	  gp 
"	  .i 	  .dx @	   0��  �f�  gexc �!>  -E�  �"-  /c ��  /�� ��   HG�  B�A           ���  bexc B!>  �n �n 4x  D@	  uo ko 4py  D@	  �o �o 4��  ET  Cp =p 4��  FT  �p �p 4 �  G	  �p �p 5WD  �yA     V�W  ߲  7vec z�  Mq Cq Nk -A       X  }��  K k Ws Ss Kk �s �s O X  M*k �s �s M6k ?t ;t   Nk TA      �X  �β  S k Sk O�X  M*k ~t zt M6k �t �t   T{A     9Us   V�V  }�  4c �	  u �t 4��  �@	  _u Uu 4��  �@	  �u �u /��  �'@	  6aA     _       �  7vec ��  )v v Nk aA      �V  ���  K k �w �w Kk �w �w O�V  M*k x x M6k Zx Vx   Nk �A      pW  ���  S k Sk OpW  M*k �x �x M6k �x �x   T�A     9Us   :�A     �  9Us  :�A     3�  9Us  :A     X�  9Us 9Ts�9Q 
�� 8�A     �� 9U~ 9T��9Q��  :!A     ��  9Us  :PA     ��  9Us  T�A     9Us   0��  �  gexc !!>  -E�   !"-  .p1 "�  .p2 "�  /d�  #@	   0��  ��  gexc �!>  -E�  �"-  /c ��  .a0 ��  .a1 ��  .b0 ��  .b1 ��  //}  �@	  /��  �@	  .dx �@	  .dy �@	  .dax �@	  .day �@	  .dbx �@	  .dby �@	  .val �@	  .R ��   0X�  �'�  gexc � !>  /c ��  /d�  �@	  1WD  � Hh�  �0A     �      �4�  bexc �!>  y y 3E�  �"-  �y ~y 4c ��  �y �y 4)�  �'	  z z 4��  �@	  �z �z 4d�  �@	  +{ '{ 4��  �@	  k{ a{ 4��  �@	  �{ �{ 4�}  �@	  -| +| 4\�  �@	  T| R| 4�� �@	  �| y| 5WD  oSA     Nf�  �A      V  "��  K��  �| �| K��  I} ?} Kx�  �} �} OV  X��    :�A     ��  9Us  ;A     ��  ��  9U}  ;,A     ��  з  9U}  :iA     �  9Us  :�A     ��  9Us  :A     �  9Us 9T}  TLA     9Us 9Ts�9Q~ 
��  0ۃ  ��  gexc �!>  -E�  �"-  /c ��  /��  �@	  /d�  �@	  /\�  �%@	  1WD  yR��  /<  T  /"<  T   E/<  #T  /"<  $T  E.vec /�     0	�  �g�  gexc �!>  -E�  �"-  /)�  �'	  /c ��  /d�  �@	  /��  �@	  /�}  �@	  1WD  �E/�� �@	    0��  K��  gexc K!>  -E�  L"-  /c N�  /��  O@	  /d�  P@	   0��   ��  gexc  !>  -E�  "-  /c �  /d�  @	   0��  `^�  gexc `!>  -E�  a"-  .dx c@	  .dy c@	  /c d�  /��  i�  1WD  � 0�}  0к  gexc 0!>  -E�  1"-  .zp 3>  /�}  4�  .dx 5@	  .dy 6@	  /��  8�  .i 8�   0�}  �i�  gexc �!>  -E�  �"-  .zp �>  /�}   �  .dx @	  .dy @	  /2 �  /�7 �  /�k �  /��  �  .i $�   0sw  �̻  gexc �!>  .zp �>  /�}  ��  .dx �@	  .dy �@	  /c ��  1WD  � 0k�  ��  gexc �#!>  -c �#�  gdx �#@	  gdy �#@	  -��  �#�   2�z  j�  �A     �      ��  bexc j/!>  �} �} bx k/�  _~ Y~ by l/�  �~ �~ 3�y  m/>  D > 3�}  n/�2  � � 7zp p>  � � 7p q�  �� �� 7d r@	  �� �� :�A     �  9Us  ;�A     �� �  9U}  8�A     �� 9U}   @	  0�~  Jm�  gexc J"!>  -E�  K""-  .I M�  .K M�  .L M�   0S�  $��  gexc $!!>  -E�  %!"-  .I '�  .K '�  .L '�   0��  ��  gexc �!>  /c ��  1WD   0�  ��  gexc �!!>  -E�  �!"-   0e�  �F�  gexc �!!>  -E�  �!"-  .A �	   0�|  k��  gexc k!!>  -E�  l!"-  .K n'	  .L n'	  .Kf n'	   0e�  H��  gexc H!>  -E�  I"-   0��  *�  gexc *!>  -E�  +"-   0��  �  gexc !>  -E�  "-   0��  �5�  gexc �!>  -E�  �"-   0�  �ܿ  gexc �!>  -E�  �"-  .A �	  .B �	  .C �	  .p1 ��  .p2 ��  /�|  ��  R��  .v1 �T  .v2 �T   E.v1 �T  .v2 �T    0�  Mq�  gexc M!>  -E�  N"-  .K P�  .L P�  .D Q@	  RE�  /<  hT  /"<  iT   E/<  pT  /"<  qT  E.vec |�     0?�  "��  gexc "!>  -E�  #"-  .K %	  .L &�   0-�  ���  gexc �!>  -E�  �"-  .L �'	  .R  @	   0{  ��  gexc �!!>  -E�  �!"-   0{�  �A�  gexc �!>  -E�  �"-   0v�  �]�  gexc �!>   0Y�  �y�  gexc �!>   0��  ���  gexc �!>   0�  ���  gexc �!>   0��  ���  gexc �!>   0�  ���  gexc �!>   0��  t�  gexc t!>  -E�  u"-   0{�  f;�  gexc f!>  -E�  g"-   í  Y0J�  La�  gexc L !>   0�  ?}�  gexc ?!>   0��  0��  gexc 0!>  -E�  1"-   0'�  "��  gexc "!>  -E�  #"-   07�  ��  gexc !>  -E�  "-   0��  !�  gexc !>  -E�  "-   0��  �J�  gexc �!>  -E�  �"-   0��  �s�  gexc �!>  -E�  �"-   0��  ���  gexc �!>  -E�  �"-   0��  ���  gexc �!>  -E�  �"-   0=|  ���  gexc �!>  -E�  �"-   0ۛ  �8�  gexc �!>  -E�  �"-  .S ��  .X �	  .Y �	   0�  ���  gexc �!>  -E�  �"-  .S ��  .X �	  .Y �	   0?{  |��  gexc |!>   0��  h��  gexc h!>  -E�  i"-   0ގ  S��  gexc S!>  -E�  T"-   0��  /1�  gexc /!>  .AA 1�  .BB 1�  /�|  3�   , �  ��  ��  gexc �!>  -�{  ��  -�{  ��  gVec ���  .A �	  .B �	  .C �	  .p1 �T  .p2 �T  /�|  ��   �	  0W}  ��  gexc �!>  -E�  �"-  .L ��  .K ��   0�|  �B�  gexc �!>  -E�  �"-  .L ��  .K ��   0r~  ���  gexc �!>  -E�  �"-  .L ��  .K ��   0	~  z��  gexc z!>  -E�  {"-  .L }�  .K }�   0��  (�  gexc (!>  -E�  )"-  .def +R  /��  ,R   0��  �i�  gexc �!!>  -E�  �!"-  .F �'	  /��  ��  .def �R  1WD  E/��  �R    0*�  r��  gexc r!>  -E�  s"-  .F u'	  /��  v�  .def wR  1WD  �E/��  �R    0�  A��  gexc A!>  /��  C�   0�  F�  gexc !>  -E�  "-  .n '	  .rec R  /��  R   0��  �o�  gexc �!>  -E�  �"-   04�  ���  gexc �!>  -E�  �"-   0�{  ���  gexc �!>  -E�  �"-   i*�  �0a�  ���  gexc �!>  /�w  �	   0��  p7�  gexc p!>  -E�  q"-  /�w  s	  .Out t�   26�  O�  �A     �       �{�  fexc O!>  U5<�  c�A      0@�  A��  gexc A!>  -E�  B"-   0��  $��  -E�  $"-  .A &	  .B &	  .C &	   0J�  
�  gexc 
!>  -E�  "-  .L 	   0��  �T�  gexc �!>  -E�  �"-  .L �	  .K �	   0ܒ  �p�  -E�  �"-   0�  ���  -E�  �"-   0F  ���  gexc �!>  -E�  �"-   0��  ���  gexc �!>  -E�  �"-   0�|  ���  gexc �!>   iˉ  �09�  v8�  gexc v!>  -E�  w"-  .I y'	   0�  _l�  gexc _!>  -E�  `"-  .I b'	   0H�  H��  gexc H!>  -E�  I"-  .I K'	   01�  1��  gexc 1!>  -E�  2"-  .I 4'	   0֗  �  gexc !>  -E�  "-  .I '	   0��  �$�  -E�  �"-   0`�  �@�  -E�  �"-   03�  �\�  -E�  �"-   0ʅ  �x�  -E�  �"-   0��  ���  -E�  �"-   0}  ���  gexc �!>  -E�  �"-   0��  ���  -E�  �"-   0�  ���  -E�  �"-   0�  ��  -E�  �"-   0��  |-�  -E�  |"-   0;�  oI�  -E�  o"-   0~�  ar�  gexc a!>  -E�  b"-   07{  S��  gexc S!>  -E�  T"-   0�  F��  -E�  F"-   0[�  9��  -E�  9"-   0P�  ,��  -E�  ,"-   0��  �  -E�  "-   0~�  '�  -E�  "-   0��  C�  -E�  "-   0ލ  �
l�  gexc �
!>  -E�  �
"-   0H�  �
��  -E�  �
"-  .L �
	   0h~  �
��  gexc �
!>   i�  �
0P�  �
��  -E�  �
"-   0�{  �
��  gexc �
!>  -E�  �
"-   0��  �
'�  gexc �
!>  -E�  �
"-   ,�  e
�  h�  gVx e
@	  gVy f
@	  gR g
��  .V i
�   H�  
�	A     �      ���  fexc 
"!>  U 2��  
@	  �	A            ���  fexc 
!>  Ufdx 
�  Tfdy 
�  Q 2��  �	@	  �	A            �5�  fexc �	!>  Ufdx �	�  Tfdy �	�  Q 2��  �	@	  p	A     8       ��  fexc �	!!>  Ubdx �	!�  3� /� bdy �	!�  p� l� c.�  p	A      p	A     5       �	Kd�  �� �� KX�  ۃ ك KL�  � 	� K@�  H� F� Lp	A     5       Mp�  q� k� M}�  Ƅ     2��  �	@	  0	A     8       ���  fexc �	!>  Ubdx �	�  � � bdy �	�  B� >� c.�  0	A      0	A     5       �	Kd�  }� {� KX�  �� �� KL�  ߅ ۅ K@�  � � L0	A     5       Mp�  C� =� M}�  �� ��    H��  _	�A     \      �L�  fexc _	"!>  U3��  `	"3	  � ӆ 3�f a	"	  Ӈ ��  0v|  '	u�  gexc '	"!>  -��  (	"�   ,��  �@	  ��  gexc �#!>  -d�  �#@	  -H�  �#@	  .val  	@	   ,r�  �@	  �  gexc � !>  -d�  � @	  -H�  � @	  .val �@	   ,,�  �@	  J�  gexc �)!>  -d�  �)@	  -H�  �)@	  .val �@	   ,�  e@	  ��  gexc e%!>  -d�  f%@	  -H�  g%@	  .val i@	   ,�  8@	  ��  gexc 8'!>  -d�  9'@	  -H�  :'@	  .val <@	   ,�  @	  �  gexc '!>  -d�  	'@	  -H�  
'@	  .val @	   ,ȇ  �@	  f�  gexc �"!>  -d�  �"@	  -H�  �"@	  .val �@	   ,{  �@	  ��  gexc �!>  -d�  �@	  -H�  �@	  .val �@	   HƑ  ��A            ��  fexc �'!>  UI�y  �'>  T3c �'�  �� �� Id�  �'@	  R H��  ��A            �q�  fexc �'!>  UI�y  �'>  T3c �'�  ۈ ׈ Id�  �'@	  R Hm�  h0A     M       ���  fexc h"!>  UI�y  i">  T3c j"�  � � Id�  k"@	  R HW�  O�A     G       �5�  fexc O"!>  UI�y  P">  T3c Q"�  U� Q� Id�  R"@	  R Hf�  )�A     �       ���  bexc )%!>  �� �� 3�y  *%>  ,� "� 3c +%�  �� �� 3d�  ,%@	  A� 5� 7v .@	  ͋ ɋ ;8A     �� ��  9U}  8nA     �� 9U}   HP�  ��A     +      ���  bexc � !>  � � 3�y  � >  �� � 3c � �  �� � 3d�  � @	  l� b� 7v �@	  � � P-A     �� 8�A     �� 9U��  ,ˎ  y�  ��  gexc y'!>  -ۚ  z'	  gaIP {'	  /x  }��   �O  ,�}  ]�  ��  gexc ] !>   HA�  D 4A     G       ���  bexc D'!>  M� G� bidx E''	  �� �� 3<v F'@	  � � ;#4A     �  u�  9Us  8.4A     � 9U}   H��  ;�A            ���  fexc ;!>  Ufidx <'	  TI<v =@	  Q H�  2P4A     0       �b�  bexc 2(!>  C� =� bidx 3('	  �� �� 3<v 4(@	  � � ;b4A     �  M�  9Us  8x4A     � 9Uv   H��  )�A            ���  fexc )!>  Ufidx *'	  TI<v +@	  Q 2ǝ  !@	  �4A     9       �g�  bexc !'!>  9� 3� bidx "''	  �� �� Nk �4A        Z  $R�  K k ِ א Kk � �� O Z  M*k t� p� M6k �� ��   8�4A     �  9Us   2Y�  @	  �A            ���  fexc !>  Ufidx '	  T 2O�  	  �4A     &       �L�  bexc +!>  �� � Nk �4A       `Z  7�  K k F� D� Kk o� i� O`Z  M*k ג Ӓ M6k � �   8�4A     �  9Us   2�~  	  �A            ��  fexc !!>  U 2]�  �	  �3A     �       �.�  bexc �"!>  [� U� L�3A     *       7x �@	  �� �� 7y �@	  �� � P�3A     ��  ;�3A     ��  �  9Uq 9Tr 0$0& P�3A     ��   ,tx  �[  ��  gax �$[  gay �$[  gbx �$	  gby �$	  /g  �.  /M  �.   28�  G[  �A            ���  fa G$[  Ubb H$	  7� 3� 7ret K.  x� p� 7tmp P.  � �  aԞ  X!>  0�A     �       �/�  3K X�M  D� @� 4ڰ  Zu  �� }� )�U [Z	  �X4BJ  ]!>  �� �� 1WD  pNK�  d�A      ��  j�  Kj�  5� 1� K]�  q� k� O��  Zw�  �\[��  ��A     ;��A     �� ��  9Uv 9T 9Q09R 9X09Y�\ 8��A     ��  9Us    8U�A     �� 9Uv 9T
P9Q�X  ,�  #Z	  O�  -BJ  ##!>   0Ɨ  ���  -BJ  �$!>  -ֳ   $KB  .i 	   2�  �Z	  0#A     7      �v�  3BJ  �$!>  Ė �� 3��  �$�5  C� 9� 3ֳ  �$KB  �� �� 7i �	  � � htmp �'	  �X4}` �Yd  }� s� 4�U �Z	  � � ;)'A     v�  U�  9T�X9Q89Rs0 8u'A     v�  9T�X9Q19Rs�  2�x  gZ	  �"A     W       �K�  3ڰ  gu  ?� ;� 3ֳ  h/  ~� x� 3��  i'	  Ι ʙ 3��  ja   � � 3�N  k'	  _� Y� )�U mZ	  �\4��  n!  �� �� 8#A     �� 9T19Rv �Q9Y�\  ,��  #Z	  ��  -BJ  #!!>  -ڰ  $!u  /�U &Z	  1;�  A `�  ��A     �       �2�  >BJ  �$!>  � �� ?ڰ  �u  h� d� ;�A     �� ��  9Uv  ;�A     �� �  9Uv  ;A     �� �  9Uv  j<A     �� 9T�U  k3  �X�  BBJ  �'!>  Bx  �'	   kǘ  ���  BBJ  �%!>  Bx  �%	  BǞ  �%a   B��  �%	   k�  ���  BBJ  �&!>  Bx  �&	  _IP �&	  C�  ���   H�  {� A     	      �5�  3��  {�5  �� �� 4ڰ  }u  � � 4E�  ~�3  4� ,� O0Y  7i �	  �� �� 4�  �	  �� �� ;� A     �� v�  9U|  ;!A     �� ��  9U|  ;!A     �� ��  9U|  ;0!A     �� ��  9U|  ;e!A     �� ��  9U|  ;�!A     �� ��  9U|  ;�!A     5�  �  9U~  ;�!A     �� �  9U|  ;�!A     �� 6�  9U|  ;�!A     �� N�  9U|  ;�!A     5�  f�  9U~  ;"A     �� ~�  9U|  ;"A     �� ��  9U|  ;-"A     �� ��  9U|  ;J"A     5�  ��  9U~  ;Z"A     �� ��  9U|  ;n"A     �� ��  9U|  ;�"A     �� �  9U|  ;�"A     �� &�  9U|  G�"A     ��   HB�  V�A     �       ��  3��  V6�5  � ݜ 3�  W6�S   � � 4ڰ  Yu  n� l� 7i Z	  �� �� ;, A     �� ��  9U}  ;G A     �� ��  9U}  ;a A     �� ��  9U}  ;� A     �� �  9U}  8� A     �� 9U}   ,e|  6Z	  o�  -��  6"�5  -�  7"R=  -Ԛ  8"�J  -��  9"�J  -;�  :"�I   2Х  �Z	   YA     �      ��  3��  �,�5  Y� O� 3x �,	  ۞ Ϟ 3Mj  �,�  m� c� 3�~  �,T  � � 30�  �,	  m� c� )�U �Z	  ��4^�  �A  � � 4ڰ  �u  �� q� 4��  �T  ~� r� 4��  �T  � � 4F�  ��  �� �� 4"	 �'	  
� � 4��  �	  �� �� 4�  �'	  B� &� 4��  �'	  � s� 4��  �'	  � � 7i �	  �� �� 7j �	  o� I� 4ܢ  �   � �� 4  �   �� �� 4͚  �   Y� M� 4E�  ��3  � � )-�  �	  ��),�  �	  ��4҅  ��2  .� � 4�|  ��2  � � 4N5  ��2  [� S� 4�  �   î �� 42�  �   P� 8� 4
�  �   p� R� 4,�  �   Ǳ �� 5}�  "#ZA     5Z  jbA     5Ob  PbA     V�`  ��  4��  	  Ҳ ʲ 4Ą  	  R� F� 4a� M	   � �� V0a  ~�  4|  \M	  b� \� 4+|  ]M	  �� �� 4|  _M	  � �� 4/|  `M	  � �� Nk peA      �a  _%3�  S k Kk �� �� O�a  M*k � �� M6k F� B�   Yk �eA       b  `%S k Kk �� �� O b  M*k ͷ ɷ M6k � �    VPb  M�  7idx ��  O� K� Nk _A      �b  � ��  S k Kk �� �� O�b  M*k �� �� M6k �� ��   ck 4_A      4_A     #       � S k Kk 8� 4� L4_A     #       M*k �� �� M6k ˹ ǹ    V`c  ��  4|  �M	  � � 4+|  �M	  �� �� 4|  ��  � � 4/|  ��  �� y�  N#�  j_A      �b  �	a�  K1�  ;� 1� K1�  ;� 1� KX�  �� �� KK�  <� 2� K>�  �� �� O�b  Me�  :� .� Mr�  Ҿ �� M�  �� �� M��  ߿ ˿ M��  �� �� M��  �� �� N��  �dA        c  4�  K�  � � K��  R� N� K��  �� �� K��  �� �� K��  � � K��  l� h� O c  X�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  Xq�  8�dA     3w 9R~ 9X��}9Yv    J��  �dA      �dA     k       B��  K��  �� �� K��  �� �� K��  �� �� K��  � � K��  :� 8� L�dA     k       M��  e� ]� X��    J��  �fA       �fA            K��  K�  �� �� K��  �� �� K��  � � K��  6� 2� K��  p� l� K��  �� �� L�fA            X�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  Xq�  8�fA     3w 9Us9T~9Qs 9R} 9X��}9Yv    Y��  �fA       0c  SK�  �� �� K��  � 	� K��  2� 0� K��  W� U� K��  ~� z� K��  �� �� O0c  X�  X�  X$�  X1�  X>�  XK�  XX�  Xe�  Xq�  8�fA     3w 9U���9T}9Qs 9R} 9X��}9Yv      ;W]A     �� y�  9U}  ;c]A     �� ��  9U}  ;�]A     �� ��  9U��~ ;�]A      ��  9U 9Ts 
��9Q��~9R��~9X��~ ;K^A     _+ ��  9U}  ;l^A     _+ �  9U}  ;EaA     �� 7�  9U��~9T��~ ;`aA     �� W�  9Us 9T��~ ;paA     �� w�  9Us 9T��~ ;�bA     �� ��  9U}  ;�bA     �� ��  9U}  ;�cA     �� ��  9U}  8�fA     �, 9U} 9Q��  ; ZA     �� �  9U| 9T@9Q09R~ 9X09Y�� ;0ZA     �� /�  9U| 9T��} ;=ZA     �� O�  9U| 9T��} ;IZA     �� n�  9U| 9Tw  ;�ZA     �� ��  9U| 9T@9Q09R~ 9X09Y�� ;�ZA     �� ��  9U| 9T19Qw 9R~ 9Xw 9Y�� ;�ZA     u� ��  9U} 9Ts  ;[A     Ă �  9U} 9Tv  ;I[A     �� D�  9U| 9T89Q09X09Y�� ;z[A     �� r�  9U| 9T89Q09X09Y�� ;�[A     �� ��  9U| 9T89Q09X09Y�� ;�[A     �� ��  9U}  ;�[A     �� ��  9U}  ;C\A     �� �  9U| 9T89Q09R~ 9X09Y�� ;s\A     �� 8�  9U| 9T89Q09R~ 9X09Y�� ;�`A     �� X�  9U| 9T��~ ;�`A     �� x�  9U| 9T��~ ;�`A     �� ��  9U| 9T��~ ;�`A     �� ��  9U| 9T��~ ;�`A     т ��  9U}  ;]bA     �� ��  9U| 9T��~ ;jbA     �� �  9U| 9T��~ ; cA     �, /�  9U} 9Q�� ;fcA     �� c�  9U| 9T89Q09R~ 9X09Y�� ;�cA     �� ��  9U| 9T89Q��~9R~ 9X��~9Y�� ;dA     �� ��  9U| 9T��~ ;*dA     �� ��  9U| 9T��~ ;EdA     �� ��  9U| 9T��~ 8OdA     �� 9U| 9T0  `  �  0P�  ��  -Mj  '�  -��  	'T  -�  
'T  -F�  '�  /�>  	  /t�  	  /ϋ  	  /z�  	  /c 	  /2 �   0r�  ���  gp1 �%S   gp2 �%S   -~�  �%S   -�|  �%S   -�  �%T  -��  �%T  .p �
S   .i �S   .out ��  .in1 ��  .in2 ��  /x  ��  /x  �"�  .d1 �(�  .d2 �,�  E/1� �M	    0d�  ���  gp1 �S   gp2 �S   gref �S   -�  �T  -��  �T  .p �S   /�� ��   2p  SZ	  =A     y      �p�  3��  S �5  � � 3^�  T A  3� !� )�U VZ	  ��4ڰ  Wu  � �� 4ah Yh  �� �� 42�  ['	  �� �� )ց  \'	  ��4��  ^	  � � 4�  _'	  �� v� 4��  a'	  �� �� 7i b	  (� � 7j b	  	� �� 4ܢ  d   :� .� 4  e   �� �� 4͚  f   Z� R� 4E�  h�3  �� �� )-�  j	  ��),�  k	  ��4҅  m�2  � �� 4�|  n�2  �� �� 4N5  o�2  �� �� 4_�  q   w� c� 4��  r   [� I� 5�  �BA     5�  �BA     V�[  ��  4��  �	  $� � 4Ą  �	  �� �� 4a� �M	  �� �� 6xCA     $       ��  48�  2M	  �� �� ck xCA      xCA            6+S k Kk  � � LxCA            M*k M� I� M6k �� ��    V \  Z�  4��  WS   �� �� 48�  XM	  �� �� Yk @AA      0\  `0S k Kk *� (� O0\  M*k W� S� M6k �� ��    ;�?A     �� r�  9U  ;@A     �� ��  9U  ;J@A     �� ��  9U~  ;k@A      ��  9U| 9Ts 
��9Q~ 9R��~9X��~ ;�@A     _+ ��  9U  ;|AA     �� �  9U��9T��~ ;�AA     �� 4�  9U��9Tv  ;�BA     �� L�  9U  ;�BA     �� d�  9U  ;�BA     �, ��  9U 9Q�� 80CA     �� 9U   :\=A     ��  9Us 9Travc9Q 9R�� ;�=A     �� ��  9Uv 9T��~ ;�=A     ��  �  9Uv 9T~  ;�=A     ��  �  9Uv 9T��~ ;�=A     �� @�  9Uv 9T��~ ;�=A     �� ^�  9Uv 9T}  ;�=A     ̃ ��  9Us�9T	`A     9Q0 ;>A     Ă ��  9U  ;->A     � ��  9U  ;E>A     т ��  9U  ;k>A     �� ��  9Uv 9T89Q09X09Y�� ;�>A     т �  9U  ;�>A     �� E�  9Uv 9T89Q09X09Y�� ;�>A     т ]�  9U  ;?A     �� ��  9Uv 9T89Q09X09Y�� ;.?A     �� ��  9U  ;<?A     �� ��  9U  ;�?A     �� ��  9Uv 9T89Q09X09Y�� ;BA     т �  9U  PZBA     т ;�CA     �, -�  9U 9Q�� ;1DA     �� [�  9Uv 9T89Q09X09Y�� 8{DA     т 9U   2��  -Z	  `A            ���  I�K  -'�
  UI�  .'a   T4ֳ  0KB  �� ��  2��  �Z	  �A     �       �Z�  3��  �#�5  � �� 3�' �#	  �� �� 4�U �Z	  H� 8� 4E�  ��3  �� �� 4;�  ��I  6� 0� 4��  �	  �� �� 5�  ̞A     6F�A     g       $�  4ڰ  �u  �� �� 4�i  �;I  �� �� 4f�  ��.  � � )�  ��  �H:v�A     ��  9Us 9Q�H ;��A     �� �  9U|  8��A     H  9Us   ;̞A     H  F�  9Us 9T09Q0 8��A     �
 9T0  2,�  �Z	  �A           �H  3��  �!�5  D� 8� 3�  �!	  �� �� 3Ԛ  �!   S� G� 4�U �Z	  �� �� 4E�  ��3  D� >� 7i �	  �� �� 7nc �	  '� !� ;ߟA     �
 $  9T0 8	�A     � 9U} 9T09Q09R1  2��  Z	  ��A     c      �� 3��  !�5  |� p� 3�  !	  � � 3Ԛ  !   b� P� )�U 
Z	  ��4E�  �3  *� &� 4;�  �I  l� d� 7i 	  �� �� 4ڰ  u  u� q� 7c    �� �� 7n    �� �� 4�     �� �� 4��  �  K� A� 5�  t�A     6@�A     L       � 4�' ;	  �� �� 4f�  <�.  � �  60�A     P       � 7a N�.  e� c�  ;��A     ��  9U| 9T89Q09X09Y�� ;ݜA     �{ + 9Ts 9R dy }  ;�A     � N 9U} 9Q 9R0 ;�A     �� l 9U| 9T  ;��A     �( � 9U}  ;��A     �
 � 9T0 8ϝA     �� 9U| 9T89Q09X09Y��  2��  �
Z	   �A           �� 3��  �
�5  �� �� 3�  �
	  #� � 3Ԛ  �
   �� �� 4�U �
Z	  0� (� 4E�  �
�3  �� �� 7i �
	  �� �� 7nc �
	  w� q� ;�A     �
 � 9T0 8�A     � 9U} 9T09Q09R1  ,e�  �
Z	  � -��  �
�5  -�  �
	  -Ԛ  �
   /�U �
Z	   2�  �	Z	  ��A     �      ��
 3��  �	�5  �� �� 3�  �		  �� {� 3Ԛ  �	   �� �� 3�  �	�  �� �� )�U �	Z	  ��4E�  �	�3  ;� 5� 4;�  �	�I  �� �� 7i �		  �� �� 4�z  �	�  �� �� 4ڰ  �	u  �� �� lZ   �	 ��   +�  p�   4��  �	� 9� 1� 5�  d
�A     Vpm  � 4��  �	�  �� �� .j �		  7c �	    � � 7n �	   �� �� LߓA     V       4�' 
	  
� �   N� ��A       �m  @
% K� z� r� K �� �� K� B� :� K� �� �� O�m  M �� �� M" v� p� M/ �� �� M: .� � ME J� @� MP �� �� ^\  n  s M] R� L� P?�A     ��  Nk ��A      `n  �� K k �� �� Kk �� �� O`n  M*k �� �� M6k 3� /�   ck ��A      ��A             �K k r� n� Kk �� �� L��A             X*k X6k     N� �A      �n  �	�	 K� �� �� O�n  M� U� M� M� �� �� M �� �� Z ��M& � � M1 q� i� Z< ��MI �� �� MV �� �� Zc ��[� ��A     ]� W�A     i       , M� '� %� ;e�A     Ă  9U��~ 8��A     � 9U��~  ]� =�A     ^       � M� U� S� ;J�A     Ă l 9U��~ 8u�A     �� 9U��~  :5�A     � 9U| 9Travg9Q��~9R�� ;K�A     [� � 9U��~ ;d�A     ؃ � 9U��~9T	��F     9Q�� ;�A     �� '	 9U��~9T89Q09X09Y�� ;�A     т A	 9U��~ ;��A     �� q	 9U��~9T89Q09X09Y�� ;��A     u� �	 9U��~ ;�A     Ă �	 9U��~ ;<�A     �� �	 9U��~ 8��A     т 9U��~   ;��A     �� �	 9T~ 9Q
s ����3$ ;��A     �� 
 9U��~ ;��A     �\  /
 9U|  ;̖A     �� I
 9U��~ ;G�A     �
 `
 9T0 ;��A     ��  x
 9U|  ;��A     �� �
 9U��~9T89Q09X09Y�� 8�A     �� 9U��~9T89Q09X09Y��  2��  �Z	  `�A     ?      �� 3��  ��5  �� �� 3�  ��I  �� �� 4^�  �A  � � 4ڰ  �u  �� |� )ց  �'	  ��~)�U �Z	  ��~4�  �'	  �� �� 7i �	  �� �� 7j �	  b� ^� 4;�  ��I  �� �� 4v�  �   [  W  7nsc �   �  �  4��  ��   
 7a ��.  � � 7c �   � � 7ns ��.  7 ' );�  �FY  ��4F�  ��  � � 4��  �	  � � 4�  �	  (  4��  ��2  � � 4E�  �t	  ] Y 4��  �t	  � � 4)�  �t	  � � 4�  �t	  C = 4�{  �t	  � � 4�  �t	    4��  ��  � � )"�  �"� 	 �F     )�   "� 	 �F     5�  �	�A     6��A     �       � )m�  ��Y  ��8�A     ؃ 9Uv 9T	 �F     9Q~   6��A     -       1 4�  �'	  � � ;��A     [� � 9Uv  ;ʑA     �(  9U}  8ՑA     u� 9Uv 9T~   Vm   4�i  :	;I  7	 3	 4�  <		  u	 m	 )��  <		  ��~)�y  <	!	  ��4cy  =		  �	 �	 :K�A     � 9U} 9TA9Q��~9R~  :l�A     � 9U} 9T29Q��~9R~  T��A     9U} 9T69Q��~9R��~  V�l  W 7n q		  <
 8
 ;,�A     �� I 9U��~9Q��~ PU�A     ��  N� ��A      @m  j	^ K� x
 t
 O@m  M� �
 �
 M� �
 �
 M�   M� M G M� � � M� � � Z ��~M U S Z ��M* ~ z M7 � � MD � � ]Q o�A            Y MR   8z�A     _ 9U} 9Tt   :	�A     � 9U} 9TRAVM9Qv 9R��~ ; �A     [� � 9Uv  ;5�A     � � 9Uv 9T��~ ;W�A     � � 9Uv 9T2 ;��A     �� � 9U~ 9T09Q��~ ;��A     �  9Uv 9T4 ;ЎA     � 9 9Uv 9T��~ ;��A     � X 9Uv 9T��~ ;�A     [� p 9Uv  ;0�A     �# � 9U} 9T��~�
����~" ;f�A     �� � 9U~ 9T@9Q09X09Y��~ ;��A     u� � 9Uv 9T��~ ;��A     Ă   9Uv  ;�A     �  9Uv  ;�A     �� 0 9Uv  ;��A     �� H 9Uv  8M�A     т 9Uv    :n�A     � 9Travg9Qv 9R��~ :��A     � 9U} 9T2FFC9Qv 9R��~ :��A     � 9U} 9Travf9Qv 9R��~ ;ωA     [� � 9Uv  ;�A     ؃  9Uv 9T	 �F     9Q�� ;�A     �� A 9U��~9T�9Q��~ ;��A     �� � 9U��~9T#| 2$| "������~"��~"��~"��~"# 9Q��~ ;��A     u� � 9Uv  ;��A     �� � 9U��~9T89Q09X09Y��~ ;ŐA     Ă � 9Uv 9T��~ ;ܐA     �� 	 9Uv  ;�A     �� ! 9Uv  ;�A     � 9 9Uv  ;G�A     �{ d 9T��~�9R| dy ��~ ;T�A     т | 9Uv  ;��A     �� � 9Uv  8��A     u� 9Uv   m$  � L    	� m$  � L    	� 0 �  Lk -��  L �5  -�  M 	  -Ԛ  N    -4�  O    /E�  Q�3  /;�  R�I  .a S�.  .i U	  .j U	  .nc U	  E.av k�R    0��  � -��  �$�5  -�  �$	  -Ԛ  �$   -�  �$   /E�  ��3  /;�  ��I  .i �	  .j �	  .a ��.  .av ��R  E/9z 
M	    2�  �M	  �A     �       �� 3E�  �"�3  5 ) 3Ą  �"�  � � 3ܢ  �"     3  �"   � � 3͚  �"   C 7 7i �	  � � 4a� �M	  i ] P5A     �� P�A     ��  ,��  �Z	  � -��  ��5  /^�  �A  /ڰ  �u  /E�  ��3  /�U �Z	  .i �	  .j �	  /ց  �'	  /Q�  �'	  /�  �'	  /b�  ��X  )��  �"� 	��F     1�  dR� /��  '	   E/��  .'	    HS�  1�A     �      �$ 3��  1�5  � � 4E�  3�3  r n 4<v 4�T  � � 4��  4�T  C = 4��  5�  � � 4�  6�  , " 4�z  7�  � � VPo  � 7p B�E    4�� C	  u o ;��A     _ � 9U| 9Tt  8��A     v| 9U d{ |   O�o  4ah gh  � � /
�  ��  jy�A     ̃ 9U�U#�9T	�A     9Q0   2w�  Z	  �A            �� 3�K  (�
    3�  (a   T P 4ֳ  KB  � � 8�A     {`  9T1  0B�  �_ -��  ��5  /^�  �A  /ڰ  �u  /E�  ��3  /�  ��S  /<v ��T  /��  ��T  /�U �Z	  /��  ��  /ց  �'	  /�) �'	  /ʰ  ��  /+�  �'	  E.p �E    2��  X�E  �A     �      �� 3��  X'�5   � I7�  Y''	  T7p [�E  � m  2��  =Z	   �A     
       �E 3��  = �5  � � 3J�  > 	  � � 3iy  ? �F  6 2 j
�A     � 9U�U9T�T9Q�Q9R1  2��  4Z	  �A            �� 3��  4 �5  s o 3J�  5 	  � � 3iy  6 �F  � � j�A     � 9U�U9T�T9Q�Q9R0  2\�  �Z	  �A           �i 3��  �!�5  0 & 3J�  �!	  � � 3iy  �!�F  � r 3<  �!�  R B 4�U �Z	    4�y  �	  � � 4"�  �	  � � 4�� �	    4�B �eT  6 2 5�  .;�A     6��A            � 7idx 	  n l  6;�A             4��  �R  � �  ;_�A     2 . 9T0 ;��A     v| U 9Us�	9Rv d{ s  8�A     2 9T1  ,A�  c	  2 -��  c+�5  -�  d+�S  -"�  e+	  -�y  f+	  /��  h�R  /�  i�E  /�  k	  .j k	  /�z  lM	  /�  mM	  /�� nM	  E/v�  zM	  /؟  {	  /�~  }>S    2�  �Z	  p�A     l      ��" 3��  ��5  � � 3<  ��  f  ^  4^�  �A  �  �  4ڰ  �u  ! ! 4E�  ��3  �! �! 4�B �eT  �! �! 4�U �Z	  " " 4��  ��  -" )" )ց  �'	  ��4�) �'	  m" c" 4ʰ  �'	  �" �" 4�  �'	  9# /# 1�  EN�" 5�A       s  9^! K�" �# �# K�" �# �# K�" �# �# K�" $ $ K�" �$ �$ O s  M�" �$ �$ M�" �$ �$ M�" `% ^% M# �% �% M# �% �% M # )& %& M-# w& s& M:# �& �& ME# 	' ' [P# ȲA     ^Y# �s  �  MZ# Z' T' Mg# �' �' Mt# �' �' m�# �s  M�# ( 
( 8R�A     �� 9U 9T��   ;I�A     u� �  9U 9Tw s " ;h�A     � �  9U 9T�� ;��A     �  ! 9U 9T�� ;ñA     �� 0! 9U��9T49Q09X09Y�� 8�A     �� 9U��9T49Q09X09Y��   :��A     �! 9U~ 9TRAVV9Qs 9R�� :�A     �! 9TRAVH9Qs 9R�� ;��A     [� �! 9Us  ;�A     � �! 9Us 9T�� ;*�A     �  " 9Us 9T2 ;S�A     � " 9Us 9T�� ;q�A     � >" 9Us 9T�� ;��A     �� c" 9U} 9T89Q�� ;��A     �# �" 9U~ 9Tw  "9Q}  P�A     ��  ,=�  uZ	  �# -��  u;�5  -�  v;'	  gmap w;+T  -�  x;�S  /^�  zA  /ڰ  {u  /�U }Z	  /��  �  /�  �	  /�  �	  /��  �	  .i �	  .j �	  1�  �E/�  �	  /"�  �	  /�y  �	  E/Kl  ��     2J�  �Z	  �EA     
      ��( 3��  �6�5  3( /( 3�  �6'	  t( l( 3�  �6�S  �( �( 4^�  �A  >) :) 4ڰ  �u  x) t) )�U �Z	  ��4��  ��  �) �) 4	�  �'	  �) �) 7i �	  M* ;* 7j �	  -+ + 7k �	  Q, O, 4zy  �	  x, v, 4E�  ��3  �, �, 4��  ��R  �, �, 4��  �/  - - 5�  m�EA     6�GA     �       �% 4�  �>S  �- �- V`\  �% 4�k  �  �- �- 4��   �  �- �- 7end   �  . �- ;�GA     � �% 9Us 9T�� ;HA     � �% 9Us 9T�� 85HA     � 9Us 9T��  8�GA     �� 9Uv 9TH9Q09X09Y��  V�\  (& 4�� V�  &. $. 8'JA     � 9Us 9T��  V�\  b& 4�� b�  K. I. 8vJA     �� 9Us 9T��  ;�EA     u� �& 9Us 9T|  ;�EA     �� �& 9Uv 9T  ;FA     � �& 9Us 9T�� ;5FA     � �& 9Us 9T�� ;OFA     � �& 9Us 9T�� ;�FA     �� )' 9Uv 9T89Q09X09Y�� ;�FA     � H' 9Us 9T�� ;�FA     u� k' 9Us 9T��| " ;GA     � �' 9Us 9T�� ;&GA     � �' 9Us 9T�� ;mGA     �� �' 9Uv 9T89Q09X09Y�� ;�HA     �� ( 9Uv 9TH9Q09X09Y�� ;�HA     u� ( 9Us  ;�HA     � <( 9Us 9T�� ;IA     � [( 9Us 9T�� ;9IA     � z( 9Us 9T�� ;yIA     �� �( 9Uv 9T49Q09X09Y�� ;�IA     � �( 9Us 9T�� 8�IA     �� 9Uv 9T29Q09X09Y��  H̖  M�:A           �_+ 3��  M�5  r. n. 4^�  OA  �. �. 4ڰ  Pu   / �. 4E�  Q�3  O/ I/ 4��  R�R  �/ �/ )�U SZ	  ��4��  T	  �/ �/ 4�  U	  /0 !0 7i V	  �0 �0 7j V	  A1 71 )ց  W'	  ��5�  ��;A     :1;A     (* 9U�U9Trava9Qs 9R�� ;];A     Ă @* 9Us  ;m;A     � X* 9Us  ;x;A     � p* 9Us  ;�;A     т �* 9Us  ;�;A     �� �* 9U} 9T@9Q09R~ 9X09Y�� ;�;A     �� �* 9Us  ;-<A     �� + 9U} 9T@9Q09X09Y�� ;W<A     �� + 9Us  ;s<A     �� 2+ 9Us  ;�<A     �� J+ 9U}  8�<A     �� 9U}   2U�      2A     x      ��, 3^�  'A  �1 �1 3ֳ  ''	  62 22 3�y  '	  y2 o2 4_�     �2 �2 4D�  		  �3 ~3 7cnt 		  �3 �3 7i 
	  &4 4 7j 
	  �4 �4 4ڰ  u  �5 �5 )�U Z	  ��;F2A     �� �, 9U��9T89Q09Rv ����9X09Y�� ;h2A     )� �, 9U~  ;�2A     )� �, 9U~  ;�2A     �� �, 9U~  8h3A     �� 9U��  <ԕ  ��2  00A     �      ��. >^�  �'A  �5 �5 >ֳ  �''	  g6 [6 >��  �'R=  �6 �6 ?N5  ��2  �7 �7 @n �	  
8  8 ?D�  �	  �8 �8 @i �	  @9 $9 @j �	  q: g: ?��  ��  �: �: ?ڰ  �u  =; 7; (�U �Z	  ��;^0A     )� �- 9U|  ;�0A     �� -. 9U} 9T29Q09R~����9X09Y�� ;�0A     )� E. 9U|  ;�0A     )� ]. 9U|  ;,1A     )� u. 9U|  ;�1A     �� �. 9U|  ;�1A     �� �. 9U|  8�1A     )� 9U|   2��  �
Z	  P�A     ,	      ��7 3ֳ  �
 KB  �; �; 3ȩ  �
 �M  �; �; 3x �
 	  `< T< 3�1  �
 [  = �< 4�U �
Z	  7> !> )��  �
�C  ��|1�  �V�  )4 /A� �
M	  4�� �
M	  !? ? 6��A     D      �1 4��  �
�5  ? }? )�C  �
�  ��|)�W  �
�  ��|)C!  �
�  ��|)�  �
�  ��|JHe ��A      ��A     '       �0 Kye �? �? Kme �? �? Kae Q@ M@ KUe �@ �@ T �A     9U��{9T09Qs 9R��|9X��|  Nk Z�A      ��  )�0 K k �@ �@ Kk �@ �@ O��  M*k 
A A M6k MA IA   Nk ��A       �  ),1 K k �A �A Kk �A �A O �  M*k �A �A M6k $B  B   Nk ��A      p�  )z1 S k Kk aB _B Op�  M*k �B �B M6k �B �B   Nk ��A      ��  )�1 S k Kk C C O��  M*k BC >C M6k �C �C   89�A     �d 9U��{9Ts 9Q09R��|9X|   NA@ ��A      `�  �
�2 KS@ �C �C Kz@ ,D $D Sm@ K`@ �D �D O`�  M�@ �D �D M�@  E �D M�@ :E 8E M�@ eE ]E Z�@ ��|T��A     9Q��{�9Rs 9Yv�   J�7 ��A      ��A            4�2 K�7 �E �E 8��A     � 9U|�9T09R0  Jk �A      �A            ;*d3 K k �E �E Kk F F L�A            M*k 8F 4F M6k {F wF   Jk D�A      D�A            >*�3 K k �F �F Kk �F �F LD�A            M*k G G M6k IG EG   ;��A     �7 4 9U| 9T} 9Qv 9Rs 9X1 8��A     �A 9U| 9T��{�9Q09R1  N�@ ��A      ��  ��6 K�@ �G �G K�@ *H H O��  M�@ �H �H MA @I :I ZA ��|MA �I �I M)A IJ =J M6A �J �J ^CA P�  A5 MHA  K K Y�Z  ��A       ��  �K�Z  cK ]K K�Z  �K �K K�Z  �K �K O��  M[  8L 2L M[  �L �L M$[  �L �L M1[  M M    ^VA ��  �6 MWA iM _M MdA �M �M ^qA  �  �5 MvA �N �N 8�A     � 9T��{  ^�A 0�  �5 M�A �N �N Z�A ��|M�A �N �N T��A     9T��{�9Q19R��|  Nk ��A      `�  ;	?6 K k 6O 4O Kk ]O [O O`�  M*k �O �O M6k �O �O   Nk ��A      ��  <	�6 K k P P Sk O��  M*k -P )P M6k eP cP   ;m�A     � �6 9T��{ 8��A     � 9T��{  8(�A     &� 9U�9T��|   J�7 �A      �A            �07 K�7 �P �P 84�A     � 9U|�9T09R0  ;��A     �7 _7 9U| 9T} 9Qv 9Rs 9X0 ;��A     �A �7 9U| 9T��{�9Q09R0 8��A     2� 9Uv�9Q0  0�  �
�7 -��  �
�:   2{�  �	Z	  �A     5      �A@ 3��  �	!�:  �P �P 3ֳ  �	!KB  &Q Q 3ȩ  �	!�M  �Q �Q 3�1  �	![  �R �R 3�  �	!�  pS ^S 4��  �	�5  =T 9T 4^�  �	A  wT sT 4�U �	Z	  �T �T 4ؘ  �	�  �T �T 4K �	�M  V V V��  @ 4BJ  �	!>  �V �V 4}~  �	�  6W &W 4)�  �	�  �W �W 4��  �	�  AX ;X 4�  �	�  �X �X Ncc  ��A      �  �	�? K�c  ZY NY Kuc   Z Z O�  M�c  QZ CZ [�c  ��A     N�c  ��A      `�  ��? K�c  �Z �Z S�c  O`�  Z�c  ��X�c  M�c  �[ �[ Md  �[ �[ Md  \ \ M d  \ }\ e-d  ^6d  ��  : M;d  �\ �\  Nv  p�A       �  r�; K;v  ] ] KGv  A] =] K/v  �] {] K#v  �] �] O �  ZSv  ��;��A     �� �: 9U��9T@9Q09R��9X09Y�� ;��A     �� �: 9U��9T@9Q09R��9X09Y�� ;�A     `v  �: 9U�� ;��A     �� /; 9U��9T@9Q09R��9X09Y�� ;��A     �� g; 9U��9T19Q09R��9X09Y�� 8�A     �� 9U��9T29Q09R09X09Y��   ^Id  ��  �; MJd  ^ ^  N�g  )�A      �  �> Kh  :^ 6^ Kh  �^ �^ O�  M+h  �^ �^ M8h  ._ (_ MEh  �_ {_ ]Rh  ��A     ?       J< MSh  �_ �_ M`h  K` C`  JX�  ��A      ��A            r�< K��  �` �` K}�  �` �` Kq�  a a Ke�  -a +a  J2�  ��A      ��A            x�< KK�  Ra Pa K?�  xa va  J2�  �A      �A            y*= KK�  �a �a K?�  �a �a  NO�  8�A      ��  �s= Kj�  �a �a K]�  b b O��  Mw�  8b 0b   J��  �A      �A     #       }�= K��  �b �b K��  �b �b K��  �b �b L�A     #       M��  c 	c   ;1�A     ��  	> 9U��9T��9Qv  TH�A     9U��   ;��A     �� 7> 9U�� ;��A     �� Q> 9U�� ;�A     �� k> 9U�� ;!�A     �� �> 9U�� PR�A     ��  ;{�A     `v  �> 9U�� P��A     ��  ;I�A     �� �> 9U��9T(9Q09X09Y�� ;��A     �� ? 9U��9T(9Q09X09Y�� ;��A     �� K? 9U��9T89Q09X09Y�� ;�A     �� {? 9U��9T89Q09X09Y�� 8B�A     ed  9Uv    m�c  ��  M�c  Qc Mc 8�A     [e  9Uv     ;K�A     ��  �? 9U��9T| 9Qv  8��A     [e  9Uv 9T����  L��A     #       4�m  �
0  �c �c 8��A     ?� 9U}    ,ar O	Z	  �@ -ֳ  O	"KB  -ȩ  P	"�M  -x Q	"	  -�1  R	"[  /��  T	�5  /�i  U	;I  /^�  V	A  /�U W	Z	  /�  X	�1   ,:�  �Z	  �A -��  �%�:  -x �%	  /��  ��5  /K ��M  /�;  �  /�� �M	  /ȩ  ��M  /ֳ  �KB  RVA /��  �   E.top ��  /� ��  R�A /��  ��   E/T�  	'D#  /�|  	'&"  /�U 	'Z	     2W�  )Z	  gA     �      ��W 3��  )#�:  �c �c 3x *#	  8e e 3�  +#	  �f �f 3��  ,#�  i �h )�U .Z	  ��}4A� /M	  {i gi 4�� /M	  Vj Rj 4�  0'	  �j �j 4��  1�5  vk Zk 4�m  20  �l �l 4<�  4�  �m �m )Z�  7{  ��~))�  8B
  ��}4�  9�  �n �n 1�  �5�  �}wA     6biA     �      �C )N5  ��W ��})�   ��W ��})H� ��W ��})Mj  �`  ��})�~  ��W ��~8_jA     o�  9T| 9Q��}9R��~9X4  V�d  uO 4ڰ  ?u  [o So 4�J A	  �o �o 4E|  B	  np dp 4bL  C'	  q q 4�K  E�
  �q �q 4~�  E�
  �q �q V i  %F 7i �A  r �q 4��  �A  's !s 4i�  ��  |s ts )Mj  �`  ��~4N5  �T  �s �s 4�   ��   2t ,t 4H� �Z  �t |t 4�~  �T  �t �t ;StA     �� 	E 9U~ 9T@9Q09R��|�#0$0&9X09Y��} ;�tA     �� 7E 9U~ 9T19Q09X09Y��} ;�tA     �� eE 9U~ 9T29Q09X09Y��} ;�tA     �� �E 9U~ 9T@9Q09X09Y��} ;evA     o�  �E 9Uv 9T| 9Q��~9R��| ;�wA     �� �E 9U~  ;�wA     �� �E 9U~  ;�wA     �� F 9U~  8�wA     �� 9U~ 9T��|  VPe  L 7n 	  �u �u 4��  	  �u �u 4i�  �  0v v 4��  	  $w 
w 4�  	  kx gx 4��  	  �x �x 4��  A  �x �x 4��  	  y sy V�f  RJ 7pp '�W !z z 4�  )	  ~{ |{ 4k�  *	  �{ �{ N\Y �zA      Pg  `/J K�Y �{ �{ K�Y U| I| K{Y } } KnY v} j} OPg  M�Y ~ �} Z�Y ��~M�Y u~ q~ M�Y �~ �~ M�Y � � ]�Y ^yA     B       H M�Y �� }� M�Y �� �� M�Y 5� /� MZ �� ~� MZ �� ��  ]@Z P{A     �       I MAZ ʁ ȁ MNZ �� � Nk X{A      �g  ��H K k � � Kk <� :� O�g  M*k c� _� M6k �� ��   Nk ~{A      �g  ��H K k � � Sk O�g  M*k � � M6k N� J�   n[Z �{A     2       M\Z �� �� MiZ �� ��   ] Z �~A     j       �I M%Z ۃ ك M2Z  � �� Nk $A       h  ��I S k Sk O h  M*k '� #� M6k j� f�   Nk LA      ph  ��I S k Sk Oph  M*k �� �� M6k � �   PA     �� P$A     ��  ;�|A     K� J 9U��~9T��|# 8�|A     2� 9U��~9T 9Qs    8HzA     �A 9U~ 9Q��}�9R0  N�X �}A      �e  t�K K�X � � K�X �� �� K�X 5� -� O�e  Z Y ��}MY �� �� MY Ն φ ^%Y f  oK M&Y %� � M3Y r� n� M@Y �� �� ZMY ��~;NmA     � K 9U| 9T��} ;�mA     v�  <K 9T��~9Q19X}  ;�mA     X� ZK 9U| 9Q}  8�~A     u� 9U|   N] 3nA      �f  y�K KM] � � K@] 5� 3� K3] e� c� K&] �� ��  ;�nA     @[ �K 9Us 9T1 8mA     e� 9U| 9Q0   8yA     q� 9U   N
X hqA      �h  SUL K)X �� �� KX � � O�h  M6X |� t�   Jk xA      xA            ��L K k ܊ ڊ Kk �  � LxA            M*k +� '� M6k n� j�   Jk &xA      &xA            �1M K k �� �� Kk ы ϋ L&xA            M*k �� �� M6k =� 9�   Nk MxA      0i  �M K k z� x� Kk �� �� O0i  M*k Ɍ Ō M6k � �   Nk yxA      `i  �M K k I� G� Kk p� n� O`i  M*k �� �� M6k ܍ ؍   Jk �xA      �xA            KN K k � � Kk ?� =� L�xA            M*k h� d� M6k �� ��   Jk �xA      �xA            �N K k � � Kk � � L�xA            M*k 8� 4� M6k {� w�   ;�qA     }� �N 9U��|9T  ;�sA     }� �N 9Us�9T  :�sA     O 9Us  :�sA      O 9Us  ;M}A     �� DO 9U~ 9TH9Q��} ;o}A     �� ^O 9U��| 8~}A     q� 9U��|  Jud -hA      -hA     �       ��P K�d �� �� K�d ݏ ۏ L-hA     �       M�d �  � M�d '� %� M�d N� J� Z�d ��}Z�d ��}Z�d ��}Z�d ��~M�d �� �� oHe �hA      �c  ��P Kye Ȑ  Kme � � Kae n� l� KUe �� �� T�hA     9U 9T09Q| 9R��}9X��}  ;ohA     [� �P 9U��| ;�hA     �d �P 9U 9T| 9R��}9X��~ 8�hA     u� 9U��|9T��|   Nk 6kA      �c  SQ K k �� �� Kk ޑ ܑ O�c  M*k � � M6k J� F�   Nk �kA      d  �Q K k �� �� Kk �� �� Od  M*k ג Ӓ M6k � �   Jk `kA      `kA            R K k W� U� Kk }� {� L`kA            M*k �� �� M6k � �   Nk �kA      pd  mR K k &� $� Kk L� J� Opd  M*k u� q� M6k �� ��   Nk �kA      �d  �R K k �� � Kk � � O�d  M*k D� @� M6k �� ��   Jk �kA      �kA            1S K k ĕ  Kk � � L�kA            M*k � � M6k W� S�   NyZ [oA      �i  1oV K�Z �� �� O�i  M�Z �� �� Z�Z ��~M�Z b� Z� M�Z Η ʗ M�Z � � M�Z z� h� [�Z qA     ^�Z �i  {U M�Z J� :� M�Z � �� M
[ ƚ �� M[ ,� $� M$[ �� �� Nk �pA      @j  JQT S k Kk �� ܛ O@j  M*k � � M6k _� [�   Jk �pA      �pA            K�T S k Sk L�pA            M*k �� �� M6k � ݜ   n1[ �rA     y       M2[ $� � Nk �rA      pj  AU S k Kk �� �� Opj  M*k  �� M6k � �   ck 'sA      'sA            BS k Sk L'sA            M*k D� @� M6k �� ��     N] |A      �j  ��U KM] Ğ  K@] Ğ  K3] � � K&] � �  ;
qA     @[ �U 9Us 9T0 ; qA     ��  V 9U  ;�qA     �� :V 9U 9T@9Q09R~  $ &9X09Y��~ ;rA     o�  `V 9Q|� 9Rw 9X~  P|A     ��   :�gA     �V 9T| 9Q��} ;�gA     o^  �V 9Uu 9T| 9Qq  PCiA     DX ;NiA     �c �V 9Us 9T|  :TlA     �V 9T��} ;�lA     �� W 9U  :�lA      W 9Us 9T|  :�lA     4W 9Us  :�lA     HW 9Us  P�nA     DX ;�nA     �c mW 9T|  : oA     �W 9Us 9T|  :CoA     �W 9Us  :[oA     �W 9Us  ;@qA     q� �W 9U��| T�qA     9Us   �  �W L    �   �W L    A  
X L    ,�  
�
  DX -�q  
!�
  gidx !	  .cur �
   Ht{  �� A     �       ��X I��  � �:  U4��  ��  >� 8� 4}~  ��  �� �� 4�  ��  � ޟ 4K ��M  T� N�  ,j�  (Z	  \Y -��  (*�:  -�J )*	  -E|  **	  /�U ,Z	  /Mj  -�  .i .	  E/^�  GA  /Z�  H�  /%�  H�  .tmp I'	    ,Q  Z	  yZ -��  0�:  -i�  �0�  -�J �0	  -��  �0	  /�m  �0  /�  �`  /��  ��  .x ��  .y ��  R Z /��  �	  .k �	  .l �	  .p1 �T  .p2 �T   R@Z /,�  �M	  /z�  �M	   E/A� �M	  /�� �M	  E/��  ��5  /K ��M     ,}  �Z	  @[ -��  �'�:  /�m  �0  /�U �Z	  /Mj  ��  /0�  �	  /ڰ  �u  /�~  �T  1�  mE.vec �T  /��  �T  /A� �M	  /�� �M	  /N�  ��  E.u <T     p{�  )Z	  P+A     i      �] 3��  )�:  �� �� 3�w  *�  ?� ;� 4��  .�5  z� x� 4K /�M  �� �� 4�y  2>  �� � 4Z�  5	  �� �� 6p-A     �      �\ 4�U cZ	  � � 4�m  e0  � � 4�  f`  D� B� NX�  �-A       �Y  i�\ K��  o� m� K}�  �� �� Kq�  �� �� Ke�  ߣ ݣ  Y/�  .A      �Y  oKA�  � � Y��  .A      �Y  %K��  )� '� K��  O� M� K��  u� s� O�Y  M��  �� ��     P�+A     �� P�/A     ��  0�y  [] -�y  ">  -" "�  -�J "	  -E|  "	   0�~  w] -��  #�5   2�  EZ	  �JA     7      �_ 3��  E'�:  Ȥ �� 4�U GZ	  4� (� 7p H  � �� 4��  I  �  � 4�m  J0  >� :� 4�  K	  x� t� 4i�  L�  �� �� 4�  M	  � �� 5WD  ��MA     1o�  �V]  �^ 7xx TM	  �� y� 7xy TM	  K� =� 7yy TM	  �� � 7yx TM	  ͫ �� 4/� U	  �� z� 8�KA     �� 9Us 9T   O`]  4^�  �A  3� 1� P�MA     [�   2Y�  [Z	  �4A     �      ��a 3" [$�:  i� W� 4�U ]Z	  5� '� 7p ^  � ή 4��  _  J� F� 4�m  `0  �� �� 4   a	  �� �� 4Mj  b�  �� �� 4Z�  c�  P� L� 40�  d	  �� �� 4~� f  � � 4��  f  � �� 7c g�  [� M� 4/� g�  �� � 7vec hT  9� /� 4��  hT  �� �� 7x i�  �� �� 7y i�  `� \� 43�  j�E  �� �� 4�  j�E  2� &� 4.�  j)�  Է ̷ Qȥ  k	   1WD  ;1M�  >V�Z  Ha htmp �'	  ��;�6A     v�  *a 9T��9Q19Xw  8�6A     �� 9Tw 9Q��  V�Z  za 4�� ��  D� 0� 7f ��  {� q�  V[  �a 4�� �  �� � 7f �   � ��  ;�8A     e� �a 9U| 9T09Q~  8�8A     e� 9U| 9T9Q0  2�  ?Z	  0 A     �       �Jb I��  ?$�:  U7p A  D� 6� 4��  B  � �  HF�  5 0A     	       ��b 3��  5%�:  � 
� 4^�  7A  K� G� G)0A     т  2��  Z	  �/A     R       ��c 3��  %�:  �� �� 3x %	  � � 3�   %'	  B� >� 3!�  !%	  �� {� 4�U #Z	  �� �� 4^�  $A  8� 4� ;�/A     u� ac 9Us 9T�Q 8�/A     Ă 9Us 9T| ����  `҉  ���@     �       �ud >��  �-�:  v� n� >x �-	  ۾ վ ?��  ��5  +� '� ?�C  ��  i� c� q�W  �"�   ?C!  ��  �� �� q�  �#�   5�   A     O�U  (�|  �"&"  �P?�U �"Z	  	� � T��@     9T�T9Q09Rw    A�  �Z	  �d B��  ��:  Bx �	  C��  ��5  C�U �Z	  C^�  �A  C�C  ��  C�W  �"�  CC!  ��  C�  �#�  Fpos �'	   kJ�  uHe B��  u �5  _idx v 	  BH  w �  _tsb x �E  _ah y �2   k��  c�e B��  c �5  _idx d 	  _lsb e �E  _aw f �2   ,̓  A  �e -K A">  -o�  B"�  /�-  Dm  /�Y  E  /֒  F>  /�i  G;I   2j�  �Z	  ��A     �       ��f 3�  � �  :� ,� 3��  � <  �� �� 3x � 	  �� �� 3�1  � [  j� Z� 4�  ��M  (� � 4ֳ  �KB  �� �� 4��  �h  �� �� )�U �Z	  Pr�A     �. �f 9U�T9T�U j+�A     �. 9U�T9T�U  ,v�  LZ	  kg -ֳ  L%<  greq M%s  /��  OKB  /�U PZ	  R[g /�H  W�5  /�i  X;I  /m Y'	   E/� p	    2n�  'Z	  PA     S       �uh 3ֳ  '<  �� �� 3m ('	  8� 0� 4�H  *�5  �� �� 4��  +KB  �� �� 4�U ,Z	  D� >� 6dA     !       Nh 4�i  :;I  �� �� 4I�  ;E  �� �� TuA     9T�T9Qs  P�A     �� 8�A     {`  9Us 9T0  Af�  �Z	  i B�H  �h  B�k �	  B/� �	  B�1  �[  B�@  �   Fnn �	  C��  ��5  R�h Ftsb ��  Fah ��   E.lsb 
�  .aw �    <8�  �Z	  P�@     3       ��i >�H  �h  )� #� >sl  �	  {� u� >�J  �	  �� �� >/�  �T  !� � ?��  ��5  �� �� ?�i  �;I  �� �� Tu�@     9U�U9T�T9Q�Q  <��  wZ	  �MA     /       ��j >ϖ w!>  '� #� >�1  x!�  _� ]� =<v y!9  Qq�U {Z	   ?K |�M  �� �� ?��  ~	  �� �� LNA            @val �R=  �� ��   A�  >Z	  k Bϖ >!>  B�1  ?!�  B<v @!9  B�h  A!�  C�U CZ	  CK D�M  EC��  M	  R�j Fs S�   EFiv [R=     AVJ  �[  Ck _a �[  _b �[  Fret �.  Ftmp �.   sf�  �A     (       ��k tx�  UK��  %� � K��  v� n� M��  �� ��  s�d  NA     |       �dl Ke � �� Ke �� |� K$e .� (� K0e �� z� K<e �� �� ^�d �]  8l Ke O� K� K<e �� �� K0e �� �� K$e �� �� Ke �� ��  u@NA     9U�U9T19Q�T9R�R9X�X  suh �NA           �8n K�h (� � K�h �� �� K�h 6� ,� K�h �� �� K�h �� �� M�h k� g� M�h �� �� 6�NA     "       -m Z�h ��Z�h ��8	OA     �d 9U| 9Ts9Q09R} 9X~   muh �]  K�h 8� 4� K�h z� t� K�h �� �� K�h � � K�h p� j� O�]  M�h �� �� X�h n�h `OA     +       Z�h ��Zi ��cHe `OA      `OA     "       	Kye �� �� Kme � � Kae E� ?� KUe �� �� T�OA     9U| 9T09Qs9R} 9X~       s�  �OA     f       ��n K-�  �� �� K:�  � � KG�  _� Y� tT�  Rta�  Xn�   PA     #       K-�  �� �� KT�  �� �� Ka�  �� �� KG�  � � K:�  A� ?�   s��  0PA     ]       �o t��  Ut��  Tt��  QM��  f� d�  s�  `QA     7       ��o t1�  Ut>�  TKK�  �� �� MX�  � � n�  �QA            K1�  �� �� KK�  �� �� K>�  � � L�QA            MX�  K� A�    s��  �QA     <       �^p t��  Ut��  TK�  �� �� M�  V� P� n��  �QA            K��  �� �� K�  �� �� K��  � � L�QA            M�  7� 3�    s��  �QA     :       ��p t��  Ut��  TK��  |� r� M��  �� �� n��   RA            K��  �� �� K��  �� �� K��  �� �� L RA            M��  *�  �    sJ�   RA     7       ��q t\�  Uti�  TKv�  �� �� M��  5� )� nJ�  @RA            K\�  �� �� Kv�  � � Ki�  C� A� L@RA            M��  p� f�    s�  `RA     7       �>r t�  Ut"�  TK/�  � � M<�  �� u� n�  �RA            K�  -� +� K/�  T� P� K"�  �� �� L�RA            M<�  �� ��    s��  �RA     P       ��r t��  Ut��  Tt��  QM��  a� W� n��  �RA            K��  �� �� K��  � � K��  >� <� L�RA            M��  m� a�    su�  �RA     U       �xs t��  Ut��  TK��  C� ;� M��  �� �� nu�  (SA            K��  �� �� K��  �� �� K��  �� �� L(SA            M��  � �    s��  PSA     �       ��s t��  Ut��  Tn��  �SA     "       K��   � �� K��  %� #�   s̻  �SA     �       �bt tڻ  UK�  N� H� t��  Qt �  Rt�  Xm̻  p^  K��  �� �� K�  �� �� K �  � � K�  L� H� Kڻ  �� ��   s4�  �TA     �      �3w KB�  �� �� SO�  M\�  +� #� Mi�  �� �� Mv�  3� +� M��  �� �� [��  �UA     ]��  �TA     $       u M��  �� �� M��  �� �� TUA     9Us   Nf�  8VA      �^  ^ju K��  "� � K��  �� �� Kx�  �� �� O�^  M��  � �   ^��  �^  �v M��  �� �� MǸ  �� �� ]Ը  �VA     ]       dv Mո  F� <� Nk �VA       _  2v K k �� �� Kk '� !� O _  M*k �� �� M6k �� ��   Nk �VA      �_  4Sv S k Sk O�_  M*k � � M6k J� F�   T�VA     9Us   Jk +WA      +WA            +�v K k �� �� Kk �� �� L+WA            M*k �� �� M6k � �   T+WA     9Us   :yUA     �v 9Us 9T  :�UA     w 9Us  T�UA     9Us 9Ts�9Q} 
��  s��  PWA     �      ��x K��  [� S� K��  �� �� K��  � �� K��  �� �� K��  [� U� K�  �� �� M�  %� � M�  t� r� M$�  �� �� M1�  � � M>�  �� �� MK�  S� I� MX�  �� �� Me�  d� Z� Mq�  4� *� m}�  `  M~�  �� �� Nk �XA      ``  �ux S k Kk 9� 5� O``  M*k x� t� M6k �� ��   8�WA     � 9Ts |    s��  �A     �      �3z K��  �� �� Kͯ  g� ]� Kٯ  �� �� K�  G� C� K�  �� �� M��  �� �� M
�  �� �� M�  c� [� M$�  �� �� M1�  � �� M>�  g� a� MK�  �� �� MX�  F� B� Me�  �� |� ^��  �j  z M��  �� �� M��  ]� Q� m��   k  M��  �� �� Nk ��A      `k  w�y K k H� F� Kk m� k� O`k  M*k �� �� M6k �� ��   8X�A     � 9Uw ��9T	����   m��  �k  M��        s�f ��A     �       ��{ K�f O  A  Kg �  �  Mg � � M!g h Z VPl  �z M3g  � M@g & $ ZMg �X:ɄA     �z 9T| 9Q�X 8u�A     kg 9Us   ]�f �A     P       �{ Kg O K K�f � � L�A     P       Xg M!g � � ][g �A     @       n{ M\g   8Q�A     �� 9T
   8�A     {`  9Us 9T0   8�A     �� 9T|   sk ��A     �      �v| K� A 9 K� � � K� ) ! Sy M� � � M� � � M�  � M� 3 ) M� � � M�  	 ^� �l  h| M� � � P'�A     � P�A     �  P8�A     ��  si 0�A     �      ��} K� 	 	 K� �	 �	 K� �	 �	 S{ M� ,
 (
 M� l
 d
 M�  �
 M� � � M�   M� y w M� � � m �n  M	 � � M � � M#   Nk j�A      o  ��} K k C A Sk Oo  M*k � � M6k � �   PѡA     �� P`�A     ��   s� 0�A     7       ��~ K�   K� Z T K� � � M� � � ]� I�A            Y~ K� 
  K� 2 0 K� W U LI�A            X�   8E�A     � 9Us 9Tv 9Q�Q9R1  s�e  �A     b       �� K�e � z K�e   X�e M�e � � X�e X�e ^�e  t  b K�e   K�e ^ X O t  M�e � � X�e M�e � � M�e � � ;a�A     Ȅ H 9T	��F      u��A     9U�U9T�T   84�A     Մ 9U	 �F     9Tv   s�j ��A     ~       ��� K�j )  K�j � � K�j 	 � K�j � ~ v�j  M�j � � m�j Pt  K�j ~ | K�j � � K�j � � K�j | r OPt  X�j X�j m�j Pt  M�j � � ]�j ϴA            o� M�j r p  n�j  �A            M�j � � 8�A     � 9U�Q9T09Q:      s'�  �A     R       �� K9�  � � KE�  > : SQ�  SQ�  Z\�  �P8-�A     � 9Uw   s1�  p�A     �       ��� KC�  � w KP�    K]�  � � Kj�  D < Mw�  � � M��  R F M��  � � M��    M��  @ 0 M��  ^ R N'�  ʵA      �t  0� KQ�  � � KQ�  { q KE�  � � K9�  [  Q  O�t  X\�  8�A     �� 9Q�R9R�R#dQ�  �R   n1�  صA            KP�  �  �  K]�  ! ! Kj�  B! >! KC�  |! x! LصA            Xw�  X��  X��  X��  X��  X��     wKS  KS  �x�I  �I  '�w@G  @G  �w�a  �a  �x�S  �S  Tw\P  \P  x�s  �s  '�w!`  !`  �x?  ?  ((w�]  �]  �w�X  �X  �w]>  ]>  �w�]  �]  �y�  �  ) w�Z  �Z  �w�?  �?  4wM  M  �we  e  �xn  n  (w-R  -R  wWN  WN  �x�`  �`  'vyBY  8Y  ) x�J  �J  *�wd  d  wHg  Hg  �ww  w  �w�k  �k  �w�[  �[  �w�M  �M  *x@  @  +�w�a  �a  +x�W  �W  `wCA  CA  +Ew�D  �D  �x�?  �?  ex�>  �>  �x\u  \u  *`x
^  
^  *sw)p  )p  vxO\  O\  �wf  f  �wR  R  �w$i  $i  -wF>  F>  kx$  $  ,.w�E  �E  H 0�   #  &  ]�  �:  ��A     �`      § ,  i   	�@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ��  
�5  ;  �s  
�H  �  	H  s&  
G   �  
N   )  A"z  �  �   ��  �  �U    ��  ��  <h ��  �I  �
   �  X�  �  U   �  n  -    �   m�  �  
  n  U    f  �    U   :  n  -   -   U    J   �"F  L  �  PH�  Ǟ  JI   ֳ  K@   pos L@     N  /[  O   �K P  (�R QV  0ڰ  Sn  8O�  TI  @��  UI  H �  �  <v �-   ��  �U    �  ��  ""  �%  +  @   I  :  @   I  @    O  �  �   c  i  t  :   v  :-   �  L�  x Nt   y Ot   �  Q�  	�  ~   w�  
  yt   �!  yt  �   zt  H  zt   "  |�  �  (�  M} N    5�  N   `�  	G   _| 
I  
!  H  ?   O  2   O  B  U     �    	�  �  (Q�     S5   0�  T5  N5  V�  �   W�   H� X�  �1  ZG     �  5  �  \�  �  �  N   �T  �!   �   pmoc�  stibu!  ltuo�  tolp :  �  �8  5"n  t  �$  �4  S�  x U5   len VH  e� WO   �#  Yy  	�  �%  {�  �  �  G   G   �  U    �  �#  �    G   !  G   G   U    �.  �.  4  I  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(  �  (�/  !  0�  U   8*  �  @ �  �  u(  
I  	�  �2  (    G     U      a  �3  ;/  5  @  a   v)  ]M  S  h  a  I  @    �3  yu  {  G   �  a  @   U    H7  ��  �  G   �  a  �   �  51  0�$  y2  �T   � ��   �@  *
 �h  / ��   $ �"  ( 2$  ��  -4  lO  +  �I  �  $8  �O  	P  \  Ab  �a    ��   	s  {"  �5  !  �H  	�  \   �G   �  �N   	�  }  �-   )$  �@   �   -   c,  +G   C*  6U   +D  C4    :   �M	  xx ��   xy ��  yx ��  yy ��   5  �
	  	M	  8  ��	  ��  �a   ��  ��   $  �_	  c   ��	  �	  �	  U    �  ��	  Kl  �U    �  ��	   s  ��	  �"  $�	   
  �   +9
  �� -�	   �W .�	  Kl  /U    %  Dd
  uR F�	   �
 G�	   }  I9
  N   $��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<3  5�  >t   ��  ?t  �"  At  �"  Bt  i!  Ct   %!  Et  (2!  Ft  0�  Gt  8   I�  �"   s�  ��  u�   5�  v�  ֳ  xt  !  zt  m  {t   v  }@  J  �#�  �  �!  �}s  ڰ  n   {3  ��  S0  ��  �/  ��  �1  ��  �1  ��$  Y/  �d
  �*  �  (�)  �s  0+:  ��$  8<8  ��$  X�*  ��  � �3  �"�  �  �(  ��  Oe �Z$   �-  ��  ڰ  �n   U  �"�  �  �  8  ah !`$   Oe "�  U1  #d
   ;+  $  0 i(  �$&  ,  l;  ���  ah �`$   Oe �m$  y2  �T   {:  �M  (�� �a  h/ ��  p�� ��  x T   � �  �  _  �q  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"  �  8�  �  @`  !�  Hd  "�  P�@  $�	  X�;  )�  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7q  ��� 8(  �K <�  �ڰ  =n  �^�  >:  �U  @d
  �t  B�	  �k  CU   ��L  Ea  � "   ~  �  1  Xm�  ��  o�   �@  p�	  �e q�  �L  r  P @  $%�  �    0\(  �-  ^�   ��  _�  �W `�  x a�  �@  b�	   �e d3  0�"  e�  pi"  f�  x� g�  ���  iT  �.a k�  ��  l�  �J  m�  �Mj  o  ��  q�  ��  r�  �M  tU    Z  u-   _"  wt  (   xt  Ud zU    �L  |Y  ( �!  F#5  ;  Z!  A�  ��  C�   T DG  �!  E�  "  F�   S  N   �G  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  �C  H;  0  `)n  t  �"  �e�  �1  gM	   H+  h�   x+  i�  0��  k�   8�)  n#"  h�'  q=  p��  rT  t�*  y�  x s  �  (  �S  I�  �  �)  %  �!  H�^  $  �U    7:  �  s4  ��   b  8H�  !  J�   m  K�  A� M�  �� N�  �  Pt  
  Qt   ��  Rt  (�  St  0 �  U^   x  t�  x   �$  
  �!  0'Y  ad  )�   �1  *�  &D  +�  2B  ,�  x� -M	     �)f  l  �"  P��  ��  �   �1  ��  �&  �1  �3  �M	  ]7  ��  0�7  �U   @�1  �T  H �  ~�  P6    tag �   Kl  �   �6  	�    �5  N   
`  i7   �&  9  F9  8%  �*   �,  
(  ./   6
�  b 8
`   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  m  �8  N   �  �:   4,  �6  $  �/  l9   �2  ��  P  �#  ��  �'  �8  >  �  M  s   �2  �Y  _  j  s   l/  �v  |     �  s  �   �   ;)  H�  �#  ��   :  ��  �5  �  F1  ��  ,8  ��   2*  ��  (�*  �,  0`1  �M  8��  �j  @   �-  ��  d)  s8  >  �  M  U    9  F#^  	M  �$  @J�  �#  L�   y2  MT  W� O.  �� PT  �,  Q�   M4  Rq  (�;  S�  0�*  T�  8 c/  X!�  �  �-  (q(  �-  s�   Oe t(  ��  uT  � v�   Y  �/  ):  @  �  T  �  �   g%  .`  f  q  �   �.  1}  �  �  �  �     Z	  73  6�  �  �  �  �   �  �8  :�  �  �  �  �  �   "3  >:  $)  Y  
  �  (    �       �6  _4  :  �  X    �  �     �3  fd  j      �  �   ;0  l�  �  �  �    �  �   �&  x�  ah �    y2  � T  H�8  � �  P�8  � (  X�'  � X  `� �   h�9  �   p $  �.  ��  P  5  @    "9  H2�  Mj  4   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :5  T%  �=  ڰ  ?n   �0  @�  q5  A�  L)  B�  )  C1  Ǟ  E�  �  F�  `Ud HU   � X+  J  �  1  $  *  �  M  :  �  �  �  "   �&  &Y  _  j  �   �1  *v  |  �  �  q   �6  -�  �  �  q   w-  1�  �  �  �  �   �;  4�  �  �  �   =;  8�  �  �    q  �   B$  <    �  2  q  �   2  @>  D  �  b  �  q  �  T   7  Gn  t  �  �  �  �  �  �   q8  N�  �  �  �  �  :   )2  S�  �  �  �  �  �  �  T  �   �  k.  ���  ah �   #,  ��  H�4  ��  P,;  ��  XEY �  `/q �M  hZ)  �j  p�#  ��  x'0  ��  �.  ��  ���  �2  �� �b  �`9  ��  ���  ��  �5  ��  �U#  �  � �/  ��  	�  �2  ��  �  U   8S  �"   �d  ��   �W  ��   C  ��  	"   �&  0��   y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  �3   *  V'�   �   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  �!  !  �  3!  �   �  3!   �	  �9  �E!  K!  [!  �   3!   A2  �g!  m!  �  �!  �   �  1  �!   �   8(  �!  ��  )!   $�  )9!  �-  )[!   )  �!  	�!  3  <"  �� >%"   ��  ?%�    �!  #  A�!  "  �U  �,,"  2"  �B  �Z"  �� �T   Oe �Z"   fP  �,f"  �"  4I  P��"  ֳ  ��   �� �#  �q �3#  R` �P#  �W �v#   P �#�#  (�U  �#�#  0�v  �#�#  8�v  �##$  @�J  �#N$  H 	l"  ��  �2"  wq  �#  #  �  3#   "  �   �J  �?#  E#  P#   "   �\  �\#  b#  �  v#   "  a   \  ��#  �#  �  �#   "  �#   a  U  ��#  �#  �  �#   "   "  a  a   �O  ��#  �#  �  �#   "  a  a   �n  �	$  $  �#  #$   "  n   ;O  �/$  5$  �#  N$   "  n  a   -k  �/$    �(  ��    �D  &�  s  �$  @    +  �$  @    �  �$  @    �$  �  �$  �   �$  �  �$  �  �  �  �   �$  �  %  �     H'  �%$  ��  8Y�%  ��  [�   ��  \�  п  ]�  �U ^�  ��  _�   �  `�  (W�  a1  0�  b�  2�  c�  4 ��  e%  �  p$�%  %  ��  ��'  ��  ��   ��  ��  *�  �P  ��  �P  	��  �P  
�  �P  .�  �'  ��  �'  (��  �'  <�  �'  X0�  ��  pY�  ��  xA�  ��  |M�  �$'  ���  �$'  ���  �P  �W�  �P  ���  �1  ��  �1  ���  �4'  �[�  �4'  ���  ��  ���  ��  ���  ��  ��  �D'  � �  '  @    �  $'  @   	 �  4'  @     �  D'  @    �  T'  @    c�  ��%  �  �#l'  �%  8�  �T'  ��  �'  ��  P   +�  �'  r�   �   �  [�  "~'  ��  "�'  ~'  0�   (�(  ��  *�   �~  +�  U�  -�(  ª  .�(  (��  /�(  �|�  1�  P�  2�  ��  4�(  ��  5�(  �n�  7�  (��  9�(  0��  A)  ���  B�  � �  �(  @    �  �(  @    �'  �(  @    �%  �(  @    `'  �(  @    �  )  @    �  )  @    p�  D�'  ��  D5)  �'  �  N   4m)  �   5�  B�  �  ��   �  <;)  c�  N   {�*  �   ��  x�  �  Q�  ��  ��  f�  ��  �  	�  
Ƹ  {�  ��  [�  l�  ��  �  p�  i�  ��  ��  ��  �  ��  ��  4�  ��  T�  �  ۳  =�  $�   ��  !e�  "4�  #�  $[�  %��  &��  '��  (7�  )�  *2�  +p�  ,��  -x�  - 
�  �z)  $�  )$�*  �*  P�  a�  ,�*  �*  �  �*  n  �*  �*   r'  �*  ;�  1+  +  4+  �*  �  �  �  �   w�  8@+  F+  Q+  �*   *�  ;�+  � =�*   �� >+  �� ?4+   M�  A�+  Q+  ��  h!�+  �+  ��  ��  u-�+  2,  ��  8V2,  �7  X�+   ��  Y7,  �R Z�,  �� [T,  �� \{,   �� ]�,  (a� ^�,  0 	�+  t�  �C,  I,  T,  �+   S�  �`,  f,  {,  �+  �  �   !�  �`,  ��  ��,  �,  �,  �+  �   e�  
�,  �,  �  �,  �+  �   |�  1�,  �,  �  -  �+  -  �*       �  �!-  -  ì  ��  �-,-  �-  �  8��-  �7  �-   ��  ��-  �R �H.  O� ��-  �  ��-   y� � .  (a� �o.  0 	2-  ��  ��-  �-  �-  -   ��  ��-  �-  �-  -  �  �  �   i�  � .  .   .  -  �  �  a   p�  &-.  3.  H.  -  �  a   !�  DU.  [.  �  o.  -  �   %�  j|.  �.  �  �.  -  -  �*     ��  ��.  ��  ��.   �� ��.  � �/   �+  �.  s   �.  �+  �.  s   �.  -  /  s   /  ��  ��.  �  � 2/  /  hG  5^/   num 7�   str 8�   *f  :8/  �_  =�/  key ?^/   Kl  @4    �K  D$�/  j/  �d  H�/  �/  �  �/  �/   ^/  �r  K�/  �/  1  �/  �/  �/   Uj  (OM0  ��  Q�   ֳ  R�  [M S�  �V  U�/  �F  V�/  �B XM0    �/  �@  \ _0  �/  N�  #q0  w0  a  �0  �   :�  )�0  �0  �  �0  �   8�  /�0  �  5�0  V 7a   x 8�   ��  :�0  ��  =$�0  �0  ��  (?.1  I_ A#   J�  B�  �m C.1    �0  f�  M@1  F1  �  Z1  �  �   �  Uf1  l1  |1  �  �   ��  Y�1  �1  �  �1  n  �0  �  41  Z1  �   r�  a�1  �1  �  �1  �0  a   ��  e�1  �1  a  2  �0  �#   ��  @ix2  4v k e0   �y m |1  v n �1  Ty o �1  hn q �0   S�  r �0  (��  s �2  0��  t �2  8 	2  q�  i�2  x2  O  �   I�2  ��  K�   ��  L�  ��  M�  R` O�2  K�  P�2   �    ��  R�2  ��  R3  �2  I�  Z)3  ��  \�    A�  ^3  !Ŀ  a�4  ��  c�%   ת  d)3  8�  eT'  @"*�  f�   "��  hm)  ("T i�2  0"��  k  P"�  l  X"��  m  `"��  o�  h"+ p�4  p"��  q�4  x"��  rS0  �"�  t�  �"�o u�4  �"�" v�4  �"C�  w�4  �"��  yP  �"��  zP  �"}�  {M	  �"	�  |�  �"j�  }�  �"[ ~�   "�  ��     �  �  ��  �53  ��  ��4  53  ��  (�5  N  ��   ��  ��  �  ��  ��  ��  A�  ��    \�  �5  �4  �  �`5  v�  ��   }�  ��  x ��  y ��   \�  �l5  "5  I�  X��5  ��  �1   o�  ��  )r  ��  (dS  ��  0"�  �5  81�  ��  @��  �`5  H'�  ��  P �  ��5  r5  ��  �!6  6  !��  x��6  ah �   �O  ��4  �"Q  ��  "g  ��  "�  ��  "�  ��6   "d  ��6  @"E�  �()  P"��  ��  X"��  ��  \"��  ��  `"f�  ��'  h"�  ��  p T  �6  @    (  �6  @    N�  �6  ��  - 7  7  ��  XZ(7  ah \�    ��  8%47  :7  !��  Pt�7  ah v�   "�� x1  0"��  y1  1"A� {�  8"�� |�  @"�0  ~�  H"q5  �  L �I  `U�8  Q  W�   �g  X�  �;  Z�  �U  [�  �B ]�   �o  ^�  "Y  `�8  (+I  a�8  8
  c�  H�!  d�  J�   e�  LH  f�  N�`  h�  P�X  i�  RO  k�  T,G  l�  V�t  m�  X �  �8  @    I  o�7  �g  8��9  ��  ��   )r  ��  dS  ��  
�B  ��  �P  ��  �p  ��  �K  ��  =  ��  me  ��  +^  ��  �]  ��  �u  ��9  
h  ��  $^K  ��  &tR  �U   (%?  �U   0 �  �9  @    �]  ��8  �S  8?�:  ��  A�   )r  B�  dS  C�  
�B  D�  �A  F�  �n  H�  �n  I�  �W  J�  me  K�  +^  L�  �]  M�  �u  O�9  
h  Q�  $�V  R�  &tR  XU   (%?  YU   0 �u  [�9  JW  �x�<  ��  z�   =  {�  �<  |�  tB  }�  �k  ~�  �m  �  
�D  ��  gJ  ��  !X  ��  �S  ��  5f  ��  ?X  ��  �a  ��  �_  ��  �a  ��  Gf  ��  �=  ��<   �E  ��  0F  ��  8�A  ��  @F  ��  H�E  ��<  P5D  ��  TH  ��  V#l  ��  X$r  ��  Z_S  ��  \'N  ��  ^?_  ��  `L  ��  b�O  ��  h�O  ��  p~e  ��  x [  ��  z0m  ��  |�M  ��  ~rM  ��  �]  ��  ��g  ��  � P  �<  @   	 =  �<  @    �X  ��:  kE  @��=  �^  ��   zp  ��  dv  ��  �i  ��  �<  ��  �F  ��   �D  ��  (�p  ��  03X  ��  8 �b  �=  K_  @��>  ��  ��   �J  ��  �<  ��  e  ��  $� ��  dk  ��  ![  ��  L^  ��  �`  ��>  yN  ��>  ,ma  ��>  4�Z  �=  :�q  �=  ;r  �P  <�u  �P  = =  �>  @    =  �>  @    =  �>  @    	l  ��=  �M  (8�?  ��  :�   �T  ;�  �P  <�  
�K  =�  B  >�  ^  ?�  �g  @�  /o  A�  %B  B�  �O  C�  �<  D�  �]  E�  *w  F�  dW  G�   �F  H�  " e=  J�>  |[  O�?  �� QP   �\  RP  red SP  q  TP   �[  V�?  �?  (�H@  `a  ��   �L  �H@  r  �H@  &W  ��  �F  �H@    �  Ik  ��?  ��  L�@  }W N�   ��  O�  ��  P�   ��  RZ@  8y  hl�@  �~  n�   ��  o�  �~  p�@   �@  �@  @    `�  r�@  ,�  0�HA  }W ��   ��  ��  def ��  ��  ��  tag ��   cy  ��  ( ˣ  ��@  ��  ��A  Ԛ  ��   cy  ��  �}  ��   	�  �TA  U�   ��A  �~  ��   ��  ��  ˧  ��  �~  ��A  i{  ��A   HA  �A  �  ��A  >i    J>B  tag  L�   ��   M�  /�  N�  �f   O>B   �  2\   Q�A  G    ��B  Tag  ��   g   ��  �=   ��  Ja   ��   mn   ��B  PB  �v    �C  �T   ��   �Y   ��  D   ��  S   ��  E]   ��  ;C   ��  �:  �   �[   ��B  DQ   RC  E]   �   ;C   �  �:     �i   C  >M  0 .�C  ��   0�   �Z   1�  vv   2�  �r  3�C  =P   4�  �Q   5�C   ^�   6:  ( C  RC  �p   8_C  CE   YD  �B   [�   b   \�   Pq   ^!D  �C  �m   x`D  ��   z�   �R   {�  Up   |D   �=   ~'D  �U   E  �   =   
    =  Sd   !P  �Q   "=  �G   #=  �v   $=  �=   %=  sD   &=  �\   '=  �X   (=  	`N   )E  
 =  &E  @    �T   +mD  >t   ��E  �>   �&E   �  �&E  !   �P  m   �P  �[   �P  SX   �P   �<   ��E  3E  x@   "�E  �   $�   �`   %�  TL   &�2  �o  '�E   �E  =  �h   )�E  �Z   <4F  �   >�   �f   ?�E   fR   A	F  # ZfF  $j  \�E  $�Y  ]4F   ms    V�F  �   X1   �r  _AF   J   afF  �t   r!�F  �F  U<  �c  ( �G  �B  �   �c   �  �y  �  �Y   ��  cC   ��   �   �1  $ 	\   ��F   L   � 3G  9G  �i  � ��K  ah  �   �u   �DB  ��v   ��  �R   ��   o   ��B  (�&  ��8  0�Q   ��9  �@   ��?  �5�   �1  �<   ��:  ��`   ��  0�a   ��C  8%os2  ��<  hF�   ��=  �j   �  0 M   ��  8w_  ��M  @�>   ��M  H�A   �KN  P^Z   �)N  X�f   �)N  `KT   �)N  h�i   �U   pQ   �U   x%mm  �U   �%var  �U   �g   �U   ��Y  �`D  �Fq  ��>  �jQ   ��  �nQ   ��E  �m   �F  ��P   N@  @   �  @B   �N  H�u   1  P�u   �?  Q�;   �  XzQ     `FN   �  hT     p!u   �  x%cvt  �N  �2i   �K  �)   )�	  ��   +�  ��j   -�  �:>   .�  ��_   01  �S?   31  �E�   4�F  ��W   6a  �XA   8�  �	K   9�  ��c   ?�  �][   @�  ��J   B�  �'<   C  �	Z   E   �q   F�  �G   G�  �T   H�  �a   I   �\   K  (�u   L�  0o   M�N  8^C   N�  <:W   O�4  @_   Q  H�@   R�  P>   S�  X}?   Ta  \m?   Ua  `%bdf  XG  h�k   \�  ��Z   ]�  �Pl   h�  �(a   i�  �i  mU   ��d  nU   � �Q   �8  �g   �"L  L  �t  x ��M  ��   �&G   ֳ   ��O  ȩ   ��  �m   �  �1   ��   x  ��  (^�   �:  0��   ��  8    ��  <�;   ��  @�C   ��  `�  ��  d"f  ��  h�I   �1  lpp1  ��  ppp2  ��  �Ǟ   �]O  ��y   �]O  �BJ   �jO  �<   �  bL   ��   Ud  �U   (�W   ��  0r�   ��  4%pp3  ��  8%pp4  ��  HO�   �  X��   �  `�k   �d
  h �^   �M  �M  �  �M  &G  �  :  >B   �D   *N  N  �  )N  L  �  �  �   �b   A6N  <N  �  KN  L   SQ   QXN  ^N  iN  L   �=  N    T�N  �G   �v  k_  <L  ok   �`   _iN  �?  T  �j  @ �]O  ڰ   �n   �0   ��  q5   ��  
0�   ��      ��  org  ��  cur  ��  "  ��   �    �  (H�  ��2  0�>   ��  8 ,L   ��N  @\   �'wO  }O  �r  �d   � �O  �O  �a  
�  @!EP  ^�  !G:   �k !H�  ��  !I�  /� !J�  T�  !KP  z�  !L�   ��  !M�  (�f  !O>B  0Vu  !P  8 �  !R�O  !��  !UzP  ��  !W�   �  !X�  /� !Z�  c�  ![zP  "= !\zP   �  �P  @   � ��  !^)P  Y�  (!a�P  ��  !d�   �  !e�  c�  !g�2  ��  !h�2  "�  !j�   �  !k�  $ ��  !m�P  -�  !r&Q  ��  !y�   ��  !z�4   8�  !|�P  9�  !�gQ  z  !��   �  !��  �  !��   �  !�2Q  �  !��Q  ّ  !��Q    gQ  ��  !�sQ  J�   !��Q  ��  !��   ��  !��Q  �  !��  ��  !��  ��  !��Q   &Q  �Q  ��  !��Q  ��  !�!R  R  U�  �!RcT  �-  !T�   ^�  !U:  ڰ  !Vn  ��  !W�  �!  !X�   �  !Y�  ${3  ![P  (S0  !\P  )G�  !]P  *��  !_�  ,�_  !a1  0�  !cP  8Y�  !dP  x�  !eP  �T !g�P  ��  !h�P  ��  !jP  89�  !kP  x��  !lP  �x�  !mP  �*�  !o�  81�  !r�4  @��  !u�  H�y !v�4  Pv�  !w  Xx�  !x�  `Ω  !zSZ  h��  !{�  0��  !|`Z  89�  !~FZ  8�  !�%/  XQ  !�}2  `��  !��  h��  !�pZ  p:�  !��  x%�  !��  ���  !��	  ���  !��Q  �ת  !�vZ  � ��  0!��T  ��  !�1   ��  !�1  �  !�R  ��  !��  3�  !��  L�  !��  ��  !��   BV !��N  ( 4�  !�cT  !a�  H!�W  ��  !��   ��  !��  ��  !��  п  !��  �U !��  ��  !��  W�  !�1  �  !��   �  !��  (�  !��  0��  !��  8[@ !��  <}�  !�M	  @�  !�1  `��  !��  h	�  !��  p��  !��  �j�  !��  ��  !�t  �	�  !��  ���  !��  ��  !��  ���  !��  ���  !��  �ɼ  !��  �=�  !��  �6�  !��  �!�  !��  �"�  !��  �6�  !��  �"��  !��   "��  !��  "�  !��  "$�  !��  "n�  !��   "��  !��  ("&�  !��  0"��  !��  4"�  !��  6"ɰ  !��  8"5�  !��  @ Z�  !��T  [�  !�$+W  1W  ��  �!/�W  �  !1W   �  !2�Y  HE�  !5�T   3�  !6�  P%NDV !7�  X��  !A  `!�  !B  h��  !C�  p��  !D�  tx�  !FP  x)�  !G�4  �.�  !Ja  � !׬  �!��Y  *�  !�P   ��  !�P  ��  !�P  �  !�P  .�  !��Y  ��  !��Y  x��  !��Y  �"�  !��Y  80�  !�  �Y�  !t  �A�  !t  �M�  !t  ���  !t  ���  !P  �W�  !P  ���  !	�Y  �[�  !
�Y   ��  !1  ��  !�  ���  !�  ���  !�  ���  !�  ���  !�  ��  !�  ���  !t  ���  !t  �y�  !�  ���  !W  � t  �Y  @    t  �Y  @   	 t  �Y  @    ��  !�W  7�   !FZ  ��  !P   �  !�  Kl  !"  ��  !#�  M�  !&�  ��  !'�  �  !(P   ׵  !*�Y  ��  !L1W  W  pZ  @   � �%  )3  ��  `",�Z  ah ".�   m "/�  X ��  "1�Z  |Z  !��  H"<
[  ah ">�   "�� "@1  0"��  "A1  1"A� "C�  8"�� "D�  @ ��  "F[  �Z  xX  h#*k[  ah #,s$   �q  #.�  8�'  #/1  <iO  #0k[  @��  #1T  ` �  {[  @    Y  #3�[  [  ��  #?-�[  �[  �  `#�/\  *�  #�   O�  #��  z�  #��  �� #��  6�  #��   ��  #��  $�K #��4  (h�  #��4  0ڰ  #�n  8�� #��\  @ ��   #Xq\  �� #[�\   �q #`�\  add #c�\  U1 #i�\   �  �\  �[  �  n   q\  �\  �[   �\  �  �\  �[  �  �  �   �\  H�  #k/\  	�\  ��  #��[  ��  #�"�\  �\  ;�  �#�W]  O�  #�   Ǟ  #�  ��  #�  �U #��  ڰ  #�n   �� #��a  ( ��  #�"c]  i]  Q�  #��]  �k #�   ��  #�  b #�x^   K�  #�"�]  	�]  �]  �  0#�A^  �  #�   ��  #L_  b #�^  ��  #X_  �  #�  ֳ  #P  C�  #�   ��  #	�  $��  #�  ( &��  N   #�x^  ��   }�  ��  ��  �  ��   I�  #�A^  ��  #�i]  &"�  N   #��^  :�   G�  ��  Z�  z�  !�  ��  d�   �  \�  	��  
��  Ѻ   ��  #��^  &��  N   #�L_  ��   ��  F�  r�  ػ  ��  ��  _�  j�  ��  	 e�  #��^  [�  #�d_  j_  z_  �  �   1�  #�]  	z_  ��  h#uQ`  �� #xk`   �q #~|`  �Y #�|`  �L #�|`  ; #��`   �> #��`  (nD #��`  0�M #��`  8�: #�a  @�[ #�3a  H�l #�Ya  P` #��a  X�9 #��a  ` k`  �\      n   Q`  |`  �\   q`  �  �`  �\   �`  �  �`  �\  �   �`  �  �`  �\    �  >B  1   �`  �  �`  �\  �  �`   �  �`  �  a  �\  �  �  �   �`  3a  �\  W]   #a  Sa  �\  W]  �  Sa   �  9a  �  �a  �\  �]  �  �  >B   _a  :�  #��_  	�a  "�  #��\  ��  #��a  ;�  p#4�b  ڰ  #6n   ��  #7�  ȩ  #8
[  ��  #9  Ǟ  #:-   �  #;-  (��  #=c  0��  #>c  8�C  #@�  @� #A�  H�;  #C�  P.�  #D1  X�� #E1  Y8�  #F1  Z��  #H1  [�  #I1  \�� #Kc  ` ��  #��b  �� #��b   �q #�c   �b  �b  U   1   �a  �b  c  �b   �b  ��  #��b  t  ��  #bZc  Ǟ  #d   ��  #e  O�  #f   Q�  #h!c  (�  #ltc  zc  �  �c  &G  �  �4  >B   ;�  #r�c  �c  �c  &G  �4  �   w�  �#w�e  �I #y�a   �� #{�e  p%top #|�  ��� #~�e   �y  #�e  �a�  #��  ��  #��  ��  #�f  �%cff #�R  ��  #�W   ��  #�f  (��  #�c  0׹  #�1  8��  #��  <P�  #��  @"�  #��  Dc�  #��  H��  #��  LT�  #��4  P0� #��4  X�o #��4  `�  #��  h;:  #�  lzd #�1  p��  #�&gc  x��  #�&�c  �Q  #�}2  ���  #��  �Z�  #��4  ���  #�S0  �}�  #�M	  �	�  #��  �E�  #�()  �f�  #��'  ���  #��  � �  �e  @   0 Zc  �e  @    Zc  �  f  @    �	  ��  #��c  �  #�#1f  7f  ��  �#<Bg  ڰ  #>n   ��  #?�  ȩ  #@�  ��  #A  Ǟ  #B-   �  #C-  (��  #Et  0��  #Ft  8�C  #H�  @� #I�  P�;  #K�  `˹  #L�h  ��� #M1  �8�  #N1  ���  #P1  �b�  #RU   ��  #SU   ��� #U�h  � ^�  #�Og  Ug  �  ig  $f  �   G�  #�vg  |g  �g  $f  t  t  P   r�  #��g  �g  �  �g  $f  t  t   h�  #��g  �g  �  �g  $f    �  #��g  ��  #��g  h  h  $f   ؽ  @#��h  �� #��h   �q #��g  VY #�$Bg  c #�$ig  f #�$�g   2 #�$�g  (�J #�$�g  0� #�$�g  8 �h  $f  �  q  �  1   �h  ��  #�h  	�h  ��  N   #��h  >�    �  /�  i�   v�  #��h  f�  #W7f  ��  #vDi  O�  #x   Ǟ  #y  ��  #z   ��  #|i  ��  #|^i  i  �  #/qi  wi  ��  �#�k  �I #��h   �� #�:l  �%top #��'  ��� #�Jl  ��y  #�Qi  x
Q  #�}2  �
�  #��  �
�o #��4  �
��  #��  �
��  #��  �
+ #��4  �
��  #��4  �
��  #�S0  �
}�  #�M	  �
	�  #��  �
a�  #��  �
�  #��  �
�  #�f  �
E�  #�()  `;:  #�  h��  #�ok  p�� #�(l  xf�  #��'  ���  #��  �zd #�1  ���  #��	  � ��  #�/k  	k  jk  �   #�jk  �� #��k   �q #��k  ;U #��k  �" #�"l   	#k  õ  #�|k  �k  �  �k  di  �   �  �k  di  �  q  �  �4  ()  1    ok   �k  �k  di   �k  �  �k  di    �   �k  �  l  l    �   f  l  '�  #�#k  	(l  �  Jl  @   � Di  Zl  @    ��  #�wi  D�  #� tl  ��  �#Tm  ڰ  #Vn   ��  #W&G  ȩ  #X
[  ��  #Y  Ǟ  #Z-   �  #[-  (��  #]t  0��  #^t  8�C  #`�  @� #a�  P�;  #c�  `.�  #e1  ��� #f1  �8�  #g1  ���  #i1  �b�  #kU   ��  #lU   ��� #n�n  � 9�  #��m  �m  �  �m  �m  �   gl  ��  #��m  �m  �m  �m  t  t  P   �  #��m  �m  �  n  �m  t  t   ��  #��m  >�  #�n  %n  0n  �m   ש  #�=n  Cn  �  Rn  �m   ��  @#��n  �� #�n   �q #n  VY #
%m  c #%�m  f #%�m   2 #%0n  (�J #%n  0� #%n  8 �n  �m  &G  �Z  
[  1   �n  �  #Rn  ^�  #�<o  Ǟ  #�   ��  #�  O�  #�   ��  #�o  ��  �#��p  �I #�gl   cff #�R  ��� #��e  �%top #��  h�� #��p  p�y  #�
q  a�  #��  �  #��  �  #�f  ��  #�t  ���  #�t  �0�  #�1  �׹  #�1  ���  #��  �f�  #�q  �P�  #��  �"�  #��  �c�  #��  ���  #��  �T�  #��4  �0� #��4  ��o #��4  ��  #��  �;:  #�  �zd #�1  ���  #�W  ���  #�&gc  ���  #�&�c  � <o  
q  @    <o  �   q  @    �  #�Io  +�  #�fq  �� #��q   �*  #��q  �" #�"l   �q  �q  &G  �Z  
[  1    gc  �c    q  fq  �  �q  �q  �Z  �   �q  �  #�-q  	�q  �  #�#�q  �q  ��  (#9r  ڰ  #n   ^�  #�r   #�5  F�  #�r  w�  # U     ӫ  #�rr  �� #��r   �q #��r  �i #��r   �  �r  �q  n       rr  �r  �q   �r  �  �r  �q   �r  ��  #�9r  	�r  ��  #�#�r  �r  ��  �  �r  �  �  U    �r  ��  #"�q  R�  #-.s  ls  ��   #/ls  f�  #1Z"   ]J #2Z"  ��  #3Z"  V #4Z"   	%s  ��  X#At  8�  #D!t   ��  #E! t  �  #F!&t  ��  #G!,t  կ  #JGt   *�  #O\t  (��  #Rwt  0��  #W�t  8�  #[s  @��  #^!�t  H�  #`"�t  P �\  �a  �h  5l  Gt    �  �   2t  a  \t  a   Mt  wt  l  U   1   bt  �t  �  `'  W   }t  �r  �q  4�  #b�t  qs  N   $��v  h�   M�  �  l�  �  j�  Ҷ  ��  ��  o�  	�  
�  ^�  ۭ  ��  ��  I�  F�  h�  �  ��  
�   (�  !��  "��  #��  $��  %��  &9�  'ظ  (��  0|�  1l�  @��  AV�  QC�  RT�  S�  Tu�  UG�  V��  Wؼ  X-�  `ڿ  a�  b@�  cN�  p%�  �Ҵ  ���  ��  ��  �M�  ���  ��  ��  ���  �4�  ���  ��  ��  ��  ��  �1�  ���  ���  �9�  ��  ���  �j�  ���  ���  �u�  �n�  ���  �%�  �3�  ���  ���  �Ψ  ��  ���  �־  ���  ���  ���  �q�  �Ƿ  ���  ���  ���  ��  �>�  ��  � 
k3  %.�  ��  �&F�w  ah &H�a   ^�  &I:  ���  &K  �I�  &L�  ��  &N  ���  &O�  �k�  &Q1  �װ  &R1  �#�  &S1  � ȯ  &Uw  ��  &U�w  w  !Q�  �'"[x  ��  '$�w   ��  '&�  �Z�  ''�\  �"�  '*�  ("�o '+�\  0"�" ',�\  �"�  '-�\  �"��  '/�  P"+ '0�\  X"��  '1S0  �"��  '21  �"�  '4�  � ��  '6�w  ��  '6sx  �w  ��  ('�x  �x  �  �x  �  �x   �@  �z  (+�x  �x  �  �x  �  �x   �x  �A  9~  (/�x  �x  �  y  �  �  �'   "�  (6y  y  �  -y  �  �  �   ��  (=�x  �  (By  ��  (GQy  Wy  �  ky  �  �   Ӏ  (K�x  ݓ  (P�y  �y  �  �y  �  �4  �y  �y  �x   �  `�  (WY  ��  (Zy  3�  (_�y  �y  �  �y  �  �4  �   >�  (dz  	�y  y  `(d�z  �~  (f"yx   -�  (g"�x  g�  (h"-y  ��  (i"ky  7�  (j"�x   Y�  (k"y  (�  (l"9y  0&�  (m"Ey  8U�  (n"�y  @A�  (o"�y  HY�  (rwy  P��  (s�y  X �A  )&�$  �V  ),�$  b�  )0�z  	�z  tG  )0{  ]o )2!�z   �  )3!�z   �d  *)�$  ��  *,{  	{  `p  *,9{  g *.{    ܨ  +!E{  K{  �  _{  �  pZ   *�  +%k{  q{  �  �{  �  vZ   ]�  +)�{  �{  �  �{  �   ��  +,�{  �{  �  �{  �  �{   T'  ��  +0�{  �{  �  |  �  �*  �  U   �   ��  +7|  	|  �  (+7g|  ��  +99{   Ъ  +:_{  �  +;�{  ݱ  +<�{  ��  +=�{    �<  ,s|  y|  �  �|  s  �  �  1   s=  ,$�|  �|  �  �|  s  �  U    �  ,)�|  	�|  #P  ,)�|  R  ,+g|   bD ,,�|   'd  - }  }  �  +}  �  �  �  �   �  -%<}  	+}  T_  -%W}  F  -'�|    '��  \)�z  	p�F     'D�  o*{  	`�F     '{�  {,z  	 �F     (�  o&|  	��F     ($�  z'7}  	��F     (��  ��|  	��F     .   �}  @    	�}  (��  �#�}  	 �F     )�v  �	`�F     �_  -~  @   . 	~  (��  �-~  	��F     *7�  �  3  +��  '�w  +g  '�t  ,^�  :  ,ڰ  	n  ,�U 
�  ,ֳ  �  -WD  -]�  U-�  -cs �.�~  ,m�  �  /tag �   0/cur O  ,��  P  ,Ь  Q�  ,�  R1  0/len ��     1��  �Y  2��  �"�w  3ڰ  �n   4|�  ��  �  2��  �!�w  2^�  �!:  2ڰ  �!n  2g  �!�t  3�U ��  5tag ��  3ֳ  ��  6�  � 4��  b�  1�  2^�  b$:  2^�  c$�  2��  d$4   3�U f�  5tag g�  3��  h�  7�  ��MB      8A�  F�   &B     n       ���  9^�  F:  �! �! 9��  G�2  !" " 9�p  H>B  �" �" '�U J�  �L:tag K�  �" �" ;ֳ  L�  :# 6# <)&B     =�  �  =Uv =T�L >]&B     J�  =Uv =T�L  ?�  ��B            �.�  @K �s  U Aı  R�  @B     x       ���  @ϖ Rs  UBK T{[  r# p# (��  Va  �t A��  3�  �[B     �      ���  C^�  3 :  �# �# C��  4 �  �# �# C�  5 �  �$ �$ C�[  6 �  % % C\  7 "  S% O% B��  9�5  �% �% B�U :�  k& M& BQ  ;}2  �' �' Bg  <�t  9( +( B�O  =�4  �( �( B�  >�%  �) �) D�  =�_B     E`�  ��  Bϖ Gs  �* �* B6e  G�  �* �* >�[B     W�  =T	׷F     =Q1  E��  ��  Bah t�  W+ O+ E�  b�  B��  ��   �+ �+ B�V ��   `, Z, F0�  B��  �1  �, �,   Fp�  (�  �t  �@<�]B     p�  ��  =Us =Tw  G�_B     d�    E��  C�  Bah ��  �, �, F �  (�� T  �@B�  s  :- 4- BOe Z"  �- �- <R^B     q�  #�  =T0=Qw =R0 >�^B     q�  =T0=Qw =R0   <�[B     ~�  b�  =T	�F      <�[B     ~�  ��  =T	P�F      >\B     �  =Us   H��  �0B     Q      ��  9��  ��  G. ?. ;��  ��5  �. �. ;ڰ  �n  / / ;�O  ��4  8/ 2/ EP�  ��  ;�  ��%  �/ �/ <�B     ��  9�  =Uv  <�B     ��  Q�  =Uv  <�B     ��  i�  =Uv  <�B     ��  ��  =Uv  >�B     ��  =Uv   <]B     ��  ��  =Uv  <zB     ��  ƅ  =Us  <B     ��  ޅ  =Uv  <0B     ��  ��  =Uv  <JB     ��  �  =Uv  <dB     ��  &�  =Uv  <~B     ��  >�  =Uv  <�B     ��  V�  =Tv  <�B     ��  n�  =Uv  <�B     ��  ��  =Uv  <�B     ��  ��  =Uv  <�B     ��  ��  =Uv  < B     ��  Ά  =Uv  <) B     ��  �  =Uv  <C B     ��  ��  =Uv  >b B     ��  =Uv   I`�  ��  �B     M       �݇  9�  �$�  �/ �/ ;��  ��5  (0 "0 ;�  �%/  u0 s0 J�B     .       ;ϖ �s  �0 �0 KB            ��  ;�� ��+  �0 �0  >�B     ��  =T	P�F        H��  �0B            �
�  L�  �$�  U 8h�  u�  PGB     C       �È  9Գ  u%q  �0 �0 Mreq v%�  :1 41 ;ֳ  x�6  �1 �1 ;�� y�+  �1 �1 <bGB     ��  ��  Nډ  s  <pGB     ��  ��  =T|  O�GB     =R0=X0  8��  ]�  �GB     H       ���  9Գ  ]q  2 2 ;ֳ  _�6  j2 d2 ;�U `�  �2 �2 ;�� a�+  �2 �2 K�GB     (       ~�  '0� f�*  �h;��  g�5  -3 +3 O�GB     =Q�h  >�GB     ��  Nډ  s   1$�  Iɉ  2Գ  Iq  3ֳ  K�6  03�� P�+    4��  9�+  �  2ֳ  9'�6  3��  ;�5  3�  <%/  3ϖ =s   A�  �	�   NB     ~      ���  C��  �	�5  f3 P3 (��  �	[x  ��yB��  �	�w  [4 U4 B�O  �	�4  �4 �4 B��  �	`'  �5 �5 (�U �	�  ��yBg  �	�t  	7 �6 D�  �
OB     E��  ��  Pi  
�  �7 �7 >8XB     ��  =U~   K ZB     @       J�  Bڰ  
n  �7 �7 >ZB     ��  =T8=Q0=X0=Y��y  E��  �  B�_ F
�  !8 8 Pidx F
�  �8 �8 B��  F
�  9 9 B��  F
(�  ]9 U9 F �  BK�  T
  �9 �9 J-YB     �       B{ ^
  �9 �9 ><YB     ��  =U} =Tv     Qǒ  &NB      `�  �	:�  R�  ^: H: RՒ  Q; M;  QY  �NB      ��  �	�  R�  �; �; R�  g< [< Rv  �< �< Rj  l= b= F��  S�  ��yS�  ��yS�  ��yT�  �QB     U�NB     ڌ  =Us =T0=Q0=R  <�NB     �  �  =U| =T	��F     =Q> <"PB     �  .�  =U| =T	̷F     =Q: <8PB     ��  K�  =U| =T0 <YPB     1�  p�  =U| =T��y=Q}  <|PB     ��  ��  =U| =T0 <�PB     ��  ��  =U  <)QB     ��  č  =U =Q��y <OQB     ��  ܍  =U|  >XB     ��  =U|    Q��  OB      p�  �
L�  R��  �= �= Fp�  V��  > > V��  Q> O> Q3  �OB      ��  �	��  R@  x> t> F��  VL  �> �> <�OB     ��  ��  =Uv  U�OB     ��  =Us  >�PB     ��  =Uv    U9OB     ʎ  =Us� UOOB     ߎ  =Us� UeOB     �  =Us� U{OB     	�  =Us� U�OB     �  =Us� <�OB     ��  6�  =Tv  >�OB     ��  =Uv    QI~  �QB      ��  �	(�  Rh~  �> �> Rh~  �> �> R[~  �? z? F��  Vu~  �? �? V�~  N@ D@ S�~  ��yS�~  ��yT�~  �TB     W�~  T�~  �TB     T�~  �RB     X�~  @�  &�  V�~  �@ �@ V�~  �A �A V  !B B V  nB lB Y"  TB     P       k�  S#  ��yO@TB     =Us =R��y=X0  URRB     �  =Us  UkRB     ��  =Us  U�RB     ��  =Us  <�RB     �  ̐  =U} =T:=Q��y <SB     �  �  =U} =T==Q| }  <2[B     �  
�  =T}  >X[B     ��  =U =Q��y  X�~  ��  �  V�~  �B �B S�~  ��y<MWB      �  a�  =U|  <�WB     ��  y�  =U|  <�WB     1�  ��  =U| =T} =Qv  <MZB     ��  ��  =U| =T��y <nZB     ��  ܑ  =U =Q��y <�ZB     ��  ��  =U|  >�ZB     1�  =U| =T} =Q   OqTB     =Q
q�   <�QB     �  F�  =U~ =Ts  <�TB     �  d�  =U~ =Ts  <'UB     ��  |�  =U~  >eUB     ��  =U~   Z��  �	ǒ  +��  �	gx  ,��  �	�w  ,ڰ  �	n   Z��  �	�  +��  �	gx  +��  �	�5   [� ��   !B     �      �2�  C��  ��5  �B �B C��  �gx  7C 'C CǞ  �  �C �C Cֳ  ��  #D D B��  ��w  lD \D B��  �  E E B��  �  wE mE B �  �1  �E �E D�  �	"B     E��  !�  Pcur �  �F vF .�  /s ��  /b  	   K�"B     C       \�  \s 	�  ��\b 	  ��>#B     £  =U =T��=Q��  E0�  �  Plen 	�  KG EG Ep�  ו  B��  (	�]  �G �G F��  B}W -	  *H &H E�  ��  B��  S	�  pH bH ]��  F$B      P�  e	&R+�  II ;I R�  �I �I R�  �J �J FP�  V8�  �J �J SE�  ��VR�  CK %K V_�  �L �L Vl�  �M �M Ty�  �$B     U�$B     y�  =U��=T  O&%B     =U =T~ =X0    <�#B     -�  ��  =U�� >$B     9�  =U| =T��=Q��   Or#B     =U   U�!B     ��  =U  U�!B     �  =U  O�"B     =U   O.!B     =U   ?�" S�'B     �      �K�  C��  S!�5  oN cN C��  T!gx  O �N B��  V�w  �O �O B��  W�[  3P P B�a  X�[  3Q Q B�  Y�[  5R R Bڰ  Zn  :S 4S B�U [�  �S �S Bg  ]�t  �S �S Pcur _  T �S B��  `  U �T Pn a�  PU JU B�  a�  �U �U B+�  b�  	V �U B
�  cP  �V �V DWD  �%,B     E��  ,�  (ֳ  ��  ��(Ǟ  �  ��E��  �  Plen ��  W W K�)B     �       ��  B�S  �  �W |W <�)B     ��  /�  =U��~=Q�� <*B     D�  G�  =U  U*B     b�  =U =Q
� UD*B     ~�  =U��=T}  >U*B     ��  =U��~=T   <)B     £  ��  =U~ =T��=Q�� U>)B     �  =U��=T} =Q=R��~�# O�+B     =U��=T}   UW(B     �  =U~  O�(B     =U~   K�*B           �  (ɲ  `%  ��U�*B     k�  =Us =T0 U�*B     ��  =Us =T1 U+B     ��  =Us =T0=Q	��F     =R8 U8+B     ԙ  =U =T0=Q��=R5 Ud+B     �  =Us =T}  O�+B     =U =T}   U�'B     �  =U~  U],B     <�  =U~�=T} =Q��~ Uy,B     _�  =U~�=T} =Q��~ U�,B     ��  =U~�=T4=Q��~ U�,B     ��  =U =T0 U	-B     ��  =U =T1 U>-B     ̚  =U =T2 Un-B     �  =U =T3 U�-B     ��  =U =Ts  U�-B     �  =Us =T��� U�-B     5�  =U =T0 O*.B     =Us =T0  ^ֲ  �@.B     :      ���  C��  ��5  �W �W C��  �gx  �X �X B��  ��w  �Y yY B�B ��[  aZ OZ Bڰ  �n  H[ @[ (�U ��  ��B��  ��  �[ �[ B/� ��  [\ U\ Bg  ��t  �\ �\ DWD  J-1B     E �  �  Pidx ��  �\ �\ (ֳ  ��  ��(Ǟ  �  ��E`�  �  B�S     d] Z] <F/B     ��  ��  =U~ =Q�� <g/B     D�  ɜ  =U}  U|/B     �  =U} =Q
� U�/B      �  =U��=Ts  >�/B     ��  =U~ =T}   U�/B     /�  =U  U�/B     C�  =U  <0B     £  i�  =U =T��=Q�� U-0B     }�  =U  U@0B     ��  =U  Ui0B     ��  =U  Up0B     ��  =U  <�0B     O�  ם  =Ts =R~  O�0B     =U��=Ts   Uj.B     �  =U  U�.B     �  =U  U�.B     ,�  =U  U/B     Q�  =U��=T���=Q~  U1B     e�  =U  <R1B     ��  ��  =U~ =T(=Q�� >l1B     [�  =T~   ?�# �PB     �      ��  C��  ��5  �] �] C��  �gx  J_ 6_ B��  ��w  <` (` Pcur �  Da a B��  �  �b �b Bg  ��t  �c �c EЋ  �  B��  ��2  (d d B/� ��  �d �d B��  ��  Ge 7e Pn �'�  f �e B	O ��[  �f �f Bڰ  �n  ]g Sg (�U ��  ��B��  �1  �g �g E �  ��  B�_ �  *h "h K3B     n       h�  Plen /�  �h �h UAB     C�  =U  O}B     =U��=T| =Q} =Rv  UHB     |�  =U  ORB     =U   U�B     ��  =U  UB     ��  =U  <4B     ��  Π  =Uw  <OB     ��  �  =Uw  UoB     ��  =U�� <�B     ��  4�  =Uw =T2=Q0=R��=X0=Y�� <�B     ��  k�  =Uw =T8=Q0=R��=X0=Y�� U�B     ��  =U�=T| =Qw  U�B     ��  =U} =Ts=Q	��F     =R8 U�B     ͡  =U  UrB     �  =U  O�B     =U   OuB     =U   ?t�  V@2B     P      ���  C��  V$�5  �h �h C��  W$gx  di Zi B��  Y�w  �i �i B�3  Z��  bj Xj B�  [�  �j �j Bah \�  ~k tk (�S  ]��  ��B��  ^�  �k �k B�Y  _�  l l Ua2B     ��  =Uv =T6=Qw =R3 <�2B     g�  �  =U
�=T|  <�2B     g�  6�  =T|  <�2B     g�  N�  =T|  <�2B     g�  f�  =T|  <�2B     g�  ~�  =T|  <�2B     g�  ��  =T|  >L3B     t�  =Us�  M	  �  £  @    Ai�  "G   �B     �       ���  C��  " �w  Jl @l Cֳ  # >B  �l �l CǞ  $ �4  Hm >m C��  % 1  �m �m Pcur '  �m �m B��  (  7n 5n K�B     ;       ��  Ps 7�  ^n Zn U�B     ��  =Us  O�B     =Us   O�B     =Us   ?ͭ  �B            ���  @��  �5  U@��  gx  T *��  ��  ��  +��  �$�5  +��  �$gx  +#` �$�]  ,�U ��  ,��  �U   ,�  ��  ,�  ��  ,E�  �()  -�   ?`�  r`B            ��  C��  r�5  �n �n C��  sgx  �n �n OsB     =U�T=T0=Q0=R0  ?v�  % B           �T�  C��  %#�5  Do 8o C��  &#gx  �o �o (M�  (T�  ��|(��  )�  ��|B�U *�  =p 3p B��  +�w  �p �p BE�  ,()  q q B�L -W]  Tq Pq Pn .�  �q �q BK�  /  �q �q B��  0  6r .r D�  j`B     U3B     !�  =Us =T��|=Q@=R��| <�B     �  >�  =Uv =Q0 O�B     =Us =T0  �^  d�  @    ?v�  ��B           �©  C��  �&�5  �r �r C��  �&gx  �r �r (�U ��  ��zB��  ��w  ms cs BE�  �()  �s �s (o�  �©  ��{Pn ��  !t t (�~  ��  ��zBK�  �  st mt B��  �  �t �t Bڰ  �n  �t �t D�  �B     K�B     �       ��  /map ��'  B6�  �W]  9u 7u (@�  �ҩ  ��{Pp ��  bu ^u (��  ��  ��zK4B     H       -�  B��  W]  �u �u UfB     �  =U  OvB     =U =T0  U�B     T�  =U =T��{=QD=R��z >�B     ��  =U��z=T8=Q0=X0=Y��z  UB     ��  =U =T��{=Q4=R��z >LB     �  =Us =T0  �^  ҩ  @    �^  �  @    ?��  N B     �      ��  C��  N,�5  �u �u C��  O,gx  Gv =v (M�  QT�  ��|(��  R�  ��{B�~  S�  �v �v B��  T�w  w w B�U V�  �w �w BE�  W()  	x x D�  ��B     E�  ë  BK�  l  Ix Ax B��  m  �x �x Pn n�  y y F@�  (o�  x©  ��{B�L yW]  �y �y B�~  z�  �y �y (�  z�  ��{Ep�  }�  Bӱ  �W]  &z "z OaB     =U =T0  U�B     ��  =U =T��{=Q4=R��{ >
B     �  =Us =Q��{�   OUB     =U =T��|=Q@=R��{  ?��  �p&B     &      ���  C��  �&�5  dz ^z C��  �&gx  �z �z (o�  �©  ��~Pn  �  2{ ,{ (�~   �  ��~B�U �  ~{ |{ BE�  ()  �{ �{ Bڰ  n  �{ �{ D�  Hu'B     E��  U�  B�L #W]  | | B}W $  �| ~| Plen %�  �| �| <'B     ��  �  =U~  <"'B     ��  @�  =U~ =Ts����=Q��~ >J'B     D�  =Qs   U�&B     |�  =U} =T��~=Q4=R��~ >�&B     �  =Us =T0  ?��  �0B           �c�  C��  ��5  } } Bڰ  �n  p} n} BE�  �()  �} �} F��  B��  ��  �} �} B�~  ��  ~ 	~ Pn ��  Q~ C~ K�B            u�  B�� ��'  �~ �~ >�B     ��  =U|   <jB     ��  ��  =U|  <�B     ��  ��  =U|  <�B     ��  ��  =U|  <�B     ��  ծ  =U|  <,B     ��  �  =U|  <bB     ��  �  =U|  <�B     ��  �  =U|  <�B     ��  5�  =U|  <�B     ��  M�  =U|  >B     ��  =U|    Aٮ  ��  �@B     �       �K�  C��  �!�5  1 + C�  �!�  � } CԚ  �!�  � � BE�  �()  j� b� (�  �K�  ��Pi ��  Ӏ ˀ Pnc ��  6� 2� <�@B     ��  6�  =Uu =Tt =Qq  > AB     ̷  =Uvh  �  [�  @    AT�  ��  PFB     c       ��  C��  �!�5  r� l� C�  �!�  ā �� CԚ  �!�  '� !� (��  ��  ��Pi ��  y� s� G�FB     d�  >�FB     ��  =U} =Tv =Qw   �  �  @    A��  ��   GB            ���  C��  ��5  ɂ ł C�' ��  � � _GB     u�  =U�U=T0=Q0  A5�  )�  �DB     �      �s�  C��  )�5  M� ?� C�  *�  � � CԚ  +�'  ]� O� B�U -�  �� �� BE�  .()  3� /� Pn /�  s� i� Pp /�  � � (��  0s�  ��~Dcs l_EB     E0�  )�  B4�  =�  {� u� B��  >�  ʆ Ć Pmap ?�'  � � B��  @�'  h� d� B��  A�  �� �� B�j  B�  � � BR  B#�  �� �� E`�  �  B��  M�  "� �  G�EB     ��   <�EB      �  I�  =Qq Nε  s  >FB      �  =U~ =T0=Qq Nε  ��~  �  ��  @    A��  �  �B     �       ��  C��  &�5  �� �� `len &�4  TCH�  &�  � �� BE�  ()  \� P� Pi �  � �  A�  ��  � B     �       ���  C��  �&�5  n� h� alen �&�  �� �� CH�  �&�  � � BE�  �()  �� �� Pi ��   �� Pn ��  �� ��  A)�  ��   @B     �       �u�  C��  ��5  !� � C�  ��  w� m� CԚ  ��  � � BE�  �()  X� R� (�  �K�  �HPi ��  �� �� Pnc ��  � 
� >J@B     ��  =Uu =Tt =Qq   *��  ��  ��  +��  ��5  +�  ��  +Ԛ  ��  ,�U ��   *d�  o�  B�  +��  o�5  +�  p�  +Ԛ  q�  ,E�  s()  /n t�  /m t�  ,��  v1  0,�Y  ��  ,��  ��    AS�  .�  �AB     �      ���  C��  .�5  w� s� C�  /�x  �� �� Bڰ  1n  H� D� B;�  2�x  �� ~� (S�  3�@  ��~(�U 4�  ��~Pi 5�  � � (�  6K�  ��~BE�  7()  i� a� D�  i�AB     <�AB     6�  D�  =U�U=Tt  <�AB     ��  ]�  =Q��~ <�BB     ��  ��  =Uu =Tt =Qq  >�BB     ̷  =Ush  Z��  ̷  +��  �  +�   �  +è   �   8P�  ��  �1B     �       �6�  9��  � �'  Ғ Ȓ Mncv � �  O� G� :j �
G   �� �� G2B     g�   8$�  ��  P B     n       ��  9��  �*�5  � � L�  �*�x  T;E�  �()  >� <� :n ��  e� a� b�U ��  Jx B     5       ;�~  ��  �� �� :map ��'  � �   �@  8��  h�  P	B     �      �,�  9��  h�5  @� .� 9��  i�  � � 9�~  j�  �� �� ;E�  l()  _� U� ;ڰ  mn  ԗ Η ;�U n�  � � 7�  ��	B     7WD  ��	B     K�	B     P      ��  :nn ��  E� C� <�	B     ��  �  =U =T8=Q0=R~ =X0=Y�� <
B     ��  :�  =U =T�=Q0=R~ =X0=Y�� </
B     ��  o�  =U =T =Q0=R~ =X0=Y�� >]
B     ��  =U =T8=Q0=R
| 1$����=X0=Y��  K�B     a       	�  :n ��  k� i� >�B     ��  =U =T8=Q0=R| v ����=X0=Y��  >rB     ��  =U =T
 =Q��  A(�  \�  @B     �      ��  CƩ  \ �  �� �� CԳ  ] q  
� �� Cx ^ �  � � C�1  _ T  Ú �� Bȩ  a(7  M� E� B�U b�  �� �� (LM cZl  ��hB��  d�5  ~� z� Bn�  e1  Ĝ �� ,��  f1  (�  g1  ��gB�O  h�4  �� �� Bg  i�t  ՝ ϝ B �  jk  2� $� (}�  lM	  ��gB	�  m�  � ܞ ()�  n�	  ��gB~�  o1  d� Z� B�  q1  � ؟ -�  HK`B     g       �  B�L  �Y  n� l� GtB     d�  G�B     d�   E`�  ��  (�'  ��  ��gB�e ��  �� �� E��  (�  Pn �  Ѡ Ϡ Pcur -   � �� Pvec �  D� :� BA� �  á �� B��  �  � �� c`�  �B      �B            ,"�  d{�  Rq�  =� ;� J�B            V��  f� b� V��  �� ��   c`�  �B      �B            -"�  d{�  Rq�  � � J�B            V��  � � V��  R� N�   Q`�  �B       �  ';  d{�  Rq�  �� �� F �  V��  ͣ ɣ V��  � �   e`�  �B      �B            (d{�  dq�  J�B            V��  O� K� V��  �� ��    Q`�  �B      ��  "~�  R{�  Ϥ ͤ Rq�  �� �� F��  V��  � � V��  b� ^�   Q`�   B      ��  
"Կ  R{�  �� �� Rq�  ƥ ĥ F��  V��  � � V��  2� .�   G[B     d�  GpB     d�  <�B     ��  �  =U} =T��g <XB     ��  1�  =U} =T =Q~  <�B     ��  P�  =U} =T��g <(B     ��  h�  =Us0 G�B     d�  G�B     d�   U/B     ��  =U��h=Tv =Q~ =Rs  <�B     N�  ��  =U��h=T =Q��g=R��g U0B     ��  =U��h U�B     �  =T��g O=B     =U��h  3  Ag�  �  �B     T      �p�  C��  �  w� m� C��  �  � � C/� �  X� P� C�1  T  �� �� C�@  �  �� �� B��  �5  z� p� (LM Zl  ��hB�O  �4  �� � Bg  �t  y� w� Pnn �  �� �� B�U  �  "� � UEB     C�  =U��h=T} =Q0=R0 <�B     p�  b�  =U��h=Tv  G�B     d�   8�  ��  �B     !      �p�  9��  �$�5  s� k� 9�  �$c  ت Ҫ ;�U ��  *� $� 'LM �Zl  ��h;x ��  w� s� ;�O  ��4  �� �� ;g  ��t  #� !� UB     ?�  =U��h=Tv =Q0=R0 <�B     p�  ^�  =U��h=Ts  O�B     =U��h  8*�  ��  `B     Q       �N�  9LM �di  L� F� 9x ��  �� �� ')�  ��	  �`'�  �1  �_;�U ��  ٬ լ K�B     +       &�  ;��  ��5  � � O�B     =T�`  >|B     N�  =Us =T�T=Q�`=R�_  8��  +�   B     =      �j�  9LM +3di  >� 6� 9x ,3�  �� �� 9��  -33!  !� � 9�  .3j�  �� �� ;��  0�5  ծ Ѯ ;�O  1�4  � � ;�U 2�  Y� K� ;g  4�t  �� � ; �  5k  2� *� '�  6f  ��u:inc 9""  �� �� K�B     �       ��  '��  iSZ  ��lU�B     ��  =U��u=Ts =Q1 UB     ��  =Uv =Tv�=Q��l U*B     ��  =U��u OWB     =U��u  K|B     |       ?�  '�e �"�   ��lG�B     d�  G�B     d�  G�B     d�  O�B     =T} =Q0=R��l  U�B     Y�  =T} =Q  O!B     =Us   1  A�  ��  P>B     �       ���  C��  ��  а ̰ Csl  ��  � 	� C�J  ��  J� F� @/�  ��  RB��  ��5  �� �� ])�  o>B       `�  �R7�  ȱ �� R7�  8� 0� R]�  �� �� R]�  �� �� RP�  � ڲ RC�  5� /� F`�  Vj�  �� �� Vw�  ĳ �� V��  � � V��  g� a� f��  ��  V��  ˴ Ŵ     A� �   �3B     
       ��  Cϖ �$s  � � C��  �$  U� Q� _�3B     ��  =U	 �F     =T�T  8��  ��  p4B     �	      ��  9��  �'�  �� �� Mkey �'�*  �� �� Midx �'�  � ζ 9<v �'U   � Ϸ 9��  �'�  �� � ;��  ��  n� �� ;
�  ��  i� [� ;��  ��5  <� &� ;�O  ��4  ?� )� E0�  �  :val ��  ]� M�  E �  0�  :val ��  � 	�  EА  ��  Pok \1  �� �� K�7B            ��  Pval b�  � � >�7B     ��  =U�Q  G8B     D�   <�5B     -�  ��  =U|  <�5B     D�  ��  =U�H=T| =Qv  <�8B     -�  ��  =U}  >�8B     D�  =U�H=T} =Q|   4   8ڱ  ��  0 B            �c�  9��  �+�  B� <� 9��  �+�{  �� ��  8�  ��    B            ���  L��  �#�  U 8ͪ  ��   B            ���  L��  �+�  UL��  �+vZ  T 8��  ��  ��A     O       ��  L��  �)�  UL�  �)pZ  T 8�  i�  ��A            �C�  L��  i�5  U 8�  I�  � B     p       ���  9��  I(�5  �� �� 9{ J(  V� J� :i L�  �� �� F��  ;��  Q�  t� r� >� B     ��  =Uv    8V�  =�   >B     %       �c�  9��  ="�5  �� �� 9x >"�  �� �� 9_| ?"�  � � 9�H  @"�  o� i� >>>B     ��  =U�Q=Q	�R����  A�  s�  �3B     �       �)�  C��  s$�  �� �� C��  t$�  � � CN  u$�  �� �� C/�  v$�  � � Pfi x�5  �� �� Pi y�  �� �� F��  Ptk �5  (� "� GJ4B     ��    Z�  J��  gfi J!�5  +0�  K!�  +�  L!�  +/�  M!�  /min O`5  /mid O`5  /max O`5  /idx P�  0,��  Y�    8Ƚ  ��  �HB     y      �9�  9L�  ��  y� q� 9^�  �:  �� �� ;g  ��t  G� ?� ;ڰ  �n  �� �� '��  �s  ��:fi ��5  �� �� '�U ��  ��;��  ��5  �� �� ;�  ��4  �� �� D�  @<IB     E��  Z�  B�k   d� \� ]9�  ,KB       �  %Rb�  �� �� Rb�  �� �� RV�  �� �� RJ�  @� :� F �  Sm�  ��Vy�  �� �� V��  %� � V��  |� r� V��  �� �� V��  �� �� V��  ]� U� V��  � � V��  �� �� V��  � � T��  �LB     <�KB     ��  ��  =U��~=T@=Q0=X0=Y�� <tLB     ��  ��  =Us  <�LB     ��  ��  =Us  <�LB     ��  �  =Us =T�� <�LB     �  )�  =Q@=R	��A      <MB     ��  C�  =U��~ >BMB     ��  =Us     <IB     ��  r�  =U|  <1IB     ��  ��  =U| =TX=Q�� <lIB     �  ��  =U  U�IB     ��  =U�� <JB     �  ��  =U  <JB     ��  ��  =U| =Tv  UFJB     �  =U�� UVJB     $�  =U�� >KB     �  =U   4��  m�  ��  2L�  m�  2^�  n:  hfi o�5  3�U q�  3ڰ  rn  3�k s  3��  t  5p u  5kp v`5  3c�  w�  3�  x(  3�� y(  5n z�  6�  � 8o? XG   ��A     )       �t�  ia X$�  Uib Y$�  T;.�  [`5  9� 7� ;��  \`5  ^� \� ;v�  ^�  �� �� ;}�  _�  �� ��  4C�  7�  ��  2}W 7�  hlen 8�  2w�  9U   3�O  ;�4  5n <�  03��  E�     H{�  (�B     P       �`�  9ڰ  ("n  �� �� Mfi )"�5  f� ^� <�B     ��  +�  =Uv  <B     ��  C�  =Uv  _0B     ��  =U�U=T�T  4VJ  �T  ��  ha �T  hb �T  5ret �"  5tmp �"   j��   ?B           � �  k��  Uk��  Tk��  Qf��  Б  R��  �� �� R��  � �� R��  =� 9�   j��  �CB           ���  R۵  }� s� k�  Qdε  V��  �� �� V�  5� )� V�  �� �� V�  [� Q� f%�   �  V&�  �� �� V3�  <� 6� e`�  DB      DB            �R{�  �� �� Rq�  �� �� JDB            V��  � � V��  r� n�     ju�  �FB     1       ���  R��  �� �� R��  � �� R��  U� Q� V��  �� �� Yu�  �FB            ��  R��  �� �� R��  �� �� R��  � � J�FB            l��    >�FB      �  =Tv =Qq Nε  s   mɉ  GB     <       �$�  dډ  V�  <� :� V�  c� _� V��  �� �� >-GB     ��  =T	P�F       n��  �GB     9       ���  R��  �� �� V��  B� :� o��  �GB     "       R��  �� �� J�GB     "       l��  o��  �GB     "       V��  �� �� >HB     ��  Nډ  s      jt�  0HB     �       ���  R��   � � R��  �� � R��  �� �� V��  +� '� l��  ot�  JHB     k       d��  d��  d��  JJHB     k       l��  V��  l� d� f��  ��  V��  �� �� <�HB     -�  ��  =Uv  >�HB     '�  =Uv =T~ =Q��     j�  `MB     �       �=�  R�  &� � R�  �� �� R�  $� � V�  �� �� S�  �VS�  �XY�  �MB     )       ��  R�  � � R�  9� 7� R�  ^� \� J�MB     )       V�  �� �� l�  l�  T �  �MB     <�MB     9�  ��  =T| =Qv  >�MB     �  =Us    <xMB     ��  ��  =Us =T0 <�MB     1�  �  =Us =T�V=Q�X <�MB     ��  "�  =Us =T0 >�MB     �  =Us =Tv   pHg  Hg  .�p�f  �f  .�p�b  �b  8p�s  �s  7p2n  2n  p�?  �?  4q�s  �s  /�qTf  Tf  hp$i  $i  -pR  R  �q�I  �I  /�q�  �  0pM  M  .�q�`  �`  /vp�D  �D  .�pw  w  .�q��  ��  0"qn  n  0p�Z  �Z  .�qNe  Ne  02r/�  %�  1 rBY  8Y  1 qMH  MH  tq
A  
A  dp\P  \P  p�[  �[  2pe  e  �pCA  CA  2Ep�a  �a  2q@  @  2�pmY  mY  �pF>  F>  kq�o  �o  ~pu  u  /yp�Q  �Q  �p�E  �E  Wq�  �  3Xp@G  @G  .�p�a  �a  .�q��  ��  0 v  �)  &  ��  �:  ``B     o      �� (\  �9   ,  i   �L   �  int �  �   @	�   �  	�    p  	 	@   �  	#	@   X  	&	@   �  	)	@    �  	,	@   (�  	-	@   0/  	2S   8�  	5S   < �   �  	�   �  	8"c   
+  	K  �   
%  	L  
�  	M  '  ��  
�A  ;  �s  
�T  �  	T  s&  
S   	`  �  
Z   )  A"�  �  �   ��  �  �a    ��  ��  <h ��  �I  �   �  X�  �  a   �    9    �   m        a    f  �'  -  a   K    9   9   a    J   �"W  ]  �  PH�  Ǟ  JZ   ֳ  KL   pos LL     N  /[  O   �K P*  (�R Qg  0ڰ  S  8O�  TZ  @��  UZ  H �  �  <v �9   ��  �a    �  ��  ""  �6  <  L   Z  K  L   Z  L    `  �  �   t  z  �  K   v  :9   �  L�  x N�   y O�   �  Q�  	�  ~   w  
  y�   �!  y�  �   z�  H  z�   "  |�  �  (�  M} Z    5�  Z   `�  	S   _| 
Z  
!  T  ?   `  2   `  B  a     �    	�  �  (Q     SA   0�  TA  N5  V  �   W�   H� X  �1  ZS     �  A  �  \�  �  �  Z   �e  �!   �   pmoc�  stibu!  ltuo�  tolp :  �'  �8  5"  �  �$  �4  S�  x UA   len VT  e� W`   �#  Y�  	�  �%  {�  �     S   S      a    �  �#  �    S   2  S   S   a    �.  �?  E  Z  S   S   a    �8  `��  .   �   �; �  �1  S   �5  �  �+  �   `(    (�/  2  0�  a   8*    @ �  �  u(  
Z  	�  �2  (    S   -  a   -   r  �3  ;@  F  Q  r   v)  ]^  d  y  r  Z  L    �3  y�  �  S   �  r  L   a    H7  ��  �  S   �  r  �     51  0�5  y2  �e   � �   �Q  *
 �y  / ��   $ �3  ( 2$  ��  -4  l`  +  �Z  �  $8  �`  	a  m  Ab  �r    ��   	�  {"  �A  !  �T  	�  \   �S   �  �Z   }  �9   	�  )$  �L   �   9   c,  +S   C*  6a   +D  C@   �]  P-    :   �k	  xx ��   xy ��  yx ��  yy ��   5  �(	  	k	  8  ��	  ��  �r   ��  ��   $  �}	  c   ��	  �	  �	  a    �  ��	  Kl  �a    �  ��	   s  ��	  �"  $
  
  �   +W
  �� -
   �W .
  Kl  /a    %  D�
  uR F
   �
 G
   }  IW
  Z   $��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<Q  5�  >�   ��  ?�  �"  A�  �"  B�  i!  C�   %!  E�  (2!  F�  0�  G�  8   I�  �"   s�  ��  u�   5�  v�  ֳ  x�  !  z�  m  {�   v  }^  J  �#�  �  �!  �}�  ڰ     {3  ��  S0  ��  �/  ��  �1  ��  �1  ��$  Y/  ��
  �*  �7  (�)  ��  0+:  ��$  8<8  �%  X�*  ��  � �3  �"�  �  �(  ��  Oe ��$   �-  ��  ڰ  �   U  �"�  �  �  87  ah !�$   Oe "4   U1  #�
   ;+  $X  0 i(  �$D  J  l;  ���  ah ��$   Oe ��$  y2  �e   {:  ��  (�� �r  h/ ��  p�� �Z  x T   � �  �  _  ��  �!  �   �  �  �  �    �  �  �   �U   (�    03"  �  8�    @`  !�  Hd  "  P�@  $�	  X�;  )  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7�  ��� 8F  �K <�  �ڰ  =  �^�  >K  �U  @�
  �t  B�	  �k  Ca   ��L  E  � "   �  �  1  Xm�  ��  o�   �@  p�	  �e q�  �L  r0  P @  $%�  �    0\F  �-  ^�   ��  _�  �W `�  x a�  �@  b�	   �e dQ  0�"  e�  pi"  f�  x� g�  ���  ie  �.a k�  ��  l�  �J  m�  �Mj  o  ��  q�  ��  r  �M  ta    Z  u9   _"  w�  (   x�  Ud za    �L  |w  ( �!  F#S  Y  Z!  A�  ��  C�   T De  �!  E�  "  F�   S  Z   �e  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  �C  HY  0  `)�  �  �"  �e  �1  gk	   H+  h�   x+  i�  0��  k�   8�)  n#l"  h�'  qN  p��  r`  t�*  y�  x �  �  F  �S  I�  �  �)=  C  �!  H�|  $  �a    7:  �+  s4  ��   b  8H�  !  J�   m  K�  A� M�  �� N�  �  P�  
  Q�   ��  R�  (�  S�  0 �  U|   x  t�  x   �$"  (  �!  0'w  ad  )�   �1  *�  &D  +�  2B  ,�  x� -k	     �)�  �  �"  P��  ��  �X   �1  ��  �&  �B  �3  �k	  ]7  ��  0�7  �a   @�1  �`  H �  ~�  P6  3  tag �   Kl  	   �6  	  3  �5  Z   
~  i7   �&  9  F9  8%  �*   �,  
F  ./   6
�  b 8
~   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  �  �8  Z   �+  �:   4,  �6  $  �/  l9   �2  ��  �\  �o  b<  ��   1S ��  p �o   a  p  �8  �#  �	  �'  ��  �  �  �  �   �2  ��  �  �  �   l/  ��  �  �  �  �  �   �   ;)  H�{  �#  ��   :  ��  �5  �{  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  ��  8��  ��  @ �  �-  ��  d)  s�  �  �  �  a    9  F#�  	�  �$  @J6  �#  L�   y2  Me  W� O�  �� P�  �,  Q(   M4  R�  (�;  S   0�*  TN  8 c/  X!B  H  �-  (q�  �-  s�   Oe t�  ��  ue  � v�   �  �/  )�  �  �  �  6  �   g%  .�  �  �  6   �.  1�  �  �  6  �  !   x	  73  6    "  6  "     �8  :4  :  �  N  6  6   "3  >�  $)  Yf  l  �  �  7  �  +  !   �6  _�  �  �  �  7  �  �  !   �3  f�  �  �  7  �  "   ;0  l�  �  �    7  �  	   �&  x�u  ah � �   y2  � e  H�8  � Z  P�8  � �  X�'  � �  `� � �  h�9  � u  p 5  �.  �  "9  H2�  Mj  4   H5  5  (�)  6  0�  7�  8�  8  @ �0  :�  T%  �=X  ڰ  ?   �0  @�  q5  A�  L)  B�  )  CB  Ǟ  E�  �  F�  `Ud Ha   � X+  Jd  �  1  v  |  �  �  K  �  �  �  @   �&  &�  �  �  �   �1  *�  �  �  �  �   �6  -�  �  �  �   w-  1    �    �   �;  4'  -  8  �   =;  8D  J  �  ^  �  �   B$  <j  p  �  �  �  �   2  @�  �  �  �  �  �  �  `   7  G�  �  �  �  �  �  �     q8  N�  �  �  
  �  K   )2  S    �  ?  �  �  �  `  ?   �  k.  ��#   ah ��   #,  ��  H�4  ��  P,;  ��  XEY �j  `/q ��  hZ)  ��  p�#  ��  x'0  ��  �.  �  ���  ��  �� ��  �`9  ��  ���  �
  �5  �8  �U#  �^  � �/  �E  	#   �2  �@   E  a   8S  �t   �d  ��   �W  ��   C  �L   	t   �&  0��   y%  �	   �/  �	  �'  �	  �6  �	  �+  �	   �6  �	  ( �7  ��   *  V'!  !  �0  �*   uN!  |#  w�   �#  x�  � y�  C4  z�   �&  |!  �'  �f!  l!  �  �!  �   �  �!   �	  �9  ��!  �!  �!  �   �!   A2  ��!  �!  �  �!  �   �  B  �!   N!  8(  "  ��  )Z!   $�  )�!  �-  )�!   )  �!  	"  3  <Y"  �� >%Y"   ��  ?%�    )"  #  A."  _"  �U  �,~"  �"  �B  ��"  �� �r   Oe ��"   fP  �,�"  N#  4I  P�N#  ֳ  ��   �� �_#  �q ��#  R` ��#  �W ��#   P �#�#  (�U  �#$$  0�v  �#O$  8�v  �#u$  @�J  �#�$  H 	�"  ��  ��"  wq  �k#  q#  �  �#  r"  	   �J  ��#  �#  �#  r"   �\  ��#  �#  �  �#  r"  r   \  ��#  �#  �  �#  r"  �#   r  U  � $  $  �  $$  r"  r"  r  r   �O  �0$  6$  �  O$  r"  r  r   �n  �[$  a$  �#  u$  r"     ;O  ��$  �$  �#  �$  r"    r   -k  ��$  *�  ��"  	�$  �  �(  ��  {  �D  &�  �  �$  L    �  %  L    �  %  L    %  �  (%  �   .%  �  L%  �  �  	  �   R%  �  f%  �  {   H'  �%5  ��  8Y�%  ��  [   ��  \  п  ]  �U ^  ��  _   �  `�  (W�  aB  0�  b�  2�  c�  4 ��  es%  �  p$&  s%  ��  ��g'  ��  ��   ��  ��  *�  �a  ��  �a  	��  �a  
�  �a  .�  �g'  ��  �w'  (��  �g'  <�  �w'  X0�  ��  pY�  ��  xA�  ��  |M�  ��'  ���  ��'  ���  �a  �W�  �a  ���  �B  ��  �B  ���  ��'  �[�  ��'  ���  ��  ���  ��  ���  ��  ��  ��'  � �  w'  L    �  �'  L   	 �  �'  L     �  �'  L    �  �'  L    c�  �&  �  �#�'  &  8�  ��'  ��  (  ��  a   +�  (  r�   ?   �  [�  "�'  0�   (�(  ��  *�   �~  +�  U�  -�(  ª  .)  (��  /)  �|�  1?  P�  2?  ��  4+)  ��  5;)  �n�  7�  (��  9K)  0��  A[)  ���  B�  �   )  L    ?  )  L     (  +)  L    &  ;)  L    �'  K)  L    "  [)  L    �  k)  L    ��  Dx)  -(  c�  Z   {�*  �   ��  x�  �  Q�  ��  ��  f�  ��  �  	�  
Ƹ  {�  ��  [�  l�  ��  �  p�  i�  ��  ��  ��  �  ��  ��  4�  ��  T�  �  ۳  =�  $�   ��  !e�  "4�  #�  $[�  %��  &��  '��  (7�  )�  *2�  +p�  ,��  -x�  - 
�  �~)  N�  #�*  �*  r  �*  �   :�  )�*  �*  �  �*  �   8�  /�*  �  5/+  V 7r   x 8�   ��  :+  ��  =$G+  M+  ��  (?�+  I_ AS#   J�  B�  �m C�+    /+  f�  M�+  �+  �  �+  	  �   �  U�+  �+  �+  	  �   ��  Y�+  �+  �  
,    ;+  �  �+  �+  	   r�  a,  ,  �  0,  ;+  r   ��  e<,  B,  r  V,  ;+  �#   ��  @i�,  4v k �*   �y m �+  v n 
,  Ty o 0,  hn q �*   S�  r �*  (��  s �,  0��  t �,  8 	V,  q�  i�,  �,  [  $�  )$�,  �,  P�  a�  ,-  -  �  +-    +-  1-   �'  �,  ;�  1C-  I-  h-  �,  �  �  �  �   w�  8t-  z-  �-  �,   *�  ;�-  � = -   �� >7-  �� ?h-   M�  A�-  �-  ��  h!�-  �-  ��  ��  u-�-  f.  ��  8Vf.  �7  X�-   ��  Yk.  �R Z�.  �� [�.  �� \�.   �� ]�.  (a� ^/  0 	�-  t�  �w.  }.  �.  �-   S�  ��.  �.  �.  �-  �  ?   !�  ��.  ��  ��.  �.  �.  �-  �   e�  
�.  �.  �  /  �-  �   |�  1/  /  �  5/  �-  5/  �,  +     �  �!H/  N/  ì  ��  �-`/  �/  �  8��/  �7  �;/   ��  ��/  �R �|0  O� ��/  �  �'0   y� �T0  (a� ��0  0 	f/  ��  ��/  �/  �/  ;/   ��  �0  0  '0  ;/  �  �  ?   i�  �40  :0  T0  ;/  �  �  r   p�  &a0  g0  |0  ;/  �  r   !�  D�0  �0  �  �0  ;/  �   %�  j�0  �0  �  �0  ;/  5/  �,  +   ��  �1  ��  �1   �� �11  � �F1   �-  1  �   1  �-  11  �   "1  S/  F1  �   71  ��  ��0  �  � f1  L1  hG  5�1   num 7�   str 8�   *f  :l1  �_  =�1  key ?�1   Kl  @@    �K  D$�1  �1  �d  H�1  �1  �  �1  �1   �1  �r  K2  2  B  %2  �1  �1   Uj  (O�2  ��  Q�   ֳ  R�  [M S�  �V  U�1  �F  V�1  �B X�2    �1  �@  \ �2  %2  �  I�  Z�2  ��  \�    A�  ^�2  o  �    ��  (�'3  N  ��   ��  ��  �  ��  ��  ��  A�  ��    \�  �33  �2  �  �w3  v�  ��   }�  ��  x ��  y ��   \�  ��3  93  I�  X��3  ��  �B   o�  �  )r  ��  (dS  ��  0"�  �'3  81�  ��  @��  �w3  H'�  ��  P �  �4  �3  
�  @E�4  ^�  GK   �k H�  ��  I�  /� J�  T�  Ka  z�  L�   ��  M�  (�f  O�4  0Vu  Po  8 �  �  R4  ��  R�4  4  !��  U	5  ��  W�   �  X�  /� Z�  c�  [	5  "= \	5   �  5  L   � ��  ^�4  ��  ^15  �4  Y�  (a�5  ��  d�   �  e�  c�  g�2  ��  h�2  "�  j�   �  k�  $ ��  m75  ��  m�5  75  -�  r�5  ��  y�   ��  z�2   8�  |�5  9�  �6  z  ��   �  ��  �  ��   �  ��5  �  �A6  ّ  �A6    6  ��  �&6  J�   ��6  ��  ��   ��  ��6  �  ��  ��  ��  ��  ��6   �5  G6  ��  �S6  ��  ��6  S6  ��  �!�6  �6  U�  �R(9  �-  T�   ^�  UK  ڰ  V  ��  W�  �!  X�   �  Y�  ${3  [a  (S0  \a  )G�  ]a  *��  _�  ,�_  aB  0�  c�4  8Y�  d�4  x�  e�4  �T g5  ��  h�5  ��  j�4  89�  k�4  x��  l�4  �x�  m�4  �*�  o  81�  r�2  @��  u�  H�y v�2  Pv�  wo  Xx�  x�  `Ω  zh?  h��  {�  0��  |u?  89�  ~H?  8�  �Y1  XQ  ��,  `��  ��  h��  ��?  p:�  �  x%�  �  ���  ��	  ���  ��6  �ת  ��?  � ��  0��9  ��  �B   ��  �B  �  ��6  ��  ��  3�  ��  L�  �?  ��  ��   BV ��9  ( `  4�  �(9  ;�  ��9  (9  !a�  H��;  ��  ��   ��  ��  ��  ��  п  ��  �U ��  ��  ��  W�  �B  �  ��   �  ��  (�  ��  0��  ��  8[@ ��  <}�  �k	  @�  �B  `��  ��  h	�  ��  p��  ��  �j�  �  ��  ��  �	�  ��  ���  ��  ��  ��  ���  ��  ���  ��  �ɼ  ��  �=�  ��  �6�  ��  �!�  ��  �"�  ��  �6�  ��  �"��  ��   "��  ��  "�  ��  "$�  ��  "n�  ��   "��  ��  ("&�  ��  0"��  ��  4"�  ��  6"ɰ  ��  8"5�  ��  @ Z�  ��9  G�  �<  �9  [�  �$<   <  ��  �/�<  �  1�;   �  2�>  HE�  5�9   3�  6�  P#NDV 7?  X��  Ao  `!�  Bo  h��  C�  p��  D�  tx�  F�4  x)�  G�2  �.�  Jr  � !׬  ���>  *�  �a   ��  �a  ��  �a  �  �a  .�  ��>  ��  ��>  x��  ��>  �"�  ��>  80�  �  �Y�  �  �A�  �  �M�  �  ���  �  ���  a  �W�  a  ���  	�>  �[�  
�>   ��  B  ��  �  ���  �  ���  �  ���  �  ���  �  ��  �  ���  �  ���  �  �y�  �  ���  <  � �  �>  L    �  �>  L   	 �  �>  L    ��  �<  ��  �>  �<  7�   H?  ��  a   �  �  Kl  "o  ��  #�  M�  &�  ��  '�  �  (a   ׵  *�>  ��  *b?  �>  ��  L <  <  �?  L   � �%  �2  -�  ��6  �I  `U�@  Q  W�   �g  X�  �;  Z�  �U  [�  �B ]�   �o  ^�  "Y  `�@  (+I  a�@  8
  c�  H�!  d�  J�   e�  LH  f�  N�`  h�  P�X  i�  RO  k�  T,G  l�  V�t  m�  X �  �@  L    I  o�?  �g  8��A  ��  ��   )r  ��  dS  ��  
�B  ��  �P  ��  �p  ��  �K  ��  =  ��  me  ��  +^  ��  �]  ��  �u  ��A  
h  ��  $^K  ��  &tR  �a   (%?  �a   0 �  �A  L    �]  ��@  �S  8?�B  ��  A�   )r  B�  dS  C�  
�B  D�  �A  F�  �n  H�  �n  I�  �W  J�  me  K�  +^  L�  �]  M�  �u  O�A  
h  Q�  $�V  R�  &tR  Xa   (%?  Ya   0 �u  [�A  JW  �x�D  ��  z�   =  {�  �<  |�  tB  }�  �k  ~�  �m  �  
�D  ��  gJ  ��  !X  ��  �S  ��  5f  ��  ?X  ��  �a  ��  �_  ��  �a  ��  Gf  ��  �=  ��D   �E  ��  0F  ��  8�A  ��  @F  ��  H�E  ��D  P5D  ��  TH  ��  V#l  ��  X$r  ��  Z_S  ��  \'N  ��  ^?_  ��  `L  ��  b�O  ��  h�O  ��  p~e  ��  x [  ��  z0m  ��  |�M  ��  ~rM  ��  �]  ��  ��g  ��  � a  �D  L   	 N  �D  L    �X  ��B  kE  @��E  �^  ��   zp  ��  dv  ��  �i  ��  �<  ��  �F  ��   �D  ��  (�p  ��  03X  ��  8 �b  ��D  K_  @�tF  ��  ��   �J  ��  �<  ��  e  ��  $� ��  dk  ��  ![  ��  L^  ��  �`  �tF  yN  ��F  ,ma  ��F  4�Z  �N  :�q  �N  ;r  �a  <�u  �a  = N  �F  L    N  �F  L    N  �F  L    	l  ��E  �M  (8�G  ��  :�   �T  ;�  �P  <�  
�K  =�  B  >�  ^  ?�  �g  @�  /o  A�  %B  B�  �O  C�  �<  D�  �]  E�  *w  F�  dW  G�   �F  H�  " e=  J�F  |[  O�G  �� Qa   �\  Ra  red Sa  q  Ta   �[  V�G  �?  (�<H  `a  ��   �L  �<H  r  �<H  &W  ��  �F  �<H    �  Ik  ��G  ��  L�H  }W N   ��  O�  ��  P�   ��  RNH  8y  hl�H  �~  n�   ��  o�  �~  p�H   �H  �H  L    `�  r�H  ,�  0�<I  }W �   ��  ��  def ��  ��  ��  tag ��   cy  ��  ( ˣ  ��H  ��  �}I  Ԛ  �?   cy  ��  �}  ��   	�  �HI  U�   ��I  �~  ��   ��  ��  ˧  ��  �~  ��I  i{  ��I   <I  }I  �  ��I  >i    J2J  tag  L�   ��   M�  /�  N�  �f   O�4   2\   Q�I  G    ��J  Tag  ��   g   ��  �=   ��  Ja   ��   mn   ��J  >J  �v    ��J  �T   ��   �Y   ��  D   ��  S   ��  E]   ��  ;C   ��  �:  �o   �[   ��J  DQ   @K  E]   �   ;C   �  �:  o   �i   K  >M  0 .�K  ��   0�   �Z   1�  vv   2�  �r  3�K  =P   4�  �Q   5�K   ^�   6K  ( �J  @K  �p   8MK  CE   YL  �B   [�   b   \�   Pq   ^L  �K  �m   xNL  ��   z�   �R   {�  Up   |L   �=   ~L  �i   ��L  ��   ��   5�   ��  �"   ��  �"   ��  i!   ��  %!   ��  
2!   ��  �   ��   W   �[L  �U   �M  �   N   
    N  Sd   !a  �Q   "N  �G   #N  �v   $N  �=   %N  sD   &N  �\   'N  �X   (N  	`N   )�M  
 N  �M  L    �T   +�L  >t   �N  �>   ��M   �  ��M  !   �a  m   �a  �[   �a  SX   �a   �<   �N  �M  x@   "jN  �   $�   �`   %�  TL   &�2  �o  'jN   pN  N  �h   )#N  �Z   <�N  �   >�   �f   ?pN   fR   A�N  $ Z�N  %j  \vN  %�Y  ]�N   ms    VO  �   XB   �r  _�N   J   a�N  �t   r!%O  +O  U<  �c  ( ��O  �B  �o   �c   �o  �y  �o  �Y   ��  cC   ��   �   �B  $ 	\   �0O   L   � �O  �O  �i  � �pT  ah  �#   �u   �2J  ��v   ��  �R   ��   o   ��J  (�&  ��@  0�Q   ��A  �@   ��G  �5�   �B  �<   ��B  ��`   ��  0�a   ��K  8#os2  ��D  hF�   ��E  �j   �o  0 M   ��  8w_  �AV  @�>   �rV  H�A   ��V  P^Z   ��V  X�f   ��V  `KT   ��V  h�i   �a   pQ   �a   x#mm  �a   �#var  �a   �g   �a   ��Y  �NL  �Fq  ��F  �jQ   ��  �nQ   �N  �m   O  ��P   BH  @   �  @B   "W  H�u   B  P�u   �G  Q�;   �  XzQ   o  `FN   �  hT   o  p!u   �  x#cvt  �9  �2i   pT  �)   )�	  ��   +�  ��j   -�  �:>   .�  ��_   0B  �S?   3B  �E�   4O  ��W   6r  �XA   8�  �	K   9�  ��c   ?�  �][   @�  ��J   B�  �'<   Co  �	Z   Eo   �q   F�  �G   G�  �T   H�  �a   Io   �\   Ko  (�u   L�  0o   MW  8^C   N�  <:W   O�2  @_   Qo  H�@   R�  P>   S�  X}?   Tr  \m?   Ur  `#bdf  X�O  h�k   \�  ��Z   ]�  �Pl   h�  �(a   i�  �i  ma   ��d  na   � �Q   ��  �g   �"�T  �T  �t  x �AV  ��   ��O   ֳ   ��W  ȩ   ��  �m   �X  �1   ��   x  ��  (^�   �K  0��   ��  8    ��  <�;   �  @�C   ��  `�  ��  d"f  ��  h�I   �B  lpp1  ��  ppp2  ��  �Ǟ   ��W  ��y   ��W  �BJ   ��W  �<   �o  bL   ��   Ud  �a   (�W   ��  0r�   ��  4#pp3  ��  8#pp4  ��  HO�   �o  X��   �o  `�k   ��
  h �^   NV  TV  �  rV  �O  �  K  �4   �D   *V  �V  �  �V  }T  �  �  �   �b   A�V  �V  �  �V  }T   SQ   Q�V  �V  �V  }T   �=  Z    TW  �G   �v  k_  <L  ok   �`   _�V  �G  �j  @ ��W  ڰ   �   �0   ��  q5   ��  
0�   ��      ��  org  �  cur  �  "  �   �    �o  (H�  ��2  0�>   ��  8 ,L   �(W  @\   �'�W  �W  �r  �d   � X  	X  �a  ��  !!�O  ��  `!,BX  ah !.   m !/�  X ��  !1NX  X  !��  H!<�X  ah !>�   "�� !@B  0"��  !AB  1"A� !C�  8"�� !D�  @ ��  !F�X  TX  !�  !Q�X  �  !S�,   ��  !T�X   �,  �X  L   � ;�  !V�X  �X  �  "$$Y  Y  ��   "&?Y  I_ "(S#   ��  ")�2   
��  ".�$  
.�  ";�$  ��  H#4�Y  �-  #6�   �k #7o  ��  #8o  O�  #9o  �� #;�2   top #<�2  (�  #=�  0��  #C�  4��  #Da   8��  #F�  @�  #G�  B ��  #IWY  �  #IZ  WY  Z   #c]Z  `�   ��  �  u�  �  ��  -�  C�  <�  �  	 H�  #siZ  oZ  �  ~Z   Z   ��   #u�Z  ��  #wS    �* #xS   �  #y�  ֳ  #za  ��  #{]Z  C�  #|�  ��  #}�   e�  #�~Z  	�Z  Z   $�;]  x�   ��  ��  ��  �  ��  }�  W�  �  ��  	�  
O�  ��  U�  g�  ��  (�  ��  ��  X�  ��  S�   k�  !*�  "!�  #��  $v�  %��  &��  'r�  (��  0D�  1��  @��  AV�  Q��  R��  SQ�  T��  U�  V3�  W��  X��  `%�  aV�  b��  c"�  p��  ���  ��  �I�  ���  ���  ��  �Y�  �5�  ���  ���  ���  ���  ���  �x�  ���  ���  �n�  ���  ���  ��  �_�  ��  �c�  ���  ���  ��  ���  �8�  ��  �X�  ��  �W�  ���  �Y�  ��  ���  �u�  ��  ���  �E�  �&�  ���  ��  ��  ���  ���  � &?Y  k	��F     &KY  �	@�F     '<  Z   %9�]  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  %V^  <v %Xa   ֳ  %Ya  �  %Z�   yK  %\�]  	^  <e  &I.^  4^  �  W^  K  �O  �  �  @   l  &s.^  Z  &�o^  u^  �^  �O   -H  &��^  �^  �  �^  �O  �  �  o  �4   �e  &2�^  �^  �  �^  �O  �  �  �  K  �^  �^   �  �L  �h  &S_  _  �  -_  �O  �  �4   �^  &p:_  @_  �  Y_  �O  �  Y_   �  eN  &�l_  r_  �  �_  �O  �  �2   Ub  &��_  �_  �  �_  �O  K  B   #K  &��_  �_  �_  �O  B  �  �_  �2   �  3l  &��_  `  �  `  �O  �   �d  &	#`  )`  B  L`  �O  �  �2  �2  L`   u  �J  &0_`  e`  �  �`  �O  �  �  �   CZ  &N�`  �`  �  �`  �O  �  �2   :=  &p�`  �`  B  �`  �O  �  �`  �`   �  �Z  &��`  �`  �  a  �O  K   �^  &�o^  GK  &�'a  -a  �  Fa  �O  �  �   N=  0&�pc  w_ &�"AV   EY &�""^  �e &�"W^  /q &�"c^  ��  &�"�   ob &�"�^  (pR &�"�`  0�^ &�"�_  8D_ &�"�`  @x` &�"�`  HPr &�"�`  P1s &�"�`  X�k &�"�`  `�S &�"a  h�O &�"�`  p�Y &�"�`  xAq &�"�`  ��b &�"�`  �ar &�"�^  ��[  &�"__  � Q  &�"a  �� &�"a  �X &�"�`  ��U &�"�_  �`H  &�"�`  ��W  &�"a  ��n &�"_  ��T &�"-_  �zi & "�`  ��d &"�`  ��Q &"a  ��] &"a  �B  &"�_   UU &"`  �p  &"R`  �[ &"�_  ]o &
"�`   4P &"�`  ( sh  &Fa  AD  &�c  pc  xX  h'*�c  ah ',�$   �q  '.�  8�'  '/B  <iO  '0�c  @��  '1`  ` �  �c  L    Y  '3�c  �c  ��  '?-d  d  �  `'��d  *�  '�o   O�  '�	  z�  '�	  �� '��  6�  '��   ��  '��  $�K '��2  (h�  '��2  0ڰ  '�  8�� '�9e  @ ��   'X�d  �� '[�d   �q '`e  add 'c3e  U1 'ie   �  �d  d  �     �d  e  d   e  �  3e  d  �  �  �   e  H�  'k�d  	9e  ��  '�"Ve  \e  ;�  �'��e  O�  '�o   Ǟ  '�o  ��  '�o  �U '��  ڰ  '�   �� '��i  ( ��  '�"�e  �e  Q�  '�f  �k '�o   ��  '�o  b '��f   K�  '�"f  	f  f  �  0'��f  �  '�   ��  '�g  b 'Mg  ��  '�g  �  '�  ֳ  'a  C�  '�   ��  '	�  $��  '�  ( '��  Z   '��f  ��   }�  ��  ��  �  ��   I�  '��f  '"�  Z   '�Mg  :�   G�  ��  Z�  z�  !�  ��  d�   �  \�  	��  
��  Ѻ   ��  '��f  '��  Z   '��g  ��   ��  F�  r�  ػ  ��  ��  _�  j�  ��  	 e�  '�Yg  [�  '��g  �g  �g  �  	   ��  h'u�h  �� 'x�h   �q '~�h  �Y '��h  �L '��h  ; '��h   �> '��h  (nD '�i  0�M '�=i  8�: '�ai  @�[ '�wi  H�l '��i  P` '��i  X�9 '��i  ` �h  Je  o  o     �h  �h  Je   �h  �  �h  Je   �h  �  �h  Je  �   �h  �  i  Je  o  	  �4  B   �h  �  =i  Je  �  �_   $i  �  ai  Je  �  ?  �   Ci  wi  Je  �e   gi  �i  Je  �e  �  �`   }i  �  �i  Je  f  F   �  �4   �i  :�  '��g  	�i  ��  '��i  ;�  p'4�j  ڰ  '6   ��  '7�  ȩ  '8�X  ��  '9X  Ǟ  ':5/   �  ';5/  (��  '=Lk  0��  '>Lk  8�C  '@  @� 'A  H�;  'C"  P.�  'DB  X�� 'EB  Y8�  'FB  Z��  'HB  [�  'IB  \�� 'K?k  ` ��  '�k  �� '�(k   �q '�9k   "k  "k  a   B   �i  k  9k  "k   .k  ��  '��j  �  ��  'b�k  Ǟ  'do   ��  'eo  O�  'fo   Q�  'hRk  (�  'l�k  �k  �  �k  �O  �  �2  �4   ;�  'r�k  �k  �k  �O  �2  �   w�  �'wn  �I 'y�i   �� '{n  p#top '|?  ��� '~n   �y  ',n  �a�  '��  ��  '��  ��  '�2n  �#cff '��6  ��  '�<   ��  '�Bn  (��  '�Lk  0׹  '�B  8��  '��  <P�  '��  @"�  '��  Dc�  '��  H��  '��  LT�  '��2  P0� '��2  X�o '��2  `�  '��  h;:  '�+  lzd '�B  p��  '�&�k  x��  '�&�k  �Q  '��,  ���  '��  �Z�  '��2  ���  '��2  �}�  '�k	  �	�  '��  �E�  '�k)  �f�  '�(  ���  '��  � �  n  L   0 �k  ,n  L    �k  �  Bn  L    �	  ��  '��k  �  '�#bn  hn  ��  �'<so  ڰ  '>   ��  '?�  ȩ  '@�  ��  'AX  Ǟ  'B5/   �  'C5/  (��  'E�  0��  'F�  8�C  'H�  @� 'I�  P�;  'K  `˹  'L"q  ��� 'MB  �8�  'NB  ���  'PB  �b�  'Ra   ��  'Sa   ��� 'U�p  � ^�  '��o  �o  �  �o  Un  �   G�  '��o  �o  �o  Un  �  �  a   r�  '��o  �o  �  �o  Un  �  �   h�  '� p  p  �  p  Un    �  '��o  ��  '�/p  5p  @p  Un   ؽ  @'��p  �� '��p   �q '�/p  VY '�$so  c '�$�o  f '�$�o   2 '�$�o  (�J '�$p  0� '�$"p  8 �p  Un  �  �  �  B   �p  ��  '�@p  	�p  ��  Z   '�"q  >�    �  /�  i�   v�  '��p  f�  'Whn  ��  'vuq  O�  'xo   Ǟ  'yo  ��  'zo   ��  '|<q  ��  '|�q  <q  �  '/�q  �q  ��  �'�<s  �I '�/q   �� '�Nt  �#top '�(  ��� '�^t  ��y  '��q  x
Q  '��,  �
�  '��  �
�o '��2  �
��  '��  �
��  '��  �
+ '��2  �
��  '��2  �
��  '��2  �
}�  '�k	  �
	�  '��  �
a�  '��  �
�  '��  �
�  '�2n  �
E�  '�k)  `;:  '�+  h��  '��s  p�� '�<t  xf�  '�(  ���  '��  �zd '�B  ���  '��	  � �   '��s  �� '��s   �q '��s  ;U '�t  �" '�6t   õ  '��s  �s  �  �s  �q  �   �  �s  �q  �  �  �  �2  k)  B  +  �s   �s  �s  �q   �s  �  t  �q  o  �   �s  �  0t  0t  o  �   Hn  t  '�  '�<s  	<t  �  ^t  L   � uq  nt  L    D�  '� {t  ��  �'T�u  ڰ  'V   ��  'W�O  ȩ  'X�X  ��  'YX  Ǟ  'Z5/   �  '[5/  (��  ']�  0��  '^�  8�C  '`�  @� 'a�  P�;  'c  `.�  'eB  ��� 'fB  �8�  'gB  ���  'iB  �b�  'ka   ��  'la   ��� 'n�v  � 9�  '��u  �u  �  �u  �u  �   nt  ��  '��u  �u  �u  �u  �  �  a   �  '��u  �u  �  v  �u  �  �   ��  '��u  >�  '�&v  ,v  7v  �u   ש  '�Dv  Jv  �  Yv  �u   ��  @'��v  �� '�v   �q '&v  VY '
%�u  c '%�u  f '%�u   2 '%7v  (�J '%v  0� '%v  8 �v  �u  �O  BX  �X  B   �v  �  'Yv  ^�  '�Cw  Ǟ  '�o   ��  '�o  O�  '�o   ��  '�
w  ��  �'�y  �I '�nt   cff '��6  ��� '�n  �#top '�?  h�� '�y  p�y  '�y  a�  '��  �  '��  �  '�2n  ��  '��  ���  '��  �0�  '�B  �׹  '�B  ���  '��  �f�  '�y  �P�  '��  �"�  '��  �c�  '��  ���  '��  �T�  '��2  �0� '��2  ��o '��2  ��  '��  �;:  '�+  �zd '�B  ���  '�<  ���  '�&�k  ���  '�&�k  � Cw  y  L    Cw  �  'y  L    �  '�Pw  ��  '�0Fy  	4y  �y  +�  '��y  �� '��y   �*  '��y  �" '�6t   	Ly  �y  �y  �O  BX  �X  B  +  �k  �k   'y  �y  �  �y  �y  BX  �   �y  �  '�Ly  	�y  �  '�#z  z  ��  (']z  ڰ  '   ^�  '�z   '�3  F�  '#{  w�  ' a     ӫ  '��z  �� '��z   �q '��z  �i '��z   �  �z  �y    o  o   �z  �z  �y   �z  �  �z  �y   �z  ��  '�]z  	�z  ��  '�#�z  {  ��  �  #{  �  	  a    
{  R�  '-.6{  �{  ��   '/�{  f�  '1�"   ]J '2�"  ��  '3�"  V '4�"   	<{  ��  X'A1|  8�  'D!1|   ��  'E!7|  �  'F!=|  ��  'G!C|  կ  'J^|   *�  'Os|  (��  'R�|  0��  'W�|  8�  '[){  @��  '^!�|  H�  '`"�|  P Ee  �i  �p  It  ^|  o  	  �   I|  r  s|  r   d|  �|  0t  a   B   y|  �|  �  �'  <   �|  �z  �y  4�  'b�|  �{  n�  (�|  �|  �  �|  �  �|  �|  �`   �  ��  ($}  }  �  *}  �  *}   B  3�  ('<}  B}  �  [}  �  �  �2   Y�  (+l}  	[}  ��  (+�}  �  (-/�|   ��  (./}  N�  (//0}   ܨ  )!�}  �}  �  �}  �  �?   *�  )%�}  �}  �  �}  �  �?   ]�  ))�}  �}  �  ~  �   ��  ),~   ~  �  4~  �  4~   �'  ��  )0F~  L~  �  o~  �  �*  �  a   �   ��  )7�~  	o~  �  ()7�~  ��  )9�}   Ъ  ):�}  �  );�}  ݱ  )<~  ��  )=:~    �d  *)%  ��  *,�~  	�~  `p  *,  g *.�~    	�~  �e  *,    V^  +9F  �L  +;�   ��  +<�   �`  +>  {V  +B^  d  �  x  F  x   F  ��  +F�  	~  �N  +F�  �  +HR    	�  ]g  +F�  �  ��  ,!�  �  �  �  �   m�  ,$�  �  �  �  �6  <  �  ?   �  ,*�  $�  a  8�  U?  �   �  ,.D�  J�  B  h�  �9  �  �  ?   d�  ,4t�  z�  �  ��  �9  �  �  ?   ��  ,:��  	��  B�  (,:��  ��  ,<$�   �  ,=$�  Y�  ,>$�  ��  ,?$8�  ��  ,@$h�    	��  ��  ,:	�  ��  
�1  -/   ��  .''�  -�  �  A�  �  A�   �H  �z  .+S�  Y�  �  m�  �  m�   s�  �I  9~  ./��  ��  �  ��  �  �  (   "�  .6��  ��  �  ρ  �  �  ?   ��  .=��  �  .B��  ��  .G�  ��  �  �  �  �   Ӏ  .K��  ݓ  .P%�  +�  �  N�  �  �2  N�  N�  m�   ?  `�  .W�  ��  .Z��  3�  ._x�  ~�  �  ��  �  �2  ?   >�  .d��  	��  y  `.dR�  �~  .f"�   -�  .g"y�  g�  .h"ρ  ��  .i"�  7�  .j"G�   Y�  .k"��  (�  .l"ہ  0&�  .m"�  8U�  .n"`�  @A�  .o"l�  HY�  .r�  P��  .sT�  X 	��  g�  .dc�  R�  �  /'u�  {�  �  ��  �  �  �`   ¦  /,u�  ۧ  /1u�  r�  /8u�  ��  /=u�  ��  /Bu�  ʍ  /Gu�  �  /N�  ֈ  /Q��  	�  ��  @/Qo�  H�  /Si�   ��  /T��  -�  /U��  ��  /W��  ݖ  /X��   p�  /Yă  (#�  /ZЃ  0��  /\܃  8 	��  ��  /Q��  o�  �A  0&(%  �V  0,L%  b�  00��  	��  tG  00ׄ  ]o 02!��   �  03!��   	��  T  00�  ׄ  �<  1��   �  �  �  �  �  �  B   s=  1$*�  0�  �  I�  �  �  a    �  1)Z�  	I�  #P  1)��  R  1+�   bD 1,�   (�  ���  	0�F     (X�  M{~  	 �F     (��  |�~  	��F     (��  ��  	��F     (��  /g}  	��F     (�  @U�  	��F     (!�  ���  	`�F     (��  ��  	 �F     (L�  ���  	��F     �   a�  L   
 	Q�  (�  	a�  	 �F     )�  d	`�F     �  ��  L   	 	��  *��  ���  	 �F     *��  ���  	��F     �Z  ��  L   L 	І  (9�  g#��  	 �F     �  �  L   � 	��  *��  +�  	 �F     �  7�  L   � 	'�  *>�  L7�  	��F     �  b�  L   V 	R�  *��  eb�  	 �F     �  ��  L   � 	}�  *��  t��  	 �F     *��  ���  	 �F     +�  �peB            ��  ,ϖ ��  U -q�  ��  �dB     x       �E�  ,ϖ ��  U.K ��c  �� �� (��  �r  �t /��  c��B     �      �  0��  c�  � � .��  eX  {� s� .ڰ  f  �� �� .�i  g}c  � �� 1ʑB     D      M�  2cff t�6  &� $� 3̳  ڑB       �  y	8�  4ڳ  K� I� 5 �  6�  p� n� 6��  �� �� 7K�  (�B       (�B            �		�  4f�  �� �� 4Y�  �� �� 85�B     ] 9U|   3S�  \�B      P�  �	��  4a�  � �  3�  ��B       ��  �	\�  48�  C� A� 4+�  h� f� 5��  6E�  �� �� 3S�  ��B      Т  }F�  4a�  �� �� 4a�  �� �� 4n�  �� �� 8��B     | 9U}   8��B     | 9U}    3K�  �B      �  �	��  4f�  �  � 4Y�  W� U� 8��B     ] 9U| 9Ts�  34�  ��B      @�  �	��  4O�  |� z� 4B�  �� �� 8�B     � 9Ts�&  :�B     ��  �  9Us� :��B     ��  *�  9Us�
 :��B     ��  B�  9Us8 :�B     ��  [�  9Us�
 :Q�B     | s�  9U|  :�B     ��  ��  9Us�'9T|  :8�B     | ��  9U|  :R�B     |   9U|  :l�B     | ڋ  9U|  :��B     | �  9U|  :��B     | 
�  9U|  :ϓB     | "�  9U|  8�B     | 9U|    8�B     | 9U~   7o�  �B      �B            ��  4}�  �� �� ;�B            6��  �� �� < �B     9Uv    <ʑB     9Uv   -��  ��  0�B     ?&      ��  0^�  �!K  J� � 0��  �!�  �� }� 0�  �!�  �� �� 0�[  �!�  �� �� 0\  �!@  k� Y� .��  �X  h� :� .�U ��  S� O� .�i  �}c  �� �� .Q  ��,  � � .�  �Y1  �� �� .g  ��|  � � .��  ���  4� *� .��  �B  �� �� .�_  �B  �� X� .j�  �B  N� B� .�-  ��  �� �� =�  ]кB     =(�  <@�B     >��  ��  .ϖ �  =� ;� .6e  	  j� `� 8��B     � 9T	׷F     9Q1  >�  ��  .ϖ �  �� �� .6e  	  � � 8שB     � 9T	��F     9Q1  > �  �  2cff \�6  �� �� .��  ]�;   � � .ڰ  ^  d� `� .�1  _`  �� �� 2i `�  O� I� 1��B     _       �  2mm �'W�  �� �� 2var �'t�  �� �� .�' ��  � �� ?��B     ܏  9U} 9T~  <ܳB     9U}   >Ь  �  .�3  ��  D� <� .�  �  �� �� 2upm ��4  .� $� .�S  ��  �� �� :4�B     � b�  9Ts  :O�B     � z�  9Ts  :j�B     � ��  9Ts  :��B     � ��  9Ts  :��B     �   9Ts  :��B     � ڐ  9Ts  8ֻB     � 9Ts   > �  ��  2sub �;  �� �� 2top �;  7� 1� .�3  �  �� �� .�    �� �� 2upm 	�4  ?  9  .�S  
�  �  �  1��B     k       ��  .�  �  �  �  :ҴB     � ő  9Uv 9T|� 9Q~  :�B     � �  9U|� 9Tv 9Q~  8��B     � 9Q~   :ݵB     � �  9T~  :�B     � /�  9T~  :�B     � G�  9T~  :�B     � _�  9T~  :%�B     � w�  9T~  :7�B     � ��  9T~  8I�B     � 9T~   >0�  Ԗ  .�  L�     12�B     F       q�  .�U q�   � � 3��  b�B      �  v$Z�  4Ӫ  � � 4ƪ  � � 5�  @�  ��6�  	  8j�B     � 9U��}9Q    8?�B     ]�  9U��}  >��  ۔  .��  ��   . , .w�  ��   _ Q .�V ��   � � 3��  нB      Э  �'�  4Ӫ  I G 4ƪ  p l 5Э  @�  ��6�  � � 8սB     � 9U��}9Q    3�  ܽB      �  �Ĕ  4:�  � � 4-�  	  5�  6G�  . , 6T�  S Q Aa�  @�  ��  6b�  � v  :�B     � ��  9Us  8�B     � 9U|    8�B     ]�  9U��}  > �  ��  .&�  ��   R P 7��  |�B      |�B            �$�  4Ӫ  w u 4ƪ  � � ;|�B            @�  ��6�  � � 8��B     � 9U��}9Q    8n�B     ]�  9U��}  >��  ˕  .��  ��   � � 8��B     ]�  9U��}  3��  I�B      p�  �!F�  4Ӫ    4ƪ  = 9 5p�  @�  ��6�  w u 8N�B     � 9U��}9T	�F     9Q    7q�  ��B      ��B     �       ��  4�  � � ;��B     �       6��    6��  � � 6��  � �   8��B     ��  9U��}9T��}�  >P�  ��  (a�  r  ��.I_ F  { s 2nn �  � � .T %5  \	 X	 >��  w�  .Oe ?�"  �	 �	 8��B     � 9U	��F     9T09Q��9R0  8ڹB     � 9U	@�F     9T09Q��9R0  3�  T�B      ��  gZ�  4b�  :
 
 4U�  � ~ 4H�  � � 4;�  "  4.�  � � 4!�  4  4�  � � 5��  @��  ��~6��  "   6��  Q G 6��  � � @��  ��~6Ǵ  ,  BԴ   �B     Bݴ  ͰB     A��   �  ��  @��  ��6�  i ] 6�   � 3��  .�B       `�  c	5�  4��  � � 4��  � � 4��  a C 4��  � � 5`�  6��  � � @��  ��6��  � � 6�  � � 6�  � � B�  _�B     A$�  Ъ  �  6%�  J D 62�  � � 6?�  � � CL�  |�B     �       w�  6Q�    C^�  ��B     �       K�  6_�  S Q 6l�  x v 6y�  � � 6��  � � :��B     � �  9Us 9T  :��B     � 0�  9Us 9T  8�B     � 9Us 9T   8��B     	 9U��}9TH9Q09X09Y   C��  @�B           :�  6��  � � :j�B      ��  9Us  :��B     " Қ  9Us 9T4 :��B     � �  9Us 9T  :��B     	 �  9U��}9T49Q09X09Y  8�B     � 9U| 9T   :��B      R�  9Us  :��B     " o�  9Us 9T2 :пB     / ��  9Us  :�B     � ��  9Us 9T  :��B     < Û  9Us 9T  :��B     � �  9Us 9T  :�B     	 �  9U��}9T89Q��}9X��}9Y  :a�B     < 4�  9U} 9T  :��B      Y�  9Us 9T	��~��~" :��B     � w�  9Us 9T  : �B     � ��  9Us 9T  :7�B     	 Ĝ  9U��}9T89Q09X09Y  8�B     	 9U��}9T@9Q09X09Y   :s�B     | �  9U��}9T��} 8P�B     ��  9U��}#�'9T��}   3��  ��B       �  �	=�  4��    4��  B < 4��  � � 4��  � � 5�  @��  ��~6�    6�  K G B!�  ��B     B*�  ��B     :�B      ޝ  9Us  :'�B     I ��  9Us 9T��~ :q�B     � �  9Us 9T��~ 8��B     V 9Us 9Q��}#�&   :��B      U�  9Us  :ڮB     q�  ��  9U 9Ts 9Q09R��~� :"�B     	 ��  9U��}9T
�9Q09X09Y��} :��B     t�  ��  9T 9R| 9X��}9Y~  8ڰB     ��  9U   C�  h�B     R       8�  6�  � � 8��B     I 9Us 9T��}  A&�  P�  ;�  6'�  � � 3e�  ��B       ��  �	G�  4��  � � 4��  ! 	! 4��  {! m! 4��  *" " 4��  �" �" 4w�  # # 5��  6��  �# �# @��  ��6��  �$ �$ B��  h�B     A��  �  O�  6��  z% p% C�  ��B     �       ��  6�  �% �% 6�  U& Q& :��B     � [�  9Us 9T  :�B     I y�  9Us 9T  Dr�B     �  :=�B      ��  9Us  :d�B     I ��  9Us 9T  :��B     	 ��  9U��}9T29Q09R| ����9X09Y  :��B     c "�  9Us 9T|����1$���� :�B     p :�  9U}  8>�B     } 9Us   :��B     	 ��  9U��}9T29Q09Rv 9X09Y�� :\�B     ��  ��  9U��}9T| 9Q��} :��B     	 �  9U��}9T29Q09Rv 9X09Y�� :��B     | ��  9U  :��B     | �  9U  8��B     	 9U��}9T29Q09Rv 9X09Y��   E8�  ��B       �  �	4��  �& �& 4~�  ' 	' 4q�  �' �' 4d�  �' �' FW�  4J�  ^( T( 5�  @��  ��6��  �( �( 6��  �) �) 6��  �* �* 6ʽ  + + B׽  9�B     B�  N�B     A6�  p�  ��  67�  �+ �+ 6D�  ], W, G|�  ��B      ��B            .F��  F��  4��  �, �, ;��B            6��  - -    C��  1�B           ��  6��  P- N- 6�  {- s- 6�  �- �- :i�B     I �  9Us 9T  8��B     I 9Us 9T   A#�  ��  l�  6(�  . . :S�B     I 3�  9Us 9T  :��B     I Q�  9Us 9T  8��B     � 9Us 9T   C�  ��B     ~       Ȥ  6�  [. Q. :�B     c ��  9Us 9Tv � 8s�B     } 9Us   :o�B     ��  �  9U��}9T|  :��B       �  9Us  :��B     I �  9Us 9T  8�B     I 9Us 9T     :��B     / S�  9Us  :׫B     � ��  9Us 9T	��F     9Q��} :'�B     � ��  9Us 9T��} :Y�B      ��  9Us  :��B     / Х  9Us  :جB     " �  9Us  :�B     q�  �  9U��~9Ts 9Q19R1 :��B     t�  d�  9U��}#�9Tv 9Q��~�9Rs 9X 9Y	�0| �0)(  �#�` :ͭB      |�  9Us  :��B     q�  ��  9U��}#�
9Ts 9Q09R��~� :��B     ��  Ʀ  9U��~ :бB      ަ  9Us  :��B     q�  
�  9U��}#89Ts 9Q09R0 :;�B     q�  2�  9Uv 9Ts 9Q09R0 :f�B     q�  [�  9U��~9Ts 9Q19R0 :��B     q�  ��  9U��~9Ts 9Q19R0 :ͲB     <�  ��  9U��~9T��}#�9Q��}#�9R��}#� :�B     ��  ا  9U��~ :��B     ��  �  9U��~ :�B     ��  
�  9U��~ :5�B     <�  9�  9U��~9T��}#�9Q09R0 8��B     ��  9U��}9T��~�   86�B     � 9U��}9T
�9Q��~  :k�B     � ��  9Uv 9T	��F      :��B     � ɨ  9Uv 9T	P�F      :��B     � �  9Uv 9T	�F      :�B      �  9Us 9T0 ?�B     <�  9Us 9T} 9Q~ 9R��}�9X��} ?O�B     d�  9U} 9Tdaeh9Qs 9R0 ?i�B     ~�  9U} 9Ts  ?��B     ��  9U} 9T2FFC9Qs 9R0 :��B      é  9Us 9T0 ?G�B     ��  9Us 9T} 9Q~ 9R��}�9X��} <l�B     9U} 9T FFC9Qs 9R0  k	  H��  �q�  I�U �#  I�  �#{  J�  �`  J)�  �#`  KLidx ��    H��  ���  I}W �%  Lidx �`  J��  �`  J��  �B   Mf�  �  ��  Iڰ  �!  I�; �!{  J�U ��  J�Y  �   N7�  e�  pfB     T       ��  0�  e �  �. �. .��  gX  8/ 2/ .�  h�6  �/ �/ .�  iY1  �/ �/ ;�fB     .       .ϖ n�  �/ �/ 1�fB            ë  .�� uS/  0 	0  8�fB     � 9T	P�F        +;�  ^�dB            ��  ,�  ^ �  U -"�  �  0|B     D      �l�  0ֳ  &�  80 .0 Oreq &�  �0 �0 .��  BX  61 ,1 .�� �-  �1 �1 >��  ��  .��  X  �1 �1 .�i  }c  2 
2 (m �  ��?_|B     �  9Ts 9Q�� 8e}B     l�  9Uv   1�|B     �       =�  .��  0X  32 12 .�  1�6  Y2 W2 .�L  2�X  ~2 |2 .��  4�  �2 �2 2i 5�  �2 �2 >�  (�  2sub ><  �2 �2 .��  ?�  23 ,3 .A� @�  �3 }3 .�� @�  �3 �3 :�|B     � �  9T| 9Q�� :}B     � �  9T| 9Q�� <}B     9R09X0  <�|B     9R09X0  :||B     � U�  9Ts  8�|B     � P��  v   Q��  ��  �zB     �       �H�  Rֳ  ��  "4 4 Rm ��  r4 n4 S��  �BX  �4 �4 S�� ��-  5 �4 1�zB     �       �  S��  �X  95 75 S�  ��6  _5 ]5 S�L  ��X  �5 �5 S��  ��  �5 �5 Ti ��  �5 �5 >p�  �  Tsub �<  �5 �5 S��  ��  86 26 SA� ��  �6 �6 S�� ��  �6 �6 :+{B     � ί  9T| 9Q�� :C{B     � �  9T| 9Q�� <_{B     9R09X0  <�zB     9R09X0  :�zB     � 1�  9T�T 8�zB     � P��  v   QH�  ��  �}B     >      ��  R��  ��  *7 "7 Sֳ  �BX  �7 �7 *�U ��  ��}S�� ��-  �7 �7 U�  ��~B     >@�  ��  S��  �X  k8 i8 S�  ��6  �8 �8 S�L  ��X  �8 �8 *��  ��'  ��}Sڰ  �  r9 p9 Ti ��  �9 �9 1Z~B     C       ��  Tsub �<  �9 �9 :l~B     �  ��  9Tt  <�~B     9T��}9Q s "  :�}B     � ��  9T
9Q��} :~B     �  ܱ  9U}�9Tt  <(~B     9T��}9Q   D�}B     �  V��  u�fB     �      �}�  R��  u'<  �9 �9 W��  v'�'  TS��  x�>  $:  : Tn y�  �: `: S/� y�  < �;  X��  R�{B     �       �~�  R��  R�  �< �< Sڰ  T  �< �< Sֳ  UBX  = = S��  VX  Z= X= S�  W�6  �= ~= S�L  X�X  �= �= 5��  S�� ]�-  > > 1�{B     -       T�  Ti c�  K> G>  :�{B     � o�  P��  �U Y|B     |   Z;�  A�-  ̳  [ֳ  A)BX  \��  CX  \�  D�6  \�  EY1  \ϖ F�   H��  �	�  I�  �	�6  Jڰ  �	  Lidx �	�   M��  ��  6�  I�-  ��  I^�  �K  I�  ��  I�  ��6  I��  �X  I��  �B  I�_  �B  (q�  �"F�  	��F     J�U ��  Jڰ  �  J��  ��  J��  ��;  J�  ��4  JJ�  ��  ]�  �	]��  �	^��  J��  �a   ^&�  J��  \	�4  Lsub ]	<  Lidx ^	�   KJl�  �	B    ^  F�  L    	6�  H��  pt�  Iڰ  p"  I��  q"<   NB�  ��  0�B     �      �B�  0��  �"<  �> �> Oidx �"�4  ? �> 0M�  �"�  @ @ 0^�  �"K  �@ �@ 0��  �"�  �@ �@ 0�* �"�  xA rA 0�  �"�6  �A �A 0��  �"X  B B .�U ��  hB >B (��  ��Y  ��~(��  �o  ��~(�  ��  ��~2top ��;  D 
D .��  ��>  bD \D .g  ��|  �D �D .�_  �B  (E $E .�  ��  vE lE =�  h,�B     1�B     A       ,�  .K 6�c  &F $F  3��  ��B       �  �'�  49�  MF IF 4-�  MF IF 4!�  �F �F 4�  �F �F 4	�  )G %G 4��  gG _G 4��  �G �G 5�  6E�  H H @Q�  ��~B]�  !�B     :�B     	 �  9U} 9T89Q09R	�0s  $0)( 
�#`9X09Y��~ 8�B     | 9U}    3\�  ٦B      ��  ��  4j�  IH EH 4j�  IH EH 4w�  �H H _��  ��B            6��  �H �H 8̨B     � 9T}    7��  ,�B      ,�B            i�  4��  �H �H 4��  �H �H ;,�B            6��  	I I D9�B     |   :æB     ��  =�  9Uv 9T��~�9Q} 9R��~ :\�B      U�  9U|  :w�B     V s�  9U| 9Q}  :��B     ��  ��  9U��~ :��B     � ��  9U| 9T}  :ԧB     B�  ӹ  9U� 9T~ 9Q09R0 :i�B      �  9U|  :��B     q�  �  9Uv 9T| 9Q19R
s  $0)� 8��B     <�  9Uv 9T~�	9Q09R0  -�  P�  0�B     �      �8�  0�  P'�6  9I /I 0��  Q'<  �I �I 03�  R'�  gJ UJ ONDV S'?  EK 1K .�U U�  8L "L (��  V�Y  ��~2top W�;  *M M .��  X�>  �M �M .^�  YK  �N �N .�  Z�  �N �N =*t  �\�B     =�  ���B     3��  +�B       p�  w
7�  49�  �N �N 4-�  :O 6O 4!�  wO sO 4�  �O �O 4	�  �O �O 4��  aP ]P 4��  �P �P 5p�  6E�  �P �P @Q�  ��~B]�  (�B     :n�B     	 !�  9U~ 9T89Q09X09Y��~ 8�B     | 9U~    7|�  ��B      ��B            �l�  4��  Q Q  7��  ݚB      ݚB            �ڼ  4��  :Q 8Q 4��  :Q 8Q ;ݚB            6��  bQ `Q D�B     |   :��B      �  9Us  :��B     c 
�  9Us  :R�B     ��  #�  9U��~ 8\�B     } 9Us   M��  Y�  S�  IT Y$%5  I�  Z$�5  I�  [$�  I^�  \$K  I��  ]$�  I�  ^$�  J�U `�  J/� a�  Lj b�  J��  c�  J��  d�  ]�  D];�  ^��  Lp �o   ^#�  J��  ��  Li ��  Lk ��   ^6�  JJ�  ��   KLsid )�  Lgid *�    H��  Po�  IT P$%5   H��  C��  I��  CX  Lmm EW�   -U�  1�  �dB     
       �e�  0��  1#X  �Q �Q 0�  2#�2  �Q �Q 0Ԛ  3#N�  R R 0��  4#N�  CR ?R 0;�  5#m�  �R |R 2mm 7W�  �R �R `�dB     9U�U9T�T9Q�Q9R�R9X�X  -��  B  �oB     ;       ��  0E�  &�9  �R �R 0y�  &�  !S S 03�  &�  ^S ZS ONDV &?  �S �S 8�oB     � 9U�R9Q�Q����3$  -��  k�  �oB     �      �_�  0E�  k&�9  �S �S 0y�  l&�  �T �T 03�  m&�  6U *U ONDV n&?  �U �U .�U p�  VV TV .ڰ  q  ~V zV 2len s�  �V �V 2vs t�6  PW JW .��  u�6  �W �W .�  v�  �W �W =�  KrB     >��  ��  2j ��  �X �X 2idx ��  �X �X J��  ��6  5К  .�~  �A6  �X �X .I�  ��  gY eY 7�
 �qB       �qB     $       ���  F�
 4�
 �Y �Y ;�qB     $       6�
 �Y �Y 6�
 �Y �Y   D"rB     �   :�pB     	 �  9U��9T19Rs 2$9Y�� :�rB     	 B�  9U��9T19Rs 9Y�� 8�rB     � 9T��9Qs   M��   �  v�  IP�   #<  I��  # Z  I��  #�  J�� �  JǞ  �  Li �  Lj �  Jֳ  �  JE�  	�9  Jڰ    J�U �  J��  �  J/� �  ]�  a^Y�  J+�  !o  J��  "o  KJ�  4	  Lp 5�2    KJ��  Fv�  Lsum Gr    m  HE�  ���  IP�  �!<   M�  a�  ��  I��  a$��  I^�  b$K  I��  c$�  I�  d$�  Jڰ  f  J�U g�  J��  i�4  Li j�  Lj j�  ]�  �KJ�  p�  J��  q�  J}�  r�  ^��  J��  ��6  KJ�~  �A6  J��  �5  J��  �5  J*�  �&5    KJKl  ��6     �6  +��  D�eB     �       �e�  0��  D$��  8Z 2Z 0ڰ  E$  �Z �Z 2i G�  �Z �Z :�eB     |  �  9U}  :fB     | 8�  9U}  :8fB     | P�  9U}  8RfB     | 9U}   M��  ��  �  I�  �"�5  I�  �"�  I^�  �"K  I��  �"�  I�  �"�  Il�  �"B  Jڰ  �  J�U ��  J��  ��  ]�  4KLj ��  KJ��  ��  Li ��     H��  wS�  I�  w"�5  I^�  x"K  Jڰ  z   H��  n|�  I�  n'�5  Iڰ  o'   M7�  `�  ��  I�  `+�5  acid a+�  J�Y  c�   -t�  ;�  �nB     �       ���  0�  ;*�5  �[ �[ 0�  <*�  \ \ 0ڰ  =*  �\ �\ (�U ?�  �\2i @�  $]  ] 2j A�  ^] \] ."�  B�  �] �] =�  Z�nB     :#oB     	 ��  9U�Q9T29Q09Rs 
��#9X09Y�\ 8�oB     	 9U�Q9T29Qs 9R19Xs 9Y�\  -U�  �a  �cB     �       ���  ,�  �$U?  U,x �$�  T2fd �a  �] �] =�  -�cB     5 �  2p 
o  q^ c^ .��  o  _ _ 2fd2 a  N_ F_ .��  �  �_ �_ .��  �  .` $`   M��  ��  4�  I�  �%U?  I�  �%�  I^�  �%K  I�  �%�  J�U ��  J��  �a  J�  ��  ]�  �]��  � H>�  �]�  I�  �%U?  I^�  �%K   M��  �  ��  I�  �'�6  asid �'�   M��  �  ��  I�  �#�6  I��  �#�   -�  c   �B     �       �\�  0�  c!�6  �` �` 0��  d!�  ba ^a 2idx f�4  �a �a .ڰ  g  �b �b (Vu  ho  �P(��  i�  �X(�U j�  �L.}W k  �b �b =�  ��B     3\�  ��B      ��  }��  4j�  hc `c 4j�  �c �c 4w�  Ld Dd _��  ��B            6��  �d �d 8��B     � 9T�P   :I�B     ��  )�  9Us89T�T9Q�P9R�X :g�B     � G�  9Uv 9Q�L 8́B     � 9Uv   Hf�  T��  aidx T(�4  I�^  U(�2  KJ^�  YK    -��  ��   B     �      �<�  Oidx �(�4  �d �d 0��  �(�  re he 0�^  �(�2  �e �e 0-�  �(�4  �f �f .�U ��  g g =�  NDB     5��  .^�  �K  9g 3g .� ��  �g �g .� ��  �g �g 18�B     �       �  2pos �  �h �h :Y�B      ��  9U  :u�B     M ��  9T} 9Q��P[�  s  8��B     M 9T} 9Q��P[�  s   :�B      �  9U  8��B     V 9U 9Tv 9Q~    -��  ��  �rB           �I�  Oidx �'�4  �h �h 0�B �'I�  ^i Ri 0}�  �'�2  �i �i 0�  �'�4  �j �j (�U ��  ��.ڰ  �  Ck ;k 2t ��2  �k �k .v�  �o  �l wl .v  ��  8m 4m =�  ��tB     >�  ��  2n ��  �m �m .��  ��  >n .n .)  ��  o �n .�  �o  �o �o 5��  .i�  ��  �o �o DtB     �   3O�  �tB      Л  ���  4a�  mp ep 5Л  @n�  ��6{�  �p �p 6��  5q -q B��  �uB     A��  0�  ��  6��  �q �q 6��   r r 6��  +s s 6��  t t 6��  �t �t :�tB     	 ��  9U| 9T89Q09Rv 9X09Y�� :?uB      ��  9U  :iuB     c ��  9U 9Tv  8�uB     } 9U   8uB     | 9U|    :DsB     	 %�  9U| 9T89Q09R}����9X09Y�� 8xsB     � 9U| 9T��9Q��  �2  MI�  V�  ��  aidx V&�4  J�U X�  J^�  YK  Jڰ  Z  ]�  �KJ	�  _a  J��  `�  Lp ao  J��  bo  J�  c�4    +:�  D`hB     a       �q�  Oidx D�4  �u �u 50�  .^�  HK  'v %v .ڰ  I  Lv Jv :�hB     � [�  9Ts8 8�hB     | 9Uv    Q��  ��  ��B     �      �J�  bidx ��4  v ov R^�  �K  Bw 0w R" �B  
x x R�_  �B  Gx Cx *�U ��  ��Sڰ  �  �x �x S/� ��  �x �x =�  ;`�B     >�  ��  .	�  	a  |y xy .ֳ  
�  �y �y :؂B     I }�  9U} 9T  :�B     " ��  9U}  :.�B     M ��  9Ts9Q P[�  s  :\�B     V ��  9U} 9Qs8 8�B     " 9U}   :5�B     / �  9U}  :I�B     < $�  9U} 9T  :��B     | <�  9Uv  D��B     �  Z��  ��  ��  cidx �%�4  [��  �%��  \�U ��  \^�  �K  dtmp ���  \�Y  ��  Kdnn ��    �  a  ��  L    Q��  ��  �cB            ���  R�_ �'�  ?z ;z  -��  ��  ЕB     T      ���  0��  � Z  �z xz 0�k �o  { { 0��  �o  W{ I{ 2p �o  %| �{ .�U ��  ?~ 7~ =��  F��B     =�  =��B     ]��  N]��  J=s�  �0�B     =cs 3P�B     5p�  2v ��  �~ �~ 5Ф  .�* �#�  7� )� .A�  �#�  � Ӏ .#` �#��  ؁ ʁ 5 �  2val ��  �� � 2q �o  � � 1�B     �       ��  .I�  �o  v� r� .Kl  ��2  ȃ ă 8J�B     � 9U} P��  ~   7��   �B       �B            �+�  4�  � �� 4�  '� %� 4��  M� K� 80�B      9U} 9Q3  7!�  p�B      p�B            ���  4@�  r� p� 43�  �� �� 8}�B      9U} 9Q0  ?��B     ��  9U}  8��B     � 9U}      �Z  -+�  �  0�B     /       �V�  0��  # Z  �� �� .��  �;  � � .Kl  �2  c� ]� .�U �  �� �� =�  )X�B     8F�B     � 9U�U  -��  ��  ��B           �)�  0��  �  Z  �� � .��  ��>  q� k� .P�  �<  �� �� .E�  ��9  �� �� .��  ��  L� J� .�U ��  u� o� =�  ��B     3_�  2�B       �  ��  4��  ć �� 4~�  �� �� 4q�  8� 4� 5 �  6��  x� n� 6��  � � 6��  � � 6��  R� J� 6��  Ӊ ˉ 6��  <� 8� 6��  |� x� @��  ��6��  �� �� 6	�  �� � B�  ��B     CY�  ��B     �       :�  6Z�  ,� &� 6g�  }� w� :ʞB     � %�  9U}  8�B     � 9U}   _�  ��B     �       6$�  ɋ ǋ 61�  �� � C>�  p�B     H       ��  6?�  )� '� 6L�  P� L�  8%�B     	 9T19X~ 9Y��    :��B     e�  ��  9Us 9Tv 9Q| 9R~  :�B     �  �  9Us 9Tv 9Q| 9R~  8%�B     � 9U}   -o�  ��  ��B     G       ���  0��  �" Z  �� �� .��  ��>  ߌ ٌ .Kl  ��2  /� )� .E�  ��9  �� � .�U ��  �� �� =�  ���B     8�B     � 9U�U  -��  ��  `�B     ^       ���  0��  �" Z  Ӎ ͍ .��  ��;  !� � .Kl  ��2  K� E� .�U ��  �� �� :��B     � s�  9Us P��  v  :��B     � ��  9Us P��  v 8��B     � 9Us P��  v  -��  i�  ��B     m       �B�  0��  i* Z  ێ Վ .��  k�;  )� '� .�U l�  O� M� 5��  .��  ~�  x� t� 8�B     � 9Us    -0�  :�  0�B     j       �"�  0��  :' Z  �� �� .��  <�;  /� -� .Kl  =�2  ]� S� .�U >�  א ѐ =WD  `0�B     5�  2tmp E�  -� %� :`�B     � �  9Us P��  v  8y�B     � 9Us P��  v   -`�  �  ��B     �       �?�  0��  $ Z  �� �� .��  �;  ߑ ݑ .�;  "  � � .Kl   �2  6� .� .�U !�  �� �� 3!�  �B       ��  (�  4@�  ݒ Ւ 43�  C� ?� 8�B      9Uv 9Q0Pk�  s   3!�  !�B      �  )\�  4@�  � y� 43�  Г Γ 8&�B      9Uv 9Q0Pk�  s  3!�  ?�B      �  *��  4@�  �� � 43�  3� 1� 8D�B      9Uv 9Q0Pk�  s  3!�  ]�B      @�  +
�  4@�  X� V� 43�  � }� 8b�B      9Uv 9Q0Pk�  s  D�B     � D.�B     � DL�B     � Dj�B     �  -�  ��  ��B     E      �u�  0��  �& Z  �� �� .��  ��;  � 	� .�3  ��  1� /� .�  �  [� Y� 2upm ��4  �� �� .Kl  ��2  �� �� =��  �B     5P�  (
Q �u�  ��~(i�  ���  ��.��  ��  �� �� .��  ��  � � 2i �S   o� m� > �  ��  .<v ��  �� �� .9�  ��  m� g� .4�  ��  Ƙ ��  3��  ��B       ��  �^�  4��  �� ~� F��  4��  R� J� A��  �  8�  6��  �� �� 6��  9� '� D��B     � :��B     ��  *�  9Uv 9Tt  D��B     �  8s�B     ��  9Uv 9Q09R�  "p  8e�B     � 9U}�    �  ��  L    �  ��  L    M��  s�  ��  I��  s( Z  ad t(�2  I�  u((  KJ3 }�  J��  ~�    M��  g�  !�  I��  g' Z  ad h'�2  I�  i'�   M��  ]�  L�  I��  ]  Z  ad ^ �2   M	�  1�  ��  I��  1 Z  ad 2�2  I�  3�  ]��  TKLval 9�    MK�  �  ��  I��   Z  ad �2   Q��  ��  �iB     �      ���  R��  � Z  � �� R�k �o  � � Rn�  ��  X� @� R�  �(  f� ^� Tp �o  ў Ş Tnib ��  c� S� S^�  ��  � � .�Y  �  Ӡ à .3 �  �� ~� .o�  �  � � .�} �   � � e��  �   .��  ,�  �� }� .�  �  ,� $� .��  �  �� �� .��  -�  � ĥ fBad =�  �BjB     ]��  �=��  �BjB     1kB     D       ��  .��  ��  4� 2� .m�  �+�  Y� W�  3��  �iB       �  ��  4��  �� |� 4��  �� �� 4��  �� �  7��  skB      skB     
       j/�  4��  ,� *� 4��  Q� O� 4��  v� t�  7��  �kB      �kB     
       C~�  4��  �� �� 4��  �� �� 4��  � �  D�lB     � DmB     � :-mB     � ��  9T: 8xmB     � 9T| 3$ �F     "  Q0�  ��   cB     �       ���  W��  �" Z  UW�k �"o  TTp �o  � � Tv ��  V� D� Tval ��  B� 0� gBad �JcB     U�  �JcB     h��   cB      ��  ���  4��  � � 4��  )� '� 4��  R� N�  i��  JcB      JcB            ���  4��  �� �� 4��  �� �� 4��  ث ֫  h��  hcB      И  �9�  4��  �� �� 4��  $� "� 4��  M� I�  j��  �cB      �cB            �4��  �� �� 4��  �� �� 4��  Ӭ Ѭ   Z�  u�  ��  [��  u) Z  [��  v)o  [��  w)o   k��  b��  [��  b  Z  \ڰ  d   Z��  *�  f�  [��  *  Z  [�* + �  [��  , a   [�-  - �  [�  . �  [��  / �  [�  0 �  \ڰ  2  \�U 3�  l�  K Q*�  ��  P�B     �
      ���  Rȩ  �!�X   � �� Rֳ  �!BX  y� _� Rx �!�  �� �� R�1  �!`  |� d� S�U ��  �� ԰ *LM �'y  ��s*�  �Hn  ��iS��  ��O  h� `� Sn�  �B  в Ĳ \��  �B  S�  �#B  s� [� Tcff ��6  � w� Sg  ��|  � ۴ S �  �Ay  O� G� *}�  �k	  ��iS	�  ��  ӵ �� ]�  �>`�  ��  S3�  �X  � � S�i  �}c  ?� 9� S^�  �K  �� �� 5��  (�e �L  ��s>��  ��  .1�  B  �� � (� �  ��i(��  �  ��i?��B     ��  9U~ 9T09Q��i�9R��i9X��i <H�B     9U~ 9T19Q��i�9R��i9X��i  <�B     9U~ 9Q��i�9Rv 9Ys�   >��  ��  .��  d�  C� A� .��  d�  j� f� .��  ea  �� �� :0�B     ��  F�  9Uu 9T��i� :��B     � f�  9T 9Q��h 8ЈB     � 9T 9Q��h  > �  ��  (9� �o  ��i(��  ��  ��i10�B     7       ��  .��  ��4  � ޸  ?.�B     
�  9U��s9T~ 9Q| 9Rs 9Yv @&? :k�B     ��  9�  9U~ 9T��i�9Q��i9R��i ?��B     ]�  9U��s9T| 9Q��i� ?��B     ~�  9U��i9T��s9Q0 ?ʆB     ��  9U��i :�B     ��  ��  9U~ 9T��i ?'�B     ��  9U��s <��B     9U��i  1C�B     i       �  (�e �"N!  ��i<��B     9T��i�9Q09R��i  1B     Y       J�  .�L  w  � �  >Р  R�  (�'  #  ��i.�e $��  /� +� .1�  %B  o� i� 1ǊB     G       ��  (�"  *�  ��i(i!  +�  ��i<��B     9U~ 9T09Q��i�9R��i9X��i  >��  J�  (2!  E�  ��i(�  F�  ��i<�B     9U~ 9T19Q��i�9R��i9X��i  >`�  /�  2n ~�  �� �� 2cur 5/  � � 2vec �  2� (� .A� ��  �� �� .�� ��  � � 7�
 `�B      `�B            �" �  F�
 4�
 %� #� ;`�B            6�
 N� J� 6�
 �� ��   7�
 ��B      ��B            �"��  F�
 4�
 λ ̻ ;��B            6�
 �� � 6�
 :� 6�   3�
 0�B      ��  ���  F�
 4�
 y� u� 5��  6�
 �� �� 6�
 �� ��   G�
 U�B      U�B            �F�
 F�
 ;U�B            6�
 7� 3� 6�
 z� v�    3�
 ��B       �  k"��  4�
 �� �� 4�
 ޽ ܽ 5 �  6�
 � � 6�
 J� F�   3�
 �B      0�  m"��  4�
 �� �� 4�
 �� �� 50�  6�
 ׾ Ӿ 6�
 � �   :��B      ��  9U| 9T��i :"�B      �  9U| 9T} 9Q~  :��B     ! =�  9U| 9T��i 8��B     - 9Us0  m|�  ��B      0�  �4��  Y� U� 4��  Y� U� 4��  �� �� 50�  6��  � ��    Q  k �  Q��  [��  Q#�O  [��  R#�2  [��  S#�  ^��  \Kl  ^�	   Kdcff k�6    Z��  -�  j�  [��  -"�O  [x ."�  [��  /"�2  [��  0"�4  ^[�  \Kl  7�	  \�U 8�   Kdcff G�6    ME�  B�  ��  IK B#�  I2*  C#�  J�-  E�  J�i  F�  J�Y  G�   +��  ��bB     
       ��  0��  �!X  S� O� 2var �#t�  �� �� `�bB     9U�U  -D�  ��  �bB     	       ���  0��  �"X  �� �� 0J�  �"�  �� �� 0iy  �"�`  1� -� 2var �#t�  l� j� `�bB     9U�U9T�T9Q�Q  -"�  ��  �bB     
       �*�  0��  �X  �� �� 0�' ��  �� �� 2mm �W�  � � `�bB     9U�U9T�T  -�  ��  �bB     
       ���  0��  �"X  6� 2� 0�  �"�  s� o� 0Ԛ  �"?  �� �� 2mm �W�  �� �� `�bB     9U�U9T�T9Q�Q  -U�  ��  �bB     
       �V�  0��  �"X  � � 0�  �"�  Q� M� 0Ԛ  �"?  �� �� 2mm �W�  �� �� `�bB     9U�U9T�T9Q�Q  -3�  �  �bB     
       ���  0��   X  �� �� 0�  � m�  /� +� 2mm �W�  j� h� `�bB     9U�U9T�T  -=�  s�  �bB     
       �f�  0��  s'X  �� �� Olen t'�2  �� �� 0H�  u'?  � 	� 2mm wW�  H� F� `�bB     9U�U9T�T9Q�Q  -Q�  g�  �bB     
       ���  0��  g'X  q� m� Olen h'�  �� �� 0H�  i'?  �� �� 2mm kW�  &� $� `�bB     9U�U9T�T9Q�Q  -��  [�  pbB     
       ���  0��  [ X  O� K� 0�  \ �  �� �� 0Ԛ  ] ?  �� �� 2mm _W�  � � `zbB     9U�U9T�T9Q�Q  -�  O�  `bB     
       �(�  0��  O X  -� )� 0�  P �  j� f� 0Ԛ  Q ?  �� �� 2mm SW�  �� �� `jbB     9U�U9T�T9Q�Q  -Q�  �  bB     A       ���  ,��  +X  U,x 	+�  Tncid 
+�2  Qe�U �   2cff �6  � � =WD  *4bB     5p�  2c �  `� X� .��  �;  � �   -��  ��  �aB     !       �g�  ,��  �X  U,��  �*}  Te�U ��   2cff ��6  J� H� ;�aB            .��  ��;  o� m�   -��  ��  @wB     �       �a�  0��  �X  �� �� 0:�  ��|  �� �� 0%�  ��|  X� N� 0&�  ��`  �� �� .�U ��  L� F� 2cff ��6  �� �� =WD  ��wB     5М  .��  ��;  �� �� :�wB     ]�  K�  9Us  8�wB     ]�  9Us    -Q�  ��  �hB     ~       ���  0�� �$F   � � 0�  �$x  �� �� .I_ �r"  r� d� e�U ��   .��  ��  � � .�-  ��  M� I� 5`�  .�i  ��  �� �� .�b  ��  �� �� :iB     � I�  9T	��F      :iB     � m�  9T	��F     9Q0 `2iB     9U�U9T�T   -��  `�  PiB     o       ���  0��  `X  �� �� 2cff b�6  u� q� .�i  c}c  �� �� 5��  .�-  k�  �  � .��  l�  (� &� .�b  m  M� K� :�iB     � L�  9T	��F      :�iB     � p�  9T	b�F     9Q0 `�iB     9U�U   -��   �  0yB            �/�  0��   ,X  x� p� 0��  ,�?  �� �� 2cff �6  Z� V� (�U �  �L=WD  H0yB     ;xyB     �       .��  	�;  �� �� .ת  
�?  �� �� .ڰ    � � .=�    F� D� >�  ��  .<�    m� i� .��    �� �� >@�  ��  2s $  �� ��  :�yB     : ��  9T	��F      8�yB     : 9U} 9T	��F       :�yB     � �  9T29Q�L 8�yB     ]�  9U|    -��  ��  �wB     6      ���  0��  �*X  !� � 0�  �*�?  �� �� 2cff ��6  �� �� (�U ��  �\=WD  ��wB     ;`xB     �       .��  ��;  &� $� .��  ��?  R� L� .ڰ  �  �� �� :vxB     �  �  9T89Q�\ :�xB     ]�  8�  9U|  :�xB     ]�  P�  9U|  :�xB     ]�  h�  9U|  :�xB     ]�  ��  9U|  8�xB     ]�  9U|    -��  ��  �aB     
       ���  ,��  �$�  U N��  ��  �mB     
      �� 0��  �)X  �� �� 0{ �){  �� �� 2cff ��6  1� -� .�  ��5  k� g� .Q  ��,  �� �� .}W �  �� �� 2sid ��  #� � 2i ��  �� �� >0�  6 .�-  ��  �� �� .��  ��  	� � .�b  �܄  .� ,� :^nB     � �  9T	��F      :mnB     �  9T	W�F     9Q0 `�nB     9U�U9T�T  1�mB            � .ϖ ��  S� Q� .6e  �	  |� x� 8�mB     � 9T	׷F     9Q1  7��  �mB       �mB            �� 4��  �� �� 4��  �� �� 4��  �� ��  8nB     F 9Us   Mq�  =�  � I��  =#X  Ix >#�  I_| ?#	  I�H  @#�  J�  B�6  J��  C  Lsid D�  J�U E�  ]�  zKJ�-  L�  J��  M�  J�b  N܄    Q��  ��  `�B     �      �] R��  � �  � �� R�k � �  �� �� R/� � �  r� f� R�1  � `  � �� R�@  � ?  �� �� Tnn ��  `� R� S�U ��  � �� S�  ��  �� x� =h�  %(�B     >�  < S�H  ��O  �� �� *��  ��  ��1؏B     .       � oah ��  ��<��B     9U| 9T19Qs9R} 9X~   ;АB     +       paw �  ��<�B     9U| 9T09Qs9R} 9X~    8z�B     ] 9U 9Qs 9R}   Q��  ��   �B     V       �b R��  �!�  g� Y� R��  �!�  � � Rx �!�  �� �� R�1  �!`  k� ]� *�U ��  PS�  ��X  � � Sֳ  �BX  �� �� q�B     f�  3 9U�U9T�T9Q�Q9R�R q'�B     f�  J 9T0 r8�B     f�  9R�R3!  QT�  p�  �aB     3       � R�H  p �  i� c� Rsl  q �  �� �� R�J  r �  � � R/�  s   a� Y� S��  u�O  �� �� S�i  v}c  � � <�aB     9U�U9T�T9Q�Q  Q��  �r  paB            �� RAq �,;+  g� c� R��  �,�#  �� �� S��  ��O  �� �� Tcff ��6  � � SQ  ��,  /� -� `�aB     9U�U9T�T  Qx�  ��  PaB            �Z RAq �-;+  _� [� R��  �-r  �� �� S��  ��O  �� �� Tcff ��6  �� �� SQ  ��,  '� %� `daB     9U�U9T�T  Vo�  ��eB     (       �� RAq �';+  Y� S� S��  ��  �� �� Sڰ  �  �� �� D�eB     |  Q��  ��  �`B     V       �� RAq �';+  �� �� R��  �'	  `� \� S��  ��O  �� �� Sڰ  �  �� �� Tcff ��6  � � S�  ��5  �� �� SQ  ��,  $� � `,aB     9T�U9R	 wB     9X0  Q��  ��   wB            �(	 R��  �#�O  s� o� bidx �#�  �� �� Tcff ��6  �� �� S�  ��5  � � Tsid ��  <� 6� Y6wB     ]�   QS�  Jr  �`B     ;       ��	 WI_ J.Y  UW��  K.�#  TS�Y  M�  �� �� S��  Nr  '� %� 5@�  S�* U�  R� J�   Qm�  <�  �`B            �
 WI_ <.Y  UR��  =.r  �� �� S�Y  ?�  �� ��  V�  5�`B     	       �/
 WI_ 5(Y  U Q��  $�  ``B            ��
 WI_ $(Y  UW��  %(	  TS��  '�O  � � Tcff (�6  =� ;� ST )%5  g� e�  ZVJ  �`  �
 ca �`  cb �`  dret �.  dtmp �.   so�  �dB            �/ 4}�  �� �� 6��  �� �� `�dB     9U�U  s]�  �vB     K       �� 4o�  &�  � 4|�  ~� r� A]�  p�  � 4|�  � 	� 4o�  H� F� E��  �vB       ��  �4��  m� k� 4��  m� k� 4��  �� ��   `�vB     9U�T  t~�  PzB     D       �M F��  6��  �� �� 6��  �� �� 6��  � � 6��  ?� ;� 8tzB     � 9T	P�F       sJ�  �~B     Q       �� 4g�  {� u� F[�  F[�  6s�  �� �� 6�  � � @��  �\6��  D� >� C��  �~B     %       � 6��  �� ��  8�~B     R 9T�\  s��  ��B     Z       �
 4�  �� �� 4�  ;� 3� 4%�  �� �� 41�  =� 1� 1��B            { @B�  �P6N�  �� �� <��B     9T�T9Qw   _��  ЃB            41�  �� �� 4%�  (� $� 4�  b� ^� 4�  �� �� _[�  ЃB            6\�  �� �� 8�B     ��  9T�T9Qs 9Rv     s��  ��B     W       �] 4��  4� ,� 4��  �� �� 4��  �  � 1�B            z @��  �`<�B     9Tw   _��  (�B            4��  n� j� 4��  �� �� 4��  �� �� _��  (�B            6��  #� !� j\�  /�B      /�B            n4j�  H� F� 4j�  H� F� 4w�  r� n� _��  9�B            6��  �� �� 8E�B     � 9T�T      sK�  �B     �       � 4Y�  �� �� 4f�  *� $� :(�B     ��  � 9Us� :7�B     | � 9Uv  :Q�B     | � 9Uv  :k�B     | � 9Uv  8��B     | 9Uv   sL�  @�B     �       �� 4^�  |� v� 4v�  �� �� Fk�  u��  A��  p�  | 6��  N� D� 8Q�B     ��  9Uu 9Tt   r��B     ��  9R0  s��  ��B     N       �� 4��  �� �� F��  q��B     ��  � 9Uu 9Tt  8ŕB     ��  9Q09R0  sj�  �B     Y       �� 4|�  � �� 4��  �� y� v��  v��  6��  � � Aj�  p�  � 4��  w� q� 4|�  �� �� 5p�  6��  �  � 6��  '� %� v��  :Q�B     � � 9T	��F      `i�B     9T�T   8$�B     _ 9U	 �F     9Tv   s� p�B     �       �| 4 Z� J� 4 � � 4& �� �� 43 �� u� 6@ Q� K� 6M �� �� 6Z �� �� vg A� ��  N 43 "� � 4& �� �� 4     4 g  _  5��  v@ vM vZ vg ut w} ��  6~ �  �  6� �  �  6�   :�B     �  9T	��F      :��B     � , 9T	W�F     9Q0 `/�B     9U�U9Q�Q9R�R    D��B     ]�  8��B     l 9U} 9Q| ����  x�s  �s  2�y!`  !`  %�y�b  �b  8y\P  \P  yXM  XM  !y�t  �t  :ye  e  �y=T  =T  2]xNe  Ne  32y2n  2n  yHg  Hg  %�x�I  �I  2�yM  M  %�yw  w  %�y�Z  �Z  %�y�[  �[  %�y�k  �k  %�y]>  ]>  %�y@G  @G  %�yKS  KS  %�y�a  �a  %�yd  d  %x�`  �`  2vy�?  �?  4y$i  $i  -yR  R  �yf  f  �z/�  %�  4 zBY  8Y  4 y�s  �s  7y�[  �[  2yCA  CA  5Ey�a  �a  5x@  @  5�ymY  mY  �x?  ?  3(x�  �  3y�D  �D  %�yF>  F>  kyu  u  2y F�   ?1  &  ��  �:  p�B     �%      N )  A"9   ?   �   ��   �  ��    ��  ��   <h ��   �I  ��    �  X�   �   �   �   -   �    	,  �   m�   �   
�   -   �    f  ��   �   �     -   �   �   �    J   �"    �  PH�  Ǟ  J   ֳ  K  pos L    N�  /[  O�   �K P�  (�R Q%  0ڰ  S-   8O�  T  @��  U  H �  ��  <v ��   ��  ��    �  ��  ""  ��  �               	�    	�  �   2  8  
C     i   �  int 	�  �   @	�  �  	�   p  	 	C  �  	#	C  X  	&	C  �  	)	C   �  	,	C  (�  	-	C  0/  	2O  8�  	5O  < �  	�  �  �  	8"]  +  	K
  �  %  	L
  �  	M
  	'  	;  	�  6  s&  
O  �  
V  v  :�   �  L�  x N\   y O\   �  Qh  �  ~   w�  
  y\   �!  y\  �   z\  H  z\   "  |�  �  (j  M} V   5�  V  `�  	O  _| 
  
!  6  ?     2     B  �     �  �  j  �  (Q�     S/   0�  T/  N5  V�  �   W�  H� X�  �1  ZO    �  /  �  \|  �  �  V  �<  �!   �   pmoc�  stibu!  ltuo�  tolp :  ��  �8  5"V  \  �$  �4  S�  x U/   len V6  e� W   �#  Ya  �  �%  {�  �  
�  O  O  �  �    �  �#  ��  �  O  	  O  O  �    �.  �    
1  O  O  �    �8  `��  .   �   �; �  �1  O  �5  �  �+  �   `(  �  (�/  	  0�  �   8*  �  @ w  �  u(  
1  �  �2  (�  �  O    �      I  �3  ;    
(  I   v)  ]5  ;  
P  I       �3  y]  c  O  |  I    �    H7  ��  �  O  �  I  �   �  51  0�  y2  �<   � ��   �(  *
 �P  / �|   $ �
  ( 2$  ��  -4  l  +  �1  	�  $8  �  8  D    ��  O  {"  �/  !  �6  l  \   �O  �  �V  }  ��   )$  �  �   �   c,  +O  C*  6�   +D  CC   :   �$	  xx ��   xy ��  yx ��  yy ��   5  ��  $	  8  �a	  ��  �I   ��  �}   $  �6	  c   �{	  �	  
�	  �    �  ��	  Kl  ��    �  �n	   s  ��	  �"  $�	  �	  �   +
  �� -�	   �W .�	  Kl  /�    %  D;
  uR F�	   �
 G�	   }  I
  V  $��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<
  5�  >\   ��  ?\  �"  A\  �"  B\  i!  C\   %!  E\  (2!  F\  0�  G\  8   I�  �"   sl  ��  u`   5�  v`  ֳ  x\  !  z\  m  {\   v  }  J  �#�  �  �!  �}J  ڰ  -    {3  �}  S0  �}  �/  �}  �1  ��  �1  �G$  Y/  �;
  �*  ��  (�)  �J  0+:  �W$  8<8  �g$  X�*  �}  � �3  �"W  ]  �(  ��  Oe �!$   �-  �y  ڰ  �-    U  �"�  �  �  8�  ah !'$   Oe "�  U1  #;
   ;+  $�  0 i(  �$�    l;  ��t  ah �'$   Oe �4$  y2  �<   {:  �$  (�� �I  h/ �|  p�� ��  x T   � �  �  _  �H  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"  }  8�  �  @`  !}  Hd  "�  P�@  $�	  X�;  )�  h�   +l  ��  ,`  �
  -`  ���  .`  �?!  0`  ��  1`  ��  3`  ��  4`  �ȩ  6�  �ֳ  7H  ��� 8�  �K <�  �ڰ  =-   �^�  >  �U  @;
  �t  B�	  �k  C�   ��L  E8  � "   U  [  1  Xm�  ��  ot   �@  p�	  �e q�  �L  r�  P @  $%�  �    0\�  �-  ^y   ��  _t  �W `�  x a�  �@  b�	   �e d
  0�"  e�  pi"  f�  x� g�  ���  i<  �.a kj  ��  l}  �J  m}  �Mj  o�  ��  q�  ��  r�  �M  t�    Z  u�   _"  w\  (   x\  Ud z�    �L  |0  ( �!  F#    Z!  AY  ��  Ct   T D  �!  El  "  Fl   S  V  �  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  Y  �C  H  0  `)E  K  �"  �e�  �1  g$	   H+  h�   x+  i}  0��  k]   8�)  n#�!  h�'  q%  p��  rB  t�*  y}  x O  l  �  �S  I�  �  �)�  �  �!  H�5  $  ��    7:  ��  s4  ��   b  8H�  !  Jl   m  Kl  A� M�  �� N�  �  P\  
  Q\   ��  R\  (�  S\  0 �  U5   x  t[  x   �$�  �  �!  0'0  ad  )}   �1  *l  &D  +}  2B  ,}  x� -$	     �)=  C  �"  P��  ��  ��   �1  ��  �&  �  �3  �$	  ]7  ��  0�7  ��   @�1  �B  H �  ~�  P6  �  tag �   Kl  �   �6  	�  �  �5  V  
7  i7   �&  9  F9  8%  �*   �,  
�  ./   6
�  b 8
7   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  D  �8  V  ��  �:   4,  �6  $  �/  l9   �2  ��  8  �#  ��  �'  �    �  $  J   �2  �0  6  
A  J   l/  �M  S  �  g  J  g   �  ;)  H��  �#  ��   :  ��  �5  ��  F1  ��  ,8  ��   2*  ��  (�*  �  0`1  �$  8��  �A  @ [  �-  �m  d)  s    �  $  �    9  F#5  $  �$  @J�  �#  L�   y2  M<  W� O  �� P+  �,  Q�   M4  RH  (�;  Su  0�*  T�  8 c/  X!�  �  �-  (q�  �-  sy   Oe t�  ��  u<  � v�   0  �/  )    �  +  �  �   g%  .7  =  
H  �   �.  1T  Z  
o  �  o  �   1	  73  6�  �  
�  �  �   �  �8  :�  �  �  �  �  �   "3  >  $)  Y�  �  �  �  �  �  �  �   �6  _    �  /  �  �  o  �   �3  f;  A  
V  �  �  �   ;0  lb  h  �  �  �  �  �   �&  x��  ah � �   y2  � <  H�8  � �  P�8  � �  X�'  � /  `� � V  h�9  � �  p   �.  ��  "9  H2K  Mj  4�   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :�  T%  �=�  ڰ  ?-    �0  @�  q5  A�  L)  B�  )  C  Ǟ  EK  �  FK  `Ud H�   � X+  J�  W  1  �  �  �      t  }  }  �   �&  &   &  
1  t   �1  *=  C  �  R  H   �6  -^  d  
o  H   w-  1{  �  �  �  �   �;  4�  �  
�  �   =;  8�  �  �  �  H  �   B$  <�  �  �  �  H  �   2  @    �  )  �  H  �  B   7  G5  ;  �  Y  t  �  �  �   q8  Ne  k  �    t     )2  S�  �  �  �  t  �  �  B  �   �  k.  ���  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q �  hZ)  �1  p�#  �R  x'0  �o  �.  ��  ���  ��  �� �)  �`9  �Y  ���  �  �5  ��  �U#  ��  � �/  ��  �  �2  ��  �  �   8S  ��  �d  �g   �W  ��   C  ��  �  �&  0�]   y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��  *  V'v   |   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  ��   �   �  �   j   �  �    a	  �9  �!  !  
"!  j   �    A2  �.!  4!  �  R!  j   �    R!   �   8(  �!  ��  )�    $�  ) !  �-  )"!   )  X!  �!  3  <�!  �� >%�!   ��  ?%j    �!  #  A�!  �!  �U  �,�!  �!  �B  �!"  �� �+   Oe �!"   fP  �,-"  �"  4I  P��"  ֳ  ��   �� ��"  �q ��"  R` �#  �W �=#   P �#i#  (�U  �#�#  0�v  �#�#  8�v  �#�#  @�J  �#$  H 3"  ��  ��!  wq  ��"  �"  �  �"  �!  �   �J  �#  #  
#  �!   �\  �##  )#  �  =#  �!  O   \  �I#  O#  �  c#  �!  c#   O  U  �u#  {#  �  �#  �!  �!  O  O   �O  ��#  �#  }  �#  �!  O  O   �n  ��#  �#  c#  �#  �!  -    ;O  ��#  �#  c#  $  �!  -   O   -k  ��#  �  �(  �]  �  �D  &�  J  W$       g$     �  w$     }$  g  �$  t   H'  �%  ��  8Y%  ��  [�   ��  \�  п  ]�  �U ^�  ��  _�   �  `�  (W�  a  0�  b`  2�  cl  4 ��  e�$  �  p$4%  �$  ��  ���&  ��  �}   ��  �}  *�  �8  ��  �8  	��  �8  
�  �8  .�  ��&  ��  ��&  (��  ��&  <�  ��&  X0�  ��  pY�  �}  xA�  �}  |M�  ��&  ���  ��&  ���  �8  �W�  �8  ���  �  ��  �  ���  ��&  �[�  ��&  ���  ��  ���  ��  ���  ��  ��  ��&  � `  �&     `  �&    	 l  �&      `  �&     `  �&     c�  �:%  �  �#�&  :%  8�  ��&  ��  @'  ��  8   +�  @'  r�   �   �  [�  "'  0�   (!(  ��  *�   �~  +�  U�  -!(  ª  .1(  (��  /A(  �|�  1�  P�  2�  ��  4Q(  ��  5a(  �n�  7�  (��  9q(  0��  A�(  ���  B�  � �  1(     �  A(     F'  Q(     (%  a(     �&  q(     �  �(     �  �(     ��  D�(  S'  ��  P\c)  �  ^�&   ��  `�  �l�  a�  ��  b\  ���  c�  ���  e8   ��  f8  }�  g$	  	�  h�  (��  j�  8@�  k�  @��  l}  H v�  n�(  ��  y%})  �(  ��  H��*  &�  ��   ��  ��  ��  �}  :�  ��  %�  ��   &�  �}  (��  �%  0j�  ��  h(�  ��  ��  �}  � ��*  ���  ��  n�  �}   ��  �}  $�  ��  (��  �}  0��  �p)  8z�  ��  @ �  �*     :�  ��)  ��  �%�*  �)  c�  V  {�+  �   ��  x�  �  Q�  ��  ��  f�  ��  �  	�  
Ƹ  {�  ��  [�  l�  ��  �  p�  i�  ��  ��  ��  �  ��  ��  4�  ��  T�  �  ۳  =�  $�   ��  !e�  "4�  #�  $[�  %��  &��  '��  (7�  )�  *2�  +p�  ,��  -x�  - 
�  ��*  $�  )$,  ,  P�  a�  ,$,  *,  �  C,  -   C,  I,   �&  ,  ;�  1[,  a,  
�,  ,  �  �  �  �   w�  8�,  �,  
�,  ,   *�  ;�,  � =,   �� >O,  �� ?�,   M�  A�,  �,  ��  h!�,  �,  ��  ��  u--  ~-  ��  8V~-  �7  X�,   ��  Y�-  �R Z�-  �� [�-  �� \�-   �� ]�-  (a� ^.  0 -  t�  ��-  �-  
�-  �,   S�  ��-  �-  
�-  �,  �  �   !�  ��-  ��  ��-  �-  
�-  �,  �   e�  
.  .  �  .  �,  �   |�  1).  /.  �  M.  �,  M.  ,  �   �  �  �!`.  f.  ì  ��  �-x.  �.  �  8��.  �7  �S.   ��  ��.  �R ��/  O� �/  �  �?/   y� �l/  (a� ��/  0 ~.  ��  �/  /  
/  S.   ��  �/  %/  
?/  S.  �  }  �   i�  �L/  R/  
l/  S.  �  �  I   p�  &y/  /  
�/  S.  �  I   !�  D�/  �/  �  �/  S.  �   %�  j�/  �/  �  �/  S.  M.  ,  �   ��  �%0  ��  �40   �� �I0  � �^0   �,  40  J   %0  �,  I0  J   :0  k.  ^0  J   O0  ��  ��/  �  � ~0  d0  hG  5�0   num 7}   str 8g   *f  :�0  �_  =�0  key ?�0   Kl  @C   �K  D$�0  �0  �d  H�0  1  �  1  1   �0  �r  K#1  )1    =1  1  1   Uj  (O�1  ��  Q�   ֳ  R�  [M S�  �V  U�0  �F  V1  �B X�1    �0  �@  \ �1  =1  N�  #�1  �1  O  �1  g   :�  )�1  �1  g  �1  �   8�  /�1  �  5'2  V 7O   x 8�   ��  :�1  ��  =$?2  E2  ��  (?z2  I_ A�"   J�  B�  �m Cz2    '2  f�  M�2  �2  g  �2  �  �   �  U�2  �2  
�2  �  g   ��  Y�2  �2  �  3  -   32  �  �2  �2  �   r�  a3  3  �  (3  32  O   ��  e43  :3  O  N3  32  c#   ��  @i�3  4v k �1   �y m �2  v n 3  Ty o (3  hn q �1   S�  r �1  (��  s �3  0��  t �3  8 N3  q�  i�3  �3  =  l  I�  Z4  ��  \l    A�  ^�3  �  �  ��  �B4  ��  �}   �* �4   o�  �N4  4  ��  (��4  N  �}   ��  ��  �  ��  ��  ��  A�  ��    \�  ��4  T4  �  ��4  v�  ��   }�  ��  x �}  y �}   \�  ��4  �4  I�  X�{5  ��  �   o�  ��  )r  ��  (dS  ��  0"�  ��4  81�  ��  @��  ��4  H'�  ��  P �  ��5  5  ��  �!�5  �5  !\  x�*6  ah ��   Q  ��   �"g  ��    #cid ��*  "ת  �4  P"+ �B4  X"�  ��   `"n�  ��  h"��  �  p �I  `U7  Q  W�   �g  X�  �;  Z�  �U  [�  �B ]l   �o  ^l  "Y  `7  (+I  a7  8
  c`  H�!  d`  J�   e`  LH  f`  N�`  hl  P�X  il  RO  k`  T,G  l`  V�t  m`  X �  %7     I  o*6  �g  8�8  ��  ��   )r  �`  dS  �`  
�B  �`  �P  �l  �p  �`  �K  �`  =  �`  me  �`  +^  �`  �]  �`  �u  �8  
h  �`  $^K  �l  &tR  ��   (%?  ��   0 `  8     �]  �17  �S  8?9  ��  A�   )r  B`  dS  C`  
�B  D`  �A  Fl  �n  H`  �n  I`  �W  J`  me  K`  +^  L`  �]  M`  �u  O8  
h  Q`  $�V  Rl  &tR  X�   (%?  Y�   0 �u  [+8  JW  �xX;  ��  zl   =  {`  �<  |l  tB  }l  �k  ~l  �m  `  
�D  �`  gJ  �`  !X  �`  �S  �`  5f  �`  ?X  �`  �a  �`  �_  �`  �a  �`  Gf  �`  �=  �X;   �E  ��  0F  ��  8�A  ��  @F  ��  H�E  �h;  P5D  �l  TH  �l  V#l  �l  X$r  �`  Z_S  �`  \'N  �`  ^?_  �l  `L  �l  b�O  ��  h�O  ��  p~e  �`  x [  �`  z0m  �l  |�M  �l  ~rM  �l  �]  �l  ��g  �l  � 8  h;    	 %  x;     �X  �'9  kE  @�<  �^  ��   zp  ��  dv  �`  �i  �`  �<  ��  �F  ��   �D  ��  (�p  ��  03X  ��  8 �b  ��;  K_  @� =  ��  ��   �J  ��  �<  �l  e  �l  $� �l  dk  �l  ![  �l  L^  �l  �`  � =  yN  �=  ,ma  � =  4�Z  �%  :�q  �%  ;r  �8  <�u  �8  = %  =     %   =     %  0=     	l  �<  �M  (8>  ��  :�   �T  ;l  �P  <l  
�K  =l  B  >l  ^  ?l  �g  @l  /o  Al  %B  Bl  �O  Cl  �<  Dl  �]  El  *w  Fl  dW  Gl   �F  Hl  " e=  J==  |[  Om>  �� Q8   �\  R8  red S8  q  T8   �[  V+>  �?  (��>  `a  �l   �L  ��>  r  ��>  &W  �l  �F  ��>    x  Ik  �y>  >i   J?  tag L�   ��  M�  /� N�  �f  O?   �  2\  Q�>  G   �p?  Tag ��   g  ��  �=  ��  Ja  ��   mn  �|?  .?  �v   ��?  �T  �l   �Y  �l  D  �l  S  �l  E]  �l  ;C  ��  �: ��   �[  ��?  DQ  0@  E]  l   ;C  �  �: �   �i  �?  >M  0.�@  ��  0l   �Z  1�  vv  2�  �r 3�@  =P  4�  �Q  5�@   ^�  6  ( �?  0@  �p  8=@  CE  Y�@  �B  [l   b  \l   Pq  ^�@  �@  �m  x>A  ��  zl   �R  {l  Up  |�@   �=  ~A  �U  �A  �  %   
   %  Sd  !8  �Q  "%  �G  #%  �v  $%  �=  %%  sD  &%  �\  '%  �X  (%  	`N  )�A  
 %  B     �T  +KA  >t  �tB  �>  �B   � �B  !  �8  m  �8  �[  �8  SX  �8   �<  ��B  B  x@  "�B  �  $l   �`  %l  TL  &�3  �o '�B   �B  %  �h  )�B  �Z  <C  �  >l   �f  ?�B   fR  A�B  $ZDC  %j \�B  %�Y ]C   ms   VoC  �  X   �r _C   J  aDC  �t  r!�C  �C  U<  �c  (��C  �B ��   �c  ��  �y ��  �Y  ��  cC  ��   �  �  $ 	\  ��C   L  � D  D  �i  ���H  ah ��   �u  �"?  ��v  ��  �R  �l   o  �p?  (�& �%7  0�Q  �8  �@  �>  �5�  �  �<  �9  ��`  �l  0�a  ��@  8&os2 �x;  hF�  �<  �j  ��  0 M  ��  8w_ ��J  @�>  ��J  H�A  �)K  P^Z  �K  X�f  �K  `KT  �K  h�i  ��   pQ  ��   x&mm ��   �&var ��   �g  ��   ��Y �>A  �Fq �0=  �jQ  ��  �nQ  �tB  �m  oC  ��P  �>  @  l  @B  �K  H�u    P�u  m>  Q�;  �  XzQ  �  `FN  �  hT  �  p!u  �  x&cvt �K  �2i  �H  �)  )�	  ��  +g  ��j  -�  �:>  .�  ��_  0  �S?  3  �E�  4|C  ��W  6O  �XA  8g  �	K  9�  ��c  ?�  �][  @�  ��J  B�  �'<  C�  �	Z  E�   �q  F�  �G  G�  �T  H�  �a  I�   �\  K�  (�u  L�  0o  MyK  8^C  N�  <:W  O4  @_  Q�  H�@  R�  P>  S�  X}?  TO  \m?  UO  `&bdf X�C  h�k  \�  ��Z  ]�  �Pl  h�  �(a  i�  �i m�   ��d n�   � �Q  �  �g  �"�H  �H  �t  x��J  ��  �D   ֳ  �`L  ȩ  ��  �m  ��  �1  ��   x ��  (^�  �  0��  �}  8   �`  <�;  ��  @�C  �}  `� �}  d"f �}  h�I  �  lpp1 ��  ppp2 ��  �Ǟ  �;L  ��y  �;L  �BJ  �HL  �<  ��  bL  ��   Ud ��   (�W  �}  0r�  �}  4&pp3 ��  8&pp4 ��  HO�  ��  X��  ��  `�k  �;
  h �^  �J  �J  �  �J  D  �    ?   �D  *�J  �J  �  K  �H  �  �  �   �b  AK  K  �  )K  �H   SQ  Q6K  <K  
GK  �H   �=  V  TyK  �G   �v  k_  <L  ok   �`  _GK  m>  B  �j  @�;L  ڰ  �-    �0  �l  q5  �`  
0�  �l     �`  org ��  cur ��  " ��   �   ��  (H� ��3  0�>  �l  8 ,L  ��K  @\  �'UL  [L  �r  �d  � mL  sL  �a  
�  @E�L  ^�  G   �k H�  ��  I�  /� J�  T�  K8  z�  L�   ��  M�  (�f  O?  0Vu  P�  8 �  RxL  !��  UXM  ��  W�   �  X�  /� Z�  c�  [XM  "= \XM   l  hM    � ��  ^M  Y�  (a�M  ��  d�   �  e�  c�  g�3  ��  h�3  "�  j�   �  k�  $ ��  mtM  -�  rN  ��  y�   ��  z4   8�  |�M  9�  �EN  z  ��   �  ��  �  ��   �  �N  �  �lN  ّ  �lN    EN  ��  �QN  J�   ��N  ��  ��   ��  ��N  �  �l  ��  ��  ��  ��N   N  rN  ��  �~N  ��  �!�N  �N  U�  �RAQ  �-  Ty   ^�  U  ڰ  V-   ��  W�  �!  X�   �  Y�  ${3  [8  (S0  \8  )G�  ]8  *��  _�  ,�_  a  0�  c�L  8Y�  d�L  x�  e�L  �T ghM  ��  h�M  ��  j�L  89�  k�L  x��  l�L  �x�  m�L  �*�  o�  81�  r4  @��  u�  H�y v4  Pv�  w�  Xx�  x�  `Ω  z1W  h��  {�  0��  |>W  89�  ~$W  8�  �q0  XQ  ��3  `��  ��  h��  �NW  p:�  ��  x%�  ��  ���  ��	  ���  ��N  �ת  �TW  � ��  0��Q  ��  �   ��  �  �  ��N  ��  ��  3�  ��  L�  ��  ��  ��   BV ��K  ( 4�  �AQ  !a�  H��S  ��  ��   ��  ��  ��  ��  п  ��  �U ��  ��  ��  W�  �  �  ��   �  ��  (�  ��  0��  �}  8[@ �}  <}�  �$	  @�  �  `��  ��  h	�  ��  p��  ��  �j�  ��  ��  �\  �	�  ��  ���  ��  ��  ��  ���  ��  ���  ��  �ɼ  ��  �=�  ��  �6�  ��  �!�  ��  �"�  ��  �6�  ��  �"��  ��   "��  ��  "�  ��  "$�  ��  "n�  ��   "��  ��  ("&�  ��  0"��  �l  4"�  �l  6"ɰ  ��  8"5�  ��  @ Z�  ��Q  [�  �$	T  T  ��  �/�T  �  1�S   �  2�V  HE�  5�Q   3�  6�  P&NDV 7�  X��  A�  `!�  B�  h��  C�  p��  D�  tx�  F�L  x)�  G4  �.�  JO  � !׬  ��vV  *�  �8   ��  �8  ��  �8  �  �8  .�  �vV  ��  ��V  x��  �vV  �"�  ��V  80�  �  �Y�  \  �A�  \  �M�  \  ���  \  ���  8  �W�  8  ���  	�V  �[�  
�V   ��    ��  �  ���  }  ���  }  ���  �  ���  �  ��  �  ���  \  ���  \  �y�  �  ���  �S  � \  �V     \  �V    	 \  �V     ��  �T  7�   $W  ��  8   �  �  Kl  "�  ��  #�  M�  &�  ��  '�  �  (8   ׵  *�V  ��  LT  �S  NW    � %  4  ��  `,�W  ah .�   m /�  X ��  1�W  ZW  !��  H<�W  ah >�   "�� @  0"��  A  1"A� C�  8"�� D�  @ ��  F�W  �W  xX  h *IX  ah  ,:$   �q   .�  8�'   /  <iO   0IX  @��   1B  ` }  YX     Y   3eX  �W  ��   ?-wX  }X  �  ` �Y  *�   ��   O�   ��  z�   ��  ��  ��  6�   �}   ��   �}  $�K  �4  (h�   �4  0ڰ   �-   8��  ��Y  @ ��    XOY  ��  [hY   �q  `yY  add  c�Y  U1  iyY   �  hY  kX  }  -    OY  
yY  kX   nY  �  �Y  kX  }  �  �   Y  H�   kY  �Y  ��   �"�Y  �Y  ;�  � �)Z  O�   ��   Ǟ   ��  ��   ��  �U  ��  ڰ   �-    ��  �N^  ( ��   �"5Z  ;Z  Q�   �pZ  �k  ��   ��   ��  b  �J[   K�   �"�Z  pZ  �Z  �  0 �[  �   g   ��   \  b  �[  ��   \  �   �  ֳ   8  C�   �   ��   	�  $��   �  ( '��  V   �J[  ��   }�  ��  ��  �  ��   I�   �[  '"�  V   ��[  :�   G�  ��  Z�  z�  !�  ��  d�   �  \�  	��  
��  Ѻ   ��   �V[  '��  V   �\  ��   ��  F�  r�  ػ  ��  ��  _�  j�  ��  	 e�   ��[  [�   �*\  0\  
@\  t  �   1�   �Z  @\  ��  h u]  ��  x1]   �q  ~B]  �Y  �B]  �L  �B]  ;  �W]   �>  �q]  (nD  ��]  0�M  ��]  8�:  ��]  @�[  ��]  H�l  �^  P`  �H^  X�9  �H^  ` 
1]  �Y  �  �  -    ]  
B]  �Y   7]  �  W]  �Y   H]  �  q]  �Y  }   ]]  �  �]  �Y  �  �  ?     w]  }  �]  �Y  }  �]   `  �]  }  �]  �Y  }  �  }   �]  
�]  �Y  )Z   �]  
^  �Y  )Z  �  ^   }  �]  �  H^  �Y  |Z  �  �  ?   %^  :�   �R\  N^  "�   ��Y  ��   �z^  ;�  p 4w_  ڰ   6-    ��   7t  ȩ   8�W  ��   9�  Ǟ   :M.   �   ;M.  (��   =�_  0��   >�_  8�C   @�  @�  A�  H�;   C�  P.�   D  X��  E  Y8�   F  Z��   H  [�   I  \��  K�_  ` ��   ��_  ��  ��_   �q  ��_   
�_  �_  �      m^  �_  
�_  �_   �_  ��   �w_  \  ��   b `  Ǟ   d�   ��   e�  O�   f�   Q�   h�_  (�   l:`  @`  �  ^`  D  �  4  ?   ;�   rk`  q`  
�`  D  4  �   w�  � w�b  �I  ym^   ��  {�b  p&top  |�  ���  ~�b   �y   �b  �a�   �}  ��   �}  ��   ��b  �&cff  ��N  ��   ��S   ��   ��b  (��   ��_  0׹   �  8��   �}  <P�   ��  @"�   ��  Dc�   �}  H��   �}  LT�   �4  P0�  �4  X�o  �4  `�   ��  h;:   ��  lzd  �  p��   �&-`  x��   �&^`  �Q   ��3  ���   �}  �Z�   �4  ���   ��1  �}�   �$	  �	�   ��  �E�   ��(  �f�   �@'  ���   ��  � �  �b    0  `  �b      `  �  �b     �	  ��   ��`  �   �#�b  �b  ��  � <d  ڰ   >-    ��   ?t  ȩ   @�  ��   A�  Ǟ   BM.   �   CM.  (��   E\  0��   F\  8�C   H�  @�  I�  P�;   K�  `˹   L�e  ���  M  �8�   N  ���   P  �b�   R�   ��   S�   ���  Uye  � ^�   �d  d  �  /d  �b  }   G�   �<d  Bd  
\d  �b  \  \  8   r�   �id  od  �  �d  �b  \  \   h�   ��d  �d  �  �d  �b    �   �id  ��   ��d  �d  
�d  �b   ؽ  @ �Te  ��  �se   �q  ��d  VY  �$d  c  �$/d  f  �$\d   2  �$�d  (�J  �$�d  0�  �$�d  8 
se  �b  t  H  �     Te  ��   ��d  ye  ��  V   ��e  >�    �  /�  i�   v�   ��e  f�   W�b  ��   v
f  O�   x�   Ǟ   y�  ��   z�   ��   |�e  ��   |$f  �e  �   /7f  =f  ��  � ��g  �I  ��e   ��  ��h  �&top  �@'  ���  ��h  ��y   �f  x
Q   ��3  �
�   ��  �
�o  �4  �
��   �}  �
��   �}  �
+  �4  �
��   �4  �
��   ��1  �
}�   �$	  �
	�   ��  �
a�   �}  �
�   �}  �
�   ��b  �
E�   ��(  `;:   ��  h��   �h  p��  ��h  xf�   �@'  ���   ��  �zd  �  ���   ��	  � �    �h  ��  �vh   �q  ��h  ;U  ��h  �"  ��h   õ   �%h  +h  �  ?h  *f  �   �  vh  *f  t  H  �  4  �(    �  h   ?h  
�h  *f   |h  �  �h  *f  �  �   �h  �  �h  �h  �  �   �b  �h  '�   ��g  �h  �  �h    � 
f  i     ��   �=f  D�   � i  ��  � T(j  ڰ   V-    ��   WD  ȩ   X�W  ��   Y�  Ǟ   ZM.   �   [M.  (��   ]\  0��   ^\  8�C   `�  @�  a�  P�;   c�  `.�   e  ���  f  �8�   g  ���   i  �b�   k�   ��   l�   ���  n�k  � 9�   �5j  ;j  �  Oj  Oj  }   i  ��   �bj  hj  
�j  Oj  \  \  8   �   ��j  �j  �  �j  Oj  \  \   ��   ��j  >�   ��j  �j  
�j  Oj   ש   ��j  �j  �  �j  Oj   ��  @ �zk  ��  �k   �q  �j  VY  
%(j  c  %Uj  f  %�j   2  %�j  (�J  %�j  0�  %�j  8 
�k  Oj  D  �W  �W     zk  �   �j  ^�   ��k  Ǟ   ��   ��   ��  O�   ��   ��   ��k  ��  � ��m  �I  �i   cff  ��N  ���  ��b  �&top  ��  h��  ��m  p�y   ��m  a�   �}  �   �}  �   ��b  ��   �\  ���   �\  �0�   �  �׹   �  ���   �}  �f�   ��m  �P�   ��  �"�   ��  �c�   �}  ���   �}  �T�   �4  �0�  �4  ��o  �4  ��   ��  �;:   ��  �zd  �  ���   ��S  ���   �&-`  ���   �&^`  � �k  �m     �k  �  �m     �   ��k  +�   �n  ��  �Cn   �*   �bn  �"  ��h   
=n  =n  D  �W  �W    �  -`  ^`   �m  n  �  bn  =n  �W  �   In  �   ��m  hn  �   �#�n  �n  ��  ( �n  ڰ   -    ^�   wo    {5  F�   �o  w�    �     ӫ   �o  ��  �9o   �q  �Jo  �i  �_o   �  9o  zn  -   �  �   o  
Jo  zn   ?o  �  _o  zn   Po  ��   ��n  eo  ��   �#�o  �o  ��  }  �o  g  �  �    �o  R�   -.�o  p  ��    /p  f�   1!"   ]J  2!"  ��   3!"  V  4!"   �o  ��  X A�p  8�   D!�p   ��   E!�p  �   F!�p  ��   G!�p  կ   J�p   *�   O�p  (��   Rq  0��   W.q  8�   [�o  @��   ^!4q  H�   `":q  P �Y  [^  �e  �h  
�p  �  �  l   �p  O  �p  O   �p  
q  �h  �      �p  
.q  t  �&  �S   q  ro  un  4�   bMq  p  O�  �!E�q  ah !G`^   ^�  !H  �F�  !J�  ���  !K�  �z�  !M�  ��  !O�  �cid !Q�*  ���  !R}  � ��  !TSq  g�  �"�q  ��  "!�q   ��  ""}  � k�  "$�q  (�  #8!r  r  ��  `#]Cr  ah #_�   ��  #`  X ��  #C&Or  Ur  !��  H#e�r  ah #g�   "�� #i  0"��  #j  1"A� #l�  8"�� #m�  @ V  $��t  ]�   ?  ��  y�  �  ��  �  -�  ��  :�  	'  
3�  ��  @�  ��  ��  o�  ��  ��  n�  )�  4�   h�  !	  "~�  #J�  $A�  %�  &a�  '��  (��  0��  1��  @��  A�  Q��  Rz�  S$�  T��  U��  V��  W��  X��  `�  a��  b[�  c"�  p�  ���  �#�  ���  ���  �z�  ���  �	�  ���  ���  �'�  ���  ���  �J�  �K�  �#�  ��  ���  � �W�  ��  ���  ��  ���  ���  ���  ���  �T�  ���  ���  ���  ���  �1�  ���  �A�  �7�  ���  ���  ���  �r�  �i  �+�  �D�  ��  �o�  �\�  �Q�  � M\  �t    4 �t  (l�  t�t  	��F     �)  %�  �d  &)w$  ��  &,Au  0u  `p  &,\u  g &.$u    ܨ  '!hu  nu  �  �u  t  NW   *�  '%�u  �u  �  �u  t  TW   ]�  ')�u  �u  }  �u  t   ��  ',�u  �u  �  �u  t  �u   �&  ��  '0v  v  �  *v  t  �+  �  �   �   ��  '7;v  *v  �  ('7�v  ��  '9\u   Ъ  ':�u  �  ';�u  ݱ  '<�u  ��  '=�u    n�  (�v  �v  �  �v  t  �v  �v  ^   g  ��  ($�v  �v  �  �v  t  �v     3�  ('�v  �v  �  w  t  �  4   Y�  (+(w  w  ��  (+]w  �  (-/�v   ��  (./�v  N�  (//�v   �<  )iw  ow  �  �w  J  g  �     s=  )$�w  �w  �  �w  J  g  �    �  ))�w  �w  #P  ))�w  R  )+]w   bD ),�w   )@�  A*<u  	��F     )��  ^&6v  	��F     )
�  �##w  	P�F     )�  ��w  	@�F     �  Yx     Ix  )�  �#Yx  	��F     *u  �	 �F     +��  ��  ��B     
       ��x  ,ϖ �#J  S O ,�  �#g  � � -��B     �  .U	��F     .T�T  +J�  ��  0�B     
       �Ly  /��  �+�5  U/x �+�  T0cid �+4  Q1�U ��    +~�  ��   �B            ��y  /��  ��5  U/��  ��v  T1�U ��    + �  p�  ��B     .       �z  /��  p�5  U/:�  q�v  T/%�  r�v  Q/&�  s^  R2cid u�*  � �  +s�  V�  ��B            �Fz  /��  V+t  U/��  W+TW  T +��  M�  ��B     O       ��z  /��  M*t  U/�  N*NW  T +�  5g  p�B            ��z  /��  5&�5  U3�Y  7g  � �  4��  �z  5��  !�z  67^�      �q  8? 9�  |  9��  9"�z  9^�  :"  9ڰ  ;"-   9g  <"@q  :�U >�  :��  ?�  :�  ?�  ::�  ?$�  ;cur @�  :��  @�  :&D  A�  :2B  A�  <�  �<]�  Z<cs �=�{  :_| o|  :f�  r�  :��  s�  ;p t�  6:��  y�    6;tmp ��    8  |  >  	 ?�  `�B            �E|  @K J  U AK�  ��  ��B     x       ��|  @ϖ �J  UBK �YX  / - (��  �O  �t C1 �  n}  5^�  !  5%�  !t  5�  !}  5�[   !}  5\  !!�  7��  #�5  7�U $�  7g  %@q  7�  &q0  D�  ���B     6Ecid e�*  7�  f(%  67��  ~�  7�V �     F��  �`�B     �      ��  ,%�  �t  Z R 3��  ��5  � � 3ڰ  �-   "   2cid ��*  K E 3�  �(%  � � G��B     w       �~  2n �}   � G��B     D       m~  3�R �B4  O M H��B      �  X~  .U}  I��B      �  .U}   I��B      �  .U}   H�B      �  �~  .U}  H)�B      �  �~  .U}  HC�B      �  �~  .U}  H]�B      �  �~  .U}  Hw�B      �  �~  .U}  H��B      �    .U}  H��B      �  *  .U}  H��B      �  B  .U}  H��B      �  Z  .U}  H�B      �  r  .U}  I-�B      �  .U}   +��  ��  @�B     4       �-�  ,ֳ  �&H  x r Jreq �&�  � � 3�� ��,    HL�B     �  �  .T�T HT�B     ��  �  Kl�  s  Lp�B     .R0.X0  +,�  ��  ��B     Y       �'�  ,��  �H  , & 3ֳ  �	r  ~ x 3�U ��  � � 3�� ��,  	  G��B     9       �  )0� �,  �h3��  ��5  C ? 3��  �p)  ~ z 3��  ��&  � � L��B     .Q�h  I��B     ��  Kl�  s   M��  p[�  9��  pH  :ֳ  r	r  6:�� w�,    8��  `�,  ��  9ֳ  `)	r  :��  b�5  :�  cq0  :ϖ dJ   N�  :�  @�B     M       �g�  ,�  : �  ( " 3��  <�5  z t 3�  =q0  � � OV�B     .       3ϖ EJ  � � Gs�B            J�  3�� L�,     In�B     �  .T	P�F        F��  3��B            ���  /�  3 �  U C��  ��  ?�  5��  ��5  5�  �}  7��  �q  7��  �z  7ڰ  -   7�U �  En }  Ecid �*  7�  	�  7�  
�  P�  �67��  Zp)    C��  ��  )�  5Kl  � �  5{<  � �  5�  � �  5��  � �5  7^�  �  7�U ��  7_| �)�  Ep ��  7��  ��  Ed ��  7-�  ��  Eval �8  7�  �  7�q �  P�  �67h�  ��  7ֳ  ��    8  9�    � 4[�  �b�  5��  �!b�  7��  ��z   �q  4�  ���  5��  �!b�  5��  �!�5   C" �  ��  5��  �5  Ecid �*  7ڰ  -   7^�    7�U �  En }  7�R 	B4  7w�  
�  7�f  ?  7g  @q  P�  rPWD  v67��  p)  7��  }  7/� �  7��  �  7{<  �  Ep �  =��  7�N  "�   =��  Elen [�   6Elen g�     C�  ��  r�  5��  � �5  5��  � b�  5Ǟ  � �  5ֳ  � �  7��  ��z  6Ecur ��  7��  ��  67��  ��  6Elen ��  67��  �pZ  67}W ��  6En ��         ?^�  X��B            ���  @��  X!�5  U@��  Y!�z  T ?��  ?p�B     I       �%�  Q��  ?(�5  : 4 Q��  @(�z  � � B��  Bp)  � � L��B     .U�T.T0  F]�  ���B     
      �j�  ,��  � �5  	 	 ,��  � �z  }	 y	 2cid ��*  �	 �	 3ڰ  �-   -
 )
 3^�  �  g
 c
 )�U ��  �L3��  ��  �
 �
 P�  5GP�B     �       X�  Rn }  �
 �
 G��B     8       &�  B��  )p)     Ij�B     &�  .Uv .T
P.Q0.Rs .X0.Y�L  L	�B     .U�T  F��  �P�B     �      ��  ,��  �'�5  Y Q ,��  �'�z  � � 3��  �p)  !  3ah �t  [ S )�S  ��  ��3��  ��  � � S�  ���B     T��  3�3  �/�  � � 3�  ��    3�Y  �}  R P U��B     q�  .Uv .T6.Qw .R3 H��B     2�  ��  .U
�.T~  H��B     2�  ��  .T~  H��B     2�  ��  .T~  H�B     2�  ؉  .T~  H�B     2�  ��  .T~  H/�B     2�  �  .T~  I��B     ?�  .Us�   �  /�     $	  8W�  G�  ��  9��  G%�5  9��  H%b�  9��  I%|Z  :�U K�  :��  L�z  :��  M�  :��  N�   ;cid O�*  <�  �6:��  qp)    8��  +�  ��  9�k +4  9	�  ,8  :�Y  .�  ;p /�   A��  Q�  ��B     �      �H�  Q��  Q&�  } u Q��  R&H  � � Qx S&�  � � Q�1  T&B  = 1 Bȩ  VCr  � � B�U W�  : & (LM Xi  ��hB��  Y�5   
 Bn�  Z  R D B��  [  � � Bg  ]@q  z r (}�  ^$	  ��gB	�  _�  � � B~�  `  a U P�  	V`�  ��  B�L  �0  � � W��B     L�  W��B     L�   V`�  я  (�'  ��  ��gB�e �H�    V �  ��  Rn �}  N L Rcur �M.  } y Rvec ��  � � BA� ��  @ < B�� ��  ~ z XS�  x�B      0�  �m�  Yn�  Zd�  � � T0�  [x�  � � [��  ; 7   \S�  ��B      ��B            �ˍ  Yn�  Yd�  O��B            [x�  z v [��  � �   \S�  ��B      ��B            � 1�  Yn�  Zd�  � � O��B            [x�  #  [��  f b   ]S�  ��B      ��B            � Yn�  Zd�  � � O��B            [x�  � � [��       XS�  ��B      ��  � �  Zn�  L J Zd�  s q T��  [x�  � � [��  � �   XS�  ��B      б  � @�  Zn�    Zd�  C A Tб  [x�  l h [��  � �   W2�B     L�  WG�B     L�  H��B     Y�  y�  .U| .T��g H�B     f�  ��  .U| .T} .Q~  H�B     s�  ��  .U| .T��g I5�B     �  .Us0  U]�B     �  .U��h.T| .Q} .Rs .X0.Y0 H��B     N�  !�  .U��h.T~  U�B     6�  .U��h L	�B     .U��h  
  +��  -�  ��B            �S�  ,LM -*f  � � ,x .�  � { 3��  0�5  � � 2cid 1�*  f \ 2p 2�  � � 39�  3�  � � 3^�  4  � � )�U 5�  ��l39� 6�  T > 3ڰ  7-   B : 3��  8�  � � 3g  9@q  � � 3�  ;      2inc >#�!  �  �  S�  �k�B     V�  x�  ))�  Ka	  ��u^��  �B      0�  T �  Zڊ  �  �  ZΊ  1! -! T0�  [�  w! q! [�  �! �!   U��B     �  .T��k�.Q��u Uq�B     3�  .T��u H{�B     ��  [�  .Uw .T��k.Q��l I��B     ��  .U} .Q��k  V��  ��  3�  l�   " �! 3� m�  :" 6" 3� m�  v" r" ^��   �B      �  v�  Zڊ  �" �" ZΊ  �" �" T�  [�  1# +# [�  �# |#   _��  [�B       [�B     1       w�  Zڊ  �# �# ZΊ  7$ 3$ O[�B     1       [�  }$ w$ [�  �$ �$   ^��  ��B       �  yԓ  Zڊ  0% .% ZΊ  W% U% T �  [�  �% % [�  �% �%   H��B     ��  �  .U��k H�B     ��  �  .U��k.T
s 1$���� H��B     ��  0�  .U��k H�B     ��  X�  .Uw .T��k.Q��l HN�B     ʦ  ��  .U��k.Q} .R��k Ig�B     ��  .U��k  V`�  ˕  3��  �p)  & & 3�  �B4  ^& Z& 3	[  ��  �& �& G��B     �       ��  )�  ��b  ��u)��  �1W  ��lU��B     1�  .U��u.Tv .Q1 U��B     L�  .Ts .Q��l U�B     o�  .U��u.T��k.Qs  LF�B     .U��u.T��k.Qs   U^�B     ��  .U} .T��k.Q
� L��B     .Uv .T��k  G��B     �       7�  )�e �"�   ��uW��B     L�  W��B     L�  W��B     L�  L �B     .T��k�.Q0.R��u  Iw�B      �  .Uw .T}   8VJ  �B  ��  `a �B  `b �B  ;ret �(  ;tmp �(   a[�   �B     <       ���  Yl�  [x�  �& �& [��  ' ' [��  Q' M' I�B     �  .T	P�F       b'�  ��B     9       ���  Z4�  �' �' [@�  �' �' c'�  ��B     "       Z4�  [( U( O��B     "       d@�  cL�  ��B     "       [M�  �( �( I��B     ��  Kl�  s      b�|   �B     �      ��  Z�|  �( �( Z�|  �) �) Z�|  �+ �+ Z�|  G, ?, Z�|  �, �, [�|  ?- - [�|   / / [
}  �/ }/ [}  0 �/ e�|  ��  ��  Z�|  [0 O0 Z�|  �0 �0 Z�|  G1 A1 Z�|  �1 �1 Z�|  2 �1 T��  d�|  [�|  ~3 r3 d
}  d}  f$}  X��  ��B       �  NQ�  Z��  4 4 Z��  �4 �4 T �  g��  ��{[͂  6 6 [ڂ  �6 �6 g�  ��{[�  �7 �7 [��  �7 �7 [�  �9 �9 [�  �9 �9 h&�  '�B     Xh�  ��B      ��  ~�  Z��  a: A: Zv�  �; �;  X�z  ��B      г  �  Z0{  �; �; Z${  6< &< Z{  �< �< Z{  �= �= Tг  [<{  t> \> [H{  ~? n? [T{  L@ 4@ [`{  SA GA [l{  �A �A [x{  nB \B [�{  ?C 3C [�{  �C �C f�{  h�{  E�B     h�{  �B     e�{  ��  )�  g�{  ��}[�{  FD <D [�{  �D �D [�{  _E OE e�{  д  �  [�{  F F Hz�B     צ  Ț  .Uv  H��B     �  �  .Uv .T| .Q  I�B     �  .U��}.T	�  "
Y.Q9  I`�B     צ  .Uv   i�{  ��B             n�  [�{  NF LF I�B     ��  .Us .T0.Q:  U��B     ��  .U~ .T0.Q0.R��{ H��B     צ  ��  .Uv  H��B     ��  ɛ  .Uv .TO H�B     ��  �  .Uv  WE�B     ��  H&�B     ��  �  .Uv .T��{ H@�B     	�  3�  .Uv .Ts .Q~� U��B     G�  .U~  U��B     [�  .U~  U��B     o�  .U~  U��B     ��  .U~  U��B     ��  .U~  U��B     ��  .U~  H'�B     �  ʜ  .Uv .T~� I3�B     ��  .Uv .Tw    \9�  '�B      '�B     )       ���  ZG�  sF qF O'�B     )       [T�  �F �F ]�z  '�B      '�B     )       �Z�z  �F �F i�z  2�B            ��  [�z  �F �F IF�B     �  .T~�  LP�B     .U~     X��  v�B        �  ݟ  Z�  	G G Z�  0G .G Z؅  eG SG Z˅  "H  H T �  [��  YH EH j�  ��  [�  CI 'I [�  yJ iJ j'�  0�  [(�  HK DK e5�  ��  ��  [6�  �K ~K jC�   �  [D�  *L L jQ�  ��  [R�  �L �L e_�   �  ��  [`�  NM HM k5�  ��B      `�  �(Z^�  �M �M ZR�  `N PN ZF�  O O T`�  [j�  �O �O [v�  �O �O [��  �P �P g��  ��}[��  Q Q h��  �B     e��  и  Z�  [��  �Q �Q  U�B     ��  .U~ .T .Q��}.R0.X0 L��B     .U} .T~     Ii�B     #�  .Us     U��B     ɟ  .U~  L��B     .U~      X?�  ��B        �  0=�  Zx�  �Q �Q Zk�  [R YR Z^�  �R ~R ZQ�  �R �R T �  [��  �R �R [��  sS kS g��  ��}[��  �S �S [��  U U [ă  U kU [σ  YV MV [܃  �V �V [�  <W *W [��  
X �W f�  e�  ��  '�  [�  �X �X [�  !Y Y H��B     צ  �  .Us  H��B     �  �  .Us .T��} I��B     צ  .Us   I�B     ��  .Us    e/�  ��  X�  [0�  {Y uY  X��  ��B      �  ���  Z��  �Y �Y T�  [��  7Z 1Z [��  �Z �Z [ʄ  [ [ gׄ  ��}[�  ~[ j[ [�  g\ _\ [��  �\ �\ [	�  �] x] [�  �^ �^ h#�  |�B     h,�  ��B     e5�  0�  c�  [6�  '_ _ [C�  �_ �_ [P�  �` �` []�  5a )a [j�  �a �a [w�  �a �a e��  ��  ˢ  [��  :b 4b I��B     &�  .Uw .T8.Q��{�����.R��{�����.X| .Y��}  X��  �B       ��  8!�  Zڊ  �b �b ZΊ  �b �b T��  [�  c c [�  `c Xc   i��  C�B            H�  [��  �c �c  i��  ��B            ��  [��  �c �c L��B     .Q
�  H��B     ��  ��  .U  H��B     ��  ��  .U  HA�B     ��  ȣ  .U  H��B     &�  �  .Uw .T8.Q0.R��{�����.X0.Y��} H��B     ��  .�  .Uw .T��{.Q��} H�B     ��  F�  .U  I4�B     �  .U .Q��{  H��B     &�  ��  .Uw .T@.Q0.X0.Y��} H*�B      �  ��  .Uw  HO�B      �  Ĥ  .Uw  Hq�B      �  ݤ  .Uw  I��B      �  .Uw .Ts    Hr�B     ��  !�  .U��{.TP.Q��{ H��B     ��  B�  .U��{.Q��{ W��B     /�    j5}  �  [6}  Zd Pd [C}  �d �d jP}  P�  [Q}  ne `e [^}  f f     Hh�B     ��  ��  .Us .T0 H��B     <�  ץ  .T	�F      I�B     <�  .T	P�F       lF>  F>  km�s  �s  *�lR  R  �l$i  $i  -m�I  �I  *�l\P  \P  l�[  �[  2l�s  �s  7lCA  CA  +El�a  �a  +m@  @  +�lmY  mY  �m�`  �`  *vnBY  8Y  / lM  M  ,�l@G  @G  ,�l�a  �a  ,�l�^  �^  ,�l�Z  �Z  ,�l�D  �D  ,�mn  n  -m$  $  ..l]>  ]>  ,�l!`  !`  ,�mNe  Ne  -2l)p  )p  ,vl�?  �?  4 �t   �7  &  ^ �:  �B     �5      o ,  i   	�@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ��  
�5  ;  �s  
�H  �  s&  
G   �  
N   )  A"u  {  �   ��  �  �U    ��  ��  <h ��  �I  �   �  X�  �  U   �  i  -    �   m�  �    i  U    f  �    U   5  i  -   -   U    J   �"A  G  �  PH�  Ǟ  JD   ֳ  K@   pos L@     N  /[  O   �K P  (�R QQ  0ڰ  Si  8O�  TD  @��  UD  H �  �  <v �-   ��  �U    �  ��  ""  �   &  @   D  5  @   D  @    J  �  �   ^  d  o  5   v  :-   �  L�  x No   y Oo   �  Q{  	�  ~   w�  
  yo   �!  yo  �   zo  H  zo   "  |�  N`  N   �G  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} N    5�  N   `�  	G   _| 
D  
!  H  ?   J  2   J  B  U     �  G  	�  �  (Q;     S5   0�  T5  N5  V;  �   W�   H� XA  �1  ZG     �  5  �  \�  �  �  N   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  �Z  �8  5"�  �  �$  �4  S�  x U5   len VH  e� WJ   �#  Y�  	�  �%  {    3  G   G   3  U      �#  �F  L  G   e  G   G   U    �.  �r  x  �  G   G   U    �8  `�  .      �;    �1  G   �5    �+     `(  9  (�/  e  0�  U   8*  �  @ �  &  u(  
�  	'  �2  (F  L  G   `  U   `   �  �3  ;s  y  �  �   v)  ]�  �  �  �  D  @    �3  y�  �  G   �  �  @   U    H7  ��  �  G   �  �  �   4  51  0�h  y2  ��   � �9   ��  *
 ��  / ��   $ �f  ( 2$  �  -4  lJ  +  ��  �  $8  �J  	�  �    ��   	�  {"  �5  !  �H  \   �G   �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U   +D  C4    :   �{	  xx �	   xy �	  yx �	  yy �	   5  �8	  	{	  8  ��	  ��  ��   ��  ��   $  ��	  c   ��	  �	  �	  U    �  �
  Kl  �U    �  ��	   s  ��	  �"  $(
  .
  �   +g
  �� -
   �W .
  Kl  /U    %  D�
  uR F
   �
 G
   }  Ig
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<a  5�  >o   ��  ?o  �"  Ao  �"  Bo  i!  Co   %!  Eo  (2!  Fo  0�  Go  8   I�  �"   s�  ��  u�   5�  v�  ֳ  xo  !  zo  m  {o   v  }n  J  �#�  �  �!  �}�  ڰ  i   {3  ��  S0  ��  �/  ��  �1  ��  �1  ��$  Y/  ��
  �*  �G  (�)  ��  0+:  ��$  8<8  ��$  X�*  ��  � �3  �"�  �  �(  ��  Oe ��$   �-  ��  ڰ  �i   U  �"�     �  8G  ah !�$   Oe "    U1  #�
   ;+  $$  0 i(  �$T  Z  l;  ���  ah ��$   Oe ��$  y2  ��   {:  �{  (�� ��  h/ ��  p�� �&  x T   � �  �  _  ��  �!  �   �  �  �  �    �  �  �   �U !  (�  !  03"  �  8�  '  @`  !�  Hd  "-  P�@  $
  X�;  )�  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7�  ��� 8V  �K <�  �ڰ  =i  �^�  >5  �U  @�
  �t  B
  �k  CU   ��L  E�  � "   �  �  1  Xm�  ��  o�   �@  p
  �e q  �L  r@  P @  $%      0\V  �-  ^�   ��  _�  �W `�  x a�  �@  b
   �e da  0�"  e	  pi"  f	  x� g�  ���  i�  �.a k�  ��  l�  �J  m�  �Mj  oG  ��  q�  ��  r%  �M  tU    Z  u-   _"  wo  (   xo  Ud zU    �L  |�  ( �!  F#c  i  Z!  A�  ��  C�   T Du  �!  E�  "  F�   S  N   �u  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  �C  Hi  0  `)�  �  �"  �e!  �1  g{	   H+  h�   x+  i�  0��  k�   8�)  n#2"  h�'  q�  p��  rO  t�*  y�  x �  �  V  �S  I�  �  �)M  S  �!  H��  $  �U    7:  �;  s4  �   b  8H  !  J�   m  K�  A� M	  �� N	  �  Po  
  Qo   ��  Ro  (�  So  0 �  U�   x  t�  x   �$2  8  �!  0'�  ad  )�   �1  *�  &D  +�  2B  ,�  x� -{	     �)�  �  �"  P�  ��  �$   �1  ��  �&  �u  �3  �{	  ]7  ��  0�7  �U   @�1  �O  H �  ~  P6  C  tag �   Kl  	   �6  	  C  �5  N   
�  i7   �&  9  F9  8%  �*   �,  
V  ./   6
�  b 8
�   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  �  �8  N   �;  �:   4,  �6  $  �/  l9   �2  �  �  �#  �	  �'  �f  l  	  {  �   �2  ��  �  �  �   l/  ��  �  N  �  �  �   �   ;)  H�G  �#  ��   :  ��  �5  �G  F1  �	  ,8  �	   2*  �   (�*  �Z  0`1  �{  8��  ��  @ �  �-  ��  d)  sf  l  	  {  U    9  F#�  	{  �$  @J  �#  L�   y2  M�  W� O\  �� P�  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!    �-  (qV  �-  s�   Oe tV  ��  u�  � v�   �  �/  )h  n  	  �    �   g%  .�  �  �     �.  1�  �  �    �  T   �	  73  6�  �  �    �   �  �8  :     	         "3  >h  $)  Y2  8  	  V  G  �  ;  T   �6  _b  h  	  �  G  �  �  T   �3  f�  �  �  G  �  �   ;0  l�  �  	  �  G  �  	   �&  x�A  ah � M   y2  � �  H�8  � &  P�8  � V  X�'  � �  `� � �  h�9  � A  p h  �.  ��  "9  H2�  Mj  4G   H5  5;  (�)  6;  0�  7�  8�  8%  @ �0  :S  T%  �=$  ڰ  ?i   �0  @�  q5  A�  L)  B�  )  Cu  Ǟ  E�  �  F�  `Ud HU   � X+  J0  �  1  B  H  	  k  5  �  �  �  P   �&  &w  }  �  �   �1  *�  �  	  �  �   �6  -�  �  �  �   w-  1�  �  	  �  �   �;  4�  �    �   =;  8    	  *  �  �   B$  <6  <  	  P  �  �   2  @\  b  	  �  �  �  �  O   7  G�  �  	  �  �  �  �  ;   q8  N�  �  	  �  �  5   )2  S�  �  	    �  �  �  O     	  k.  ���  ah �M   #,  ��  H�4  ��  P,;  ��  XEY �6  `/q �k  hZ)  ��  p�#  ��  x'0  ��  �.  ��  ���  �P  �� ��  �`9  ��  ���  ��  �5  �  �U#  �*  � �/  �  	�  �2  �     8S  �:   �d  ��   �W  �    C  �   	:   �&  0��   y%  �	   �/  �	  �'  �	  �6  �	  �+  �	   �6  �	  ( �7  �K   *  V'�   �   �0  �*   u!  |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  �,!  2!  	  K!  �   �  K!   �	  �9  �]!  c!  s!  �   K!   A2  �!  �!  	  �!  �   �  u  �!   !  8(  �!  ��  ) !   $�  )Q!  �-  )s!   )  �!  	�!  3  <"  �� >%"   ��  ?%�    �!  #  A�!  %"  �U  �,D"  J"  �B  �r"  �� ��   Oe �r"   fP  �,~"  #  4I  P�#  ֳ  ��   �� �%#  �q �K#  R` �h#  �W ��#   P �#�#  (�U  �#�#  0�v  �#$  8�v  �#;$  @�J  �#f$  H 	�"  ��  �J"  wq  �1#  7#  	  K#  8"  	   �J  �W#  ]#  h#  8"   �\  �t#  z#  �  �#  8"  \   \  ��#  �#  �  �#  8"  �#   \  U  ��#  �#  �  �#  8"  8"  \  \   �O  ��#  �#  �  $  8"  \  \   �n  �!$  '$  �#  ;$  8"  i   ;O  �G$  M$  �#  f$  8"  i  \   -k  �G$  *�  ��"  	r$  M  �(  ��  G  �  �$  @    Y  �$  @    �  �$  @     H'  �%h  � lF&  �  \   ��  !�  x "�  G�  #�    %�  R &�  � (�  T )\  I *\   ? ,\  $� -\  (Q .\  ,j
 0�  0� 1\  4 2\  8' 4�  < 5�  @�	 6�  D� 8�  Ha 9�  L� ;\  P}	 <\  Ty	 =\  X� ?�  \�
 @�  `	 A�  d$ B�  h � D�$  ; D^&  �$  � 0N�&  ֳ  P\   �  Q\  �3  S�&  � T�  o U�  � V�    WO  $� Y\  (i Z\  , O  �&  @    z \d&  h \'  d&  � vJ'  ��  x�   � y�  � z\   � |V'  '  � (��'  � ��   � ��  �1  ��  � �\  � �\  �	 �\  W �\  � ��  � �J'    � �\'  W ��'  \'   �?(  ��  ��   � ��  � ��  � �\   t �K(  �'  � ��(  f�  ��   � ��  	 ��(   �  m �Q(  � �%�(  �(  �  � )  �W ��(   � ��  �1  ��  	� ��  
� ��  �  �+	  .�  �\  ��  �\    ���*  ڰ  �i   �  �\  * ��  � ��  � ��  �;  ��  �1  ��  8* ��  <�G ��  @�H ��  D�* ��  H�Q  ��(  P<  ��(  `[ �!  p�U �!  x�  �!  �cC  ��  �� ��  �gC  ��*  �*�  ��  �.�  ��(  �A�  ��  �0�  ��  ���  ��  �) �+	  �Cc �?(  �Y ��  �% ��(  ��
 ��*  �W ��  �O�  �H  � �'  �(  � � )  � ��*   )  6  N+  A�  	   �� !	  � "�  q	 #�  � $\  � %�   a	 '�*  �
 'h+  �*  � 80�+  ��  2�   � 8�   9�+  � :�+  ' =�  � >�  + ?,   ��  A$  (.�  Bu  0 o  N+  > Dn+  � D!,  n+  �	 (\,  I_ #   ��   �  Cc !?(    � #h,  ',  
� &-~$  D !�,  �,  !� �"�,  ah $3   �& %F&  �"N &�&  d"M	 '�*  � � !�,  �,  k X,�,  ah .    ^ !
-  -  !� h3:-  ah 5   "ȩ  6,  0 N   �}/  �  X N
 d 5	 �	 � F �	 � 	� 
 |  � � x * d �
 � y  � !� "� #~ $!
 %� &� '� (. 0� 1b @ A�	 Qc RG Sw
 T# U� V Wa X? ` a� b� c: p� �� �� �� �� �j � � �� �7 �x �I �� �) �� �� �g �$ � �\ � �� �E �� �[ �\ �< �� �� �b �+ ��
 �� �M �� �� �C �� �� �� �� �/ � �s � �� �� � #n,  �	@�F     <  N   90  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  VC0  <v X�   ֳ  Y�  �  Z�   yK  \0  	C0  d !`0  f0  	  �0  �  �0  �0       �  
 (�  � .�0  �0  	  �0  �  �  �+   � 3�0  	�0  u 31  �[ 5T0   � 6�0  � 7�0   
�8  .�  $� �#�0  	�F     F   >1  @    	.1  $� �#>1  	��F     #1  �	 �F     � 6w1  }1  	  �1  H  H  	   � :�1  b <�   ��  =k1   	�1  �
 ?�1  	�1  � A,�1  �1  O0  �1  @    	�1  $( �!�1  	��F     �1  !2  @    	2  % �"!2  	@�F     � &�2  � (H   `�  )�  5�  *�  M} +�  X$ ,�   =
 .=2  N .�2  =2  &� C	  4  'ȩ  C#�,  'ֳ  D#�,  'x E#�  '��  F#u  (�U H	  (��  Iz,  (^�  J5  (� K�*  (� L�  (� M�  (�  N?(  (�n O�'  )� h)�  #)�  *�3  +n W�   *�3  (� l�   ,(n ��  (; ��  (� �%�  (> ��  (� ��  (��  �'�  +p �H  ,+len �     &� 	  n4  -p %H  '��  %H  '��  %�  '> %u  '.  %n4  (�U 	  (.	 �2   �  &K �	  5  '7 �'5  '��  �'H  '| �'�  'm �'�5  ': �'�5  '= �'�0  '� �'�0  '� �'�5  '> �'�0  (�U �	  (�1  ��  +b ��  +p �H  (n ��  (; ��  (� ��  (> ��  (� ��  )� )�  
 H  �  .� �6  'Ǟ  &H  '��  &H  '/� &�  '�1  &�0  '��  &�  ' &�6  ' &�6  +min �  +max �  (� �  +two u  (� H  )WD  w)@ }*6  +p ,H  +lim -H  (�* .�  ( /�   ,+mid d�  (�* d�    �  /� �.7  0.	 �-�2  1p �-H  0��  �-H  2^�  ��  2/� ��  3n ��  2� ��  2�  ��  3cur �H  2�� ��  3c ��   /� {�7  0.	 {-�2  1p |-H  0��  }-H  2^�  �  2/� �  2� �7  3n ��  2� ��  2�  ��  3cur �H  2�� ��  3c ��  ,3v ��    �  �7  @    / Eb8  0.	 E.�2  1p F.H  0��  G.H  3n I�  2� I�  2�  J�  3cur KH  2�� L�  3val M�  3c N�   /� 2�8  0.	 2&�2  0.  3&n4  0> 4&u   4� �	  ��B     #      �2;  5Q �%�  ^f Vf 50�  �%�  �f �f 5�  �%�  eg Ug 5/�  �%;  "h h 6��  �z,  �h �h 6�U �	  0i $i 6M	 ��*  �i �i 6�t �\  3j +j 6�v �\  �j �j 6S � \   k k 7�  S��B     7� ��B     7cs F	��B     8@�  6� ��(  Zk Vk 6^�  �5  �k �k 9��  �:  6/� �  �k �k 6ֳ  �  Il El 6 	�  �l l 6
 
�  4m 0m 6)  �  tm jm 6Ǟ  H  ln dn 6 u  �n �n 6c u  o o :p H  to \o 6� \  xp lp ;��B     %       6<v C�  �p �p   <��B     �s  ;  =U}  <��B     �s  ;  =U}  >��B     �s  =U}    4 7	  �C     '      ��F  5� 7 �  -q q 5�	 8 �  �q �q 5J�  9 �  �r �r 5�1  : O  Ct +t 6�  <�,  Tu Fu 6ֳ  =�,  v �u 6�U >	  �v �v 6��  ?z,   w w 67 @?(  �w �w 6Mj  A�F  �w �w 6� B�  �x {x 7�  �C     9��  �>  %�'  n�  ��6�e o�F  �x �x 6� po  y y 6� q�  ]y [y 6F q&�  �y �y 6�  ru  �y �y ?[C     �       t>  :n ��  �y �y 6A� �	  z z 6�� �	  ;z 9z :vec �;  ez _z @�o  �C      ��  ��=  A�o  B�o  �z �z 8��  C�o  �z �z Cp  3{ /{   D�o  �C      �C            ��=  A�o  A�o  ;�C            C�o  r{ n{ Cp  �{ �{   @�o  �C       �  � 1>  A�o  B�o  �{ �{ 8 �  C�o  | | Cp  \| X|   E�o  �C      @�  � A�o  A�o  8@�  C�o  �| �| Cp  �| �|    F!C     �s  >%C     �s  =Us�=T��  @\  YC       P�  i:?  BT\  } } BG\  W} U} B:\  ~} z} B-\  �} �} B \  �} �} F^C     �s  >�C     b\  =Us�=Tw =Q��=R| =X��~  E�2  pC      ��  SB�2  V~ F~ B�2  k Y B�2  b� V� B�2  �� � 8��  C�2  �� �� C�2  �� �� C
3  � � C3  ;� 5� C$3  �� �� C13  ׃ σ C>3  =� ;� CK3  u� o� GX3  �C     Ha3  Gj3  �C     Is3  pC     O       8@  Cx3  Ą   J�3  ��  �A  C�3  � � @�5  \C      p�  |�A  B�5  z� t� B�5  ؅ ҅ B�5  6� 0� B�5  �� � B�5  �� ܆ A�5  B�5  � � 8p�  C�5  k� e� C6  �� �� C6  5� -� C6  �� �� C(6  � � G56  C     G>6  �C     JG6  ��  bA  CL6  �� �� CW6  � �� Cd6  >� 8� Cq6  �� ��  K6   �  C�6  � � C�6  �� ��    <C     �s  �A  =Uw  <)C     �s  �A  =Uw  >C     �s  =Uw   K�3  P�  C�3  � ؋ C�3  ]� S� C�3  � Ԍ C�3  �� �� C�3  K� ?� C�3  � ю C�3  ԏ �� @t4  �C       ��  �JC  B�4  G� C� B�4  �� �� B�4  ϑ ˑ B�4  � � B�4  W� S� B�4  �� �� B�4  � ے B�4  W� G� B�4  � � 8��  C�4  W� S� C5  �� �� C5  �� �� C 5  t� <� C+5  Ę �� C85  �� �� CE5  �� �� CR5  V� B� C_5  =� )� Hl5  Hu5    J�3  ��  CF  L�3  @4  �C      �  .F  BF4  � � B94  �� �� B,4  � �� A4  B4  q� c� 8�  CS4  � � C`4  �� `� Db8  �C      �C     *       !D  B�8  O� M� B{8  �� ~� Bo8  á ��  M�6  ��  .	�D  A�6  B�6  � � A�6  8��  C�6  )� %� C�6  c� _� C�6  �� �� C�6  ۢ Ӣ C�6  H� <� C7  ң ̣ C7  )� � C#7  Ԥ ʤ   D�7  �C      �C     �       &	iE  A8  B�7  K� E� B�7  �� �� ;�C     �       C8  ĥ �� C8  �� �� C'8  +� � C38  �� �� C?8  �� � CK8  �� �� CW8  �� �   N.7  `�  *	AQ7  BG7  �� {� A;7  8`�  C]7  � � Ci7  w� q� Cu7  ȩ �� C�7  6� 4� C�7  _� Y� C�7  �� �� C�7  ,� (� C�7  p� b� C�7  � � O�7  �C            C�7  �� ��      >wC     t  =Us   <�C     �s  \F  =Uw  FHC     �s  FjC     �s  <�C     �s  �F  =U|  <�C     �s  �F  =U| =T�� >�C     �s  =Uw      G  a  P� -��B     �       ��G  5� - �  � � 6�  /�,  ^� X� E�j  ��B      ��  2B�j  �� �� 8��  C�j  � � <��B     t  jG  =Uv  >��B     t  =Uv     4@  	   �B     [       �H  5�   �  � � 6�  "�,  g� a� 6��  #$  �� �� E�j  8�B      �  &Bk  ڮ خ Ak  Ft�B     �s    Q� D	  �C     J      ��Q  R^�  D!5  � �� RQ E!�  6� � R�  F!�  M� ?� R�[  G!�  � � R\  H!P  ,� (� S��  Jz,  }� e� S�U K	  �� �� 7�  �'C     9��  �I  S�!  a�  �� �� TZ  6C      ��  dB�Z  � � B�Z  1� +� B�Z  �� |� 8��  U�Z  ��C�Z  �� �� C�Z  2� ,� H�Z  <HC     �s  I  =Uv =T}  >aC     $t  =Uv =T��    9��  
K  SM	 ��*  �� �� 9 �  �I  Vnn ��  ǵ õ  ?�&C     �       �J  Vn ��   � �� S/� ��  &� $� Sֳ  �'  O� I� S�n ��'  �� �� Sڰ  �i  � � >�&C     1t  =T =Q0=Rv ����=X0=Y��  9��  �J  Vmax ��  � � S/� ��  n� f� S7 �?(  ҷ η  80�  %�� �  ��>@&C     =t  =U	@�F     =T0=Q��=R0   W[  �C      p�  T�K  B3[  � � B'[  ]� W� 8p�  C?[  �� �� <�C     �s  mK  =Uv =T0 >�C     Jt  =Uv =T	��F     =Qs�   X�Z  C      C     /       X�K  B�Z  � � ;C     /       C[  >� <�   W�Y  �C        �  x�N  B�Y  f� b� B�Y  �� �� A�Y  B�Y  չ ѹ B�Y  � � 8 �  C�Y  M� K� CZ  z� v� CZ  �� �� C"Z  �� �� U/Z  ��G<Z  �!C     GEZ  �!C     GNZ  �!C     JWZ  p�  �M  CXZ  �� l� CcZ  #� � CpZ  e� Y� @�[  � C      ��  ��M  B\  � � B�[  � � YL[  � C      � C     8       �B�[  >� <� Bt[  >� <� Bh[  d� b� B][  �� �� ;� C     8       C�[  �� �� C�[  � ׾ C�[  i� g� C�[  �� �� C�[  ؿ Կ H�[  H�[     <�C     �s  �M  =Uv  >�C     �s  =Uv =T|   <�C     �s  N  =Uv  <�C     $t  .N  =Uv =T�� <"C     Wt  TN  =Uv =T
 5���� <;C     $t  sN  =Uv =T�� <XC     dt  �N  =Uv =T�� >�!C     �s  =Uv    T R  �!C       ��  �BYR   � � BLR  ^� V� B?R  �� �� B2R  �� �� 8��  UfR  ��CsR  �� �� C�R  .� $� C�R  �� �� C�R  �� �� C�R  �� �� G�R  T$C     G�R  *$C     G�R  2$C     J�R  `�  �O  C�R  �� i� C�R  �� � K�R  ��  C�R  �� �� C�R  �� �� >$C     �S  =Qw    IS  �'C     �       .P  CS  �� �� CS  9� 5� >(C     1t  =Uw =T4=Q0=R| =X0=Y��  J$S  ��  �P  C%S  u� q� C0S  �� �� C=S  �� �� JJS   �  }P  CKS  &�  �  >H)C     1t  =Uw =T@=Q0=R} 
��=X0=Y��  @L[   *C      @�  f�Q  Bt[  s� o� B�[  �� �� Bh[  w� m� B][  �� �� 8@�  C�[  0� *� C�[  �� {� C�[  ;� 5� C�[  �� �� C�[  �� �� H�[  H�[  K�[  ��  C�[  D� >� Z�*C     =T} =Q|     <"C     �s  �Q  =Uv =T�� <%"C     �s  �Q  =Uv =T|  <:$C     �s  �Q  =Uv  >B$C     qt  =Uv     /0 , R  0Q ,�  2��  .z,  2ڰ  /i   &� 6	  [S  'M	 6#�*  '^�  7#5  '�  8#\  'ֳ  9#\  (�U ;	  (ڰ  <i  (�1  =�  (� >�  +p ?H  (��  @H  )�  )� )WD  *S  +q uH  +q2 vH  ,(��  ~�  (b ~�    *$S  +n ��  (/� ��   ,+n ��  (/� ��  (�m  ��  ,+cur �?(     . 
�S  'M	 
#�*  'ڰ  #i  ,(� #�(  (�W #�(    4 �	  ��B     �       ��T  [p �#H  �� �� [len �#�  ;� 3� 5ڰ  �#i  �� �� 5� �#�T  7� +� %�U �	  �L6�Y  �!  �� �� :n ��  m� e� :ok ��  �� �� 7�  � C     <��B     t  �T  =U}  <U C     ~t  �T  =U} =Ts����=Q�L >n C     �t  =Tv =Qs   !  4K s	  ��B     �      �.V  [p s3H  $� � 5��  t3H  � �� 5M	 u3�*  �� �� 6� w�(  4� $� 6�U x	  �� �� 6ڰ  yi  � � 7�  ��B     7� ���B     9�  �U  6� ��  h� T� 6� ��  � �� :q �H  �� ��  <��B     ~t  V  =U} =T =Q�L <��B     t  V  =U}  > �B     t  =U}   4� F	  �B     �       �YW  [p F0H  �� �� 5��  G0H  �� �� 5M	 H0�*  � � 6/� J�  �� r� 6� J�  =� 7� 65 J!�  �� �� 6	 K�(  �� �� %�U L	  �L6ڰ  Mi  �� �� 7�  eN�B     7� hN�B     >��B     1t  =T4=Q0=R} ����=X0=Y�L  4G ,	  P�B     u       �CX  [p ,-H  � � 5��  --H  �� �� 5M	 .-�*  �� �� %�U 0	  �\6ڰ  1i  o� i� :len 2�  �� �� 7�  ?P�B     <��B     ~t  (X  =Tv����=Q�\ >��B     �t  =T| =Qv   4% �	  ��B     �      ��Y  [p �1H  �� l� 5��  �1H  �� �� 5M	 �1�*  m� e� 6ڰ  �i  �� �� 6�n ��'  � � 6� ��  �� �� :n ��  ,� *� 6/� ��  T� P� 6� ��  �� �� 6�U �	  �� �� 7� 0�B     7�  *�B     ;H�B     O       6�N  ��  �� �� >j�B     1t  =T(=R�������=Y��   &� G	  Z  'N G#'  '^�  H#5  -idx I#�  ' J#\  '� K#u  (� M�  (�1  N�  (�  O\  (ֳ  P\  (�U Q	  )�  �)� �)WD  �,+p fH  (��  gH  ( h�    &� !	  �Z  '^�  !"5  ' ""\  'u #"�5  (�U %	  (/� &�  (�Y  '�  )�  @ &� u  [  '�& !R&  (�Y  u   \} �	  L[  0�& � R&  0^�  � 5  2�U �	   \ �	  �[  1pp �*5  0��  �*H  0� �*�1  0� �*	  2�U �	  3p �H  2� ��  2~ ��  2Kp  �%�  ]� �]�  �,2)  ��1    \B ~	  \  1pp ~$5  0��  $H   &/ C	  b\  'ȩ  C,  '^�  D5  '� E�  '�  F�  'ֳ  G�   4 �	  0C     �      ��f  5ȩ  �",  /� '� 5^�  �"5  �� �� 5� �"�  � �� 5�  �"�  �� �� 5ֳ  �"�  +� � 6�U �	  E� � :p �H  � �� 6��  �H  	� � 7�  =xC     9��  va  :n ��  T� R� 6N ��  �� x� 6/� �%�  m� g� 6��  �$  �� �� 6Ǟ  ��F  "� � 9��  _  :i ��  ~� z� 6� ��  �� �� 6��  �&�  4� *� 6i�   [+  �� �� ?C     v       �^  :vec ;  �� {� @�o  �C      ��  w^  A�o  A�o  8��  C�o  �� �� Cp  � �   E�o  �C       �  A�o  B�o  R� N� 8 �  C�o  �� �� Cp  �� ��    ?@C     8       �^  :vec ";  � �  >=C     b\  =U =T~ =Q��~  @�f  �C      0�  �1a  B�f  A� 1� B�f  !� �� B�f  ]� M� 80�  U�f  ��C�f  � � C
g  ]� W� Cg  �� �� C$g  Y� Q� C1g  �� �� C<g  !� � CIg  � � CVg  �� �� Ccg  �� �� Hpg  Hyg  G�g  �C     J�g  ��  .`  C�g  �� �� >�C     1t  =T =R} ����=Y��  @�[  C      �  Ha  B\  �� �� B�[  �� �� YL[  C      C     _       �B�[  � � Bt[  � � Bh[  <� :� B][  a� _� ;C     _       C�[  �� �� C�[  �� �� C�[  �  �  C�[  / % C�[  � � H�[  H�[     K�g  @�  C�g  � �    <�C     �s  Ia  =U~  <�C     �s  aa  =U~  >�C     �s  =U~   @�g  �C      ��  8zf  B�g    B�g  � � B�g     8��  U�g  ��~C�g  � � C�g  B 8 Ch  � � Ch  �	 �	 Ch  g
 _
 C'h  �
 �
 C3h  � � C?h  (  GJh  �C     GSh  �C     G\h  �C     Heh  Gnh  C     @�[  ]	C      P�  U9c  B\  � � B�[  � � TL[  ]	C      `�  �B�[    Bt[    Bh[  X T B][  � � 8`�  C�[  � � C�[  $  C�[     C�[  � ~ C�[  j \ H�[  H�[     @Wj  �	C      ��  Zbc  Bdj  @ 8  J�h  ��  ,f  U�h  ��C�h  � � K�h  0�  C�h  ,  C�h  � � C�h  � � C�h  V J C�h  � � J�h  ��  �c  C�h  L @ C�h  � �  Di  $C      $C            
_d  B!i  ~ | <0C     p  Qd  =Uu =Tt ^~j    F9C     �t   @.i  CC      п  %e  BKi  � � B?i    8п  CVi  J H Cbi  r n <TC     p  �d  =Uu =Tt ^~j    <�C     �q  e  =Q��^j   ^j  �� ><C     �t  =U��~=T1=Q1   @oi  �C       �  f  B�i  � � B�i  � � B�i  � � B�i  U O B�i  � � 8 �  C�i   � C�i  W Q C�i  � � G�i  �C     J�i  P�  �e  C�i    C�i  < :  >eC     �t  =U��~=T3=Q0   >C     �q  =Q��^j   ^j  ��   Owh  �C     H       C|h  c _ >C     1t  =T8=R��~�����=Y��~    <[C     �s  �f  =U~ =T��~�R" >�C     �s  =U~ =T}   &{ /	  �g  'ȩ  /',  -p 0'H  '��  1'H  (�U 3	  (��  4$  (ڰ  5i  (i�  6[+  (�1  7�  +i 7�  (/� 7�  (� 7&�  (ϋ 8�  (= 8�  )� �) �)�  �*�g  (�N  Y�   ,(��  p�    \� �	  i  0ȩ  �%,  1p �%H  0��  �%H  2�U �	  2ڰ  �i  2�1  ��  2*p ��  2� � �  3i �)�  2/� �,�  2�� �3�  +x  �  )� &) %)�  ") �	)V	 	*�h  (�N  (�   ,+pos ^i  +cur _;  ,(��  g�  ($ g�  (� g&�  (�Z g7�  +n gC�  ,+idx ��  (�� ��      �  i  @    /� �.i  0ȩ  �,   \ �	  oi  0ȩ  �",  1to �";  2��  �$  2�U �	   \� �	  �i  0ȩ  �#,  0� �#;  0� �#;  1to �#;  2��  �$  2Mj  ��F  2�U �	  ]�  �,3vec �;  3tag �H    \# 	  Wj  0ȩ  ",  1to �";  2��  �$  2Mj  ��F  2�U �	  ]�  �,3n ��    /	 xqj  0ȩ  x,   /� O�j  0ȩ  O',  2��  Q$  2Mj  R�F  2��  S�  2��  S�  ,3p1 c;  3p2 d;    /� 5�j  0ȩ  5,  2ڰ  7i   /0 (k  0ȩ  (#,  0��  )#$   QK �N  � C     
       ��k  Rϖ �&�  � � R�E  �&G  � � _� C     �t  =U	��F     =T�T  Qw c	  � C     �       ��l  RQ c�    R� d�0  � | R� e�0  � � R� f  (   R� g  � � S��  iz,  � � S� j�*  ] U SA� k	  � � S�� k	  8 2 Sֳ  l�  � � FC     �t  F4C     �t   Q� B	  ��B     5       �Bm  `Q B�  URJ�  C�  � � ` D�+  QS��  Fz,    S�U G	  > : a�  ]��B     ;��B            S� S�*  x v   \D 	  �m  0Q  �  0�    �  0c� ! �  04 " ;  2��  $z,  2� %�*   Q� c\  ��B     �       �yn  `I_ c#\,  U`��  d#�#  TS�Y  f�  � � S��  g\  �  �  a j��B     a�  ���B     8�  Vmin l�  
!  ! Vmax m�  �! |! Vmid n�  " " S7 o?(  �" �"   Q� F�  ��B     h       �o  `I_ F#\,  U`��  G#\  TVmin I�  $ $ Vmax J�  T$ J$ 8��  S7 O?(  �$ �$ Vmid P�  �% �%   b� >p�B            �;o  `I_ >\,  U Q! 	  �B     V       ��o  `I_ \,  UR��  	  h& d& S�U 	  �& �& S��   z,  �& �& a�  8`�B     8��  Vn +�  ' '   \VJ  �O  p  1a �O  1b �O  3ret �"  3tmp �"   cqj  pC     �       ��p  A~j  A~j  C�j  @' >' C�j  e' c' C�j  �' �' C�j  �' �' K�j  @�  C�j  0( ,( C�j  j( f(   cBm   C     t       ��q  BSm  �( �( B_m  8) 4) Bkm  u) q) Bwm  �) �) C�m  N* B* C�m  �* �* JBm  p�  Tq  B_m  �+ |+ Bkm  �+ �+ Bwm  4, ,, BSm  �, �, 8p�  L�m  L�m  FqC     �s    <1C     �8  �q  =Us =T�T=Q�Q=Rv  F�C     �s   c�i  �C     �       �,r  Aj  Aj  Aj  Cj  - �, C*j  f- ^- C6j  �- �- GBj  �C     IJj  �C     )       r  CKj  �- �-  >C     �t  =T1=Q0  c�Q  �C     �      ��s  B�Q  +. #. CR  �. �. LR  K�Q  ��  B�Q  �. �. 8��  LR  CR  E/ C/ W[S  /C      ��  <�s  BvS  j/ h/ BiS  �/ �/ J�S  0�  s  C�S  �/ �/ C�S  40 20 >CC     t  =Uv   <7C     t  s  =Uv  <QC     t  3s  =Uv  <kC     t  Ks  =Uv  <�C     t  cs  =Uv  <�C     t  {s  =Uv  <�C     t  �s  =Uv  >C     t  =Uv   >wC     t  =U}     dM  M  �d@G  @G  �d�a  �a  �de  e  �e@  @  �e�W  �W  `d�<  �<  �e�s  �s   �dHg  Hg  �e�I  �I   �d2n  2n  dd  d  dw  w  �d�=  �=  �d�Z  �Z  �e�`  �`   vfBY  8Y  ! e�>  �>  �e�?  �?  edF>  F>  kd\P  \P   (�   �=  &  �$ �:  �*C     �%      � ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  	0  s&  G   �  N   )  A"b  h  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  V  -    �   m�  �  �  V  U    f  ��    U   "  V  -   -   U    J   �".  4  �  PH�  Ǟ  J1   ֳ  K@   pos L@     N�  /[  O�   �K P  (�R Q>  0ڰ  SV  8O�  T1  @��  U1  H �  ��  <v �-   ��  �U    �  ��  ""  �    @   1  "  @   1  @    7  �  �   K  Q  \  "   v  :-   �  L�  x N\   y O\   �  Qh  	�  ~   w�  
  y\   �!  y\  �   z\  H  z\   "  |�  �  (j  M} N    5�  N   `�  	G   _| 
1  
!  0  ?   7  2   7  B  U     �  �  	j  �  (Q�     S)   0�  T)  N5  V�  �   W�   H� X�  �1  ZG     �  )  �  \|  �  �  N   �<  �!   �   pmoc�  stibu!  ltuo�  tolp :  ��  �8  5"V  \  �$  �4  S�  x U)   len V0  e� W7   �#  Ya  	�  �%  {�  �  �  G   G   �  U    �  �#  ��  �  G   	  G   G   U    �.  �    1  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(  �  (�/  	  0�  U   8*  �  @ w  �  u(  
1  	�  �2  (�  �  G     U      I  �3  ;    (  I   v)  ]5  ;  P  I  1  @    �3  y]  c  G   |  I  @   U    H7  ��  �  G   �  I  �   �  51  0�  y2  �<   � ��   �(  *
 �P  / �|   $ �
  ( 2$  ��  -4  	l7  +  	�1  �  $8  	�7  	8  D    	��   	O  {"  	�)  !  	�0  	l  \   	�G   �  	�N   }  	�-   )$  	�@   �   	-   c,  	+G   C*  	6U   +D  	C4    :   	�$	  xx 	��   xy 	��  yx 	��  yy 	��   5  	��  	$	  8  	�a	  ��  	�I   ��  	�}   $  	�6	  c   	�{	  �	  �	  U    �  	��	  Kl  	�U    �  	�n	   s  	��	  �"  	$�	  �	  �   	+
  �� 	-�	   �W 	.�	  Kl  	/U    %  	D;
  uR 	F�	   �
 	G�	   }  	I
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @
<
  5�  
>\   ��  
?\  �"  
A\  �"  
B\  i!  
C\   %!  
E\  (2!  
F\  0�  
G\  8   
I�  �"   
sl  ��  
u`   5�  
v`  ֳ  
x\  !  
z\  m  
{\   v  
}  J  
�#�  �  �!  �}J  ڰ  V   {3  �}  S0  �}  �/  �}  �1  ��  �1  � 0  Y/  �;
  �*  ��  (�)  �J  0+:  �00  8<8  �@0  X�*  �}  � �3  
�"W  ]  �(  ��  Oe ��/   �-  �y  ڰ  �V   U  
�"�  �  �  8�  ah ! 0   Oe "z  U1  #;
   ;+  $+,  0 i(  
�$�    l;  ��t  ah � 0   Oe �0  y2  �<   {:  ��(  (�� �I  h/ �|  p�� �-*  x T   
� �  �  _  �
H  �!  
�   �  
�  �  
�    
�  �  
�   �U 
�  (�  
�  03"  
}  8�  
�  @`  
!}  Hd  
"�  P�@  
$�	  X�;  
)�  h�   
+l  ��  
,`  �
  
-`  ���  
.`  �?!  
0`  ��  
1`  ��  
3`  ��  
4`  �ȩ  
6�  �ֳ  
7H  ��� 
8�  �K 
<�  �ڰ  
=V  �^�  
>"  �U  
@;
  �t  
B�	  �k  
CU   ��L  
E8  � "  
 U  [  1  X
m�  ��  
ot   �@  
p�	  �e 
q�  �L  
r�  P @  
$%�  �    0
\�  �-  
^y   ��  
_t  �W 
`�  x 
a�  �@  
b�	   �e 
d
  0�"  
e�  pi"  
f�  x� 
g�  ���  
i<  �.a 
kj  ��  
l}  �J  
m}  �Mj  
o�  ��  
q�  ��  
r�  �M  
tU    Z  
u-   _"  
w\  (   
x\  Ud 
zU    �L  
|0  ( �!  
F#    Z!  
AY  ��  
Ct   T 
D  �!  
El  "  
Fl   S  N   
�  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  
Y  �C  
H  0  
`)E  K  �"  �e�  �1  g$	   H+  h�   x+  i}  0��  kN'  8�)  n#�-  h�'  q%  p��  r<  t�*  y}  x O  l  �  �S  
I�  �  
�)�  �  �!  H�5  $  �U    7:  �p  s4  ��   b  8
H�  !  
Jl   m  
Kl  A� 
M�  �� 
N�  �  
P\  
  
Q\   ��  
R\  (�  
S\  0 �  
U5   x  
t[  x   
�$�  �  �!  0'0  ad  )}   �1  *l  &D  +}  2B  ,}  x� -$	     
�)=  C  �"  P��  ��  �+,   �1  ��  �&  �  �3  �$	  ]7  ��  0�7  �U   @�1  �<  H �  
~�  P6  
�  tag 
�   Kl  
�   �6  
	�  c  @
Kx  �1  
M�   %_  
NI  c  
O�  /[  
P�  ^�  
Q"   K 
RJ  (�[  
S}  0\  
Tx  8 �  �e  
V�  �5  N   

�  i7   �&  9  F9  8%  �*   �,  

�  ./   
6
%  b 
8
�   5�  
9
�  ��  
:
�  5  
;
�  Q(  
<
�    -  
I
(2  �  �8  N   
�p  �:   4,  �6  $  �/  l9   �2  
�8  8  �#  ��  �'  ��  �  �  �  J   �2  ��  �  �  J   l/  ��  �  �  �  J  �   �   ;)  H�|  �#  ��   :  ��  �5  �|  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  ��  8��  ��  @ [  �-  ��  d)  s�  �  �  �  U    1  �  �  �  �  "  t  }  }  x   �&  &�  �    t   �1  *    �  #  H   �6  -/  5  @  H   w-  1L  R  �  a  �   �;  4m  s  ~  �   =;  8�  �  �  �  H  %   B$  <�  �  �  �  H  �   2  @�  �  �  �  �  H  �  <   7  G    �  *  t  �  �  �   q8  N6  <  �  P  t  "   )2  S\  b  �  �  t  �  �  <  �   �  k.  ��i  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q ��  hZ)  �  p�#  �#  x'0  �@  �.  �a  ���  ��  �� ��  �`9  �*  ���  �P  �5  �~  �U#  ��  � �/  ��  	i  �2  ��  �  
�4  .u  ��  8Y  ��  [�   ��  \�  п  ]�  �U ^�  ��  _�   �  `�  (W�  a  0�  b`  2�  cl  4 ��  e�  �  p$3  �   |  ��  ���  ��  �}   ��  �}  *�  �8  ��  �8  	��  �8  
�  �8  .�  ��  ��  ��  (��  ��  <�  ��  X0�  ��  pY�  �}  xA�  �}  |M�  ��  ���  ��  ���  �8  �W�  �8  ���  �  ��  �  ���  ��  �[�  ��  ���  ��  ���  ��  ���  ��  ��  ��  � `  �  @    `  �  @   	 l  �  @     `  �  @    `  �  @    c�  �E  �  �#   E  8�  ��  ��  K  ��  8   +�  K  r�   �   �  [�  "  0�   (,   ��  *�   �~  +�  U�  -,   ª  .<   (��  /L   �|�  1�  P�  2�  ��  4\   ��  5l   �n�  7�  (��  9|   0��  A�   ���  B�  � �  <   @    �  L   @    Q  \   @    '  l   @    �  |   @    �   �   @    �  �  �   @    ��  D�   ^  �  N   4�   �   5�  B�  �  ��   �  <�   c�  N   {""  �   ��  x�  �  Q�  ��  ��  f�  ��  �  	�  
Ƹ  {�  ��  [�  l�  ��  �  p�  i�  ��  ��  ��  �  ��  ��  4�  ��  T�  �  ۳  =�  $�   ��  !e�  "4�  #�  $[�  %��  &��  '��  (7�  )�  *2�  +p�  ,��  -x�  - 
�  ��   $�  )$;"  A"  P�  a�  ,R"  X"  �  q"  V  q"  w"     /"  ;�  1�"  �"  �"  /"  �  �  �  �   w�  8�"  �"  �"  /"   *�  ; #  � =F"   �� >}"  �� ?�"   M�  A#  �"  ��  h!#  $#  ��  ��  u-5#  �#  ��  8V�#  �7  X#   ��  Y�#  �R Z#$  �� [�#  �� \�#   �� ]$  (a� ^J$  0 	;#  t�  ��#  �#  �#  #   S�  ��#  �#  �#  #  �  �   !�  ��#  ��  �$  $  #$  #  �   e�  
0$  6$  �  J$  #  �   |�  1W$  ]$  �  {$  #  {$  /"  p   �  �  �!�$  �$  ì  ��  �-�$  %  �  8�%  �7  ��$   ��  �"%  �R ��%  O� �@%  �  �m%   y� ��%  (a� ��%  0 	�$  ��  �/%  5%  @%  �$   ��  �M%  S%  m%  �$  �  }  �   i�  �z%  �%  �%  �$  �  �  I   p�  &�%  �%  �%  �$  �  I   !�  D�%  �%  �  �%  �$  �   %�  j�%  �%  �  &  �$  {$  /"  p   ��  �S&  ��  �b&   �� �w&  � ��&    #  b&  J   S&  )#  w&  J   h&  �$  �&  J   }&  ��  �&  �  � �&  �&  8S  ��&  �d  ��   �W  ��   C  ��&  	�&  �&  0�N'  y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��&  hG  5�'  num 7}  str 8�   *f  :['  �_  =�'  key ?�'   Kl  @4    �K  D$�'  �'  �d  H�'  �'  �  �'  �'   �'  �r  K�'   (    (  �'  �'   Uj  (Op(  ��  Q�   ֳ  R�  [M S�  �V  U�'  �F  V�'  �B Xp(    �'  �@  \ �(  (  9  F#�(  	�(  �$  @J)  �#  L�   y2  M<  W� Oi)  �� P�)  �,  Q�)   M4  R�)  (�;  S�)  0�*  T!*  8 c/  X!)  !)  �-  (qc)  �-  sy   Oe tc)  ��  u<  � v�   �(  �/  )u)  {)  �  �)  )  �   g%  .�)  �)  �)  )   �.  1�)  �)  �)  )  �)  �   1	  73  6�)  �)  �)  )  �    �8  :*  *  �  !*  )  )   "3  >u)  $)  Y9*  ?*  �  ]*  �  �  p  �   �6  _i*  o*  �  �*  �  �  �)  �   �3  f�*  �*  �*  �  �  �    ;0  l�*  �*  �  �*  �  �  �   �&  x�H+  ah � �   y2  � <  H�8  � -*  P�8  � ]*  X�'  � �*  `� � �*  h�9  � H+  p   �.  ��*  "9  H2�+  Mj  4�   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :Z+  T%  �=+,  ڰ  ?V   �0  @�  q5  A�  L)  B�  )  C  Ǟ  E�+  �  F�+  `Ud HU   � X+  J7,  �+  U   *  V'O,  U,  �0  �*   u�,  |#  w�   �#  x�  � y�  C4  z�   �&  |Z,  �'  ��,  �,  �  �,  C,  �  �,   a	  �9  ��,  �,  �,  C,  �,   A2  �-  -  �  +-  C,  �    +-   �,  8(  j-  ��  )�,   $�  )�,  �-  )�,   )  1-  	j-  3  <�-  �� >%�-   ��  ?%C,   w-  #  A|-  �-  �U  �,�-  �-  �B  ��-  �� �+   Oe ��-   fP  �,.  �.  4I  P��.  ֳ  ��   �� ��.  �q ��.  R` ��.  �W �/   P �#B/  (�U  �#r/  0�v  �#�/  8�v  �#�/  @�J  �#�/  H 	.  ��  ��-  wq  ��.  �.  �  �.  �-  �   �J  ��.  �.  �.  �-   �\  ��.  /  �  /  �-  I   \  �"/  (/  �  </  �-  </   I  U  �N/  T/  �  r/  �-  �-  I  I   �O  �~/  �/  }  �/  �-  I  I   �n  ��/  �/  </  �/  �-  V   ;O  ��/  �/  </  �/  �-  V  I   -k  ��/  �  �(  �]  N+  �D  &�  J  00  @    �  @0  @    �  P0  @    V0  �  e0  t   k0  �  �0  t  �  �  �   �0  �  �0  t  |    H'  �%  N�  #�0  �0  I  �0  �   :�  )�0  �0  �  �0  �   8�  /�0  �  5&1  V 7I   x 8�   ��  :�0  ��  =$>1  D1  ��  (?y1  I_ A�.   J�  B�  �m Cy1    &1  ! ED1  f�  M�1  �1  �  �1  �  �   �  U�1  �1  �1  �  �   ��  Y�1  �1  �  2  V  21  �  �1  �1  �   r�  a2  2  �  32  21  I   ��  e?2  E2  I  Y2  21  </   ��  @i�2  4v k �0   �y m �1  v n 2  Ty o 32  hn q �0   S�  r �0  (��  s �2  0��  t �2  8 	Y2  q�  i�2  �2  7  �   I;3  ��  K}   ��  L}  ��  M}  R` O;3  K�  PA3   l  |  ��  R�2  ��  R_3  �2  I�  Z�3  ��  \l    A�  ^e3  !Ŀ  a�4  ��  c   ת  d�3  8�  e�  @"*�  f�   "��  h�   ("T iG3  0"��  k}  P"�  l}  X"��  m}  `"��  o}  h"+ p�4  p"��  q�4  x"��  rv(  �"�  t}  �"�o u�4  �"�" v�4  �"C�  w�4  �"��  y8  �"��  z8  �"}�  {$	  �"	�  |�  �"j�  }�  �"[ ~�   "�  ��   }  �  �  ��  ��3  ��  �5  �3  ��  (�g5  N  �}   ��  ��  �  ��  ��  ��  A�  ��    \�  �s5  5  �  ��5  v�  ��   }�  ��  x �}  y �}   \�  ��5  y5  I�  X�?6  ��  �   o�  ��  )r  ��  (dS  ��  0"�  �g5  81�  ��  @��  ��5  H'�  ��  P �  �K6  �5  +  a6  @    �  q6  @    !  �!
7  ah #�   �O  $�4  �"Q  %�  "g  &�  "<! *}  "� +�   "� ,t  ("�  -Q6  0"d  .a6  P": /1  ` �# 17  q6  �  `%D7  ah '�   ��  (H  X u *P7  7  !� 8.�7  ah 0�   "�  1�  0 x 3�7  V7   @7�7  ah 90    :z  8 � <�7  �7  N   �:  �!  �  H � ' �" � $ � 	u 
� � e � 
 � � A# �$ �  �  ` !Z! "Y #�% $�! %� &� '� (K  0g# 1� @� A" Q� R S$ Td  U& VD W� X�" `�! a� b� cx! p2" �I" �% ��  �E! �~ �. �� ��! �� �'# �d �B% �a% � �
# ��# �� �� �� �- �� �#% �'! �� �: �� �� �� �c" ��  �� �� �� �5  �0 ��% �n � ��$ �H ��# �� � ��  ��" �[# � �A  &e0  �V  ,�0  b�  08:  	':  tG  0`:  ]o 2!:   �  3!:   �d  )P0  ��  ,}:  	l:  `p  ,�:  g .`:    ܨ  !�:  �:  �  �:  t  �:     *�  %�:  �:  �  �:  t  �:   �3  ]�  )�:  ;  }  ;  t   ��  ,;  #;  �  7;  t  7;   �  ��  0I;  O;  �  r;  t  ""  �  U   �   ��  7�;  	r;  �  (7�;  ��  9�:   Ъ  :�:  �  ;�:  ݱ  <;  ��  ==;    #N \)3:  	��F     #� p*x:  	��F     #T �&~;  	��F     �&  $<  @    	<  #� �#$<  	`�F     $�  �	��F     �I  `U<=  Q  W�   �g  X�  �;  Z�  �U  [�  �B ]l   �o  ^l  "Y  `<=  (+I  a<=  8
  c`  H�!  d`  J�   e`  LH  f`  N�`  hl  P�X  il  RO  k`  T,G  l`  V�t  m`  X �  L=  @    I  oQ<  �g  8�6>  ��  ��   )r  �`  dS  �`  
�B  �`  �P  �l  �p  �`  �K  �`  =  �`  me  �`  +^  �`  �]  �`  �u  �6>  
h  �`  $^K  �l  &tR  �U   (%?  �U   0 `  F>  @    �]  �X=  �S  8?A?  ��  A�   )r  B`  dS  C`  
�B  D`  �A  Fl  �n  H`  �n  I`  �W  J`  me  K`  +^  L`  �]  M`  �u  O6>  
h  Q`  $�V  Rl  &tR  XU   (%?  YU   0 �u  [R>  JW  �xA  ��  zl   =  {`  �<  |l  tB  }l  �k  ~l  �m  `  
�D  �`  gJ  �`  !X  �`  �S  �`  5f  �`  ?X  �`  �a  �`  �_  �`  �a  �`  Gf  �`  �=  �A   �E  ��  0F  ��  8�A  ��  @F  ��  H�E  ��A  P5D  �l  TH  �l  V#l  �l  X$r  �`  Z_S  �`  \'N  �`  ^?_  �l  `L  �l  b�O  ��  h�O  ��  p~e  �`  x [  �`  z0m  �l  |�M  �l  ~rM  �l  �]  �l  ��g  �l  � 8  �A  @   	 %  �A  @    �X  �N?  kE  @�9B  �^  ��   zp  ��  dv  �`  �i  �`  �<  ��  �F  ��   �D  ��  (�p  ��  03X  ��  8 �b  ��A  K_  @�'C  ��  ��   �J  ��  �<  �l  e  �l  $� �l  dk  �l  ![  �l  L^  �l  �`  �'C  yN  �7C  ,ma  �GC  4�Z  �%  :�q  �%  ;r  �8  <�u  �8  = %  7C  @    %  GC  @    %  WC  @    	l  �FB  �M  (8ED  ��  :�   �T  ;l  �P  <l  
�K  =l  B  >l  ^  ?l  �g  @l  /o  Al  %B  Bl  �O  Cl  �<  Dl  �]  El  *w  Fl  dW  Gl   �F  Hl  " e=  JdC  |[   O�D  ��  Q8   �\   R8  red  S8  q   T8   �[   VRD  �?  ( ��D  `a   �l   �L   ��D  r   ��D  &W   �l  �F   ��D    x  Ik   ��D  >i   !JCE  tag !L�   ��  !M�  /� !N�  �f  !OCE   �  2\  !QE  G   !��E  Tag !��   g  !��  �=  !��  Ja  !��   mn  !��E  UE  �v   !�F  �T  !�l   �Y  !�l  D  !�l  S  !�l  E]  !�l  ;C  !��  �: !�}   �[  !��E  DQ  !WF  E]  !l   ;C  !�  �: !}   �i  !F  >M  0!.�F  ��  !0l   �Z  !1�  vv  !2�  �r !3�F  =P  !4�  �Q  !5�F   ^�  !6"  ( F  WF  �p  !8dF  CE  !YG  �B  ![l   b  !\l   Pq  !^&G  �F  �m  !xeG  ��  !zl   �R  !{l  Up  !|G   �=  !~,G  �U  !H  �  !%   
  ! %  Sd  !!8  �Q  !"%  �G  !#%  �v  !$%  �=  !%%  sD  !&%  �\  !'%  �X  !(%  	`N  !)H  
 %  +H  @    �T  !+rG  >t  !��H  �>  !�+H   � !�+H  !  !�8  m  !�8  �[  !�8  SX  !�8   �<  !��H  8H  x@  !"�H  �  !$l   �`  !%l  TL  !&;3  �o !'�H   �H  %  �h  !)�H  �Z  !<9I  �  !>l   �f  !?�H   fR  !AI  %!ZkI  &j !\I  &�Y !]9I   ms   !V�I  �  !X   �r !_FI   J  !akI  �t  !r!�I  �I  U<  �c  (!�J  �B !�}   �c  !�}  �y !�}  �Y  !��  cC  !��   �  !�  $ 	\  !��I   L  !� 8J  >J  �i  �!��N  ah !��   �u  !�IE  ��v  !��  �R  !�l   o  !��E  (�& !�L=  0�Q  !�F>  �@  !�ED  �5�  !�  �<  !�A?  ��`  !�l  0�a  !��F  8'os2 !��A  hF�  !�9B  �j  !�}  0 M  !��  8w_ !��P  @�>  !��P  H�A  !�PQ  P^Z  !�.Q  X�f  !�.Q  `KT  !�.Q  h�i  !�U   pQ  !�U   x'mm !�U   �'var !�U   �g  !�U   ��Y !�eG  �Fq !�WC  �jQ  !��  �nQ  !��H  �m  !�I  ��P  !�D  @  !l  @B  !�Q  H�u  !  P�u  !�D  Q�;  !�  XzQ  !}  `FN  !�  hT  !}  p!u  !�  x'cvt !�Q  �2i  !�N  �)  !)�	  ��  !+�  ��j  !-�  �:>  !.�  ��_  !0  �S?  !3  �E�  !4�I  ��W  !6I  �XA  !8�  �	K  !9�  ��c  !?�  �][  !@�  ��J  !B�  �'<  !C}  �	Z  !E}   �q  !F�  �G  !G�  �T  !H�  �a  !I}   �\  !K}  (�u  !L�  0o  !M�Q  8^C  !N�  <:W  !O�4  @_  !Q}  H�@  !R�  P>  !S�  X}?  !TI  \m?  !UI  `'bdf !XJ  h�k  !\�  ��Z  !]�  �Pl  !h�  �(a  !i�  �i !mU   ��d !nU   � �Q  !��  �g  !�"O  O  �t  x!��P  ��  !�+J   ֳ  !��R  ȩ  !��  �m  !�+,  �1  !��   x !��  (^�  !�"  0��  !�}  8   !�`  <�;  !��  @�C  !�}  `� !�}  d"f !�}  h�I  !�  lpp1 !��  ppp2 !��  �Ǟ  !�bR  ��y  !�bR  �BJ  !�oR  �<  !�}  bL  !��   Ud !�U   (�W  !�}  0r�  !�}  4'pp3 !��  8'pp4 !��  HO�  !�}  X��  !�}  `�k  !�;
  h �^  !�P  �P  �  �P  +J  �  "  CE   �D  !*
Q  Q  �  .Q  O  �  �  �   �b  !A;Q  AQ  �  PQ  O   SQ  !Q]Q  cQ  nQ  O   �=  N   !T�Q  �G   �v  k_  <L  ok   �`  !_nQ  �D  <  �j  @!�bR  ڰ  !�V   �0  !�l  q5  !�`  
0�  !�l     !�`  org !��  cur !��  " !��   �   !�}  (H� !�;3  0�>  !�l  8 ,L  !��Q  @\  !�'|R  �R  �r  �d  !� �R  �R  �a  
�  @"E"S  ^�  "G"   �k "H�  ��  "I�  /� "J�  T�  "K8  z�  "L�   ��  "M�  (�f  "OCE  0Vu  "P}  8 �  "R�R  !��  "US  ��  "W�   �  "X�  /� "Z�  c�  "[S  "= "\S   l  �S  @   � ��  "^.S  Y�  ("a�S  ��  "d�   �  "e�  c�  "g;3  ��  "h;3  "�  "j�   �  "k�  $ ��  "m�S  -�  "r+T  ��  "y�   ��  "z�4   8�  "|T  9�  "�lT  z  "��   �  "��  �  "��   �  "�7T  �  "��T  ّ  "��T    lT  ��  "�xT  J�   "��T  ��  "��   ��  "��T  �  "�l  ��  "��  ��  "��T   +T  �T  ��  "��T  ��  "�!U  U  U�  �"RhW  �-  "Ty   ^�  "U"  ڰ  "VV  ��  "W�  �!  "X�   �  "Y�  ${3  "[8  (S0  "\8  )G�  "]8  *��  "_�  ,�_  "a  0�  "c"S  8Y�  "d"S  x�  "e"S  �T "g�S  ��  "h�S  ��  "j"S  89�  "k"S  x��  "l"S  �x�  "m"S  �*�  "o�  81�  "r�4  @��  "u�  H�y "v�4  Pv�  "w}  Xx�  "x�  `Ω  "zX]  h��  "{�  0��  "|e]  89�  "~K]  8�  "��&  XQ  "��2  `��  "��  h��  "��:  p:�  "��  x%�  "��  ���  "��	  ���  "� U  �ת  "��:  � ��  0"��W  ��  "�   ��  "�  �  "�U  ��  "��  3�  "��  L�  "��  ��  "��   BV "��Q  ( 4�  "�hW  !a�  H"�Z  ��  "��   ��  "��  ��  "��  п  "��  �U "��  ��  "��  W�  "�  �  "��   �  "��  (�  "��  0��  "�}  8[@ "�}  <}�  "�$	  @�  "�  `��  "��  h	�  "��  p��  "��  �j�  "��  ��  "�\  �	�  "��  ���  "��  ��  "��  ���  "��  ���  "��  �ɼ  "��  �=�  "��  �6�  "��  �!�  "��  �"�  "��  �6�  "��  �"��  "��   "��  "��  "�  "��  "$�  "��  "n�  "��   "��  "��  ("&�  "��  0"��  "�l  4"�  "�l  6"ɰ  "��  8"5�  "��  @ Z�  "��W  [�  "�$0Z  6Z  ��  �"/�Z  �  "1Z   �  "2�\  HE�  "5�W   3�  "6�  P'NDV "7�  X��  "A}  `!�  "B}  h��  "C�  p��  "D�  tx�  "F"S  x)�  "G�4  �.�  "JI  � !׬  �"��\  *�  "�8   ��  "�8  ��  "�8  �  "�8  .�  "��\  ��  "��\  x��  "��\  �"�  "��\  80�  "�  �Y�  "\  �A�  "\  �M�  "\  ���  "\  ���  "8  �W�  "8  ���  "	�\  �[�  "
�\   ��  "  ��  "�  ���  "}  ���  "}  ���  "�  ���  "�  ��  "�  ���  "\  ���  "\  �y�  "�  ���  "$Z  � \  �\  @    \  �\  @   	 \  �\  @    ��  "�Z  7�   "K]  ��  "8   �  "�  Kl  ""}  ��  "#�  M�  "&�  ��  "'�  �  "(8   ׵  "*�\  ��  "L6Z  $Z  u]  @   � ��  `#,�]  ah #.�   m #/�  X ��  #1�]  u]  !��  H#<^  ah #>�   "�� #@  0"��  #A  1"A� #C�  8"�� #D�  @ ��  #F^  �]  ��  $?-!^  '^  �  `$��^  *�  $�}   O�  $��  z�  $��  �� $��  6�  $�}   ��  $�}  $�K $��4  (h�  $��4  0ڰ  $�V  8�� $�M_  @ ��   $X�^  �� $[_   �q $`#_  add $cG_  U1 $i#_   �  _  ^  }  V   �^  #_  ^   _  �  G_  ^  }  �  �   )_  H�  $k�^  	M_  ��  $�'^  ��  $�"v_  |_  ;�  �$��_  O�  $�}   Ǟ  $�}  ��  $�}  �U $��  ڰ  $�V   �� $�d  ( ��  $�"�_  �_  Q�  $�&`  �k $�}   ��  $�}  b $� a   K�  $�"7`  	&`  =`  �  0$��`  �  $�   ��  $�a  b $ya  ��  $�a  �  $�  ֳ  $8  C�  $�   ��  $	�  $��  $�  ( (��  N   $� a  ��   }�  ��  ��  �  ��   I�  $��`  ��  $��_  ("�  N   $�ya  :�   G�  ��  Z�  z�  !�  ��  d�   �  \�  	��  
��  Ѻ   ��  $�a  (��  N   $��a  ��   ��  F�  r�  ػ  ��  ��  _�  j�  ��  	 e�  $��a  [�  $��a  �a  b  t  �   1�  $=`  	b  ��  h$u�b  �� $x�b   �q $~c  �Y $�c  �L $�c  ; $�c   �> $�3c  (nD $�\c  0�M $��c  8�: $��c  @�[ $��c  H�l $��c  P` $�
d  X�9 $�
d  ` �b  j_  }  }  V   �b  c  j_   �b  �  c  j_   
c  �  3c  j_  }   c  �  \c  j_  }  �  CE     9c  }  {c  j_  }  {c   `  bc  }  �c  j_  }  �  }   �c  �c  j_  �_   �c  �c  j_  �_  �  �c   }  �c  �  
d  j_  2`  =,  �  CE   �c  :�  $�b  	d  "�  $�|_  ��  $�<d  ;�  p$49e  ڰ  $6V   ��  $7t  ȩ  $8^  ��  $9+,  Ǟ  $:{$   �  $;{$  (��  $=�e  0��  $>�e  8�C  $@�  @� $A�  H�;  $C�   P.�  $D  X�� $E  Y8�  $F  Z��  $H  [�  $I  \�� $K�e  ` ��  $�de  �� $�e   �q $��e   ye  ye  U      /d  de  �e  ye   �e  ��  $�9e  \  ��  $b�e  Ǟ  $d}   ��  $e}  O�  $f}   Q�  $h�e  (�  $l�e  f  �   f  +J  �  �4  CE   ;�  $r-f  3f  Hf  +J  �4  �   w�  �$wch  �I $y/d   �� ${ch  p'top $|�  ��� $~sh   �y  $�h  �a�  $�}  ��  $�}  ��  $��h  �'cff $�U  ��  $�$Z   ��  $��h  (��  $��e  0׹  $�  8��  $�}  <P�  $��  @"�  $��  Dc�  $�}  H��  $�}  LT�  $��4  P0� $��4  X�o $��4  `�  $��  h;:  $�p  lzd $�  p��  $�&�e  x��  $�& f  �Q  $��2  ���  $�}  �Z�  $��4  ���  $�v(  �}�  $�$	  �	�  $��  �E�  $��   �f�  $�K  ���  $��  � �  sh  @   0 �e  �h  @    �e  �  �h  @    �	  ��  $�Hf  �  $�#�h  �h  ��  �$<�i  ڰ  $>V   ��  $?t  ȩ  $@�  ��  $A+,  Ǟ  $B{$   �  $C{$  (��  $E\  0��  $F\  8�C  $H�  @� $I�  P�;  $K�  `˹  $Lyk  ��� $M  �8�  $N  ���  $P  �b�  $RU   ��  $SU   ��� $U;k  � ^�  $��i  �i  �  �i  �h  }   G�  $��i  j  j  �h  \  \  8   r�  $�+j  1j  �  Jj  �h  \  \   h�  $�Wj  ]j  �  lj  �h    �  $�+j  ��  $��j  �j  �j  �h   ؽ  @$�k  �� $�5k   �q $��j  VY $�$�i  c $�$�i  f $�$j   2 $�$Jj  (�J $�$lj  0� $�$yj  8 5k  �h  t  H  �     k  ��  $��j  	;k  ��  N   $�yk  >�    �  /�  i�   v�  $�Mk  f�  $W�h  ��  $v�k  O�  $x}   Ǟ  $y}  ��  $z}   ��  $|�k  ��  $|�k  �k  �  $/�k  �k  ��  �$��m  �I $��k   �� $��n  �'top $�K  ��� $��n  ��y  $��k  x
Q  $��2  �
�  $��  �
�o $��4  �
��  $�}  �
��  $�}  �
+ $��4  �
��  $��4  �
��  $�v(  �
}�  $�$	  �
	�  $��  �
a�  $�}  �
�  $�}  �
�  $��h  �
E�  $��   `;:  $�p  h��  $��m  p�� $��n  xf�  $�K  ���  $��  �zd $�  ���  $��	  � �   $��m  �� $�8n   �q $�In  ;U $�hn  �" $��n   õ  $��m  �m  �  n  �k  �   �  8n  �k  t  H  �  �4  �     p  �m   n  In  �k   >n  �  hn  �k  }  �   On  �  �n  �n  }  �   �h  nn  '�  $��m  	�n  �  �n  @   � �k  �n  @    D�  $� �n  ��  �$T�o  ڰ  $VV   ��  $W+J  ȩ  $X^  ��  $Y+,  Ǟ  $Z{$   �  $[{$  (��  $]\  0��  $^\  8�C  $`�  @� $a�  P�;  $c�  `.�  $e  ��� $f  �8�  $g  ���  $i  �b�  $kU   ��  $lU   ��� $nTq  � 9�  $��o  �o  �  p  p  }   �n  ��  $�p  p  7p  p  \  \  8   �  $�Dp  Jp  �  cp  p  \  \   ��  $�Dp  >�  $�}p  �p  �p  p   ש  $��p  �p  �  �p  p   ��  @$�/q  �� $Nq   �q $}p  VY $
%�o  c $%
p  f $%7p   2 $%�p  (�J $%cp  0� $%pp  8 Nq  p  +J  �]  ^     /q  �  $�p  ^�  $��q  Ǟ  $�}   ��  $�}  O�  $�}   ��  $�aq  ��  �$�Xs  �I $��n   cff $�U  ��� $�ch  �'top $��  h�� $�Xs  p�y  $�hs  a�  $�}  �  $�}  �  $��h  ��  $�\  ���  $�\  �0�  $�  �׹  $�  ���  $�}  �f�  $�ns  �P�  $��  �"�  $��  �c�  $�}  ���  $�}  �T�  $��4  �0� $��4  ��o $��4  ��  $��  �;:  $�p  �zd $�  ���  $�$Z  ���  $�&�e  ���  $�& f  � �q  hs  @    �q  �  ~s  @    �  $��q  +�  $��s  �� $��s   �*  $�t  �" $��n   �s  �s  +J  �]  ^    p  �e   f   ~s  �s  �  t  �s  �]  �   �s  �  $��s  	t  �  $�#<t  Bt  ��  ($�t  ڰ  $V   ^�  $,u   $?6  F�  $]u  w�  $ U     ӫ  $��t  �� $��t   �q $��t  �i $�u   �  �t  /t  V  }  }   �t  �t  /t   �t  �  u  /t   u  ��  $��t  	u  ��  $�#9u  ?u  ��  }  ]u  �  �  U    Du  R�  $-.pu  �u  ��   $/�u  f�  $1�-   ]J $2�-  ��  $3�-  V $4�-   	vu  ��  X$Akv  8�  $D!kv   ��  $E!qv  �  $F!wv  ��  $G!}v  կ  $J�v   *�  $O�v  (��  $R�v  0��  $W�v  8�  $[cu  @��  $^!�v  H�  $`"�v  P Y_  d  Hk  �n  �v  }  �  l   �v  I  �v  I   �v  �v  �n  U      �v  �v  t  �  $Z   �v  'u  *t  4�  $bw  �u  " �%Ww  ah %"d   ^�  % "  ���  %"}  �I�  %#�  �װ  %%  � F %'w   %'ow  w  !� @%*�w  ��  %,Ww   ��  %.}  �Z�  %/^_  �"�  %2}  "�o %3^_   "�" %4^_  �"�  %5^_  �  %7uw  ] %7�w  uw  b  x  @    	x  #$ 7x  	��F     v N   
Rx  h  8$   � ,x  )� �x  *��   �w  +��  cw   )� ��x  *��  � �w  *��  � 
7   ,� y�  �y  *��  y
7  *��  z�w  *Ǟ  {}  *ֳ  |�  +��  ~cw  +��  }  +�# �}  -�  �./cur �}  0Wy  +΀  �}  .+�L �a    ./len ��  ./i �G   .+��  �&`  +}W �}       ,�  B�  z  *��  B!
7  *��  C!�w  *#` D!&`  +�U F�  +��  GU   +�  H=,  +�  I�  -�  s 1�" �6C     
      �~  2��  &
7  [0 W0 2��  &�w  �0 �0 3��  cw  1 �0 3��  ^  j1 b1 3�a  ^  �1 �1 3�  ^  P2 H2 3ڰ  V  �2 �2 3�U �  &3 
3 3g  �v  F4 @4 4cur }  �4 �4 3��  }  d5 ^5 4n }  �5 �5 3+�   }  #6 6 3
�  !8  �6 �6 5WD  <�9C     6�9C     b       �{  3/� H}  27 .7 7�9C     �{  8U~  7�9C     �{  8U~  7:C     �{  8U~  9*:C     8U~   6O:C     k      �|  4len ��  w7 i7 3� �  8 8 7�:C     /|  8U| 8T��� 7�:C     C|  8U~  7;C     W|  8U~  7;C     k|  8U~  9B;C     8Uv 8T���8R���#  7�6C     �|  8U~  7�6C     �|  8U~  7`7C     �|  8Uv 8Q}  7�7C     �|  8U| 8Q}  7�7C     }  8U��8T48Q}  7�7C     !}  8U~  78C     5}  8U~  :?8C     ��  M}  8Uu  7�8C     f}  8U 8T0 7�8C     }  8U 8T1 7�8C     �}  8U 8T2 7%9C     �}  8U 8T3 7L9C     �}  8U| 8Ts  7u9C     �}  8Uv 8Ts  7�9C     �}  8U| 8T0 9�9C     8Uv 8T0  1*  0C           ���  2��   
7  B8 68 2��   �w  �8 �8 3��  cw  j9 ^9 3ڰ  V  �9 �9 4cur }  Y: C: 3��  }  L; D; ;�U �  ��3�R  }  �; �; 3/� �  �< n< 4n �  �= �= 3r$ �  �> y> 3n$ !�  �? �? ;� 2�  ��3�   }  �@ }@ 38T !  �A �A 3V #Rx  �B �B 5WD  �3C     5�  
�3C     <��  P�  3ֳ  E�  �C �C <`�   �  4tmp s�  <D 8D 7�0C     �  8U�� 9�0C     8U��  <��  ��  4i �G   vD rD 4len ��  �D �D <��  N�  4p �}  E �D  =�1C     ��  8Uw 8T18Q���4$# $ &8Y��  7a1C     ��  8U�� :�2C     ��  ր  8Uw 8T18Q<8R���4$# $ &8Y�� 714C     �  8U�� :�4C     ��  %�  8Uw 8T18Q��8R| 8Xs 8Y�� 9�4C     8U��8Ts 8Q| 8R��8X1  7.0C     d�  8Us  7P0C     x�  8Us  =�3C     ��  8Uw 8T   1�# .�;C     �      ��  2��  .#
7  �E qE 2��  /#�w  �F �F 3��  1cw  �G �G 4cur 2}  �H �H 3��  3}  MJ ?J 3g  5�v  �J �J <��  ��  3��  ES3  �K qK 3/� F}  YL SL 4n F}  �L �L 3	O G^  �M �M 3ڰ  HV  
N �M ;�U I�  ��3��  J  �N �N <P�  m�  3�_ �}  �N �N 6�?C     e       H�  4len ��  LO HO 7�?C     #�  8U~  9�?C     8U��8T| 8Q} 8Rv  7>C     \�  8U~  9>C     8U~   7_<C     ��  8U~  7y<C     ��  8U~  :�<C     ��  ��  8Uw  :�<C     ��  ǃ  8Uw  7�<C     ݃  8U�� :=C     ��  �  8Uw 8T28Q08R��8X08Y�� :>=C     ��  K�  8Uw 8T88Q08R��8X08Y�� 7e=C     m�  8U~�8T| 8Qw  7�=C     ��  8U} 8Ts8Q	��F     8R8 7�=C     ��  8U~  72>C     ��  8U~  7i>C     Մ  8U~  7Q?C     �  8U~  =@C     ��  8Uu   9�;C     8U~   >� � 5C     0      �{�  ?��  �&
7  �O �O ?��  �&�w  P P @��  �cw  �P �P @�3  �{�  	Q �P @�  ��  �Q �Q #�S  ���  ��@��  ��  R R @�Y  �}  ER CR 7>5C     �  8Uv 8T68Qw 8R0 :u5C     ��  �  8T|  :�5C     ��  �  8T|  :�5C     ��  5�  8T|  :�5C     ��  M�  8T|  :�5C     ��  e�  8T|  =6C     ɝ  8Us�  $	  �  ��  @    A! �G   ��  Bc �8   CP �ӆ  D��  � cw  Eڰ  �V   Az" ��  5�  D��  �#cw  D^�  �#"  Dڰ  �#V  Dg  �#�v  E�U ��  Eֳ  ��  F�  � ,~$ �  ��  *ȩ  %�  *ֳ  �%H  *x �%�  *�1  �%<  +�U ��  +�  ��7  +F �D7  + �
7  + �z   )Z$ fه  *�  f&�   1"  \�,C            �0�  2�  \%�  lR hR 3�  ^�7  �R �R G�,C     ֝   H C�  �,C     Q       ��  2�  C%�  �R �R 3�  E�7  QS IS 3��  Ft  �S �S 3 G
7  T  T ;�  H�  �h3�U I�  VT PT =�,C     �  8T�h  )�# 11�  *F 1H  +ֳ  3D7  +��  4t  + 5
7  +�K  6�	   H� �  �+C     t       �߉  2F H  �T �T 2m �  �T �T 3ֳ   D7  KU EU 3��  !
7  �U �U 3�U "�  �U �U I�+C     �  =�+C     ��  8T|   HI$ 
�   ,C     t       ���  2F 
&H  �U �U Jreq &%  9V 3V 3ֳ  D7  �V �V 3��  
7  �V �V 3�U �  �V �V I6,C     �  =E,C     	�  8T|   Hh ��  -C     6       �O�  2ֳ  �H  'W !W 3F �D7  yW sW 3��  �t  �W �W 3 �
7  �W �W ;��  �H  �X3�U ��  X X :--C     �  A�  8T�X I=-C     �   1�# ��+C            �~�  Kϖ �J  U H� ��  0/C     /       ���  2ϖ �J  jX `X 3K ��7  �X �X 3�! �J  bY ^Y =B/C     "�  8T	��F       1*$ �P-C     �      ���  2 �t  �Y �Y 3��  �
7  Z �Y 3�O  �5  lZ fZ 3�  �'  �Z �Z 3ڰ  �V  [ [ Iz-C     /�  :�-C     ��  ��  8Uv  :�-C     ��  ��  8Uv  :�-C     ��  ٌ  8Uv  :�-C     ��  �  8Uv  :�-C     ��  	�  8Uv  :.C     ��  !�  8Uv  :%.C     ��  9�  8Uv  :?.C     ��  Q�  8Uv  :Y.C     ��  i�  8Uv  :s.C     ��  ��  8Uv  :�.C     ��  ��  8Uv  :�.C     ��  ��  8Uv  :�.C     ��  ɍ  8Uv  :�.C     ��  �  8Uv  =�.C     ��  8Uv   L� ��  pCC           ���  ?^�  �!"  E[ A[ ? �!t  �[ ~[ ?�  �!}  o] k] ?�[  �!}  �] �] ?\  �!x  �] �] @��  �
7  I^ ^ @�U ��  "` ` @Q  ��2  	a a @g  ��v  ]a Aa @ah �t  �b �b @�O  �5  �d pd @�  �'  �f �f 5�  ��JC     < �  k�  @ϖ �J  �h �h @6e  ��  	i i =�CC     <�  8T	׷F     8Q1  <��  ��  @��  ��   Oi Ai @�V ��   �i �i  <��  ��  ;E�   ~  ��{:�FC     "�  ֏  8T	��F      =GC     I�  8Tv 8Q08Rs�  <0�  |�  ;�� V+  ��{3�  Wcu  ;j 7j 3Oe X�-  �j qj :'HC     V�  ]�  8T08Qv 8R0 =�HC     V�  8T08Qv 8R0  M��  �CC      `�  �j�  N��  Sk -k O`�  P��  ��{Q��  �l �l Q̗  �m �m Qؗ  �o �o P�  ��zQ�  Vp >p R��  0DC     M�x  DC      ��  +0�  N�x  ~q Vq N�x  2s .s  M_x  0DC       �  ��  Nmx  ls hs O �  Qzx  �s �s S��  �DC      P�  Ƒ  N��  �s �s OP�  QƆ  t t 7�DC     ��  8Uv  I]FC     ��    7FDC     ۑ  8Uv� 7\DC     �  8Uv� 7rDC     �  8Uv� 9�DC     8Uv�   Mӆ  �EC      ��  8��  N�  jt Tt N��  cu Wu N��  �u �u N�  hv ^v O��  P�  ��zQ �  �v �v R,�  �IC     7�EC     ��  8Uv 8T08Q08R~  :FC     c�  ϒ  8U 8T0 :�HC     p�  �  8U 8TA :0IC     }�  �  8U  :HIC     c�  !�  8U 8T0 :sIC     ��  F�  8U~ 8T| 8Q��z :�IC     ��  d�  8U 8Q|  : KC     ��  |�  8U~  =PC     ��  8U 8T|    M�x  �IC       �  ?��  N�x  w w N�x  :w 8w N�x  qw _w N�x  <x ,x O �  Q�x  y �x Qy  �y �y Qy  �y �y Ry  :LC     T'y  `�  ��  Q(y  �z lz TWy  ��  ��  QXy  u{ k{ Tey   �  ��  Qfy  �{ �{ Uqy  `�  Qry  ^| H| Qy  ~ ~ S�y  �LC      ��  �$m�  N�y  "  N�y  >� 2� N�y  ƀ �� O��  Q�y  � � P�y  ��zQ�y  n� d� Q�y  � � R�y  JMC     7JMC     S�  8Uv 8Ts  $ &34$��F     "8Q��z8R08X0 9bPC     8U��z8Tv    :�LC     ��  ��  8U}  =�LC     ��  8U��z8T} 8Q    96JC     8Uv   V5y  pKC     �       {�  Q:y  :� 8� VGy  �KC     ,       .�  PHy  ��z7�KC     �  8Uv  9LC     8Uv 8T��z  7uKC     B�  8Uv  7KC     V�  8Uv  7�KC     j�  8Uv  9�KC     8Uv   7rJC     ��  8Uv  9�JC     8Uv   9�IC     8Uv    T�  0�  H�  Q�  m� ]� Q�  3� +� Q�  �� �� Q)�  � �� U5�  p�  Q6�  �� }� WB�  �NC     x       QC�  � � =�NC     Ǟ  8U| 8Ts     =DC     ��  8U~ 8T<8Q��z   :�CC     Ӟ  ��  8T	�F      I0GC     ��   A`  �  S�  D��   
7  E��  "�w  E��  #cw  E�O  $5  Eڰ  %V  E�U &�  Eg  (�v  F�  �.E�_ e}  Xidx e}  E��  e}  E��  e(}  .EK�  t|  .E{ ~|      Y� ��  P6C     
       ���  ?ϖ �(J  4� 0� ?� �(|  q� m� ZZ6C     �  8U	`�F     8T�T  Yh ��  p+C            ��  ?��  �,t  �� �� ?��  �,7;  � ��  Y� �}  `+C            �<�  [��  �$t  U Y�" ��  P+C            �{�  [��  �,t  U[��  �,�:  T Y� }�   +C     O       ���  [��  }*t  U[�  ~*�:  T Yc j�  �*C            ��  [��  j#
7  U Y�! H�  `/C     �       ���  ?��  H)
7  r� f� ?{ I)|  � �� \i K}  �� �� O��  @��  P�  ̇ ʇ :�/C     Ǟ  x�  8U}  =�/C     ��  8T08Q:   YC <�  `6C     %       �'�  ?��  <#
7  � � ?x =#�  0� ,� ?_| >#�  o� i� ?�H  ?#�  �� �� =~6C     �  8U�Q8Q	�R����  ]��  �6C            �m�  ^��  UW��  �6C            N��  � �   ]5�  p@C     �      ���  NG�  8� 2� NT�  �� �� Na�  ܉ ։ Nn�  .� (� Q{�  |� z� Q��  �� �� Q��  �� � Q��  E� C� Q��  k� i� S��  �@C      ��  �:�  Nˇ  �� �� =�@C     �  8Us   V5�  �AC     =      ��  NT�  �� �� _a�  Nn�  ڋ ؋ NG�  �� �� `�AC     =      a{�  a��  a��  a��  a��    :�@C     ��  ǜ  8T08Q: 9�AC     8Q} 8R| 8!  ]�  0CC     6       ���  N�  (� "� Q��  z� t� Q	�  Ȍ ƌ Q�  � � Q#�  � � V�  SCC            ��  N�  9� 7� `SCC            a��  a	�  a�  a#�  I\CC     ��    INCC     �   b�I  �I  &�b�s  �s  &�c\P  \P  
c�[  �[  '2cMc  Mc  �cIY  IY  {bno  no  (�c6U  6U  
�	c�q  �q  
q
b�B  �B  (dc$i  $i  -c�Z  �Z  
�	c�b  �b  8c�S  �S  
2	c2n  2n  cM  M  )�c@G  @G  )�c�a  �a  )�b�`  �`  &vc�D  �D  )�cw  w  )�bNe  Ne  *2d/�  %�  - b�  �  *c�?  �?  4b�t  �t  (ycF>  F>  kb$  $  +.cu  u  &yc�o  �o  �b\u  \u  ,` ;E   �C  &  p( �:  �PC     �      y� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �s  �<  �  s&  G   �  N   )  A"i  o  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  ]  -    �   m�  �  �  ]  U    f  �    U   )  ]  -   -   U    J   �"5  ;  �  PH�  Ǟ  J8   ֳ  K@   pos L@     N�  /[  O�   �K P  (�R QE  0ڰ  S]  8O�  T8  @��  U8  H �  ��  <v �-   ��  �U    �  ��  ""  �    @   8  )  @   8  @    >  �  �   R  X  c  )   v  :-   �  L�  x Nc   y Oc   �  Qo  	�  ~   w�  
  yc   �!  yc  �   zc  H  zc   "  |�  N`  N   �;  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} N    5�  N   `�  	G   _| 
8  
!  <  ?   >  2   >  B  U     �  ;  	�  �  (Q/     S)   0�  T)  N5  V/  �   W�   H� X5  �1  ZG     �  )  �  \�  �  �  N   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  �N  �8  5"�  �  �$  �4  S�  x U)   len V<  e� W>   �#  Y�  	�  �%  {    '  G   G   '  U    �  �#  �:  @  G   Y  G   G   U    �.  �f  l  �  G   G   U    �8  `�  .      �;   �1  G   �5  �  �+  �   `(  -  (�/  Y  0�  U   8*  �  @ �    u(  
�  	  �2  (:  @  G   T  U   T   �  �3  ;g  m  x  �   v)  ]�  �  �  �  8  @    �3  y�  �  G   �  �  @   U    H7  ��  �  G   �  �  �   (  51  0�\  y2  ��   � �-   �x  *
 ��  / ��   $ �Z  ( 2$  ��  -4  l>  +  ��  �  $8  �>  	�  �    ��   	�  {"  �)  !  �<  \   �G   �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U   +D  C4    :   �o	  xx ��   xy ��  yx ��  yy ��   5  �,	  	o	  8  ��	  ��  ��   ��  ��   $  ��	  c   ��	  �	  �	  U    �  �
  Kl  �U    �  ��	   s  ��	  �"  $
  "
  �   +[
  �� -
   �W .
  Kl  /U    %  D�
  uR F
   �
 G
   }  I[
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<U  5�  >c   ��  ?c  �"  Ac  �"  Bc  i!  Cc   %!  Ec  (2!  Fc  0�  Gc  8   I�  �"   s�  ��  u�   5�  v�  ֳ  xc  !  zc  m  {c   v  }b  J  �#�  �  �!  �	}�  ڰ  	]   {3  	��  S0  	��  �/  	��  �1  	��  �1  	��&  Y/  	��
  �*  	�;  (�)  	��  0+:  	��&  8<8  	��&  X�*  	��  � �3  �"�  �  �(  	��  Oe 	��&   �-  	��  ڰ  	�]   U  �"�  �  �  8	;  ah 	!�&   Oe 	"�!  U1  	#�
   ;+  	$  0 i(  �$H  N  l;  �	��  ah 	��&   Oe 	��&  y2  	��   {:  	�u  (�� 	��  h/ 	��  p�� 	�   x T   � �  �  _  ��  �!  �   �  �  �  �    �  �  �   �U   (�    03"  �  8�    @`  !�  Hd  "!  P�@  $
  X�;  )�  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7�  ��� 8J  �K <�  �ڰ  =]  �^�  >)  �U  @�
  �t  B
  �k  CU   ��L  E�  � "   �  �  1  Xm�  ��  o�   �@  p
  �e q�  �L  r4  P @  $%�       0\J  �-  ^�   ��  _�  �W `�  x a�  �@  b
   �e dU  0�"  e�  pi"  f�  x� g�  ���  i�  �.a k�  ��  l�  �J  m�  �Mj  o;  ��  q�  ��  r  �M  tU    Z  u-   _"  wc  (   xc  Ud zU    �L  |n  ( �!  F#W  ]  Z!  A�  ��  C�   T Di  �!  E�  "  F�   S  N   �i  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  �C  H]  0  `)�  �  �"  �	e  �1  	go	   H+  	h�   x+  	i�  0��  	k�"  8�)  	n#,$  h�'  	qu  p��  	rC  t�*  	y�  x �  �  J  �S  I�  �  �)A  G  �!  H	��  $  	�U    7:  	�  s4  	��   b  8H�  !  J�   m  K�  A� M�  �� N�  �  Pc  
  Qc   ��  Rc  (�  Sc  0 �  U�  x   �$    �!  0
'n  ad  
)�   �1  
*�  &D  
+�  2B  
,�  x� 
-o	     �){  �  �"  P	��  ��  	�   �1  	��  �&  	�i  �3  	�o	  ]7  	��  0�7  	�U   @�1  	�C  H P6    tag �   Kl  	   �6  	�    �5  N   
h  i7   �&  9  F9  8%  �*   �,  
0  ./   6
�  b 8
h   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  u  �8  N   �  �:   4,  �6  $  �/  l9   �2  ��  �  �) ��
  ��  ��   �>  ��  ��  �
  �+ ��  L�' ��  N�, ��  P�* ��  R�G ��  T�* ��  V�+ ��  X�' ��  Z'- ��  [?( ��  \��  ��  ^�  ��  `�@  ��  bp  ��  d�& ��  fL* ��  hSd  ��  jp& ��  l�& ��  m* ��  n�, ��  o�& ��  p+ ��  x@- ��  ��+ ��  �& ��  �Y  ��  ��1  ��  �{& ��  ��' ��  ��) ��  ��) ��  �s, �  � �    @   ; �  *  @    �' �(  �, �)B  (  �#  �	  �'  �`  f  	  u  �   �2  ��  �  �  �   l/  ��  �  H  �  �  �   �   ;)  H�A  �#  ��   :  ��  �5  �A  F1  ��  ,8  ��   2*  �  (�*  �T  0`1  �u  8��  ��  @ �  �-  ��  d)  s`  f  	  u  U    9  F#�  	u  �$  @J�  �#  L�   y2  M�  W� OV  �� P|  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!    �-  (qP  �-  s�   Oe tP  ��  u�  � v�   �  �/  )b  h  	  |  �  �   g%  .�  �  �  �   �.  1�  �  �  �  �  H   |	  73  6�  �  �  �  �   �  �8  :�     	    �  �   "3  >b  $)  Y,  2  	  P  ;  �    H   �6  _\  b  	  �  ;  �  �  H   �3  f�  �  �  ;  �  �   ;0  l�  �  	  �  ;  �  	   �&  x�;  ah � G   y2  � �  H�8  �    P�8  � P  X�'  � �  `� � �  h�9  � ;  p \  �.  ��  "9  H
2�  Mj  
4;   H5  
5/  (�)  
6/  0�  
7�  8�  
8  @ �0  
:M  T%  �
=  ڰ  
?]   �0  
@�  q5  
A�  L)  
B�  )  
Ci  Ǟ  
E�  �  
F�  `Ud 
HU   � X+  
J*  �  1  <  B  	  e  )  �  �  �  *   �&  &q  w  �  �   �1  *�  �  	  �  �   �6  -�  �  �  �   w-  1�  �  	  �  �   �;  4�  �  �  �   =;  8
      	  $   �  �   B$  <0   6   	  J   �  �   2  @V   \   	  z   �  �  �  C   7  G�   �   	  �   �  �  �  /   q8  N�   �   	  �   �  )   )2  S�   �   	  !  �  �  �  C  !   �  k.  ���!  ah �G   #,  ��  H�4  ��  P,;  ��  XEY �0  `/q �e  hZ)  ��  p�#  ��  x'0  ��  �.  ��  ���  �J   �� �z   �`9  ��   ���  ��   �5  ��  �U#  �$   � �/  �!  	�!  �2  �"  !  8S  �4"  �d  ��   �W  �   C  �"  	4"  �&  0��"  y%  �	   �/  �	  �'  �	  �6  �	  �+  �	   �6  �	  ( �7  �E"  *  V'�"  �"  �0  �*   u#  |#  w�   �#  x�  � y�  C4  z�   �&  |�"  �'  �&#  ,#  	  E#  �"  �  E#   �	  �9  �W#  ]#  m#  �"  E#   A2  �y#  #  	  �#  �"  �  i  �#   #  8(  �#  ��  )#   $�  )K#  �-  )m#   )  �#  	�#  3  <$  �� >%$   ��  ?%�"   �#  #  A�#  $  �U  	�,>$  D$  �B  	�l$  �� 	�v   Oe 	�l$   fP  	�,}$  	l$  %  4I  P	�%  ֳ  	��   �� 	�$%  �q 	�J%  R` 	�g%  �W 	��%   P 	�#�%  (�U  	�#�%  0�v  	�#&  8�v  	�#:&  @�J  	�#e&  H 	�$  ��  	�D$  wq  	�0%  6%  	  J%  2$  	   �J  	�V%  \%  g%  2$   �\  	�s%  y%  �  �%  2$  P   \  	��%  �%  �  �%  2$  �%   P  U  	��%  �%  �  �%  2$  2$  P  P   �O  	��%  �%  �  &  2$  P  P   �n  	� &  &&  �%  :&  2$  ]   ;O  	�F&  L&  �%  e&  2$  ]  P   -k  	�F&  *�  	��$  	q&  G  �(  	��  A  �  �&  @    S  �&  @    �  �&  @     H'  	�%\  <  N   9W'  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  V�'  <v X�   ֳ  Y�  �  Z�   yK  \W'  	�'  '&  �'  �  "�   - $�   �& &�'  �% )(  �  +�   #* -�  ) .�   C+ 0�'  '  3{(  �  5�   - 6�  �, 7�  
�* 9�  �' ;�  �& =�  �+ >�   �) A(  �(  D�(  }W F�(   �& H�  �, I�  _, J�   �  �(  @    r' M�(  `* PA)  �( R�   �) S�  �+ T�  -, U�  <) V�  7* W�   +) Y�(  8& \u)  }W ^�   �  _�   �% aM)  a+  d�)  + f�   ֳ  g�  �* h�  Y  i�   r* k�)  �* ��*  �  ��   �& �*  V* �"  �}, ��  ��U �  � - �**  �)  !y+  �Y*  ah �'   �  �*  � - �e*  0*  
!1  �.�!  N   ��,  �U  3Z Ik k hp q �P R eY u[ 	<b 
Y %n �c �] �d �_ �U �l �r �i QR  �O !�\ "�g #Sh $�P %�R &�e '�j (-m 0�o 1�h @�n A:o Q�Z R�[ S�T T�c U�Y V(^ W�p X�g `:] aRl b�\ c�l p�d ��f ��U �?V ��d �0f �YQ ��O �s^ �^T �e �`e ��Q ��f �` ��_ ��b ��k �Y[ ��m �#V ��r ��s ��l ��s �kl ��q ��S ��i �<s �Hj ��X �,b �on �7U ��n �j ��h ��_ ��V ��T ��R �pq ��Q �W ��X ��j � '(  �,  �,  	  �,  �  �,   *  9' $�,  	�,  q) $-  �, &�,    �'  "-  @    	-  "( + "-  	 �F     �'  M-  @    	=-  " ' 7 M-  	 �F     �'  x-  @    	h-  "\' D x-  	��F     �'  �-  @    	�-  "�' X �-  	��F     ") g �-  	��F     �'  �-  @    	�-  "�% v �-  	`�F     "T) � M-  	@�F     �'  %.  @   % 	.  ";, � %.  	��F     ,+  [y.  I_ ]%   ��  ^P  /� _P   �' a�.  @.  #, �"}&  	@�F     $P, �x$  #* i&�,  	0�F     @"  �.  @    	�.  #�* s#�.  	 �F     %k*  �	@�F     &�+ |H  PTC     
       �v/  'ϖ |)�  `� \� '�E  })A  �� �� (ZTC     ZD  )U	 �F     )T�T  &�, ]	  �PC            ��/  '��  ],�  ڍ ֍ '�& ^,�,  � � *�  `*  �� z�  &�, �	  `QC     q      ��1  '�  �!�  � � 'ֳ  �!�  g� c� 'x �!�  �� �� '�1  �!C  � � *��  �Y*  �� �� *�  �*  �  � *�U �	  Q� O� +p �"  �� u� +len ��  C� ?� *.a ��1  �� {� *�  ��  � � *.' �i  �� � ,�  W�QC     -`�  �1  *ڰ  5]  �� �� *`�  6�  � ߓ *'' 7"  2� 0� *�  8"  Y� U� .�SC     1       �1  *��  M"  �� ��  /ZSC     gD  )T~ ����)Q0)X0)Y�L  /�RC     sD  )Uv0  �  0�) �	  C2  1ֳ  �&�  2req �&�  $��  �Y*  $�& �6  $�d  �  $�U �	  $��  ��   &�& �	  QC     L       ��2  'ֳ  ��  �� �� 'm ��  
� � *��  �Y*  E� C� *�& �6  j� h� /*QC     �D  )T0  &N' �	  �UC     k      �f=  '^�  �!)  �� �� '�% �!�  �� �� '�' �!�  �� ^� '�[  �!�  � � '\  �!*  X� T� *��  �Y*  �� �� #�U �	  ��*ڰ  �]  � �� *�  ��  � � ,�  �-XC     ,WD  ��WC     .�XC     �       14  *�  �*  � � 3�XC     �D  4  )U} )T�)Q�� /�XC     �@  )Tw   - �  6  *ah �  � � *�  *  y� q� *!, �  ۛ ՛ -P�  5  *�d    (� $� #�(  �  \*:-  !�  `� ^� 30WC     �D  �4  )T~ )QH 3`WC     �D  �4  )T| )QH /�YC     �D  )TH)Q~   .lWC     S       e5  #�� Hv  ��/�WC     �D  )U	@�F     )T0)Q��)R0  3�VC     gD  �5  )U} )T )Q0)R1)X0)Y��} 3�YC     �D  �5  )U} )Tv)Q~  3)ZC     �D  �5  )Qv  3CZC     �D  �5  )U|  /]ZC     gD  )U} )T1)Qv )X| )Y~   4�>  VC      ��  ��<  5?  �� �� 6�>  7��  8?  ��}9?  :� $� 9,?  3� � 89?  ��}9F?  G� /� :S?  �XC     :\?  �YC     :e?  �]C     ;n?  ��  n<  8o?  ��};|?   �  �8  9�?  =� ;� 9�?  �� y� 9�?  � �� 9�?  �� {� ;�?  @�  d7  9�?  آ ΢ 9�?  K� G� <[C     �D  3;[C     �D  O7  )U|  /�\C     �D  )U|   3�ZC     �D  |7  )U|  3�ZC     �D  �7  )U|  3�ZC     �D  �7  )U|  3J[C     �D  �7  )U|  3�\C     �D  �7  )U|  3]C     �D  8  )U} )T�)Q��} 3']C     �D  &8  )U| )T	~ <��}" 3@]C     �D  C8  )U| )T< 3T]C     �D  [8  )U|  3u]C     �D  s8  )U|  3�]C     �D  �8  )U|  /�]C     �@  )T|   ;�?  ��  -<  8�?  ��~8�?  ��8�?  ��~8�?  ��~8@  ��~8@  ��}8!@  ��}8.@  ��~8;@  ��9H@  �� �� 9U@  
� � 9b@  t� l� 9o@  � ֤ 9z@  ʥ ĥ 9�@  � � 3}[C     �D  d9  )U|  3�[C     E  �9  )U| )T	��F     )Q��~ 3H\C     E  �9  )U| )T	��F     )Q��} 3�]C     �D  �9  )U|  3�]C     E  :  )U| )T	��F     )Q��~ 3Q^C     �D  5:  )U| )T��}�
��3$ $ &��}"# 3o^C     E  a:  )U| )T	`�F     )Q��} 3�^C     �D  �:  )U| )T��} 3�^C     E  �:  )U| )T	��F     )Q��~ 3_C     �D  �:  )U| )T} 
��3$ $ &��}"# 38_C     E  
;  )U| )T	`�F     )Q��} 3z_C     �D  (;  )U| )Ts  3�_C     E  T;  )U| )T	��F     )Q��~ 3�_C     �D  �;  )U| )Tv 
��3$ $ &s " 3`C     E  �;  )U| )T	`�F     )Q��~ 3/`C     �D  �;  )U|  3L`C     E  �;  )U| )T	@�F     )Q�� 3�`C     �D  <  )U��})T�)Q��} /aC     �@  )T|   3=YC     �D  E<  )U|  /[YC     E  )U| )T	 �F     )Q��}  3VC     �D  �<  )U| )T0 3RXC     E  �<  )U| )T	 �F     )Q��} /wXC     �@  )U    =f=  �WC      ��  �5t=  d� b� 7��  9�=  �� �� >�=  ?f=  ��  5t=  �� �� 7��  >�=  9�=  Ӧ Ѧ 3
XC     �@  M=  )U  /XC     E  )Us       @X& ��=  1�% ��  $��  �Y*  $ڰ  �]   &J( �P  �PC     /       �>  AI_ �#y.  UA��  �#�%  T*J�  ��  �� �� *�Y  �P  f� \� *��  �P  � ק  &�+ v�  �PC            �z>  AI_ v#y.  U'��  w#P  ]� Y� *J�  y�  �� ��  &S+ e	  �PC             ��>  AI_ ey.  UA��  f	  T*��  hY*  �� �� *�  i*  � ߨ  0�+ 	  �@  1��  $Y*  1�' $�  $�U 	  $^�  )  $ڰ  ]  $9+ �'  $�  �  B�  VBWD  RB]( �C$f& &(  D�?  $, 3�  $�& 5�  $� 6�  $	�  7�  C$�* T�  $/� T�    C$�& �!{(  $�* �!�(  $O& �!A)  $�) �+A)  $1- �5A)  $�* �!u)  $& �-u)  $& �9u)  $�, �!�)  $�( ��  $�) �%�  $�( �6�  Ei ��  Ej ��  Ek ��     F�' �	  �@  G�  �*  G^�  �)  H�U �	  H�& �6  H.' �i  Hֳ  ��  ,�  	�UC      I�' ��SC     l       ��A  J��  �Y*  $� � Kڰ  �]  r� p� K^�  �)  �� �� K�  �*  © �� 3TC     $E  �A  )Tv� 3&TC     E  �A  )U|  /<TC     E  )U| )Tv   L�1  `TC     �       ��B  5�1  �� �� 5�1  Q� K� 92  �� �� 92  ۪ ת 92  !� � M(2  952  c� [� N�1  �TC            5�1  ū �� 5�1  � �� O�TC            >2  >2  >2  >(2  >52  (�TC     C2  )U�U)T0    L�@   UC     �       ��C  5�@  K� ;� 5�@  � �� 9�@  ƭ �� 9�@  � � >�@  9�@  � � ;�@  ��  �C  5�@  %� � 5�@  w� q� 7��  9�@  ȯ Ư >�@  >�@  >�@  P�@  3�UC     �D  cC  )Uv  (�UC     1E  )U�T)Q�U#�   3UC     �D  �C  )Uv  /9UC     E  )Uv )T	��F     )Qs  Lf=  @aC     A       �ZD  5t=  � � 9�=  Z� R� >�=  ?f=  ��  5t=  �� �� 7��  >�=  9�=  � � 3ZaC     �@  CD  )Us  /faC     E  )Uv     QF>  F>  kR�I  �I  �QmY  mY  	�Qf  f  	�R�`  �`  vQe  e  �Q2n  2n  	SBY  8Y   RNe  Ne  2Q�c  �c  �Q�Z  �Z  �QM  M  �Q@G  @G  �Q�a  �a  �Qd  d  R�s  �s  �Q!`  !`  �Q]>  ]>  � A[   0H  &  < �:  �aC     u#      l� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �s  �<  �  s&  G   �  N   )  A"i  o  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  ]  -    �   m�  �  �  ]  U    f  �    U   )  ]  -   -   U    J   �"5  ;  �  PH�  Ǟ  J8   ֳ  K@   pos L@     N�  /[  O�   �K P  (�R QE  0ڰ  S]  8O�  T8  @��  U8  H �  ��  <v �-   ��  �U    �  ��  ""  �    @   8  )  @   8  @    >  �  �   R  X  c  )   X�  W;  v  :-   �  L�  x Np   y Op   �  Q|  	�  ~   w�  
  yp   �!  yp  �   zp  H  zp   "  |�  N`  N   �H  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} N    5�  N   `�  	G   _| 
8  
!  <  ?   >  2   >  B  U     �  H  	�  �  (Q<     S)   0�  T)  N5  V<  �   W�   H� XB  �1  ZG     �  )  �  \�  �  �  N   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  �[  �8  5"�  �  �$  �4  S�  x U)   len V<  e� W>   �#  Y�  	�  �%  {    4  G   G   4  U      �#  �G  M  G   f  G   G   U    �.  �s  y  �  G   G   U    �8  `�  .      �; !  �1  G   �5    �+     `(  :  (�/  f  0�  U   8*  �  @ �  '  u(  
�  	(  �2  (G  M  G   a  U   a   �  �3  ;t  z  �  �   v)  ]�  �  �  �  8  @    �3  y�  �  G   �  �  @   U    H7  ��  �  G      �      5  51  0�i  y2  ��   � �:   ��  *
 ��  / ��   $ �g  ( 2$  �  -4  	l>  +  	��  �  $8  	�>  	�  �    	��   	�  {"  	�)  !  	�<  \   	�G   �  	�N   }  	�-   )$  	�@   �   	-   c,  	+G   C*  	6U   +D  	C4    :   	�|	  xx 	�	   xy 	�	  yx 	�	  yy 	�	   5  	�9	  	|	  8  	��	  ��  	��   ��  	��   $  	��	  c   	��	  �	  �	  U    �  	�
  Kl  	�U    �  	��	   s  	��	  �"  	$)
  /
  �   	+h
  �� 	-
   �W 	.
  Kl  	/U    %  	D�
  uR 	F
   �
 	G
   }  	Ih
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @
<b  5�  
>p   ��  
?p  �"  
Ap  �"  
Bp  i!  
Cp   %!  
Ep  (2!  
Fp  0�  
Gp  8   
I�  �"   
s�  ��  
u�   5�  
v�  ֳ  
xp  !  
zp  m  
{p   v  
}o  J  
�#�  �  �!  �}�  ڰ  ]   {3  ��  S0  ��  �/  ��  �1  ��  �1  ��$  Y/  ��
  �*  �H  (�)  ��  0+:  ��$  8<8  ��$  X�*  ��  � �3  
�"�  �  �(  ��  Oe �j$   �-  ��  ڰ  �]   U  
�"�    �  8H  ah !p$   Oe "�  U1  #�
   ;+  $  0 i(  
�$U  [  l;  ���  ah �p$   Oe �}$  y2  ��   {:  �b  (�� ��  h/ ��  p�� �  x T   
� �  �  _  �
�  �!  
�   �  
�  �  
�    
�  �  
�   �U 
"  (�  
"  03"  
�  8�  
(  @`  
!�  Hd  
".  P�@  
$
  X�;  
)�  h�   
+�  ��  
,�  �
  
-�  ���  
.�  �?!  
0�  ��  
1�  ��  
3�  ��  
4�  �ȩ  
6�  �ֳ  
7�  ��� 
8W  �K 
<�  �ڰ  
=]  �^�  
>)  �U  
@�
  �t  
B
  �k  
CU   ��L  
E�  � "  
 �  �  1  X
m�  ��  
o�   �@  
p
  �e 
q  �L  
rA  P @  
$%      0
\W  �-  
^�   ��  
_�  �W 
`�  x 
a�  �@  
b
   �e 
db  0�"  
e	  pi"  
f	  x� 
g�  ���  
i�  �.a 
k�  ��  
l�  �J  
m�  �Mj  
oH  ��  
q�  ��  
r  �M  
tU    Z  
u-   _"  
wp  (   
xp  Ud 
zU    �L  
|{  ( �!  
F#d  j  Z!  
A�  ��  
C�   T 
Dv  �!  
E�  "  
F�   S  N   
�v  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  
�  �C  
Hj  0  
`)�  �  �"  �e"  �1  g|	   H+  h�   x+  i�  0��  k�   8�)  n#"  h�'  q�  p��  rC  t�*  y�  x �  �  W  �S  
I�  �  
�)N  T  �!  H��  $  �U    7:  �"  s4  �   b  8
H  !  
J�   m  
K�  A� 
M	  �� 
N	  �  
Pp  
  
Qp   ��  
Rp  (�  
Sp  0 �  
U�  x   
�$&  ,  �!  0'{  ad  )�   �1  *�  &D  +�  2B  ,�  x� -|	     
�)�  �  �"  P��  ��  �   �1  ��  �&  �v  �3  �|	  ]7  ��  0�7  �U   @�1  �C  H P6  
*  tag 
�   Kl  
	   �6  
	�  *  �5  N   

u  i7   �&  9  F9  8%  �*   �,  

=  ./   
6
�  b 
8
u   5�  
9
�  ��  
:
�  5  
;
�  Q(  
<
�    -  
I
(�  �  �8  N   
�"  �:   4,  �6  $  �/  l9   �2  
��  �  �#  �	  �'  �M  S  	  b  �   �2  �n  t    �   l/  ��  �  5  �  �  �   �   ;)  H�.  �#  ��   :  ��  �5  �.  F1  �	  ,8  �	   2*  �!  (�*  �A  0`1  �b  8��  �  @ �  �-  ��  d)  sM  S  	  b  U    9  F#s  	b  �$  @J�  �#  L�   y2  M�  W� OC  �� Pi  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!�  �  �-  (q=  �-  s�   Oe t=  ��  u�  � v�   n  �/  )O  U  	  i  �  �   g%  .u  {  �  �   �.  1�  �  �  �  �  U   �	  73  6�  �  �  �  �   �  �8  :�  �  	    �  �   "3  >O  $)  Y    	  =  H  �  "  U   �6  _I  O  	  m  H  �  �  U   �3  fy    �  H  �  �   ;0  l�  �  	  �  H  �  	   �&  x�(  ah � 4   y2  � �  H�8  �   P�8  � =  X�'  � m  `� � �  h�9  � (  p i  �.  ��  "9  H2�  Mj  4H   H5  5<  (�)  6<  0�  7�  8�  8  @ �0  ::  T%  �=  ڰ  ?]   �0  @�  q5  A�  L)  B�  )  Cv  Ǟ  E�  �  F�  `Ud HU   � X+  J  �  1  )  /  	  R  )  �  �  �  7   �&  &^  d  o  �   �1  *{  �  	  �  �   �6  -�  �  �  �   w-  1�  �  	  �  �   �;  4�  �  �  �   =;  8�  �  	    �  �   B$  <  #  	  7  �  �   2  @C  I  	  g  �  �  �  C   7  Gs  y  	  �  �  �  �  <   q8  N�  �  	  �  �  )   )2  S�  �  	  �  �  �  �  C  �   	  k.  ���  ah �4   #,  ��  H�4  ��  P,;  ��  XEY �  `/q �R  hZ)  �o  p�#  ��  x'0  ��  �.  ��  ���  �7  �� �g  �`9  ��  ���  ��  �5  ��  �U#  �  � �/  ��  	�  �2  ��  �  8S  �!   �d  ��   �W  �!   C  ��  	!   �&  0��   y%  �	   �/  �	  �'  �	  �6  �	  �+  �	   �6  �	  ( �7  �2   *  V'�   �   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  �!  !  	  2!  �   �  2!   �	  �9  �D!  J!  Z!  �   2!   A2  �f!  l!  	  �!  �   �  v  �!   �   8(  �!  ��  )!   $�  )8!  �-  )Z!   )  �!  	�!  3  <"  �� >%"   ��  ?%�    �!  #  A�!  "  �U  �,+"  1"  �B  �Y"  �� ��   Oe �Y"   fP  �,e"  �"  4I  P��"  ֳ  ��   �� �#  �q �2#  R` �O#  �W �u#   P �#�#  (�U  �#�#  0�v  �#�#  8�v  �#"$  @�J  �#M$  H 	k"  ��  �1"  wq  �#  #  	  2#  "  	   �J  �>#  D#  O#  "   �\  �[#  a#  �  u#  "  P   \  ��#  �#  �  �#  "  �#   P  U  ��#  �#  �  �#  "  "  P  P   �O  ��#  �#  �  �#  "  P  P   �n  �$  $  �#  "$  "  ]   ;O  �.$  4$  �#  M$  "  ]  P   -k  �.$  *�  �k"  	Y$  4  �(  ��  .  �  �$  @    @  �$  @    �  �$  @     H'  �%i  <  N   9?%  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  Vt%  <v X�   ֳ  Y�  �  Z�   yK  \?%  	t%  p: N   J�%  �:  �0 �; 9  �9 Q�%  �- v�%  b x�%   u ~�%   !y&  ;G z�  :�  {C  �: |P   : ��%  B0  '^&  b )�   ��  *�  ֳ  +�  �  ,�   +6 .&  X= .v&  &  �3 1�&  ��  3�   /� 4�  �R  5j&   �5 7|&  �/ 7�&  |&  �0 :'  }W <�   52 =�  <v >�   �- @�&  �- @'  �&  !HM'  ;G J"  "l K�  "ul L�   �= C�'  }W E"   52 F�  <v N"'   A7 P�'  M'  : S�'  �: U�   '9 V�  �: W�  �G X�  �H Y�   �4 [�'  O8 ^X(  �: `�   '9 a�  �: b�  �G c�  �H d�  v; e�  
c� g�   �> i�'  ?> ip(  �'  �0 l�(  �4 n�   �; o�  �5 p�  �< q�  b4 r�  �  t�(   �  R1 vv(  �. v�(  v(  n4 �y�)  �> {�   �> |�  �3 }�  �0 ~�  �1 �  �5 ��  n- ��  �5 ��   . ��  �< ��  �7 �X(   �/ �X(  8�7 �X(  P�/ �X(  h �= ��(  �; ��)  �(  #6 8��*  ah �4   J> �c  �$�; �)  H$�7 ��   P$o/ ��   X%toc ��&  `$,8 ��)  x$w. �G   �$�  ��'   $�: ��  $�e �d(  %enc ��(  $W9 ��  0 �5 ��*  �)  
2  %.�  N   ��,  P0  �2 �= �> >2 e9 ?= �. H3 �: 	�7 
�> �9 �6 #0 �7 Z; �4 ]< �= �5 �;  E. !)4 "�8 #�2 $�0 %q= &3? 'e> (�> 0�< 1�0 @4 A�6 Q�8 R1 S�- T�. U�/ VN5 W�1 X= `�6 a�5 b"7 cp2 p�< �j5 �[0 ��. �33 ��1 �T/ ��3 �2 ��< �V2 ��6 �s3 �,5 ��7 �Q- �|4 ��4 �]1 �B: ��1 �/; �5/ �89 ��1 �> ��8 �? �5 ��= ��2 ��3 �V6 �86 �
. ��5 �e6 �G4 ��/ �/ ��/ �^8 ��9 ��6 ��9 ��8 ��; � ;  -  -  	  '-  �  '-  '-   �  �6 %9-  ?-  	  X-  �  �  X-   &  ? *o-  	^-  �< *�-  �= ,�,   bD ---   �<  �-  �-  	  �-  �  �  !  v   s=  $�-  �-  	  �-  �  �  U    �  ).  	�-  #P  )+.  R  +�-   bD ,�-   }8  FS.  ah H #   enc I�(   r0 K_.  +.  &�> �e$  	��F     '�. �#j-  	��F     '�3 ��-  	��F     -   �.  @    	�.  '�; �#�.  	@�F     (�*  (	��F     �%  �.  @    	�.  &�7 C�.  	`�F     �%  #/  @    	/  &�- P#/  	@�F     �%  N/  @    	>/  ''1 N/  	 �F     '�< N/  	 �F     �%  �/  @    	�/  '28 /�/  	��F     �%  �/  @    	�/  '3 ��/  	��F     '3 ��/  	��F     '�- ��/  	��F     ']: ��/  	`�F     �%  .0  @    	0  '�4 {.0  	 �F     '*= �.0  	��F     )E1 U�0  *buf U!8  +�0 V!4   ,-c Z>    )91 B�0  *buf B 8  +�0 C 4   ,-c G>    )N7 ,�0  *buf ,#8  +�0 -#4   ,-val 1N     .�. �	  �mC     ?      ��A  /^�  �)  n� 0� /��  ��*  � � /�  ��  	� � 0ah ��  8� � 0�U �	  � � 0ڰ  �]  9� 1� 0�1 �v  �� �� 1�  ��}C     2��  �6  0Cp ��'  ӹ �� 20�  �3  0�d  &(  �� �� 0M; '�  ,� � 0
6 ',�  
� �� 3�{C     #X  Y2  4U| 4T} 4Q	F�F     5SG  s  3
|C     #X  �2  4U| 4T} 4Q	��F     5SG  s  3F|C     #X  �2  4U| 4T} 4Q	��F     5SG  s  3�|C     #X  �2  4U| 4T} 4Q	w�F     5SG  s  3�|C     #X  %3  4U| 4T} 4Q	��F     5SG  s  33}C     �Y  C3  4U 4QH 3i}C     �Y  [3  4U  3x�C     �Y  ~3  4T�;$4QN  6�C     �Y  4U 0$0&4T24Q3  20�  o4  0o/ ��'  �� �� '�7 �)�'  P3�}C     #X  4  4U| 4T} 4Q	��F     5SG  s  3�}C     #X  64  4U| 4T} 4Q	��F     5SG  s  3�C     �Y  T4  4U 4Q~  61�C     �Y  4U 4Q~   7�A  �xC      ��  �^6  8�A  L� F� 9��  :�A  ��~;�A  �� �� ;�A  '� #� ;�A  e� ]� :�A  ��:B  ��;B  Ǿ �� ;B  � � <)B  ��  �5  ;*B  �� �� <5B   �  h5  ;6B  ڿ ؿ =CB  �}C     &       S5  ;DB  �� ��  6�zC     �Y  4Qv   6bzC     �Y  4U| 4Q}   3�xC     #X  �5  4Uv 4T~ 4Q	<�F     5SG  s  3MyC     #X  �5  4Uv 4T~ 4Q	B�F     5SG  s  3�yC     #X  6  4Uv 4T~ 4Q	N�F     5SG  s  3�yC     #X  O6  4Uv 4T~ 4Q	\�F     5SG  s  >zC     �Y    3�zC     #X  �6  4Q	k�F     5SG  s  38{C     Z  �6  4Uw 4T 4Q04R14X04Y~  6��C     �Y  4Uw 4Q~   7NI  �mC      ��  �`8  8kI  1� #� 8_I  �� �� 9��  :wI  ��;�I  �� ~� ;�I  D� 6� ;�I  �� �� ;�I  �� �� ;�I  �� �� ?�I  �nC     <�I  @�  �7  ;�I  ?� ;� ;�I  }� u� @�I  p�  ;�I  �� ��   3�mC     Z  �7  4Uv 4T0 3�mC     Z  �7  4Uv 4T	`�F     4Qs� 3JnC     Z  8  4Uw 4T 4Q04X04Y�� 3�nC     Z  I8  4Uv 4T	@�F     4Q}  6�nC     *Z  4Uw    7`F  �nC      `�  ��;  8F  }� c� 8rF  �� �� 9`�  ;�F  h� J� ;�F  �� �� ;�F  p� ^� ;�F  G� 9� ;�F   � �� :�F  ��:�F  ��:�F  ��~;�F  � � ;�F  �� �� ;G  e� M� ?G  VpC     <"G  ��  �9  ;#G  c� a� =0G  _C     5       }9  A1G  6�C     �Y  4U| 4Q}   6�C     �Y  4U| 4Q}   3oC     �G  �9  4Uv 4R14X��4Y�� 36oC     6Z  �9  4Uv 4T}  3eoC     6Z  �9  4Uv 4T}  3�oC     Z  4:  4U| 4TH4Q~ 4R 4X~ 4Y}  35pC     Z  L:  4Uv  3apC     *Z  j:  4U| 4T  3lpC     *Z  �:  4U| 4T~  >�sC     CZ  3:~C     PZ  �:  4Uv 4T��~��~9 3j~C     CZ  �:  4Uv 4T}  3�~C     Z  ;  4U| 4T14Q~ 4R��~#4X~ 4Y}  3�~C     ]Z  9;  4Uv 4T~ 4Q��~ 3	C     Z  n;  4U| 4TH4Q04R��~4X04Y}  3R�C     PZ  �;  4Uv 4T��~	� >��C     6Z  6K�C     PZ  4Uv 4T4��~3   7�G  �pC       @�  �<  8�G  �� �� 8�G  �� �� 8�G  �  � 9@�  ;�G  >� :�   7�E  �pC      ��  ��=  8�E  }� u� 8�E  �� �� 9��  :�E  ��~;�E  �� �� :
F  ��:F  ��;$F  � 
� ;1F  �� �� ;>F  �� �� ;KF  L� H� ?VF  �rC     3qC     �G  �<  4Uv 4R44X��4Y�� 3'qC     6Z  =  4Uv 4T}  3oqC     jZ   =  4Uv 4T}  3�qC     Z  M=  4U~ 4TH4Q04X04Y}  3�rC     �H  k=  4Uv 4Q  3�rC     *Z  �=  4U~  >�sC     CZ  >�uC     wZ  >�uC     6Z    7�D  �rC      ��  �X?  8E  �� �� 8E  � �� 9��  :(E  ��~A5E  :BE  ��:OE  ��;\E  :� 2� ;iE  �� �� ;vE  �� �� ;�E  B� 4� ;�E  �� �� B�E  <�E  0�  �>  ;�E  V� P� >�sC     CZ  6�sC     6Z  4Uv 4T}   3�rC     �G  �>  4Uv 4R84X��4Y�� 3�rC     �Z  �>  4Uv 4T8 3sC     �Z  �>  4Uv  3&sC     �Z  ?  4Uv  31sC     �Z  ?  4Uv  3�uC     CZ  <?  4Uv 4T}  >�}C     6Z  >~C     �Z    7D  )vC      p�  �^A  8*D  �� �� 8D  �� �� 9p�  :7D  ��~;DD  �� �� :QD  ��:^D  ��;kD  �� �� ;xD  i� e� ;�D  �� �� ;�D  �� �� ;�D  7� /� ;�D  �� �� ;�D  �� �� ;�D  � � ;�D  T� N� ;�D  �� �� ?�D  hxC     ?�D  G�C     35vC     �G  �@  4Uv 4R 4X��4Y�� 3LvC     6Z  �@  4Uv 4T}  3�vC     Z  �@  4Uv  3wC     Z  �@  4U~ 4T24Q04R 4X04Y}  3,wC     �Z  A  4Uv 4T 1$ >%xC     �Z  3ZxC     �Z  0A  4Uv  3dxC     �Z  HA  4Uv  6V�C     *Z  4U~    3�pC     tB  �A  4Uv 4Ts 4Q2 6�C     tB  4Uv 4Ts 4Q
   C.: 	  TB  Dpcf "�*  E�U 	  E��  �  Eڰ  ]  ECp !�'  E�y #TB  Eh�  $dB  Fnn $4   Flen $"4   ,Fs Z�   ,Fsrc d�  ,Fmm v4       �  dB  @    4   tB  @    .$8 �	  �kC     �      �D  /^�  �)  L� D� /��  ��*  �� �� /b ��  � � '��  ��  �P'ֳ  ��  �X0�U �	  f� d� 0,8 ��)  �� �� 1�4 �lC     3�kC     �G  \C  4Uv 4R�Q4X�P4Y�X 3�kC     6Z  zC  4Uv 4T�L 3#lC     Z  �C  4Uv  3�lC     �H  �C  4Uv 4Qs� 3�lC     �H  �C  4Uv 4Qs� 3UmC     �H  �C  4Uv 4Qs� 6xmC     �H  4Uv 4Qs�  C8 �	  �D  G^�  �!)  G��  �!�*  E�U �	  Eڰ  �]  E��  ��  Eֳ  ��  Fenc ��(  E�9 ��  E�  ��(  EV> ��  E�; �!�  Eb= ��  Ep7 �!�  Fi ��  Fj ��  Fpos �/  H�4 uH�  r CM< .	  �E  G^�  .)  G��  /�*  E�U 1	  E7 2�E  E��  3�  Eֳ  3�  Fpos 3�  Ew? 4�  Er? 4�  Fi 4(�  E�1 4+�  H�4 �,E�  u�    �  �E  @    C�2 �	  `F  G^�  �)  G��  ��*  E�U �	  Eڰ  �]  E��  ��  Eֳ  ��  E�e �d(  E�: ��  E�: ��  Fi �*�  H�4 ( C]7 �	  AG  G^�  �")  G��  �"�*  E3g �'  E�  ��'  Ew. ��  Er. � �  Fi �-�  E��  ��  Eֳ  � �  E�U �	  Eڰ  �]  Er$ ��  E�y �"  H�4 �,EE- r�  ,E�[ ��     C�3 ��'  �G  G��  �(�*  GCp �(.  E�  ��'  E�  �v  Fi �G    C�; �v  �G  G�R  �"j&  G0 �"�  Gb �"�  Fi ��   .0 u	  �gC     �       ��H  /^�  u&)  � �� /�R  v&j&  �� {� /0 w&�  �� �� /b x&�  k� a� /> y&�H  �� �� /�p  z&�H  �� �� 0�U |	  Z� L� Ii }�  �� �� 1WD  ��gC     6.hC     PZ  4U�U  �  C�: ?	  HI  G^�  ?)  G��  @�  G�: Ad(  E�U C	  1�  oSkC     J8I  E�k HHI   ,E�? U!�'    �%  K,. _	  �I  +^�  _)  +��  `�*  L�U b	  -toc c�&  L�R  dj&  Lڰ  f]  -n g�  Lֳ  i�  H�  ,-i ��  L�9 ��  ,-tmp �^&     M{0 !0cC            �J  Nϖ !�  U .�3 	   cC            �OJ  Nϖ �  U .^3 5  phC     
       ��J  /ϖ &�  G� C� /}W &�  �� �� OzhC     �Z  4U	@�F     4T�T  .a? �	  cC            �K  Nϖ �"�  UN�1  �"�  TN<v �"!  Q .P? �	   cC            �vK  Nϖ �"�  UN�1  �"�  TN<v �"!  Q/�h  �"v  �� ��  .�= w	  �bC            ��K  N��  w%�*  UN�7 x%'-  TNn/ y%'-  Q .*> N	  �jC     U       �]L  /��  N+�*  �� �� /M9 O+�  =� 7� /�9 P+X-  �� �� 0Cp R�'  � � 6�jC     #X  4Q�T5SG  �U  .; �	  �dC     -      ��N  /�  �!�  L� B� /ֳ  �!�  �� �� /x �!�  0� (� /�1  �!C  �� �� 0��  ��*  ]� S� 0^�  �)  �� �� 0�U �	  =� 1� 0.a ��N  �� �� 0�: �d(  T� L� 0Vu  ��  �� �� H�  BPa0  ofC       ofC     A       =	�M  8z0  � � 8n0  Z� T� @�0  ��  ;�0  �� ��   P�0  gC       gC     d       .N  8�0  �� �� 8�0  � � @�0   �  ;�0  m� W�   P�0  �gC       �gC     4       9	fN  8�0  �� �� 8�0  �� �� @�0  P�  ;�0  ?� =�   3�eC     �Z  ~N  4Us0 3�eC     �Z  �N  4Us 4T}  3fC     Z  �N  4U|  6fC     ]Z  4U| 4Q}   �  .�2 �	  �cC     �       ��O  /ֳ  �&�  j� b� Qreq �&�  �� �� 0��  ��*  )� � 0�d  �(  �� �� R�U �	  0��  ��  �� x� S�O  dC      dC     ;       �8P  �� �� 8�O  � � TdC     ;       ;P  +� )� 6dC     �Z  4Us 4T0    C�2 �	   P  Gֳ  ��  Gm ��  E,8 ��)   U�7 �	  ��C     E      ��S  V^�  �!)  ]� Q� V�/ �!�  �� �� V�  �!�  �� �� V�[  �!�  � � V\  �!7  H� D� W��  ��*  �� �� W�U �	  R� B� 1WD  ���C     H�  �2��  ?Q  0P  	  � �� 3�C     [  $Q  4U~ 4T|  6�C     [  4U~ 4T|   X��C            �Q  0$6 	  M� K� 6��C     [  4U~ 4T|   20�  7R  0o/ `"  v� p� 0�7 a"  �� �� 0�k  bv  �� �� Xp�C     �       �Q  Is g�   <� :�  9`�  '�� }�  �@6��C     [  4U	��F     4T04Q�@4R0   7�S  �C      ��  �R  8�S  a� _� 9��  ;�S  �� �� A�S  6��C     =V  4Us    7�S  @�C      ��  Z�R  8�S  �� �� 9��  ;�S  � � A�S  6V�C     =V  4Us    P�S  ��C      ��C            �NS  8�S  9� 5� T��C            ;�S  v� r� A�S  6ĄC     =V  4Us    3��C     �0  rS  4U| 4Ts 4Qv  63�C     �0  4U~ 4Ts 4Qv   )d. ��S  +�/ ��  L��  ��*  Lڰ  �]  ,-i ��  ,LCp ��'     U�: ��   bC     �       ��T  V|- �""  �� �� Y9 �#�#  TWI_ �S.  �� �� Zenc ��(  +� )� W�_ �P  V� N� W~. ��  �� �� W9. ��  �� �� W�Y  ��  -� '�  U/ i�  �aC     c       �7U  V|- i#"  {� w� V�_ j#P  �� �� WI_ lS.  
� � Zenc m�(  E� C� W~. n�  n� h� W9. o�  �� ��  [�4 _�aC     	       �xU  Y|- _"  UWI_ aS.  � �  Ux1 O	  �aC            ��U  Y|- O"  UY�h  P	  TWI_ RS.  ;� 9� W��  S�*  `� ^�  \�O  @cC     N       �=V  8�O  �� �� 8P  �� �� ;P  � � 6TcC     �Z  4Uv 4T�T  \�S  �hC     �      ��W  8�S  E� ;� A�S  ;�S  �� �� =�S  �hC            W  ;�S  �� �� =�S  �hC     E       �V  ;�S  _� [� 3iC     *Z  �V  4U}  62iC     *Z  4U}   6HiC     *Z  4U}   3�hC     *Z  W  4U}  3�hC     *Z  5W  4U}  3biC     *Z  MW  4U}  3yiC     *Z  eW  4U}  3�iC     *Z  }W  4U}  3�iC     *Z  �W  4U}  3�iC     *Z  �W  4U}  3�iC     *Z  �W  4U}  >jC     +[   \�S   jC            �#X  8�S  �� �� ;�S  �� �� A�S  O*jC     =V  4U�U  \AG  @jC     h       ��X  8`G  E� 9� ]SG  ]SG  ;mG  �� �� ;zG  7� 1� ;�G  �� �� 6ojC     8[  4T|   \�H  kC     �       ��Y  8�H  �� �� 8�H  _� W� 8�H  �� �� ;I  [ 	 U 	 X kC            CY  ;*I  � 	 � 	 66kC     Z  4U�U4T! �F      �F     �T4 $0.( 4Qs   @�H  ��  8�H  	 	 8�H  D	 >	 8�H  �	 �	 9��  ;I  �	 �	 BI  @8I  ��  :9I  �k6OkC     Z  4U�U4T	��F     4Q�k     ^e  e  
�^=T  =T  ]_BY  8Y   `�`  �`  v`Ne  Ne  2`�I  �I  �^M  M  �^d  d  `�s  �s  �^�f  �f  �^�[  �[  �^w  w  �^�D  �D  �^Hg  Hg  �^�G  �G  �^@G  @G  �^�s  �s  �^�]  �]  �^�a  �a  �^KS  KS  �^�c  �c  �^F>  F>  k^mY  mY  �^�<  �<  �^f  f  �`w< w< [`�- �- Y^2n  2n  ^~l  ~l  |`�  �   �p   �M  &  �@ �:  �C     �@      �� (\  �9   ,  i   �L   �  L   int �  �   @�   �  �    p   	@   �  #	@   X  &	@   �  )	@    �  ,	@   (�  -	@   0/  2X   8�  5X   < 	�   �  �   �  8"h   
+  K  	�   
%  L  
�  M  '  ;  �  s&  X   �  _   )  A"n  	t  �   ��  �  �f    ��  ��  <h ��  �I  ��   �  X�  	�  f   �  b  9    �   m�  	�  �  b  f    f  �
  	  f   .  b  9   9   f    J   �":  	@  �  PH�  Ǟ  J=   ֳ  KL   pos LL     N  /[  O   �K P  (�R QO  0ڰ  Sb  8O�  T=  @��  U=  H �  �  <v �9   ��  �f    �  ��  ""  �  	  L   =  .  L   =  L    	C  �  C  �   \  	b  m  .   v  :9   �  L�  x Nm   y Om   �  Qy  �  ~   w�  
  ym   �!  ym  �   zm  H  zm   "  |�  N`  _   �E  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} _    5�  _   `�  	X   _| 
=  
!  A  ?   C  2   C  B  f     �  E  �  �  (Q9     S:   0�  T:  N5  V9  �   W�   H� X?  �1  ZX     	�  	:  �  \�  	�  �  _   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  �X  �8  5"�  	�  �$  �4  S�  x U:   len VA  e� WC   �#  Y�  �  �%  {  	  1  X   X   1  f    	�  �#  �D  	J  X   c  X   X   f    �.  �p  	v  �  X   X   f    �8  `�  .      �;   �1  X   �5    �+     `(  7  (�/  c  0�  f   8*  �  @ 	�  	$  u(  
�  %  �2  (D  	J  X   ^  f   ^   	�  �3  ;q  	w  �  �   v)  ]�  	�  �  �  =  L    �3  y�  	�  X   �  �  L   f    H7  ��  	�  X   �  �  �   	2  51  0�f  y2  ��   � �7   ��  *
 ��  / ��   $ �d  ( 2$  �  -4  lC  +  ��  �  $8  �C  �  	�    ��   �  {"  �:  !  �A  \   �X   �  �_   }  �9   )$  �L   �   9   c,  +X   C*  6f   +D  C@    :   �y	  xx �	   xy �	  yx �	  yy �	   5  �6	  y	  8  ��	  ��  ��   ��  ��   $  ��	  c   ��	  	�	  �	  f    �  �
  Kl  �f    �  ��	   s  ��	  �"  $&
  	,
  �   +e
  �� -
   �W .
  Kl  /f    %  D�
  uR F
   �
 G
   }  Ie
  _   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @	<_  5�  	>m   ��  	?m  �"  	Am  �"  	Bm  i!  	Cm   %!  	Em  (2!  	Fm  0�  	Gm  8   	I�  �"   	s�  ��  	u�   5�  	v�  ֳ  	xm  !  	zm  m  	{m   v  	}l  J  	�#�  	�  �!  �
}�  ڰ  
b   {3  
��  S0  
��  �/  
��  �1  
��  �1  
�z$  Y/  
��
  �*  
�E  (�)  
��  0+:  
��$  8<8  
��$  X�*  
��  � �3  	�"�  	�  �(  
��  Oe 
�a$   �-  
��  ڰ  
�b   U  	�"�  	�  �  8
E  ah 
!g$   Oe 
"�  U1  
#�
   ;+  
$  0 i(  	�$R  	X  l;  �
��  ah 
�g$   Oe 
�t$  y2  
��   {:  
�Y  (�� 
��  h/ 
��  p�� 
�  x T   	� �  	�  _  �	�  �!  	�   �  	�  �  	�    	�  �  	�   �U 	  (�  	  03"  	�  8�  	%  @`  	!�  Hd  	"+  P�@  	$
  X�;  	)�  h�   	+�  ��  	,�  �
  	-�  ���  	.�  �?!  	0�  ��  	1�  ��  	3�  ��  	4�  �ȩ  	6�  �ֳ  	7�  ��� 	8T  �K 	<�  �ڰ  	=b  �^�  	>.  �U  	@�
  �t  	B
  �k  	Cf   ��L  	E�  � "  	 �  	�  1  X	m�  ��  	o�   �@  	p
  �e 	q	  �L  	r>  P @  	$%  	
    0	\T  �-  	^�   ��  	_�  �W 	`�  x 	a�  �@  	b
   �e 	d_  0�"  	e	  pi"  	f	  x� 	g�  ���  	i�  �.a 	k�  ��  	l�  �J  	m�  �Mj  	oE  ��  	q�  ��  	r  �M  	tf    Z  	u9   _"  	wm  (   	xm  Ud 	zf    �L  	|x  ( �!  	F#a  	g  Z!  	A�  ��  	C�   T 	Ds  �!  	E�  "  	F�   S  _   	�s  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  	�  �C  	Hg  0  	`)�  	�  �"  �
e  �1  
gy	   H+  
h�   x+  
i�  0��  
k�   8�)  
n#"  h�'  
q  p��  
rH  t�*  
y�  x 	�  	�  	T  �S  	I�  �  	�)K  	Q  �!  H
��  $  
�f    7:  
�  s4  
�	   b  8	H	  !  	J�   m  	K�  A� 	M	  �� 	N	  �  	Pm  
  	Qm   ��  	Rm  (�  	Sm  0 �  	U�  x   	�$#  	)  �!  0'x  ad  )�   �1  *�  &D  +�  2B  ,�  x� -y	     	�)�  	�  �"  P
��  ��  
�   �1  
��  �&  
�s  �3  
�y	  ]7  
��  0�7  
�f   @�1  
�H  H P6  	'  tag 	�   Kl  		   �6  		�  	'  �5  _   	
r  i7   �&  9  F9  8%  �*   �,  	
:  ./   	6
�  b 	8
r   5�  	9
�  ��  	:
�  5  	;
�  Q(  	<
�    -  	I
(�  	  �8  _   	�  �:   4,  �6  $  �/  l9   �2  	��  �#  �	  �'  �D  	J  	  Y  �   �2  �e  	k  v  �   l/  ��  	�  ,  �  �  �   	�   ;)  H�%  �#  ��   :  ��  �5  �%  F1  �	  ,8  �	   2*  �  (�*  �8  0`1  �Y  8��  �v  @ 	�  �-  ��  d)  sD  	J  	  Y  f    9  F#j  Y  �$  @J�  �#  L�   y2  M�  W� O:  �� P`  �,  Q�   M4  R}  (�;  S�  0�*  T�  8 c/  X!�  	�  �-  (q4  �-  s�   Oe t4  ��  u�  � v�   	e  �/  )F  	L  	  `  �  �   g%  .l  	r  }  �   �.  1�  	�  �  �  �  R   	�	  73  6�  	�  �  �  �   	�  �8  :�  	�  	  �  �  �   "3  >F  $)  Y  	  	  4  E  �    R   �6  _@  	F  	  d  E  �  �  R   �3  fp  	v  �  E  �  �   ;0  l�  	�  	  �  E  �  	   �&  x�  ah � +   y2  � �  H�8  �   P�8  � 4  X�'  � d  `� � �  h�9  �   p 	f  �.  ��  "9  H2�  Mj  4E   H5  59  (�)  69  0�  7�  8�  8  @ �0  :1  T%  �=  ڰ  ?b   �0  @�  q5  A�  L)  B�  )  Cs  Ǟ  E�  �  F�  `Ud Hf   � X+  J  	�  1     	&  	  I  .  �  �  �  4   �&  &U  	[  f  �   �1  *r  	x  	  �  �   �6  -�  	�  �  �   w-  1�  	�  	  �  �   �;  4�  	�  �  �   =;  8�  	�  	    �  �   B$  <  	  	  .  �  �   2  @:  	@  	  ^  �  �  �  H   7  Gj  	p  	  �  �  �  �  9   q8  N�  	�  	  �  �  .   )2  S�  	�  	  �  �  �  �  H  �   		  k.  ���  ah �+   #,  ��  H�4  ��  P,;  ��  XEY �  `/q �I  hZ)  �f  p�#  ��  x'0  ��  �.  ��  ���  �.  �� �^  �`9  ��  ���  ��  �5  ��  �U#  �  � �/  ��  �  �2  ��  	�  8S  �   �d  ��   �W  �   C  ��     �&  0��   y%  �	   �/  �	  �'  �	  �6  �	  �+  �	   �6  �	  ( �7  �)   *  V'�   	�   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  �
!  	!  	  )!  �   �  )!   	�	  �9  �;!  	A!  Q!  �   )!   A2  �]!  	c!  	  �!  �   �  s  �!   	�   8(  �!  ��  )�    $�  )/!  �-  )Q!   )  �!  �!  3  <�!  �� >%�!   ��  ?%�    	�!  #  A�!  	"  �U  
�,""  	("  �B  
�P"  �� 
��   Oe 
�P"   fP  
�,\"  	�"  4I  P
��"  ֳ  
��   �� 
�#  �q 
�)#  R` 
�F#  �W 
�l#   P 
�#�#  (�U  
�#�#  0�v  
�#�#  8�v  
�#$  @�J  
�#D$  H b"  ��  
�("  wq  
�#  	#  	  )#  "  	   �J  
�5#  	;#  F#  "   �\  
�R#  	X#  �  l#  "  U   \  
�x#  	~#  �  �#  "  �#   	U  U  
��#  	�#  �  �#  "  "  U  U   �O  
��#  	�#  �  �#  "  U  U   �n  
��#  	$  �#  $  "  b   ;O  
�%$  	+$  �#  D$  "  b  U   -k  
�%$  *�  
�b"  P$  	+  �(  
��  	%  �  �$  L    7  �$  L    �  �$  L     H'  
�%f  hG  5�$  !num 7�  !str 8�   *f  :�$  �_  =%  key ?�$   Kl  @@    �K  D$%  	�$  �d  H/%  	5%  �  D%  D%   	�$  �r  KV%  	\%  s  p%  D%  D%   Uj  (O�%  ��  Q�   ֳ  R�  [M S�  �V  U#%  �F  VJ%  �B X�%    	%   M Zp%  �@  \ �%  	p%  (@ N2&  �D PX    cF QX   RA RX   aN SX    nL U�%  2&  	2&  	�   "sz&  ;G u�   !l v9   !ul wL    G n�&  }W p�   ��  qX   M rX   <v yO&   �? {z&  �&  �A �)'  5�  �A   ��  �A  XC �:  y�  �:  �G �:  �H �:  
 �L ��&  }C 8��'  }W ��    T �L   |L �A  ZN �A  bbx �)'  .a �=   bpr �L   (Vu  �A  0 �G �5'  �M ��$)  }W ��    bbx �)'  �' �L   M; �L    
6 �L   (�C �X   0�E �A  4* �L   8G �9   @�H �9   H�A �L   PNN �L   X4x �$)  `zN �L   hQM �L   phF �$)  xiH �L   ��B �L   �3g �*)  �WA ��   �&G �L   ��L  �f   �bpp �A  �ڰ  �b  �CC �*)  �BC �L   �tH ��%  � 	�'  	�&  XF ��'  _   �+  8E  �F cG @G tD 1N H �L �B s@ 	)D 
�K �L \K �I �L O �B �G �F CJ AD  K !�@ "(B #2H $�K %lJ &�G '�I (�B 0�F 1L @@F A�I Q�M RC SaC T_B U�J VCE W�G X�@ `)L a:A blA c�K pEK ��K �,J �_E ��A ��D �6O �oM ��K ��C ��D ��M ��H �@ ��? ��A ��B ��I �NH ��H ��L �+M ��C �rF ��G �F ��D �DB �J �BL �N ��J ��N �
B ��F ��M ��J �-I ��? �$F ��N �J@ �I ��F ��A ��E ��E � #E >>&  �&  �+  L   R �+  $
D P �+  	��F     %D �S   S�N ��+  	�+  	  �+  �   L   L   f   f    uE  �:,  #` �I&   ֳ  �L   [M �L   ڰ  �b   tI ��+  �N x�2-  �1  �L    cnt �L   row  L   |H :  �N :  �J :  �A :  XD :   �O :  "{ 
�   (
N 9   0�  2-  8E C&  @�q  :,  Hڰ  b  hֳ  L   p 	0)  xK F,  �   U-  L     E-  &?K oU-  	��F     J  �-  L    q-  'a2i ��-  	 �F     J  �-  L    �-  &G ��-  	 �F     &�I ��-  	��F     J  �-  L    �-  &�B ��-  	��F     p: _   J7.  �:  �0 �; 9  �9 Q.  �- vi.  b x7.   u ~i.   "y�.  ;G z�  :�  {H  �: |U   : �C.  ;  �.  	�.  	  �.  �  �.  �.   	�  �6 %�.  	�.  	  �.  �  �  �.   	�.  ? */  /  �< *>/  �= ,�.   bD -�.   O (f/  enc *�   ȩ  +�   �C ->/  (�F  0�/  ah 21   �7 4�   �)o/ 5�    ).O 72-  )�M 9�/  )�E ;�   	f/  �J =�/  	r/  
g+  @.�  �H (6,0  I_ 8�"   �@ 9�  �@ :�/    7@ <80  	�/  $�E �\$  	��F     &�E �#/  	p�F     $   {0  L    k0  &L �#{0  	@�F     *�/  �	��F     +�? �,  ��C     
       �1  ,ϖ �&�  �	 �	 ,}W �&�  3	 /	 -�C     �o  .U	@�F     .T�T  +�G �	  p�C            �k1  /��  �%�/  U/�7 �%�.  T/n/ �%�.  Q +YL r	  0�C     �       �F2  ,��  r+�/  p	 l	 ,M9 s+�  �	 �	 ,�9 t+�.  	 �	 0Cp v*)  &	 	 1WD  �~�C     2�H  7�C       ��  {3I  �	 �	 3I  $	  	 4��  5'I  6i�C     �j  .T�T    +�C 	  ��C     �      �r3  ,�  !�  f	 Z	 ,ֳ  !�  �	 �	 ,x !�  [	 U	 ,�1  !H  �	 �	 7bdf �/  	 	 0��  �  L	 H	 8�U 	   0.a r3  �	 �	 0ȩ  �'  7	 %	 7bpp X   �		 �		 1�  f��C     9k�C     �o  ]3  .Us  6�C     �o  .Us0  	�  :�D �	  �3  ;ֳ  �&�  <req �&�  =��  ��  =�d  �%  =.O �2-  =�U �	  =��  ��   +�H �	  ��C     G       �^4  ,ֳ  ��  �		 �		 ,m ��  3
	 /
	 0.O �2-  n
	 l
	 6��C     �o  .T�T  +aI ]	   �C     �      �=D  ,^�  ]!.  �
	 �
	 ,�L ^!�  s	 O	 ,�  _!�  �	 �	 ,�[  `!�  :	 6	 ,\  a!4  w	 s	 0�U c	  �	 �	 =��  d�/  0ڰ  eb  �	 �	 0�  g2-  �	 �	 &Ũ h2&  ��~1�  �&�C     1WD  ���C     > �  �?  0Cp �*)  W	 =	 >��  �8  0�d  �%  o	 a	 0M; ��  	 	 0
6 �,�  ,	 	 0<v �9   ,	 	 ?�H  ��C      P�  �F6  3I  �	 �	 3I  	 	 4P�  5'I  6��C     �j  .Uv .T	F�F        @�H  ӣC      ӣC            ��6  3I  @	 >	 3I  n	 l	 AӣC            5'I  6�C     �j  .Uv .T	��F        @�H  �C      �C            :7  3I  �	 �	 3I  �	 �	 A�C            5'I  64�C     �j  .Uv .T	��F        @�H  Z�C      Z�C            %�7  3I  �	 �	 3I  	 	 AZ�C            5'I  6w�C     �j  .Uv .T	w�F        @�H  ��C      ��C            :.8  3I  9	 7	 3I  g	 e	 A��C            5'I  6̤C     �j  .Uv .T	��F        9��C     �o  F8  .QH 9��C     �o  p8  .T} 0$0&.Q~ 0$0& 9H�C     �o  �8  .T2.Q3 6$�C     �o  .T�;$.QN   B��C     �       9  7cur _$)  �	 �	 7n `L   �	 �	 6�C     �o  .Uw .T@.Q0.X0.Y��~  >��  �;  0o/ z*)  	 �	 0�7 z-*)  g	 c	 0�k  {s  �	 �	 >`�  �:  7s ��  		 	 >��  �9  &�� ��  ��6z�C     �o  .U	��F     .T0.Q��.R0  9��C     �o  �9  .U~ .Q��~ 9��C     �o  �9  .U~ .Q��~ 9��C     p  #:  .Uv .T	��F      9�C     p  H:  .Uv .T	��F      9 �C     p  g:  .T	4�F      91�C     p  �:  .Uv .T	��F      6F�C     p  .T	��F       >0�  �:  &�� ��  ��6�C     �o  .U	��F     .T0.Q��.R0  ?�H  ��C      ��  Q;  3I  A	 ?	 3I  o	 m	 4��  5'I  6��C     �j  .Uv .T	��F        2�H  §C       �  �3I  �	 �	 3I  �	 �	 4 �  5'I  6ѧC     �j  .Uv .T	��F         ?�H  y�C      ��  �<  3I  �	 �	 3I  U	 O	 4��  5'I  6��C     �j  .Uv .T	�F        @�H  ��C      ��C            ��<  3I  �	 �	 3I  �	 �	 A��C            5'I  6ǠC     �j  .Uv .T	k�F        ?�E  �C      ��  �Y?  3�E  �	 �	 4��  C�E  ��~D�E  g	 U	 D�E  (	 "	 D�E  s	 q	 D�E  �	 �	 CF  ��CF  ��DF  V	 P	 D$F  �	 �	 E�H  I�C      I�C     %       ��=  3I  	 	 3I  H	 F	 AI�C     %       5'I  6n�C     �j  .U| .T	<�F        E�H  }�C      }�C            �>  3I  o	 m	 FI  A}�C            5'I  6��C     �j  .U| .T	B�F        G�H  ��C       �  �e>  3I  �	 �	 FI  4 �  5'I  6��C     �j  .U| .T	N�F        G�H  ˡC      P�  ��>  3I  �	 �	 FI  4P�  5'I  6�C     �j  .U| .T	\�F        H0F  ��  J?  D1F  7	 3	 H<F  ��  .?  D=F  o	 m	 IJF  ��C     <       ?  DKF  �	 �	  6��C     p  .Q~   6j�C     p  .U} .Q��~  J�C     +p    9�C     �o  y?  .Uw .Q��~ 6�C     �o  .Uw .T .Q0.R1.X0.Y��~  ?�I  ��C      @�  x�C  3�I  �	 �	 3�I  �	 ~	 3�I  � 	 z 	 3�I  �!	 x!	 4@�  D�I  _"	 Q"	 D�I  #	 �"	 D�I  �$	 i$	 C�I  ��~KJ  �C     K
J  �C     ?tb  �C      ��  ��B  3�b  �%	 �%	 3�b  z&	 n&	 3�b  *'	 '	 3�b  �'	 �'	 4��  C�b  ��D�b  �(	 �(	 D�b  )	 �(	 D�b  �)	 �)	 D�b  �*	 �*	 D�b  ,+	 (+	 Dc  g+	 e+	 Dc  �+	 �+	 D!c  �+	 �+	 D.c  �,	 �,	 D;c  [-	 W-	 DHc  �-	 �-	 DUc  �.	 �.	 Cbc  ��Koc  �C     Hxc  ��  �A  Dyc  ~/	 z/	 6�C     �o  .U��~.T1.Q} .Rs .X .Y��~  9(�C     �o  �A  .U��~.T1.Q0.R
 .X0.Y��~ 9��C     7p  B  .U��~.T } ".Q��}}  9�C     Dp  (B  .U��~ LQ�C     [B  .U��~.Tv .Q��~.R��.X��~ L��C     �B  .Tv .Q��~.R��.X��~ 6�C     Pp  .U .Q}    ?3f  �C       ��  ��B  3Nf  �/	 �/	 3Af  �/	 �/	  @;I  �C      �C            	GC  3II   0	 �/	 A�C            5VI  5cI  5nI  5{I  6�C     �g  .Uv    9��C     p  lC  .Uv .Tx.Q��~ 9�C     �o  �C  .T1.Y��~ 9 �C     Dp  �C  .Uw  9�C     �e  �C  .U��~ 9"�C     Dp  �C  .Uw  65�C     Dp  .Uw .T    9:�C     \p  D  .U~ .T0 9�C     =D  (D  .Us  6ШC     =D  .Us   M^J B��C     �       ��E  ,�L B�  ,0	 $0	 0��  D�/  �0	 �0	 0ڰ  Eb  �0	 �0	 @;I  ��C       ��C     
       ME  3II  1	 1	 A��C     
       5VI  5cI  5nI  5{I  J�C     �g    9��C     Dp  E  .Uv  9�C     Dp  3E  .Uv  9-�C     Dp  KE  .Uv  9D�C     Dp  cE  .Uv  9X�C     Dp  {E  .Uv  9l�C     Dp  �E  .Uv  6��C     Dp  .Uv   N�I �	  [F  Obdf �"�/  #�U �	  #��  ��  #ڰ  �b  #�  �2-  #Cp �*)  #�y �[F  #h�  �kF  Pnn �@   Plen �#@   QRs �   QRsrc �  QRmm 0@       �  kF  L    @   {F  L    S E ��  ��C     �       �vG  T�N �#"  @1	 <1	 U9 �#�#  TVI_ �,0  }1	 y1	 V�@ ��/  �1	 �1	 Wmin ��  �1	 �1	 Wmax ��  32	 +2	 Wmid �!�  �2	 �2	 V�Y  ��  S3	 I3	 V�_ ��  �3	 �3	 X�  � �C     4 �  V�* ��  b4	 \4	   S�N [�   �C     {       �SH  T�N [#"  �4	 �4	 T�_ \#U  �4	 �4	 VI_ ^,0  )5	 %5	 V�@ _�/  d5	 b5	 Wmin `�  �5	 �5	 Wmax `�  �5	 �5	 Wmid `!�  46	 &6	 V�Y  a�  �6	 �6	 4��  V�* j�  (7	 "7	   YlO P �C            ��H  U�N P"  UVI_ R,0  s7	 q7	  SC @	  ��C             ��H  U�N @"  UU�h  A	  TVI_ C,0  �7	 �7	 V��  D�/  �7	 �7	  :PO b	*)  5I  ;�  b	'2-  ;}W c	'�  =\G e	5I   	@   Z�@ 	�I  ;�  	2-  =Cp 	*)  Ri 	L   =4x 	$)  =ڰ   	b   :�@ �	  J  ;^�  �".  ;NC �"b  ;E �"C&  ;�  �"J  =HI �L   Rp �J  =ڰ  �b  =�U �	  [�  	[WD  	 	2-  	8-  +�E N	  �C     �      �R  ,� N$�   �7	 �7	 ,�H O$L   Z8	 08	 ,HI P$L   :	 :	 ,D Q$f   f:	 L:	 ,`A R$f   �;	 ;	 &�H TL   ��}0�W UR   <	 �;	 Rp VJ  0�  W2-  !=	 =	 7s X�   �=	 �=	 0ڰ  Zb  (>	 >	 0�U [	  �>	 �>	 1�  t>�C     >��  �K  7i �@   �?	 �?	 0Cp �*)  �?	 �?	 9?�C     ip  �K  .U~ .T  6��C     up  .Tv .Q~ .R   B��C     L       �K  7bpp 0A  @	 @	 J��C     da   B%�C     �       �L  &oD MR  ��}9Q�C     �p  4L  .U��}.T	4�F      9d�C     3k  cL  .T	�F     .Q��}\�]  �Q 9��C     �p  �L  .U��}.T	4�F      6��C     3k  .T	�F     .Q��}\�]  �Q  @Kb  �C       �C            �&M  3]b  >@	 <@	 A�C            5hb  J*�C     \f    ?�a  ݳC       ��  �OM  3�a  c@	 a@	 4��  5�a  J�C     �f    @�a  ��C      ��C            ��M  3�a  �@	 �@	 A��C            5�a  J�C     �f    ?�^  .�C       ��  O  3�^  �@	 �@	 3�^  �@	 �@	 3�^  0A	 *A	 4��  D	_  }A	 yA	 C_  ��}C#_  ��}D0_  �A	 �A	 D=_  �A	 �A	 KJ_  ޵C     ]S_  ?3f  X�C      @�  �pN  3Nf  �B	 �B	 3Af  �B	 �B	  9��C     +p  �N  .Us  9��C     p  �N  .U��}.Ts .Q|  9��C     �c  �N  .U��}.T	{�F     .Q��}.R|  9޵C     �e  �N  .U��} 6��C     �e  .U��}   ?Kb  }�C       ��  )QO  3]b  �B	 �B	 4��  5hb  J��C     \f    @Kb  ��C      ��C            *�O  3]b  C	 C	 A��C            5hb  J��C     \f    @Kb  ��C      ��C            +P  3]b  AC	 ?C	 A��C            5hb  J��C     \f    J��C     m_  9
�C     p  5P  .U .T�.Q��} 9��C     �c  iP  .U}� .T	N�F     .Q�U.R�T 9��C     �c  �P  .U}� .T	N�F     .Q�U.R�T J�C     da  J&�C     da  9��C     �c  �P  .U| .T	N�F     .Q�U.R�T 9��C     no  Q  .U|  9��C     �n  Q  .Tt  9شC     Dp  2Q  .Uv  9�C     �o  `Q  .Uv .T1.Q0.X0.Y��} 9*�C     p  xQ  .T|  9a�C     �c  �Q  .U}� .T	N�F     .Q�U.R�T 9�C     �o  �Q  .Uv .TH.Q0.X0.Y��} 9^�C     p  �Q  .U .T(.Q��} 6��C     ip  .T   	�+  �   *R  L    +�J �	  ��C     $      ��V  ,� �)�   hC	 dC	 ,�H �)L   �C	 �C	 ,HI �)L   	D	 D	 ,D �)f   \D	 BD	 ,`A �)f   �E	 uE	 &�B �L   ��~0�W �R  �F	 �F	 7p �J  �G	 �G	 0}W ��   *I	 I	 0<v ��   �I	 �I	 &oD �R  ��~0�U �	  iJ	 MJ	 1�  G��C     @�H  #�C       #�C     !       �S  3I  �K	 �K	 3I  �K	 �K	 A#�C     !       5'I  6D�C     �j  .T	�F        @�H  Q�C       Q�C     !       8T  3I  �K	 �K	 3I  L	 L	 AQ�C     !       5'I  6r�C     �j  .T	�F        ?L^  ٮC       ��  2NU  3�^  8L	 0L	 3�^  �L	 �L	 3x^  M	 M	 3k^  �M	 �M	 3^^  �M	 �M	 4��  D�^  �N	 �N	 D�^  ;O	 !O	 D�^  VP	 BP	 D�^  *Q	 &Q	 2Q`  �C      �  #	3p`  iQ	 aQ	 3c`  �Q	 �Q	 4�  D}`  -R	 )R	 9"�C     �p  /U  .U| .T� 6?�C     �p  .U| .T�     9�C     3k  oU  .T| \�]  �Q 9o�C     �p  �U  .Uw .T	4�F      9��C     3k  �U  .T	�F     .Qw \�]  �Q 9��C     �p  �U  .Uw .T	4�F      9��C     3k  V  .T	�F     .Qw \�]  �Q 9��C     �c  FV  .U~ .T	N�F     .Q| .Rv  9��C     no  ^V  .U~  9��C     �n  vV  .Tw  9��C     3k  �V  \�]  �Q 6�C     3k  .T| .Qs \�]  �Q  +�A 	  ��C     I      �M]  ,� %�   gR	 cR	 ,�H %L   �R	 �R	 ,HI 	%L   ]S	 US	 ,D 
%f   �S	 �S	 ,`A %f   JV	 BV	 7c X   �V	 �V	 0�M X   1W	 -W	 7s �   �W	 �W	 7bp =  X	 
X	 7i L   �X	 �X	 &�H L   ��0)N !L   4Y	 ,Y	 0�W R  �Y	 �Y	 7p J  
\	 \	 0ȩ  $)  }\	 i\	 0�  2-  []	 K]	 0ڰ  b  ^	 ^	 &�U 	  ��1�  �o�C     1�E �p�C     B��C     >       �X  7sw �A  @^	 >^	 6��C     �o  .T@   >P�  �X  0nN �L   g^	 c^	 6p�C     �o  .U| .T1.Q0.X0.Y��  ?Kb  g�C       ��  ?$.Y  3]b  �^	 �^	 4��  5hb  J~�C     \f    ?�a  ?�C      ��  ~oY  3�a  �^	 �^	 4��  5�a  JV�C     �f    @Kb  �C       �C            W'�Y  3]b  �^	 �^	 A�C            5hb  J��C     \f    @Kb  ��C       ��C            d'!Z  3]b  #_	 !_	 A��C            5hb  J��C     \f    ?�a  �C        �  }bZ  3�a  J_	 F_	 4 �  5�a  J3�C     �f    9S�C     �c  �Z  .Uv� .T	N�F     .Qs .R  9h�C     m_  �Z  .U}  9�C     Dp  �Z  .U|  94�C     �o  �Z  .U| .T8.Q0.X0.Y�� 9ϽC     �p  [  .Q8.R	��C      9 �C     Dp  0[  .U|  9�C     �c  a[  .U} .T	N�F     .Qs .R  9/�C     no  y[  .U}  99�C     �n  �[  .Tt  9e�C     �o  �[  .U| .T1.Q0.X0.Y�� 9��C     p  �[  .Ts  9��C     �c  	\  .Uv� .T	N�F     .Qs .R  JվC     �a  9׿C     �c  H\  .Uv� .T	N�F     .Qs .R  9��C     �c  z\  .Uv� .T	N�F     .Qs .R  9�C     �c  �\  .Uv� .T	N�F     .Qs .R  Jg�C     da  Jx�C     da  9��C     �o  �\  .U| .T8.Y�� J��C     �a  9�C     �o  ]  .U| .T8.Y�� 9=�C     Dp  5]  .U|  6Y�C     �o  .T@   +�M �	  ІC            ��]  /� �"�   U/�H �"L   T/HI �"L   Q/D �"f   R/`A �"f   X :OI L	  L^  ;�  L%2-  ;}W M%�  ;<v N%�   ;HI O%L   =\G Q5I  =Cp R*)  Rfp R*)  =ڰ  Sb  =�U T	  [�  � :3G X   �^  ;�  �   ;�H  L   ;}W  I&  ;<v  I&  ;�   2-  =�8 X   Rsp �   Rep �   Rp *)   :�C �	  ]_  ;�  �-2-  ;E �-C&  ;HI �-L   Rlen �@   =}W �]_  =�q  �:,  =ڰ  �b  =�U �	  [�  [WD   �   m_  L   � +�C �	  P�C     �       �Q`  ,�  �$2-  �_	 �_	 ,�C �$�   �_	 �_	 ^len �$L   ,`	 $`	 7cp ��   �`	 �`	 0ڰ  �b  �`	 �`	 &�U �	  �L1�  �͋C     9��C     �o  6`  .T1.Y�L 6��C     p  .T} .Qv   :^D r*)  �`  ;}W r"�   ;�  s"2-  =\G u5I   :M @	  �`  ;}W @%�  ;��  A%X   ;�  B%2-  Rn D@   Rp E*)  =ڰ  Fb  =�U G	  [�  l +�J ,X   ��C            �da  _a ,  U_b -  T7c1 /$)  �`	 �`	 7c2 /$)  �`	 �`	  +i@ :  ��C     �       ��a  ^s �  +a	 !a	 7v :  �a	 �a	 7neg :  %b	 b	  :%E �A  �a  <s ��  Rv �A   +@@ �9   �C     �       �Kb  ^s ��  �b	 �b	 7v �9    c	 c	 7neg �9   �c	 �c	  :K �L   tb  <s ��  Rv �L    :�? 	  �c  ;^�  &.  ;L�  &�+  ;`A 	&f   <lno 
&�c  Rcb �+  =HI L   =�@ L   =z# X   =�8 X   =�N %X   =Vu  -   =�k -   Rend %-   =O�  *-   =fO 2-   Rbuf �   =ڰ  b  =�U 	  [�  �Q=v  P�    	L   :�B �	  ?d  ;�q  �#?d  ;7C �#�  ;� �#�   ;�H �#L   =9K �L   =]� �X   Rsp ��  Rend ��  Rep ��   =oI �Ed  =�U �	  1�  �	�C      	:,  �   Ud  L    :`M s�   �d  ;�q  s#?d  <c t#X   ;$D u#�c  Ri wL   Rj wL   Rdp x�   QRfp ��     Z�? X�d  ;�q  X#?d  <n Y#L   Ri [L   Ru [L    +�H 6	  ��C     �       ��e  ,�q  6$?d  3d	 +d	 ,� 7$L   �d	 �d	 &�U 9	  �\1�  R��C     4`�  0E >L   �d	 �d	 0zO ?L   (e	 e	 00E @L   �e	 �e	 0ڰ  Ab  �e	 �e	 6܊C     �o  .T8.Y�\   M�H (�C     6       �3f  ,�q  (!?d  Ef	 ?f	 0ڰ  *b  �f	 �f	 J%�C     Dp   Z�O \f  ;�q  !?d  ;ڰ   !b   `Kb  ��C     y       ��f  3]b  �f	 �f	 Dhb  g	 g	  `�a  p�C     g       ��f  3�a  sg	 mg	 D�a  �g	 �g	  `x3  ��C     �       ��g  3�3  *h	 $h	 3�3  |h	 vh	 D�3  �h	 �h	 D�3  i	 i	 D�3  Di	 @i	 a�3  D�3  �i	 ~i	 bx3  P�C            3�3  �i	 �i	 3�3  %j	 !j	 AP�C            5�3  5�3  5�3  5�3  5�3  -W�C     �3  .U�U.T0    `;I  ��C     @      ��i  3II  dj	 ^j	 DVI  �j	 �j	 DcI  �j	 �j	 DnI  l	 l	 D{I  �l	 �l	 9��C     Dp  !h  .Uv  9��C     �p  9h  .Tv  9ɍC     Dp  Qh  .Uv  9�C     Dp  ih  .Uv  97�C     Dp  �h  .Uv  9[�C     Dp  �h  .Uv  9��C     Dp  �h  .Uv  9��C     Dp  �h  .Uv  9ԎC     Dp  �h  .Uv  9�C     Dp  �h  .Uv  9�C     Dp  i  .Uv  9�C     Dp  )i  .Uv  93�C     �p  Hi  .Us�.Tv  9m�C     Dp  `i  .Uv  9��C     Dp  xi  .Uv  6��C     Dp  .Uv .T|   `�c  ��C     G      ��j  3�c  �l	 �l	 3�c  Om	 Km	 3�c  �m	 �m	 3�c  n	 n	 5�c  5�c  5�c  5�c  5d  5d  a d   c�c  ��  3�c  an	 Yn	 3�c  �n	 �n	 3�c  ho	 `o	 3�c  �o	 �o	 4��  D�c  9p	 1p	 D�c  �p	 �p	 D�c  Fq	 (q	 D�c  }r	 wr	 Dd  �r	 �r	 Cd  ��D d  �s	 �s	 K-d  ~�C     90�C     �d  �j  .U|  6L�C     �d  .U|     `�H  �C     4       �3k  3I  �t	 zt	 3I  �t	 �t	 D'I  Ou	 Ku	 6�C     �p  .U�T  `�]  �C           ��n  3�]  �u	 �u	 3�]  Xv	 Fv	 3�]  "w	 w	 3�]  �w	 �w	 D^  �w	 �w	 D^  �x	 �x	 D^  �x	 �x	 D(^  �y	 �y	 C5^  ��KB^  �C     @Kb  ��C      ��C            s,l  3]b  �y	 �y	 A��C            5hb  6��C     \f  .U|    @Kb  ЗC      ЗC            ��l  3]b  z	 z	 AЗC            5hb  6�C     \f  .U|    ?�`  0�C      �  ��m  3�`  9z	 5z	 3�`  uz	 qz	 3�`  �z	 �z	 4�  D�`  �z	 �z	 D�`  @{	 <{	 D�`  {{	 w{	 C�`  ��K�`  O�C     9J�C     �p  .m  .Uv .T~  9�C     �o  Rm  .U .TH.Y�� 94�C     +p  jm  .Uv  9W�C     �o  �m  .U .T1.Q0.R��.X0.Y�� 9}�C     p  �m  .Tv .Q�� 6��C     up  .Q~ .R    9%�C     �p  �m  .Uv  9��C     �p  n  .Uv .T~  9��C     Dp  *n  .U}  9ؖC     �o  On  .U} .T| .Q�� 9)�C     �o  ln  .U} .TH 9��C     �o  �n  .U} .T| .Q�� 9�C     up  �n  .R}  9(�C     �a  �n  .U|  9�C     �a  �n  .U|  6j�C     �p  .Uv .T~   `Ud  �C     �       �no  dgd  Udd  TD�d  �{	 �{	 D�d  |	 |	 D�d  U|	 S|	 etd   b�d  �C     E       D�d  z|	 x|	   `�d  p�C     I       ��o  d�d  U5�d  5�d  e�d   fF>  F>  kf[l  [l  
�fmY  mY  
�ff  f  
�fe  e  	�g�I  �I  �f2n  2n  
f=T  =T  ]g�  �  hBY  8Y   g�`  �`  vgNe  Ne  2f�h  �h  �g�s  �s  �gn  n  fM  M  �g2A  2A  `gV@  V@  ngIM IM ggt  t  zg�  �  XgTf  Tf  h �.  �S  &  �^ �:  ��C     W�      � ,  i   �@   �  int G   �  S   �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < 	�   �  �   �  8"a   
+  K  	�   
%  L  
�  M  '  �M  ?  -   O  @    ��  �[  ;  �s  �n  �  n  s&  G   �  S   �  )  A"�  	�  �   ��  �  �_    ��  ��  <h �  �I  �5   �  X�  	�  _     �  -    �   m  	%  5  �  _    f  �A  	G  _   e  �  -   -   _    J   �"q  	w  �  PH  Ǟ  Jt   ֳ  K@   pos L@     N8  /[  O8   �K PD  (�R Q�  0ڰ  S�  8O�  Tt  @��  Ut  H �  �8  <v �-   ��  �_    �  �  ""  �P  	V  @   t  e  @   t  @    	z  �  z  �   �  	�  �  e   v  :-   �  L�  x N�   y O�   �  Q�  �  ~   w'  
  y�   �!  y�  �   z�  H  z�   "  |�  N`  S   �|  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} S    5�  S   `�  	G   _| 
t  
!  n  ?   z  2   z  B  _     �  |  �  �  (Qp     S[   0�  T[  N5  Vp  �   W�   H� Xv  �1  ZG     	�  	[  �  \  	�  �  S   ��  �!   �   pmoc�  stibu!  ltuo�  tolp :  ��  �8  5"�  	�  �$  �4  S)  x U[   len Vn  e� Wz   �#  Y�  )  �%  {H  	N  h  G   G   h  _    	6  �#  �{  	�  G   �  G   G   _    �.  ��  	�  �  G   G   _    �8  `�O  .   O   �; U  �1  G   �5  ;  �+  ;   `(  n  (�/  �  0�  _   8*  '  @ 	  	[  u(  
�  \  �2  ({  	�  G   �  _   �   	�  �3  ;�  	�  �  �   v)  ]�  	�  �  �  t  @    �3  y�  	�  G     �  @   _    H7  �  	   G   4  �  4   	i  51  0��  y2  ��   � �n   ��  *
 ��  / �   $ ��  ( 2$  �:  -4  lz  +  ��  �  $8  �z  �  	�  Ab  ��    ��   �  {"  �[  !  �n  		  \   �G   �  �S   &	  }  �-   )$  �@   �   -   c,  +G   \	  C*  6_   +D  C4    :   ��	  xx �O	   xy �O	  yx �O	  yy �O	   5  ��	  �	  8  �
  ��  ��   ��  �	   $  ��	  c   �"
  	(
  3
  _    �  �^
  Kl  �_    �  �
   s  �3
  �"  $x
  	~
  �   +�
  �� -k
   �W .k
  Kl  /_    %  D�
  uR Fk
   �
 Gk
   }  I�
  S   %�2  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<�  5�  >�   ��  ?�  �"  A�  �"  B�  i!  C�   %!  E�  (2!  F�  0�  G�  8   I2  �"   s  ��  u�   5�  v�  ֳ  x�  !  z�  m  {�   v  }�  J  �#-  	3  �!  �}�  ڰ  �   {3  �	  S0  �	  �/  �	  �1  �&	  �1  �
%   Y/  ��
   �*  ��  ( �)  ��  0 +:  �%  8 <8  �*%  X �*  �	  � �3  �"�  	  �(  �=  Oe ��$   �-  �   ڰ  ��   U  �"J  	P  �  8�  ah !�$   Oe "s   U1  #�
   ;+  $�  0 i(  �$�  	�  l;  ��  ah ��$   Oe �%  y2  ��   {:  ��  (�� ��  h/ �  p�� ��  x T   � (  	.  _  ��  �!  7	   �  7	  �  7	    7	  �  7	   �U q  (�  q  03"  	  8�  w  @`  !	  Hd  "}  P�@  $^
  X�;  )'  h�   +		  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6I  �ֳ  7�  ��� 8�  �K <=  �ڰ  =�  �^�  >e  �U  @�
  �t  B^
  �k  C_   ��L  E�  � "   �  	  1  XmI  ��  o   �@  p^
  �e q[  �L  r�  P @  $%V  	\    0\�  �-  ^    ��  _  �W `I  x a&	  �@  b^
   �e d�  0�"  eO	  pi"  fO	  x� g�  ���  i�  �.a k�  ��  l	  �J  m	  �Mj  o|  ��  q&	  ��  rh  � M  t_     Z  u-    _"  w�   (   x�   Ud z_     �L  |�  ( �!  F#�  	�  Z!  A   ��  C   T D�  �!  E		  "  F		   S  S   ��  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �     �C  H�  0  `)�  	�  �"  �eq  �1  g�	   H+  h�   x+  i	  0��  k!!  8�)  n#�"  h�'  q�  p��  rz  t�*  y	  x 	�  	  	�  �S  I.  �  �)�  	�  �!  H��  $  �_    7:  �q  s4  �[   b  8H[  !  J		   m  K		  A� MO	  �� NO	  �  P�  
  Q�   ��  R�  (�  S�  0 �  U�  x   �$u  	{  �!  0'�  ad  )	   �1  *		  &D  +	  2B  ,	  x� -�	     �)�  	�  �"  P�N  ��  ��   �1  �&	  �&  ��  �3  ��	  ]7  ��  0�7  �_   @�1  �z  H P6  y  tag C	   Kl  n	   �6  	N  	y  �5  S   
�  i7   �&  9  F9  8%  �*   �,  
�  ./   6
&  b 8
�   5�  9
7	  ��  :
7	  5  ;
&	  Q(  <
&	    -  I
(3  	�  �8  S   �q  �:   4,  �6  $  �/  l9   �2  �9  �\  ��  b<  �&	   1S �&	  p ��   	�  �  p  �~  �#  �n	  �'  ��  	�  \	  �  �   �2  �  	    �   l/  �#  	)  �  =  �  =   	�   ;)  H��  �#  �C	   :  �7	  �5  ��  F1  �O	  ,8  �O	   2*  �U  (�*  ��  0`1  ��  8��  �  @ 	�  �-  �C  �  d)  s�  	�  \	  �  _    9  F#  �  �$  @J�  �#  L7	   y2  M�  W� O�  �� P  �,  Qx   M4  R#  (�;  SP  0�*  T�  8 c/  X!�  	�  �-  (q�  �-  s    Oe t�  ��  u�  � v�   	  �/  )�  	�  \	    �  I   g%  .  	  #  �   �.  1/  	5  J  �  J  �   	�	  73  6\  	b  r  �  r   	'  �8  :�  	�  \	  �  �  �   "3  >�  $)  Y�  	�  \	  �  �  I  q  �   �6  _�  	�  \	  
  �  I  J  �   �3  f  	  1  �  I  r   ;0  l=  	C  \	  \  �  C	  n	   �&  x��  ah � �   y2  � �  H�8  � �  P�8  � �  X�'  � 
  `� � 1  h�9  � �  p 	�  �.  �\  "9  H2&  Mj  4|   H5  5p  (�)  6p  0�  7&	  8�  8h  @ �0  :�  T%  �=�  ڰ  ?�   �0  @&	  q5  A&	  L)  B&	  )  C�  Ǟ  E&  �  F&  `Ud H_   � X+  J�  	2  1  �  	�  \	  �  e    	  	  �   �&  &�  	       �1  *  	  \	  -  �   �6  -9  	?  J  �   w-  1V  	\  \	  k  I   �;  4w  	}  �  I   =;  8�  	�  \	  �  �  &   B$  <�  	�  \	  �  �  C	   2  @�  	�  \	    I  �  &	  z   7  G  	  \	  4    &	  &	  p   q8  N@  	F  \	  Z    e   )2  Sf  	l  \	  �    &	  &	  z  �   	O	  k.  ��s   ah ��   #,  �7	  H�4  �7	  P,;  �7	  XEY ��  `/q ��  hZ)  �  p�#  �-  x'0  �J  �.  �k  ���  ��  �� �  �`9  �4  ���  �Z  �5  ��  �U#  ��  � �2  �   	�  8S  ��   �d  �=   �W  �U   C  ��   �   �&  0�!!  y%  �n	   �/  �n	  �'  �n	  �6  �n	  �+  �n	   �6  �n	  ( �7  ��   *  V':!  	@!  �0  �*   u�!  |#  w7	   �#  x7	  � y7	  C4  z7	   �&  |E!  �'  ��!  	�!  \	  �!  .!  &	  �!   	
  �9  ��!  	�!  �!  .!  �!   A2  ��!  	�!  \	  "  .!  &	  �  "   	�!  8(  U"  ��  )�!   $�  )�!  �-  )�!   )  "  U"  3  <�"  �� >%�"   ��  ?%.!   	b"  #  Ag"  	�"  �U  �,�"  	�"  �B  ��"  �� ��   Oe ��"   fP  �,�"  	�#  4I  P��#  ֳ  �C	   �� ��#  �q ��#  R` ��#  �W �$   P �#-$  (�U  �#]$  0�v  �#�$  8�v  �#�$  @�J  �#�$  H �"  ��  ��"  wq  ��#  	�#  \	  �#  �"  n	   �J  ��#  	�#  �#  �"   �\  ��#  	�#  &	  $  �"  �   \  �$  	$  &	  '$  �"  '$   	�  U  �9$  	?$  &	  ]$  �"  �"  �  �   �O  �i$  	o$  	  �$  �"  �  �   �n  ��$  	�$  '$  �$  �"  �   ;O  ��$  	�$  '$  �$  �"  �  �   -k  ��$  *�  ��"  	�  �(  �  	�  �  %  @    �  *%  @    �  :%  @    	@%  =  O%     	U%  \	  s%    &	  n	  &	   	y%  &	  �%    �   !H'  �%�  <  S   9&  �?   Mm  2a  �=  	2r  �u  0@  �>  gd  �e  Lo  s  �Y  �^  �f  �l  E  �M   _c  VN&  <v X�   ֳ  Y�  �  Z		   yK  \&  N&  �I  `UJ'  Q  WO	   �g  XO	  �;  Z7	  �U  [7	  �B ]		   �o  ^		  "Y  `J'  (+I  aJ'  8
  c�  H�!  d�  J�   e�  LH  f�  N�`  h		  P�X  i		  RO  k�  T,G  l�  V�t  m�  X C	  Z'  @    I  o_&  �g  8�D(  ��  �O	   )r  ��  dS  ��  
�B  ��  �P  �		  �p  ��  �K  ��  =  ��  me  ��  +^  ��  �]  ��  �u  �D(  
h  ��  $^K  �		  &tR  �_   (%?  �_   0 �  T(  @    �]  �f'  �S  8?O)  ��  AO	   )r  B�  dS  C�  
�B  D�  �A  F		  �n  H�  �n  I�  �W  J�  me  K�  +^  L�  �]  M�  �u  OD(  
h  Q�  $�V  R		  &tR  X_   (%?  Y_   0 �u  [`(  JW  �x�+  ��  z		   =  {�  �<  |		  tB  }		  �k  ~		  �m  �  
�D  ��  gJ  ��  !X  ��  �S  ��  5f  ��  ?X  ��  �a  ��  �_  ��  �a  ��  Gf  ��  �=  ��+   �E  �C	  0F  �C	  8�A  �C	  @F  �C	  H�E  ��+  P5D  �		  TH  �		  V#l  �		  X$r  ��  Z_S  ��  \'N  ��  ^?_  �		  `L  �		  b�O  �C	  h�O  �C	  p~e  ��  x [  ��  z0m  �		  |�M  �		  ~rM  �		  �]  �		  ��g  �		  � �  �+  @   	 �  �+  @    �X  �\)  kE  @�G,  �^  �O	   zp  �O	  dv  ��  �i  ��  �<  �C	  �F  �C	   �D  �C	  (�p  �C	  03X  �C	  8 �b  ��+  K_  @�5-  ��  �O	   �J  �C	  �<  �		  e  �		  $� �		  dk  �		  ![  �		  L^  �		  �`  �5-  yN  �E-  ,ma  �U-  4�Z  ��  :�q  ��  ;r  ��  <�u  ��  = �  E-  @    �  U-  @    �  e-  @    	l  �T,  �M  (8S.  ��  :O	   �T  ;		  �P  <		  
�K  =		  B  >		  ^  ?		  �g  @		  /o  A		  %B  B		  �O  C		  �<  D		  �]  E		  *w  F		  dW  G		   �F  H		  " e=  Jr-  m<  S   m�.  nA   ZY  TE  �U  �R  {H  b  �c   �`  y`.  |[  O�.  �� Q�   �\  R�  red S�  q  T�   �[  V�.  �?  (�N/  `a  �		   �L  �N/  r  �N/  &W  �		  �F  �N/    		  Ik  ��.  	7	  ��   L�/  }W  Nq   ��   O7	  ��   P7	   ��   Rf/  8y  h l�/  �~   n&	   ��   o&	  �~   p�/   �/  �/  @    `�   r�/  ,�  0 �T0  }W  �q   ��   �O	  def  �O	  ��   �O	  tag  �C	   cy   �&	  ( ˣ   ��/  ��   ��0  Ԛ   ��   cy   �&	  �}   �&	   	�   �`0  U�    ��0  �~   �&	   ��   �&	  ˧   �&	  �~   ��0  i{   ��0   	T0  	�0  �   ��0  >i   !JJ1  tag !LC	   ��  !MO	  /� !N7	  �f  !OJ1   	C	  2\  !Q1  �k !l�1  �v  !nC	   �R  !o		  ei !p		  
�f !q		  j !r		  �  !tC	   �` !v\1  ad !v�1  	\1  G   !�2  Tag !�C	   g  !�C	  �=  !�C	  Ja  !�C	   b !��1  mn  !�02  	�1  �v   !��2  �T  !�		   �Y  !�		  D  !�		  S  !�		  E]  !�		  ;C  !�C	  �: !��   �[  !�62  M  !��2  	62  DQ  !�2  E]  !		   ;C  !C	  �: !�   �i  !�2  hh  !3  	�2  >M  0!.�3  ��  !0		   �Z  !1&	  vv  !2&	  �r !3�3  =P  !4&	  �Q  !5�3   ^�  !6e  ( 	�2  	�2  �p  !83  �a !8�3  	3  CE  !Y�3  �B  ![		   b  !\		   Pq  !^�3  	�3  �m  !x*4  ��  !z		   �R  !{		  Up  !|�3   �=  !~�3  �i  !��4  ��  !�		   5�  !�		  �"  !��  �"  !��  i!  !�		  %!  !��  
2!  !��  �  !�		   W  !�74  l !��4  	74  �U  !5  �  !�   
  ! �  Sd  !!�  �Q  !"�  �G  !#�  �v  !$�  �=  !%�  sD  !&�  �\  !'�  �X  !(�  	`N  !)5  
 �  �5  @    �T  !+�4  			  >t  !�6  �>  !��5   � !��5  !  !��  m  !��  �[  !��  SX  !��   �<  !�6  	�5  x@  !"_6  �  !$		   �`  !%		  TL  !&�5  �o !'_6   	e6  	�  �h  !)6  qo !)�6  	6  �Z  !<�6  �  !>		   �f  !?e6   fR  !A�6  |o !A�6  	�6  "!Z�6  #j !\k6  #�Y !]�6   ms   !V&7  �  !X�   �r !_�6   J  !a�6  rk !a@7  	�6  �t  !r!S7  	Y7  U<  �c  (!��7  �B !��   �c  !��  �y !��  �Y  !�C	  cC  !�&	   �  !��  $ 	\  !�^7  �s !��7  	^7   L  !� �7  	�7  �i  �!��<  ah !��   �u  !�P1  � �v  !�C	   �R  !�		    o  !�$2  ( �& !�Z'  0 �Q  !�T(  � @  !�S.  � 5�  !��  � <  !�O)  � �`  !�		  0 �a  !��3  8$os2 !��+  h F�  !�G,  � j  !��  0  M  !�C	  8 w_ !��>  @ �>  !��>  H �A  !�?  P ^Z  !��>  X �f  !��>  ` KT  !��>  h �i  !�_   p Q  !�_   x$mm !�_   �$var !�_   � g  !�_   � �Y !�*4  � Fq !�e-  � jQ  !�C	  � nQ  !�6  � m  !&7  � �P  !T/   @  !		  @ B  !c?  H �u  !�  P �u  !�.  Q �;  !C	  X zQ  !�  ` FN  !C	  h T  !�  p !u  !C	  x$cvt !i?  � 2i  !�<  � )  !)^
  � �  !+=  � �j  !-C	  � :>  !.C	  � �_  !0�  � S?  !3�  � E�  !4F7  � �W  !6�  � XA  !8=  � 	K  !9&	  � �c  !?C	  � ][  !@C	  � �J  !BC	  � '<  !C�  � 	Z  !E�    �q  !FC	   �G  !G&	   �T  !HC	   �a  !I�    �\  !K�  ( �u  !LC	  0 o  !MV?  8 ^C  !N&	  < :W  !Oo?  @ _  !Q�  H �@  !RC	  P >  !S&	  X }?  !T�  \ m?  !U�  `$bdf !X�7  h �k  !\C	  � �Z  !]C	  � Pl  !hC	  � (a  !iC	  � i !m_   � �d !n_   � �Q  !��  �g  !�"�<  	�<  �t  x!��>  ��  !��7   ֳ  !�C@  ȩ  !�I  �m  !��  �1  !�C	   x !�&	  (^�  !�e  0��  !�	  8   !��  <�;  !�'  @�C  !�	  `� !�	  d"f !�	  h�I  !��  lpp1 !��  ppp2 !��  �Ǟ  !�@  ��y  !�@  � BJ  !�+@   �<  !��   bL  !�C	    Ud !�_   ( �W  !�	  0 r�  !�	  4$pp3 !��  8$pp4 !��  H O�  !��  X ��  !��  ` �k  !��
  h �^  !�>  	�>  \	  �>  �7  C	  e  J1   �D  !*�>  	�>  \	  �>  �<  &	  C	  &	   �b  !A�>  	�>  \	  ?  �<   SQ  !Q?  	?  $?  �<   �=  S   !TV?  �G   �v  k_  <L  ok   �`  !_$?  	�.  	z  	&	  �j  @!�@  ڰ  !��   �0  !�		  q5  !��  
0�  !�		     !��  org !�p  cur !�p  " !�p   �   !��  (H� !��5  0�>  !�		  8 ,L  !�u?  @\  !�'8@  	>@  �r  �d  !� P@  	V@  �a  �p X"-A  � "/C	   9g "0C	  ��  "1C	  �R  "2		  Y  "3		  �X "4C	   ��  "5		  (@g "6		  *f] "7C	  0ER "8C	  8�m "9C	  @ W ":C	  H�^ ";C	  P �] "=[@  �g 0"^zA  Tag "`C	   �=  "aC	  fo "bC	  �m "cC	  g  "dC	   �q "fC	  ( �k "h�A  	A  <e  #I�A  	�A  \	  �A  e  �7  	  	  �   l  #s�A  Z  #��A  	�A  �A  �7   -H  #��A  	�A  \	  B  �7  C	  7	  �  J1   �e  #2,B  	2B  \	  _B  �7  C	  &	  &	  e  _B  eB   	�  	�4  �h  #SxB  	~B  \	  �B  �7  &  J1   �^  #p�B  	�B  \	  �B  �7  C	  �B   	[  eN  #��B  	�B  \	  �B  �7  &	  �B   	q  Ub  #�C  	C  \	  'C  �7  e  �   #K  #�4C  	:C  YC  �7  �  &	  YC  �5   	�  3l  #�lC  	rC  \	  �C  �7  &	   �d  #	�C  	�C  �  �C  �7  &	  o?  o?  �C   	�  �J  #0�C  	�C  \	  �C  �7  &	  I  I   CZ  #N D  	D  \	  D  �7  		  �B   :=  #p,D  	2D  �  PD  �7  		  PD  PD   		  �Z  #�cD  	iD  \	  }D  �7  e   �^  #��A  GK  #��D  	�D  	  �D  �7  &	  &	   N=  0#��F  w_ #�"�>   EY #�"�A  �e #�"�A  /q #�"�A  ��  #�"   ob #�"�A  (pR #�"VD  0�^ #�"�B  8D_ #�"VD  @x` #�"VD  HPr #�"VD  P1s #�"VD  X�k #�"VD  `�S #�"}D  h�O #�"VD  p�Y #�"VD  xAq #�"VD  ��b #�"VD  �ar #�"B  ��[  #�"�B  � Q  #�"}D  �� #�"�D  �X #�"VD  ��U #�"�B  �`H  #�"VD  ��W  #�"}D  ��n #�"kB  ��T #�"�B  �zi # "VD  ��d #"VD  ��Q #"}D  ��] #"}D  � B  #"_C    UU #"�C   �p  #"�C   �[ #"'C   ]o #
"�C    4P #"D  ( sh  #�D  �F  AD  #�F  	�F  
�7  $�  S   %�TI  �U  2Z Hk k gp q �P R dY t[ 	;b 
Y $n �c �] �d �_ �U �l �r �i PR  �O !�\ "�g #Rh $�P %�R &�e '�j (,m 0�o 1�h @�n A9o Q�Z R�[ S�T T�c U�Y V'^ W�p X�g `9] aQl b�\ c�l p�d ��f ��U �>V ��d �/f �XQ ��O �r^ �]T �e �_e ��Q ��f �` ��_ ��b ��k �X[ ��m �"V ��r ��s ��l ��s �jl ��q ��S ��i �;s �Gj ��X �+b �nn �6U ��n �j ��h ��_ ��V ��T ��R �oq ��Q �W ��X ��j � p: S   &JI  �:  �0 �; 9  �9 &QTI  �- &v�I  b &xI   u &~�I   %&y�I  ;G &z=  :�  &{z  �: &|�   : &��I  ; ' �I  	�I  \	  J    J  J   	=  �6 '%(J  	.J  \	  GJ    =  GJ   	�I  ? '*^J  MJ  �< '*�J  �= ',�I   bD '-J   �u  (*.�J  	�J  �R  X(X�J  �Y  (Z3   Ǟ  (\�  @��  (]�  HgY  (^K  P�U (_\	  T �J  �G  S   (FK  X   �t  *u   �k  (L�J  �r (a�J  V^  )9QK  �L  );C	   ��  )<7	   �`  )>)K  {V  )BiK  	oK  \	  �K  �  �K   	QK  ��  )F�K  �K  �N  )F�K  �  )H]K    LQ (*"�K  I_ *$�#   Kl  *%�  �1  *&	    W *(�K  Q *(L  	�K  Ss **,L  L  L  	fL  �T h*1fL  Oe *3�$   ��  *4&	  P�r *5kL  X�  *6]K  ` $L  �c *.wL  	}L  \	  �L  �  �J   %U *8$L  �L  p `*^�L  a *`K   �  *a&	  X �m *c�L  �L  Za *c�L  	�L  
.k *j-�L  �A  +&O%  �V  +,s%  b�  +0"M  M  tG  +0JM  ]o +2!�L   �  +3!M   �d  ,):%  ��  ,,gM  VM  `p  ,,�M  g ,.JM    �g  -(�M  	�M  \	  �M    C	  7	  �  J1   3?  -2�M  	�M  _   �M    �.   �K  -:�M  	�M  \	  N    &	  J1  J1  J1   �o -A#N  N  6q  -AXN  �s  -C�M   I  -D�M  Y -E�M   ��  .'dN  	jN  \	  ~N    ~N   	�/  �z  .+�N  	�N  \	  �N    �N   	�N  	�0  9~  ./�N  	�N  \	  �N    &	  `/   "�  .6�N  	�N  \	  O    &	  �   ��  .=�N  �  .B�N  ��  .G0O  	6O  \	  JO    &	   Ӏ  .K�N  ݓ  .PbO  	hO  \	  �O    o?  �O  �O  �N   	�  `�  .W�  ��  .Z�N  3�  ._�O  	�O  \	  �O    o?  �   y  `.d~P  �~  .f"XN   -�  .g"�N  g�  .h"O  ��  .i"JO  7�  .j"�N   Y�  .k"�N  (�  .l"O  0&�  .m"$O  8U�  .n"�O  @A�  .o"�O  HY�  .rVO  P��  .s�O  X �O  g�  .d�P  	~P  &BW �N  	�G     &�p �M  	�G     �  �P  @    �P  &] ��P  	pG     �a ��P  	�P  G   Q  G    �   Q  @    Q  '�h Q  	`G     'o BbM  	XG     '�n L�K  	PG     '�e yYJ  	@G     �   �Q  @    Q  'YZ ��Q  	�G     '@P ��F  	�G     (G  	@G     N�  /#�Q  	�Q  �  �Q  =   :�  /)R  	R  =  R  &	   8�  //R  �  /5JR  V /7�   x /8&	   ��  /:"R  ��  /=$bR  	hR  ��  (/?�R  I_ /A�#   J�  /B&	  �m /C�R    	JR  f�  /M�R  	�R  =  �R  n	  &	   �  /U�R  	�R  �R  n	  =   ��  /Y�R  	�R  \	  %S  �  VR  &	  �R  �R  n	   r�  /a1S  	7S  &	  KS  VR  �   ��  /eWS  	]S  �  qS  VR  '$   ��  @/i�S  4v /k �Q   �y /m �R  v /n %S  Ty /o KS  hn /q �Q   S�  /r R  (��  /s �S  0��  /t �S  8 qS  q�  /i�S  	�S  	u  �  0'T  	T  \	  /T    &	  PD   ¦  0,T  ۧ  01T  r�  08T  ��  0=T  ��  0BT  ʍ  0GT  �  0N�  ��  @0Q�T  H�  0ST   ��  0T/T  -�  0U;T  ��  0WGT  ݖ  0XST   p�  0Y_T  (#�  0ZkT  0��  0\wT  8 �T  ��  0Q
U  	�T  
S }U  	"U  q  6U  �2  �   )�R ��L  	�G     * [ T�L  	@G     nW P��U  I_ ��K   �_ ��  (�P �&	  ,�  �&	  0py  �&	  4e_ �&	  8�\ �&	  <z�  �	  @�l ��  H �U ��U  	cU  *D^ �L  	�G     *P ��L  	@G     *�j ��L  	�G     *h ��L  	@G     �q P��V  I_ ��K   ��  ��  (�_ �C	  0�P �&	  8�S �C	  @1X �C	  H uV ��V  	_V  *�a �	�L  	�G     VY P
OW  I_ 
�K   ��  
�  (�_ 
C	  0�P  
&	  8�S !
C	  @1X "
C	  H ZW $
\W  	�V  *�_ *�L  	@G     �o H��W  I_ ��K   qr �C	  (>n ��  0�s �'$  8ڰ  ��  @ dW ��W  	yW  *QS $�L  	�G     +�L  �	@G     L  X  @   	 X  '�n �X  	�G     �a 0lX  gid 2		   �r 3		  b<  4		   �p 67X  �h (9�X  ��  ;		   �X <		  b<  =		  �X ?�  �]  @�  �B C_   �@  DC	    �U FxX  [d (0IY  ��  2		   \p 3		  `p 5�  Zq 6�  �B :_   �@  ;C	    �O =�X  �P X�Z  ��  ��7   ^�  �e  .a �_B  �e ��4  �` ��   1T ��  !�] ��  "Pl  �C	  ((a  �C	  0[f �C	  8p �C	  @ [ ��  Hr ��  P }Z �UY  �s �4Z  	UY  �Y �GZ  	MZ  \	  uZ  'Z  �  �  	  	  &	   ,Yr :\	  pqD           �N_  -��  :1�7  �|	 �|	 -m ;1C	  }	 }	 -x <1&	  ~}	 n}	 -�1  =1&	  9~	 /~	 -^�  >1e  �~	 �~	 .map ?1_B  �	 �	 /�e @1eB  � 0�U B\	  u�	 ]�	 1�sD           f\  'LM JN_  ��~2Qm  �sD      �sD     �       M1\  3�m  q�	 o�	 3}m  ��	 ��	 3pm  	�	 �	 3cm  .�	 ,�	 4�sD     �       5�m  \�	 T�	 5�m  ��	 ��	 6�m  �tD     7�m  ItD     S       \  5�m  �	 �	  8�sD     �, 9U|    8�tD     d`  9U��~9T} 9Q09R09X09Y~ F%1  :�
 ]  '�[ r�  ��~0�-  s   ��	 ��	 ;�tD     �, �\  9U��~ ;uD     �, �\  9U| 9T 9Q��~9R1 ;uD     �, �\  9U| 9T��~ <duD     �,  =^_  �qD      P
 ]3�_  ��	 �	 3�_  �	 �	 3�_  M�	 C�	 3�_  τ	 ��	 3�_  o�	 g�	 3}_  х	 ˅	 3p_  7�	 +�	 >P
 5�_  ��	 ��	 5�_  χ	 Ň	 5�_  B�	 >�	 ?�_  ?�_  5`  ��	 x�	 5`  �	 ܈	 5&`  ��	 ��	 53`  ��	 ��	 6>`  sD     ;"rD     �, ^  9U|  ;9rD     �, #^  9U| 9T8 ;KrD     �, ;^  9U|  ;VrD     �, S^  9U|  ;arD     �, k^  9U|  ;�rD     �, �^  9U|  ;�rD     �, �^  9U| 9T ���� ;�rD     �, �^  9U|  ;�rD     �, �^  9U|  ;�rD     �, �^  9U|  ;sD     �, _  9U|  ;sD     �, _  9U|  ;XsD     �, 7_  9U|  8�sD     �, 9U|     Z  ^_  @     @q] �\	  d`  A��  �1�7  Am �1C	  Ax �1&	  A^�  �1e  Bmap �1_B  A�e �1eB  A��  �1�  C9j �&	  C"	 �&	  C� �+&	  CdU �	  CrU �	  C�W ��  C�V �	  C�U �\	  Dp ��  E)f �FC�j )�  C� *		    ,-h �\	  �D     (      �je  -LM �/'Z  0�	 �	 -x �/&	  ,�	 �	 -ϋ �/	  =�	 /�	 -= �/	  �	 ؍	 -�  �/&	  ��	 ��	 -��  �/�  �	 ��	 Gp ��  ��0��  ��  �	 �	 0�  �C	  6�	 ,�	 0�k �&	  ��	 ��	 Hend �&	  ��	 ~�	 0�p �&	  [�	 Q�	 05W �)&	   �	 �	 0�k �C	  �	 ޔ	 0�k � C	  ݕ	 ŕ	 0W^ �/C	  �	 ۖ	 E �I{c _D     IOP �D     :��  ;b  '�Z -C	  R8ID     "l  9Uu 9Tt 9Q 9Rr   :��  �b  Hmm KC	  ��	 ��	 '�  KC	  T>�  0J�  Z&	  ��	 �	   :��  c  C�Z oC	  Hmm oC	  �	 �	 0�  o#C	  9�	 5�	 :��  �b  0J�  �&	  }�	 o�	  8�D     "l  9Uu 9Tt 9Q 9Rr   =je  VD      `�  �3�e  ��	 ��	 3�e  ��	 ��	 3�e  M�	 G�	 3�e  ��	 ��	 3�e  �	 �	 J�e  J�e  3|e  .�	 $�	 >`�  5�e  ��	 ��	 5�e  a�	 Y�	 K�e  ��5	f  ĝ	 ��	 Kf  ��6#f  _D     6,f  D     L5f  ��  �d  56f  �	 �	 LCf  0�  +d  5Df  y�	 s�	 5Qf  ў	 Ϟ	 5^f  ��	 ��	 5kf  ��	 ��	  M�l  �D      `�  ��d  3�l  ̟	 ȟ	 3�l  �	 �	 >`�  5�l  D�	 <�	 5�l  ��	 ��	 5m  ��	 ��	 5m  (�	 "�	 5m  t�	 r�	 6+m  D     <HD     �,   N�D     9Uv 9Qs 9R} 9X~ 9Y|   ;�D     �, e  9U  ;�D     	- (e  9U 9Ts 9Q�� ;�D     - Ge  9U 9T�� 8�D     "l  9Uu 9Tt 9Qs     @Z Q\	  {f  ALM Q0'Z  Ay2  R0&	  A"	 S0C	  A�#  T0C	  Aϋ U0	  A= V0	  A�  W0&	  A��  X0�  C�U Z\	  C^�  [e  Dp \�  C��  ]�  CKl  ^�  E�  �EWD  �FC��  � :Z  FC5�  �&	  C��  �&	  C�i �&	  C�[ �&	     ,c �\	  �D     K      �ah  -LM �2'Z  ��	 ��	 .p �2�  �	 ��	 -��  �2�  ��	 ��	 -ϋ �2	  �	 �	 -= �2	  S�	 K�	 -�  �2&	  ��	 ��	 0�U �\	  #�	 �	 0BT �&	  ��	 ��	 Hnn �&	  ��	 ��	 0�"  ��  ��	 ��	 0�"  ��  "�	  �	 0i!  ��  K�	 I�	 0%!  ��  t�	 r�	 02!  ��  ��	 ��	 0�  ��  Ʀ	 Ħ	 IWD  �D     I�  �D     4mD     =       0J�  �&	  �	 �	 Gdx ��  QHdy ��  �	 �	 8�D     d`  9Us 9Xv 9Y0   ,i Q\	  ��C     �      �3j  -LM Q5'Z  @�	 8�	 .p R5�  ��	 ��	 -��  S5�  h�	 ^�	 -ϋ T5	  �	 ۨ	 -= U5	  ��	 ��	 -�  V5&	  �	 �	 O�U X\	   0� Y�  `�	 R�	 0`�  Z	  �	 ��	 05�  Z	  ��	 x�	 0��  Z	  �	 ��	 0�k Z'	  �	 �	 Hh Z2	  ��	 ��	 0g Z5	  T�	 B�	 0md [&	  �	 �	 0�h [&	  R�	 L�	 0.a \_B  ��	 ��	 0oh ]		  �	 ֯	 I�  �&�C     >��  0�W ��  ˰	 ��	 Hw �	  ��	 ��	   ,�m �\	  ��C     -      �"l  -LM �6'Z  $�	 �	 .p �6�  ��	 ��	 -��  �6�  4�	 (�	 -ϋ �6	  ϳ	 ��	 -= �6	  ��	 ��	 -�  �6&	   �	 �	 O�U �\	   0� ��  g�	 Y�	 0`�  �	  �	 ��	 05�  �	  @�	 :�	 0��  �	  ��	 ��	 0�k �'	  ��	 �	 Hh �2	  M�	 ?�	 0md �&	  �	 �	 0�h �&	  (�	 "�	 0.a �_B  w�	 q�	 I�  &��C     :��  �k  0�W ��  Ƹ	 ��	 Hw �	  �	 �	  >��  0�W 	�  J�	 @�	 Hw 
	  ��	 ��	 0�S &	  ��	 �	   ,�e �\	  ��C     �       ��l  /LM �1'Z  UPpp �1�l  T-��  �1�  �	 ݺ	 Pbig �1�  RHp ��  9�	 /�	 0�e ��4  ��	 ��	 EWD  � 	�  @a 1\	  5m  ALM 11'Z  A��  21�  C�U 4\	  C5�  5&	  C��  5&	  Dmap 6_B  Cֳ  7C	  E�  z QMg *Qm  ALM *)'Z   @C[ �\	  �m  ALM �.'Z  A��  �.�7  Am �.C	  A�e �.eB  C�U �\	  C^�  �e  E�  $FDp �    ,�T  \	  @ D     )      �kp  -��   2�7  ݻ	 ջ	 -m !2C	  D�	 <�	 -�e "2�B  ��	 ��	 :p�  �n  0�n :�  7�	 1�	 0�R ;�  ��	 ��	 0~P <�  �	 �	 ;�!D     #- �n  9T@B$ 8�!D     #- 9T@B$  >@�  0^�  �e  l�	 b�	 C�  �&	  0�e �		  ߾	 ݾ	 0� �		  �	 �	 C� �%		  0�>  �kp  >�	 <�	 0ab ��  f�	 d�	 0�U �\	  ��	 ��	 Hp ��  �	 �	 ;� D     �, io  9U}  ;� D     �, �o  9U} 9T4 ;p"D     �, �o  9U}  ;{"D     �, �o  9U}  <�"D     �, ;�"D     #- �o  9T} 9Q~  ;�"D     #- �o  9T} 9Q~  ;�"D     #- p  9T} 9Q~  ;#D     #- ;p  9T} 9Q~  ;!#D     #- Tp  9T@B$ 8:#D     #- 9T@B$   	T(  ,�n \	  p#D     
       ��p  -��  -�7  Z�	 V�	 .req -&  ��	 ��	 -m -J1  ��	 ��	 Rz#D     0- 9U�U9T�T9Q09R�Q  S�m 
��C     /       �[q  -��  
�7  (�	 "�	 0^�  e  v�	 t�	 8��C     - 9Ts�
  TrT 2\	  �#D     �      �u  U��  2!�7  ��	 ��	 U^�  3!e  �	 �	 V�U 5\	  ��	 ~�	 &�@  6C	  ��V2�  7C	  �	 �	 W�  �:��  Wr  Xp b�  f�	 \�	 V��  cO	  ��	 ��	 VcC  dC	  ��	 ��	 V/� e&	  !�	 �	 8�%D     	- 9Uv 9Q|   :��  �s  V��  �		  J�	 D�	 V�1  �		  ��	 ��	 VcC  �C	  ��	 ��	 V/� �&	  5�	 1�	 ;h$D     �, �r  9Uv 9T8 ;x$D     �, �r  9Uv  ;�$D     �, �r  9Uv  ;�$D     �, s  9Uv  ;�$D     �, -s  9Uv  ;�$D     =- Es  9Uv  ;�$D     �, ]s  9Uv  8%D     	- 9Uv 9T~ 2$#����9Qs�
  :�  5t  &(a  �C	  ��Y�&D     �s  9Us 9TTDBC9Qv 9R�� Y�&D     �s  9Us 9TTDBE9Qv 9R�� Y'D      t  9Us 9Ttadb9Qv 9R�� 8H'D     =- 9Uv   Y�#D     _t  9Us 9TCLBC9Qv 9R�� ;$D     - }t  9Uv 9T|  ;8$D     =- �t  9Uv  YF%D     �t  9Us 9TCLBE9Qv 9R�� Y~%D     �t  9Us 9Tcolb9Qv 9R�� N�%D     9Us 9Txibs9Qv 9R��  @�^ �\	  �u  A��  �%�7  Bidx �%&	  A{W �%�B  C�U �\	  C�r �37  C��  �O	  CQ  ��S  ZEnd 6[�u  C�B x6  FC�  		    FC�B &�6    S
[ � D           ��v  -��  �#�7  s�	 k�	 0ڰ  ��  ��	 ��	 0�r �37  �	 ��	 0��  �O	  r�	 l�	 1PD     �       �v  0�B �x6  ��	 ��	 Hn �		  ��	 ��	 ;_D     J- �v  9U}  ;�D     J- �v  9U}  8�D     J- 9U}   4�D     (       0�B ��6  J�	 H�	 8�D     J- 9U}    ,�S ~\	  �QD     n      ��}  -��  ~�7  ��	 p�	 0^�  �e  ��	 ��	 0�U �\	  o�	 ]�	 0��  �O	  0�	 *�	 '7S �C	  ��0�V �C	  ��	 y�	 I�  �_RD     M1~  pRD      � ��{  3Z~  I�	 A�	 3N~  ��	 ��	 3B~  Y�	 I�	 >� 5f~  �	 �	 Kr~  ��5~~  f�	 ^�	 5�~  ��	 ��	 5�~  ��	 ��	 5�~  _�	 =�	 6�~  �RD     6�~  �UD     \�~  L�~    �x  5�~  ��	 ��	 ;�RD     V- �x  9U~ 9T29Q09R 9X09Y�� ;�RD     �, �x  9Uv 9T 1$ ;,SD     �, �x  9Uv  ;QSD     �, �x  9Uv  87VD     �, 9Uv   L�~  P 8y  5�~   �	 ��	 ]�~  `SD     %       5�~  >�	 8�	   L�~  � �z  5�~  ��	 ��	 L  � ?z  5  <�	 .�	 L  0 �y  5  ��	 ��	 8�TD     =- 9Uv   ;�SD     =- �y  9Uv  ;$TD     V- �y  9U~ 9T19Q09R}����9X09Y�� ;ETD     b- z  9Uv 9Q}  ;uTD     =- #z  9Uv  8�TD     o- 9Uv 9T��  ;�SD     V- zz  9U~ 9T89Q09R	���
��9X09Y�� ;PVD     V- �z  9U~ 9T89Q09R09X09Y�� 8�VD     V- 9U~ 9T19Q09R19X09Y��  74  VD            {  55  )�	 '�	 8 VD     J- 9U~   7!  gVD     0       ?{  5&  O�	 M�	  ;�RD     |- ^{  9Uv 9T�� ;�UD     J- ~{  9U~ 9T�� 8�UD     J- 9U~ 9T��   M�}  �TD      p �%}  3�}  w�	 u�	 3�}  ��	 ��	 3�}  ��	 ��	 >p 5�}  �	 �	 K�}  ��5�}  S�	 M�	 5�}  ��	 ��	 6�}  �TD     6�}  �UD     7~  cUD     G       k|  5~  :�	 6�	 ^~  � 5~  y�	 q�	   7!~  �VD            �|  5"~  ��	 ��	  ;�TD     |- �|  9Uv 9T�� ;+UD     V- �|  9U} 9T19Q09R��~9X09Y�� ;SUD     b- }  9Uv 9T��~9Q�� 8�UD     J- 9U}    Y�QD     O}  9Us 9Ttsop9Qv 9R�� ; RD     =- g}  9Uv  8<RD     �- 9Uv 9T   @�Y ;\	  1~  A��  ;�7  A^�  <e  A�V =C	  Cڰ  ?�  C�U @\	  C�  B	  C�p Ce6  E�  xEWD  u[!~  Dn Z	  FDidx _7	    FC�B l�6    _zj �\	  B  `��  ��7  `^�  �e  `�V �C	  aڰ  ��  a�U �\	  a�  �	  a�`  �		  aTL  ��5  aDl �_6  E�  5EWD  1E}�  ([�~  bn �	   [�~  bn �	  Fbidx �	    [!  bn �		  Fblen �&	  Fbd �	     [4  C�B x6   FDn *		    c�[ 
�p�C     �      ��  U��  
�$�7  �	 �	 U<  
�$�  ��	 ~�	 UJ�  
�$&	  ��	 ��	 U�j 
�$YC  *�	 "�	 U� 
�$�5  ��	 ��	 &�U 
�\	  ��V^�  
�e  F�	 D�	 V�& 
�kp  m�	 k�	 VHh 
�C	  ��	 ��	 V�@  
� C	  ��	 ��	 V�c  
�,C	  ��	 ��	 Xk 
�		  s�	 k�	 Xvar 
�#�T  ��	 ��	 IOY 
0 �C     :��  ��  dv 
�_   P : �  �  Hf 
8  �	 	�	 Ga 
9	  ��Gb 
:	  ��Y?�C     ��  9Us 9T 9Q�� YU�C     �  9Us 9T 9Q�� N��C     9Us 9T 9Q��  ;��C     �, A�  9U��9T�� ;�C     |- b�  9U��9T�� ;a�C     �, |�  9U�� ;��C     |- ��  9U��9T�� ;��C     |- ��  9U��9T�� ;��C     �, ׁ  9Uw  8�C     |- 9T��  T�^ 
�\	  p,D     t       ��  U��  
�!�7  M�	 C�	 U^�  
�!e  ��	 ��	 U<  
�!�  Z�	 V�	 V�U 
�\	  ��	 ��	 V�& 
�kp  ��	 ��	 &�m 
�")�  	�
G     eWD  
��,D     :��  ڂ  Xv 
�_    �	 �	 N�,D     9Us�|9Taehv9Qv 9R0  ;�,D     �- �  9Uv 9T	�
G     9Qs  N�,D     9Taehh  Z&  )�  @    �  T�U 
I\	  ��C     u       �1�  U��  
I!�7  a�	 Y�	 U^�  
J!e  ��	 ��	 U<  
K!�  B�	 <�	 V�U 
M\	  ��	 ��	 Xtag 
NC	  ��	 ��	 &�@  
NC	  �HVd^ 
OJ1  :�	 6�	 V` 
PJ1  t�	 p�	 eWD  
gC�C     Y(�C     �  9U�U9Qv 9R�H 8?�C     =- 9Uv   ,{Y x\	  �D     B      ��  -��  x!�7  ��	 ��	 -^�  y!e  d�	 V�	 0�U {\	  �	 ��	 0ڰ  |�  +�	 %�	 Hj ~&	  v�	 t�	 0�  ~&	  ��	 ��	 0l �3  ��	 ��	 I�  ��D     Y�D     �  9Uv 9Tpsag9Qs 9R0 ;�D     �, ;�  9Us 9T4 ;�D     �, S�  9Us  ;�D     �, k�  9Us  ;�D     �, ��  9Us  ;BD     V- ��  9U| 9T49Q09R} 9X09Y�L ;eD     �, օ  9Us 9T} 2$ ;�D     �, �  9Us  ;�D     �, �  9Us  8�D     �, 9Us   ,9q 9\	  �'D     J       ��  -��  9!�7  "�	 �	 -^�  :!e  ��	 ��	 'vg <"�  	�G     0�U T\	  X�	 V�	 0Fq U$�  ��	 {�	 I�  `�'D     Y�'D     �  9Us 9TTLCP9Qv 9R0 R�'D     �- 9U�T9T	�G     9Q�U#�  Z&  �  @    �  	e-  ,)s �\	  0+D     J       ��  -��  �!�7  *�	 �	 -^�  �!e  ��	 ��	 0�U �\	  `�	 ^�	 06s ��  ��	 ��	 '^ "#�  	`G     YL+D     ��  9Us 9Ttsop9Qv 9R0 Rz+D     �- 9U�T9T	`G     9Q�U#�  	G,  Z&  #�  @   
 �  @Hr Y\	  ܈  A��  Y �7  A^�  Z e  C�U \\	  Dos2 ]܈  '�k _"�  	�G     'Jn �"�  	�G     '\n �"�  	`G     '�k �"�  	PG     I�  �X_D      	�+  Z&  �  @   + �  Z&  �  @    ��  Z&  �  @    �  @<_ 3\	  l�  A��  3!�7  A^�  4!e  C�U 6\	  I�  @�QD      SxS �D     
      ���  -��  ��7  ,�	 &�	 0ڰ  ��  z�	 x�	 0�B ��3  ��	 ��	 14D     X       <�  0�, �2  ��	 ��	 0��  �2  K�	 I�	 ;`D     J- !�  9Uv  8�D     J- 9Uv 9Ts   4�D     S       0�, 3  t�	 n�	 0��  3  ��	 ��	 ;�D     J- ��  9Uv  8�D     J- 9Uv 9Ts    ,�k 8\	  �'D     Z      �=�  -��  8!�7  ��	 ��	 -^�  9!e  U�	 K�	 '�U ;\	  ��0ڰ  <�  ��	 ��	 0Hh =C	  �	 �	 'ց  =C	  ��0�S >C	  V�	 P�	 0�j >"C	  ��	 ��	 0�B ?�3  3�	 +�	 '<e A"M�  	�G     '!l M"�  	�G     '�j \"b�  	�G     I�  �G(D     :��  4�  0�, �3  ��	 ��	 0��  �3  ��	 ��	 8�*D     �- 9Us 9T	�G     9Q   :@�  ��  0�, ��2  �	 ��	 0/� �&	  p�	 b�	 ;�(D     �- ��  9Us 9T	�G     9Q  8�)D     V- 9U| 9T 9Y��  Y(D     ތ  9U~ 9Teman9Qs 9R�� ;((D     =- ��  9Us  ;?(D     �- "�  9Us 9T	�G     9Q~� ;�(D     V- Q�  9U| 9T 9Q09X09Y�� ;�(D     �, i�  9Us  ;�)D     �, ��  9Us  ;�)D     �, ��  9Us 9T}  ;�)D     |- ��  9Us 9T�� ;*D     V- �  9U| 9TH9Q09R 9X09Y�� ;6*D     �, 
�  9Us  ;�*D     �, "�  9Us  8�*D     �, 9Us 9Tv  Z&  M�  @    =�  Z&  b�  @    R�  ,p` �\	  �+D     �       ���  -��  �!�7  �	 �	 -^�  �!e  ��	 v�	 0�U �\	   �	 ��	 0�S ���  ��	 ��	 '�` �"�  	@G     '�g �"��  	 G     I�   `,D     Y�+D     E�  9Us 9Tpxam9Q| 9R0 ;�+D     �- p�  9U| 9T	@G     9Q}  8,D     �- 9U| 9T	 G     9Q}   	S.  Z&  ��  @    ��  ,�b �\	  @^D            �&�  -��  �!�7  �	 �	 -^�  �!e  I�	 E�	 RG^D     ��  9U�U9T�T9Qdehb  ,hR �\	  P^D            ���  -��  �!�7  ��	 ��	 -^�  �!e  ��	 ��	 RW^D     ��  9U�U9T�T9Qdaeh  @�i n\	  �  A��  n+�7  A^�  o+e  Btag p+C	  C�U r\	  C�& s�  'd' u"+�  	@G     I�  �^D      	Z'  Z&  +�  @    �  ,gb *\	  �D     �       ���  -��  * �7  �	 ��	 .tag + C	  n�	 f�	 -�  , 7	  ��	 ��	 -_| - �  )�	 �	 -��  . J1  ��	 ��	 '�U 0\	  P0^�  1e  �	 �	 0�B 2$2  F�	 D�	 0ֳ  3C	  s�	 i�	 E�  VMY�  �D       @�  9v�  3j�  ��	 ��	 3j�  ��	 ��	 3v�  �	 �	 >@�  5��  E�	 A�	 5��  }�	 {�	   fWD     �- f�D     �-  ,X X\	   ZD     �      �f�  -��  X%�7  ��	 ��	 -^�  Y%e  �	 �	 '�i  [�1  ��'�U \\	  ��0ڰ  ]�  v�	 n�	 Hnn ^		  ��	 ��	 0+] ^		  8�	 "�	 '�e `"v�  	�G     I�  ��]D     :� 	�  0�, �2  8�	 "�	 Hi �		  ��	 ��	 0�Y ��  ��	 ��	 ;b[D     �, ē  9Us  ;m[D     �, ܓ  9Us  ;y[D     �, ��  9Us  8�[D     �, 9Us   M{�  �[D       ���  3��  ��	 ��	 3��  ��	 ��	 3��  �	 �	 3��  q�	 k�	 > 5��  ��	 ��	 5��  ��	 ��	 5ǖ  M�	 G�	 5Ӗ  ��	 ��	 5ߖ  !�	 �	 5�  ��	 ��	 5��  ��	 ��	 \�  L"�  ` r�  K#�  ��L/�  � I�  ?0�  ;�\D     �, ��  9Us  ;]D     �- �  9Us 9T�� 83]D     �, 9Us 9Tv 
��#4$ $ &w "  8�\D     �- 9Us 9T	�G     9Q��  8\D     �, 9Us 9Tw    ;@ZD     =- ��  9Us  ;RZD     �- ƕ  9Us 9T�� ;�ZD     �- �  9Us 9T	�G     9Q�� ;�ZD     V- !�  9U~ 9T 9Q09X09Y�� ;�ZD     �, 9�  9Us  ;[D     �, Q�  9Us  8�]D     �, 9Us   Z&  v�  @    f�  _3[ �\	  ?�  `�i  �!�1  `^�  �!e  `��  �!�5  a�U �\	  bnn �		  a+] �		  a�R �&	  aps �&	  a�l �,&	  a�  �C	  &�a �"v�  	�G     E�  9Fa�B �2  Fa�  ��     To_ �\	  ��C     V       �Y�  U��  �"�7  U�	 O�	 gtag �"C	  ��	 ��	 U^�  �"e  ��	 ��	 U��  �"J1  K�	 E�	 V�B �$2  ��	 ��	 a�U �\	  e�  �'�C     hY�  ��C       ��  �C�  3j�  ��	 ��	 3j�  �	 �	 3v�  d�	 `�	 >��  5��  ��	 ��	 5��  ��	 ��	   R;�C     �, 9U�Q  _�l :$2  ��  `��  :#�7  itag ;#C	  a�, =$2  a��  >$2   T�V �	  ��C           �Ě  j��  �!�7  UUsl  �!&	  �	 �	 U�J  �!&	  f�	 `�	 V�Y  �	  ��	 ��	 V/� �&	  L 
 B 
 V�� �&	  � 
 � 
 Xp ��  .
 
 V��  ��  m
 i
 I�Z . �C     Ics (��C     >��  VǞ  ��  �
 �
 V�W ��  "
  
 V��  �&	  O
 E
 V��  �&	  7
 '
 Ve� �&	  �
 }
 VzR �&	  g
 _
 V<v �	  �
 �
 >P�  a�e �C	  : �  ��  Xmin �&	  _
 [
 Xmax �&	  �
 �
 >P�  Xmid �&	  
 �
 Xq ��  ~
 r
 Xkey �C	  	
 	
   >��  0�Q 
&	  �	
 �	
 >��  Hkey C	  �	
 �	
      krm ��  `��  ��7  a^�  �e   T�O ,\	  p�C     E      ��  U��  ,!�7  �

 �

 U^�  -!e  %
 
 V�U /\	  �
 �
 &�@  0C	  ��Xp 1�  $
 �
 V��  2�  �
 �
 Xnn 3&	  �
 �
 V�R  3&	  D
 @
 VfO 4�  �
 �
 V  4�  �
 �
 e�  ���C     e�Z �p�C     :p�  Ϝ  VzR X&	  (
 "
 V��  X&	  {
 w
 Ve� X%&	  �
 �
 V��  X/&	  �
 �
 V�_ Y�  (
  
 V�� Z�  �
 �
 4%�C     [       V/� �C	  �
 �
 VS �C	  +
 %
 4:�C     /       Vn ��  �
 
    Y��C     ��  9Us 9Tnrek9Qv 9R�� 8��C     	- 9Uv 9Qs�
  ,sQ \	   �C     �       �ם  /��  !�7  U-@  !&	  
 
 0i 	ם  q
 m
 0�  �  �
 �
 Hp �  �
 �
 Hq c?  �
 �
 0��  c?  �
 �
 0�e  		  
 �
  	IY  c�Q ��D     G       �q�  U��  ��7  �
 �
 V^�  �e  
 
 Vڰ  ��  B
 @
 Vi �ם  o
 g
 ;�D     - c�  9Ts f�D     J-  Tri K\	  �D     =      �D�  U��  K!�7  �
 �
 U^�  L!e  >
 4
 &�U N\	  ��Vڰ  O�  �
 �
 &�B Q�  ��Xp R�  
 �
 Vi Tם  �
 y
 VFm VC	  
 

 &�@  WC	  ��e�O ��D     eIc ��D     :�  S�  V�P �C	  5
 /
 &$X � C	  _&X �.C	  _V; ��5  �
 �
 V��  ��5  �
 �
 Xq ��5  G
 ;
 ;�D     V- ��  9U~ 9T29Q09X09Y�� ;wD     V- (�  9U~ 9T29Q09X09Y�� 8{D     V- 9U~ 9T29Q09X09Y��  Y�D     }�  9Us 9TLAPC9Qv 9R�� ;D     - ��  9Uv 9T|  ;D     J- ��  9U~ 9T}  ;@D     	- נ  9Uv 9Q|  ;wD     �- ��  9U~ 9T(9Q�� ;D     V- *�  9U~ 9T49Q09X09Y�� 8+D     �  9Uu 9T0  ,S \	  D     -      �Ф  -��  +�7  �
 �
 -�e  +&	  f
 Z
 -�h +I  �
 �
 -Q +I  7
 -
 '�U \	  ��Hx &	  �
 �
 Hy &	  
 
 Hb �  �
 �
 Hg �  
 
 Hr �  b
 \
 0q  �  �
 �
 0ֳ  C	  
 �
 Hsrc �  �
 {
 Hdst �  �
 �
 :��  ݣ  0�� 5	  �
 �
 0� 5	  w 
 o 
 0�Z 5	  7!
 1!
 0G�  5$	  �!
 �!
 4�D     I      0ڰ  E�  "
 "
 05�  G&	  A"
 ="
 0M} H&	  }"
 y"
 0`�  I&	  �"
 �"
 Hbuf K�  �"
 �"
 Hp L�  C#
 A#
 Hq M�  j#
 f#
 ;D     �- ��  9T���| ����9Q�� ;�D     �- ��  9T}  8�D     �, 9Us 9T��   : �  ��  Haa �G   �#
 �#
 Hfa �G   $
 $
 Dfb �G   Dfg �G   Dfr �G   Hba2 �G   <$
 8$
 Hbb �G   {$
 w$
 Hbg �G   �$
 �$
 Hbr �G   �$
 �$
 Hba �G   <%
 :%
  ;�D     �, ��  9U~ 9Ts  8�D     �- 9T09Qs   TMU ��  ��C     i      �#�  j��  �.�7  UUOq �.&	  k%
 _%
 j�j  �.o?  QU�e  �.o?   &
 �%
 j��  �.�C  XV�d �#�  {&
 u&
 VX_ �lX  �&
 �&
 >��  V�  �C	  *(
 &(
 l)�  ��C       �  �3^�  d(
 `(
 3R�  �(
 �(
 3F�  �(
 �(
 3:�  D)
 @)
 > �  5j�  �)
 z)
 5v�  �)
 �)
 ^��  p�  5��  *
 *
 5��  �*
 z*
 5��  +
 +
      	�X  _N_ ��  ��  `�` �-�  `Kq �-	  `�W �-&	  `w� �-��  bmin �	  bmax �	  Fbmid �	  bp ��  bgid �		    	lX  c�] �`D     G       �A�  U��  ��7  �+
 �+
 V^�  �e  �+
 �+
 Vڰ  ��  ,
 ,
 V�d �#�  <,
 4,
 ;�D     - 3�  9Ts f�D     J-  T�d T\	  �D     �      ��  U��  T!�7  �,
 �,
 U^�  U!e  "-
 -
 &�U W\	  ��Vڰ  X�  �-
 �-
 &�B Z�  ��Xp [�  
.
 �-
 V�d ]#�  �.
 �.
 V�Q _C	  {/
 y/
 V�l _"C	  �/
 �/
 &�@  `C	  ��e�U �(D     eIc � D     YD     g�  9Us 9TRLOC9Qv 9R�� ;3D     - ��  9Uv 9T}  ;>D     J- ��  9U| 9T~  ;hD     	- ��  9Uv 9Q}  8�D     �- 9U| 9T(9Q��  ,@S \	  ��C            �s�  -�� #�  �/
 �/
 -�  #�K  0
 0
 0I_  �"  m0
 g0
 0Oe !L  �0
 �0
 m��C     9U�U9T�T  ,Qi �\	  �,D           �;�  -��  �!�7  �0
 �0
 0�B ��  1
 u1
 0��  ��   2
 �1
 '�s �2	  ��~Gp ��  ��~0�-  �   w2
 s2
 >��  '�� ��  ��0�  ��  �2
 �2
 >0�  'I_ �(�  ��~'��  �(2	  ��~'Ne �(A�  ��~'Oe �(L  ��~>p�  '��  �'�L  ��'�U �'i	  ��~1�/D     +       �  '�` ��"  ��~8�/D     �- 9Q��9R��~  ;Q/D     �- �  9U��9Qw 9R0 ;n/D     �- &�  9U�� N�/D     9T��     	L  ;�  ,�Y ��  ��C            �֫  -Aq �+VR  �2
 �2
 -��  �+'$  73
 33
 0��  ��7  r3
 p3
 0Q  ��S  �3
 �3
 m��C     9U�U9T�T  ,?a z&	  p�C            �f�  -Aq z,VR  �3
 �3
 -��  {,�  4
 �3
 0��  }�7  <4
 :4
 0Q  ~�S  b4
 `4
 m}�C     9U�U9T�T  S�c n�D     (       �Ҭ  -Aq n&VR  �4
 �4
 0��  p  �4
 �4
 0ڰ  q�  5
 5
 <�D     J-  ,�b W\	  0�C     6       ���  -Aq W&VR  45
 ,5
 -��  X&n	  �5
 �5
 0��  Z�7  �5
 �5
 0ڰ  [�  6
 
6
 0Q  \�S  J6
 D6
 m[�C     9T�U9R	`YD     9X0  ,U J=  `YD     ?       �`�  -��  J�7  �6
 �6
 .idx K&	  �6
 �6
 '{W Mq  �h=u  mYD      0 P3<u  A7
 ;7
 3/u  �7
 �7
 3"u  �7
 �7
 >0 ?Iu  ?Vu  ?cu  ?pu  \}u  8�YD     r 9U�U9T�T9Q�h    ,$_ �'$  ��C     P      ���  -I_ �'�K  H8
 28
 -ڰ  �'�  K9
 59
 -�I  �'�  ;:
 5:
 Hp ��  �:
 �:
 Hi �	  I<
 '<
 0�g �C	  �=
 �=
 0�g �C	  �=
 �=
 :p�  ��  0�o ��W  C>
 9>
 0�R  ��  �>
 �>
 0�` ��   ?
 ?
 0�e ��  @
 @
 0�o ��  �@
 t@
 0�_ ��  "A
 A
 Hdp ��  �A
 �A
 Hdi �&	  >B
 <B
 Hni �&	  jB
 bB
 Hk �&	  �B
 �B
 Hret �'$  �C
 �C
 MԲ  ��C      ��  �F�  3�  D
 D
 >��  5�  oD
 kD
 5��  �D
 �D
   ;?�C     O�  e�  9U 9Q�T no�C     ��  ��  9U�U9Q�T R��C     ��  9U�U  8��C     K�  9Uu 9Tt   ,�S '$  ��C     �       ���  -I_ +�K  LE
 @E
 .p �+�  �E
 �E
 -ڰ  �+�  �F
 �F
 0�o ��W  G
 G
 C�` ��  Hi �&	  �G
 �G
 Hret �'$  �G
 �G
 8�C     O�  9U| 9Ts9Q�Q  ,1c Z'$  �C     �       �Բ  -I_ Z'�K  H
 H
 .p ['�  �H
 �H
 -ڰ  \'�  �I
 �I
 0�o ^�W  J
 �I
 0�R  _�  �J
 �J
 Hcnt `&	  pK
 jK
 Hq a'$  �K
 �K
 1p�C     6       _�  Huni l�  @L
 >L
  MԲ  �C      0�  d��  3�  qL
 cL
 >0�  5�  M
 M
 5��  �M
 �M
   ;_�C     O�  ��  9U|  8��C     O�  9T1  @vX H&	  �  Bp H'�  C�R  J�  Dtot K&	   ,�h "'$  ��C           �a�  -I_ "'�K  �M
 �M
 -ڰ  #'�  PN
 JN
 -�W $'�  �N
 �N
 0�o &�W  _O
 WO
 0/� '�  �O
 �O
 Hp (�  P
 �O
 Hq )'$  �P
 �P
 :0�  ?�  0gZ 1�  NQ
 JQ
 0�g 2C	  �Q
 �Q
 0�g 3C	  R
 R
 ;^ D     ߸  $�  9Uu 9Tt  8� D     �  9Uu 9Tt   8��C     O�  9U| 9T}9Q�T  ,5r '$  � D     �       �5�  -I_ "�K  rR
 fR
 -ڰ  	"�   S
 �R
 0�o �W  XS
 LS
 0/� �  �S
 �S
 Hp �  =T
 /T
 0�Y  '$  �T
 �T
 Hi �  U
 U
 8� D     O�  9U| 9Tv9Q�T  ,]j �	  ��C     x       �+�  -I_ �,�K  VU
 RU
 -�_ �,�  �U
 �U
 -�I  �,�  ?V
 5V
 Hp ��  �V
 �V
 0�g �C	  "W
 W
 0�g �C	  nW
 hW
 ;��C     K�  �  9Uu 9Tt  ;��C     �  �  9Uu 9Tt  8�C     ߸  9Uu 9Tt   ,P �&	   �C     �       �K�  -I_ �(�K  �W
 �W
 -�n  �(�K  X
 X
 -�_ �(�  �X
 �X
 -�I  �(�  �Y
 �Y
 Hp ��  Z
 
Z
 0�g �C	  aZ
 ]Z
 0�g �C	  �Z
 �Z
 ;>�C     K�  ��  9Uu 9Tt  ;t�C     ߸  �  9Uu 9Tt  o��C     0�  9U�T R��C     �  9Uu 9Tt   ,�o ��  ��C     �       ��  -Ǟ  �'�  [
 [
 /QT �'�  T0�Q ��  L[
 J[
 Hmax ��  �[
 �[
 Hmin ��  `\
 \\
 >��  Hmid ��  �\
 �\
 Hp ��  ]
 ]
 0gZ �C	  �]
 �]
   ,�Z �&	  ��C     �       �߸  -Ǟ  �1�  D^
 @^
 /��  �1�  T0�` ��  ~^
 |^
 Hmax ��  �^
 �^
 Hmin ��  h_
 d_
 >p�  Hmid ��  �_
 �_
 Hp ��  $`
 `
 Huni ��  �`
 �`
   ,�` f&	   �C     �       ���  -Ǟ  f.�   a
 a
 /��  g.�  T0�R  i�  Za
 Xa
 Hmax j�  �a
 �a
 Hmin j�  nb
 jb
 >0�  Hmid u�  �b
 �b
 Hp v�  0c
 c
 0�k wC	  3d
 -d
 Hcnt x&	  �d
 �d
   ,Tm X\	   �C            � �  /I_ X%�K  U/�  Y%�K  T ,�] L�  ��C     	       �B�  /I_ L$�K  U/��  M$'$  T ,�T @&	  ��C            ���  /I_ @$�K  U/��  A$�  T ,Z �\	  LD           ��  -�B �%�  �d
 �d
 -��  �%�J  Ye
 Qe
 Hp ��  �e
 �e
 0��  �C	  �f
 �f
 0qr �C	  g
 �f
 :��  н  Hn �C	  &g
 $g
 0�O �C	  Xg
 Jg
 >��  0gZ �C	  �g
 �g
 0�g �C	  bh
 Zh
 0�g �C	  �h
 �h
 :  �  0#r ��  hi
 Ti
 0�R  �C	  mj
 ej
 Hi �C	  �j
 �j
 0�j �C	  Pk
 Hk
 :P  H�  0Ǟ  C	  �k
 �k
 Hcnt C	  �k
 �k
 ;ND     . .�  9Us 9T8 8ND     . 9Us 9T8  ;�OD     . e�  9Us 9T8 8PD     . 9Us 9T8  :�  ��  Hndp �  Nl
 >l
 0�` C	  m
 �l
 Hi C	  �m
 vm
 0i C	  n
 n
 :�  a�  Huni 'C	  tn
 nn
 Hgid (C	  �n
 �n
 ;!OD     . *�  9Us 9T8 ;AOD     . G�  9Us 9T8 8yOD     . 9Us 9T@  ;�OD     . ~�  9Us 9T8 8�OD     . 9Us 9T8  ;AMD     . ��  9Us 9T8 8]OD     . 9Us 9T8   ;�LD     . �  9Us 9T8 8PD     . 9Us 9T8  ,V �\	  ��C     !       �O�  /I_ ��W  U-�B ��  o
 o
  ,�g �\	  ��C     X       ���  -I_ � �W  _o
 Wo
 -�s � �  �o
 �o
 -ڰ  � �  Dp
 :p
 0-Q  ��  �p
 �p
 '�U �\	  �\8��C     V- 9U�Q9T49Rv 9Y�\  S�q �PD     1       �T�  -I_ ��W  �p
 �p
 0ڰ  ��  ^q
 Zq
 <uD     J-  ,�f \	  ��C            ���  /I_ %�K  U/�  %�K  THp  �  �q
 �q
  @�r �  �  AI_ $�K  A��  $'$  C�o OW  CJ�  &	   ,b\ �
&	  p�C            �^�  -I_ �
$�K  �q
 �q
 -��  �
$�  r
 r
 8��C     ^�  9U�U9T�t9Q0  ,] �
&	  `�C     	      ���  -I_ �
*�K  ]r
 Mr
 -��  �
*'$  s
 s
 -�W �
*�  �s
 �s
 0J�  �
&	  �s
 �s
 Hp �
�  �t
 �t
 01X �
�  Vu
 Ru
 0��  �
�  �u
 �u
 0�k �
�  ,v
 &v
 Hend �
�  �v
 �v
 Hmax �
�  �w
 �w
 Hmin �
�  �x
 �x
 Hmid �
�  �x
 �x
 > �  0��  �
  �y
 �y
 0�o �
OW  z
 z
 8��C     ��  9Uu    Ss q
��C     �       ���  /I_ q
OW  U0��  s
  �z
 �z
 Hp t
�  �z
 �z
 0�k u
C	  L{
 B{
 Hend u
C	  G|
 A|
 0�W u
C	  �|
 �|
 0��  u
%C	  j}
 h}
 Hn v
C	  �}
 �}
 0J�  w
&	  �}
 �}
 IWD  �
P�C      ,S] 7
\	  �JD     2      �5�  -�B 7
%�  z~
 p~
 -��  8
%�J  �~
 �~
 Hp :
�  x
 h
 0��  ;
C	  2�
 ,�
 01X <
C	  ��
 ��
 1@KD     �       ��  Hn P
C	  �
 ��
 0�k P
C	  d�
 `�
 Hend P
C	  ��
 ��
 0�W P
 C	  ց
 ԁ
 0��  P
*C	  .�
 $�
 ;gKD     . ��  9U 9T8 ;�KD     . ��  9U 9T8 8�KD     . 9U 9T@  ;@KD     . �  9U 9T8 8�KD     . 9U 9T8  ,as (
\	  ��C            �}�  /I_ (
OW  U-�B )
�  ��
 ��
  ,]` �	\	  ��C            ���  /I_ �	%�K  U/�  �	%�K  THp �	�  ��
 ܂
  @b �	�  �  AI_ �	$�K  A��  �	$'$  C�o �	�V  CJ�  �	&	   ,-d �	&	  p�C            ���  -I_ �	$�K  !�
 �
 -��  �	$�  ^�
 Z�
 8��C     ��  9U�U9T�t9Q0  ,g S	&	  @�C     !      ���  -I_ S	*�K  ��
 ��
 -��  T	*'$  Z�
 P�
 -�W U	*�  Ԅ
 ̄
 0J�  W	&	  @�
 6�
 Hp X	�  ��
 ��
 01X Y	�  ��
 ��
 0��  Z	�  �
 �
 0�k [	�  e�
 ]�
 Hend [	�  ��
 ��
 0e [	�  $�
 "�
 Hmax \	�  ��
 ��
 Hmin \	�  X�
 R�
 Hmid \	�  ��
 ��
 >��  0��  �	  ��
 ��
 0�o �	�V  �
 ڌ
 8��C     ��  9Uu    S�W 	0�C     	      ���  /I_ 	�V  U0��  	  l�
 h�
 Hp 	�  ��
 ��
 0�k 	C	  )�
 %�
 Hend 	C	  c�
 _�
 0e 	C	  ��
 ��
 0��  	%C	  �
 ӎ
 Hn 	C	  z�
 v�
 0J�  	&	  ��
 ��
 IWD  M		�C     E]�  -	 ,!Q �\	  `ID     j      ���  -�B �%�  :�
 0�
 -��  �%�J  ��
 ��
 Hp ��  8�
 (�
 0��  �C	  �
 �
 01X �C	  m�
 g�
 1�ID     �       j�  Hn �C	  ��
 ��
 0�k �C	  ��
 ��
 Hend �C	  4�
 .�
 0e � C	  ��
 ��
 0��  �*C	  ߓ
 ד
 1JD     -       3�  Hd  	�  D�
 >�
 89JD     . 9U~ 9T@  ; JD     . P�  9U~ 9T8 8�JD     . 9U~ 9T8  ;�ID     . ��  9U~ 9T8 8�JD     . 9U~ 9T8  ,�W �\	  �C            ���  /I_ ��V  U-�B ��  ��
 ��
  ,eS v\	  ��C            �>�  /I_ v%�K  U/�  w%�K  THp y�  ה
 Ӕ
  ,�W M�  @�C     �       ��  -I_ M$�K  �
 �
 /��  N$'$  T0�B P�  W�
 Q�
 0��  Q�  ��
 ��
 0J�  R&	  ��
 ��
 Hp S�  G�
 5�
 C�k T�  C/� U�  Hidx V�  �
 �
  ,H` 2&	   �C     3       ���  /I_ 2$�K  U-��  3$�  ��
 ��
 0�B 5�  ͚
 ɚ
 0�Y  6&	  �
 �
 Hp 7�  2�
 *�
 0�k 8�  ��
 ��
 0/� 9�  (�
 $�
 Hidx :�  ��
 ��
  ,�r \	  �HD     �       ���  -�B %�  b�
 V�
 -��  %�J  �
 �
 Hp �  ��
 x�
 0��  C	  D�
 >�
 0/� C	  ��
 ��
 :P�  ��  0J�  "&	  '�
 �
 8ID     . 9U| 9T@  ;�HD     . ��  9U| 9T8 8UID     . 9U| 9T8  ,�i �\	  ��C            ��  /I_ �$�K  U/�  �$�K  THp ��  ֠
 Ҡ
  ,�R ��  ��C     �       �*�  -I_ �#�K  �
 �
 /��  �#'$  T0��  �  i�
 e�
 0�Y  ��  ��
 ��
 0��  ��  <�
 2�
 0J�  �&	  Ǣ
 ��
 0�B ��  ��
 ��
 Hp ��  �
 �
 01X ��  Ӥ
 Ϥ
 C�k ��  Dend ��  0e ��  g�
 c�
 E]�  � ,Gf f&	  p�C     e       ���  -I_ f#�K  �
 �
 -��  g#�  (�
 $�
 0�B i�  e�
 a�
 O�Y  j&	   Hp k�  ��
 ��
 01X l�  N�
 L�
 C�k m�  Dend m�  0e m�  ��
 ��
  ,�Q \	  �ED     �      �q�  -�B $�  j�
 \�
 -��  $�J  �
 �
 Hp �  ��
 ��
 04o �  �
 �
 0��  �  c�
 _�
 01X �  �
 �
 :p�  �  Hn �  ��
 w�
 0�k �  �
 
�
 Dend �  0e !�  ��
 ��
 0/� +�  9�
 1�
 0��  2�  ��
 ��
 >��  Hhi !&	  �
 �
 Hlo !&	  ��
 ��
 : �  ��  Hd 0�  >�
 4�
 ;�FD     . t�  9U} 9T@ ;`GD     . ��  9U} 9T8 ;�GD     . ��  9U} 9T8 ;9HD     . ��  9U} 9T8 8QHD     . 9U} 9T8  ;�FD     . �  9U} 9T8 8�GD     . 9U} 9T8   ;uGD     . :�  9U} 9T8 ;mHD     . W�  9U} 9T8 8�HD     . 9U} 9T8  ,�m �\	  @�C     $       ���  /I_ �$�K  U/�  �$�K  THp ��  ��
 ��
  ,�h x�  p�C     �       ���  -I_ x#�K  �
 �
 /��  y#'$  T0�B {�  ,�
 "�
 0�Y  |�  ��
 ��
 0��  }�  ,�
  �
 0J�  ~&	  �
 ֲ
 Hp ��  ?�
 +�
 0�k �&	  *�
 �
 0/� �&	  `�
 T�
 Hidx �&	  ��
 ��
  ,xb b&	   �C     I       �x�  /I_ b#�K  U-��  c#�  ݷ
 ٷ
 0�B e�  �
 �
 0�Y  f&	  S�
 Q�
 Hp g�  �
 w�
 0�k h&	  �
 �
 0/� i&	  ��
 ��
 Hidx j&	  z�
 x�
  ,h <\	   ED     �       �}�  -�B <$�  ��
 ��
 -��  =$�J  Q�
 E�
 Hp ?�  �
 ֻ
 0��  @&	  r�
 n�
 0/� @&	  ��
 ��
 1mED     E       F�  0J�  R&	  �
 �
 8�ED     . 9Uv 9T@  ;�ED     . c�  9Uv 9T8 8�ED     . 9Uv 9T8  ,�b �\	  ��C     $       ���  /I_ �$�K  U/�  �$�K  THp ��  ��
 ��
  @�d ��  �  AI_ �#�K  A��  �#'$  CJ�  �&	  FC�Z ��U    ,ys �&	  ��C     :       ���  -I_ �#�K  ʽ
 ½
 -��  �#�  2�
 ,�
 ;��C     �  ��  9U�U9T�t9Q0 <��C     ��   ,w\ �&	  `�C     P      ��  -I_ �)�K  ��
 }�
 -nf �)'$   �
 �
 -�W �)�  ��
 ��
 0��  ��7  �
 �
 0��  ��  =�
 ;�
 0�j �&	  q�
 o�
 0�k �&	  ��
 ��
 Hend �!&	  ��
 ]�
 0�  �&&	  ��
 ��
 0�� �	  !�
 ��
 Hmax �&	  ��
 ��
 Hmin �&	  5�
 -�
 Hmid �&	  ��
 ��
 0<R �&	  h�
 ^�
 0�_ �&	  ��
 ��
 0J�  �&	  ��
 l�
 Hp ��  ��
 ��
 :��  ��  Hi 
&	  ��
 ��
 :P�  p�  0PZ &	  ��
 ��
 0�q �  �
 �
  >��  0�j D&	  x�
 p�
 0gm D"&	  ��
 ��
   >p�  0�Z ��U  ��
 ��
 ;R�C     ��  ��  9Uu  ;��C     ��  ��  9Uu  8��C     m�  9Us    ,f ?&	  ��C     �      ���  -I_ ?)�K  ��
 ��
 -nf @)'$  *�
 &�
 -�W A)�  n�
 b�
 0��  C�7  ��
 ��
 0��  D�  �
 �
 C�j G&	  0�k G&	  T�
 P�
 Hend G"&	  ��
 ��
 0�  G'&	  ��
 ��
 0�� H	  H�
 @�
 Hi I&	  N�
 @�
 0<R I&	  ��
 ��
 0�_ J�  b�
 X�
 0J�  K&	  ��
 ��
 Hp L�  m�
 i�
 Hq M�  ��
 ��
 E]�  o>0�  Hr r�  ��
 ��
   ,�[ }\	  �>D     	      �m�  -�B }$�  W�
 A�
 -��  ~$�J  U�
 A�
 Hp ��  X�
 ,�
 0��  �&	  I�
 7�
 0�  ��  �
 �
 0�[ ��  ��
 ��
 0�f  � �  )�
 #�
 0_�  �*�  x�
 r�
 0
\ �3�  ��
 ��
 0<R �&	   �
 �
 0�U �\	  ��
 ��
 :��  �  0ei �&	  P�
 D�
 0�f �&	  ��
 ��
 0j �&	  d�
 \�
 ;�?D     . ��  9U~ 9T8 8�DD     . 9U~ 9T8  : �  ��  0�k �&	  ��
 ��
 Hend �&	  e�
 U�
 0�  �&	  ?�
 3�
 Hn �%&	  ��
 ��
 02\ �&	  ��
 ��
 0�Q �!&	  ]�
 S�
 0�� �	  ��
 ��
 0�r ��  o�
 a�
 0��  ��  0�
 "�
 0�z  ��  ��
 ��
 0�  ��  ��
 ��
 :@�  I�  Hi &	  d�
 b�
 Hidx &	  ��
 ��
 8CD     . 9Uv 9T@  ;AD     . h�  9U��9T8 ;�AD     . ��  9U��9T8 ;;BD     . ��  9U��~9T8 8dCD     . 9U��9T8  ;�CD     . ��  9U~ 9T8 ;�CD     . ��  9U~ 9T8 ;DD     . �  9U~ 9T8 ;-DD     . 6�  9U~ 9T8 ;EDD     . S�  9U~ 9T8 8�DD     . 9U~ 9T8  Sth  �C     W      ���  -I_ �U  .�
 �
 0��  �7  ��
 ��
 0��  �  �
 �
 0�_ &	  [�
 I�
 IWD  v��C     I�[ m`�C     >��  0
Q (�  2�
  �
 Hend )&	  �
 ��
 0�� *	  l�
 d�
 :��  ~�  Hp 1�  ��
 ��
 > �  0J�  :&	  ��
 ��
   :`�  ��  0J�  M&	  z�
 r�
  8o�C     ��  9Uu    ,d �	  ��C     '      ���  /I_ �!�U  U-�\ �!&	  ��
 ��
 0�B ��  �
 �
 Hp ��  U�
 7�
 0�  �&	  �
 �
 >@�  0�  �&	  C�
 9�
 4��C     0       0��  ��7  ��
 ��
 0��  ��  ��
 ��
    ,�g �\	  ��C     (       ���  /I_ ��U  U/�B ��  THp ��  '�
 %�
  ,�S G\	  ��C     $       �9�  /I_ G$�K  U/�  H$�K  THp J�  N�
 L�
  ,T ��  0�C     ]      ���  -I_ �#�K  w�
 s�
 -nf �#'$  ��
 ��
 0�B ��  ��
 ��
 0J�  �&	  �
 �
 0�Y  ��  ��
 ��
 0�_ ��  ��
 ��
 0�p ��  t�
 j�
 I�  ?��C     I{e 8��C     :��  ��  Hp ��  ��
 ��
 0�k  &	  ��
 ��
 0/� &	  �
 �
 0�� 	  w�
 o�
 0�  &	  7�
 /�
 0DQ &	  ��
 ��
 Hpos &	  g�
 e�
 Hidx &	  ��
 ��
  ;[�C     -�  ��  9Uy 9Tx  8��C     -�  9Uy 9Tx   ,_ �&	  ��C     �       �-�  -I_ �#�K  ��
 ��
 -��  �#�  9�
 3�
 0�B ��  ��
 ��
 0�Y  �&	  ��
 ��
 0�p ��      1��C     z       �  Hp ��  l  `  Hidx �&	    �  0�k �&	  � � 0/� �&	  n d 0�� �	  B < 0�  �&	  � �  8��C     -�  9Tx   ,�p ��  0�C     `       ��  -�B �&�    -��  �&�  a [ O�Y  ��   I�  ���C     >��  0DQ �&	  � � 0s �&	    Hp ��  � � 0+ ��   	 Hsub ��  2 .   ,�o '\	  p<D     v      �k�  -�B '$�  | h -��  ($�J  e Y Hp *�   � 0��  +&	  4	 ,	 Hn -&	  �	 �	 0� -&	  C
 9
 0�Q .�  �
 �
 0+ /�  @ < 0
\ 0�  � v :0�  �  Hidx C&	   � 8=D     . 9U~ 9T8  :`�  �  0=` Z&	  � � 0�b Z&	  � � 0�  Z(&	  ] [ 0�� [	  � � :��  ��  Hids q�  - + :��  ��  0��  {�  R P Hidx |&	   u 8�>D     . 9U~ 9T@  8>D     . 9U~ 9T9  8�=D     . 9U~ 9T8  ;(=D     . 4�  9U~ 9T8 ;�>D     . Q�  9U~ 9T8 8�>D     . 9U~ 9T8  TP\ �\	   �C     $       ���  jI_ �$�K  Uj�  �$�K  TXp ��  = ;  T�b ��  ��C     3       �K�  jI_ �#�K  Uj��  �#'$  TV�B ��  f b V�_ ��  � � V�Y  ��  � � VJ�  �&	      T=i �&	  ��C            ���  jI_ �#�K  Uj��  �#�  TV�B ��  � ~  _ \ `\	  ��  `�B `$�  `��  a$�J  bp c�  a��  d&	  Fbn s&	  bidx s&	    T(r ?\	  ��C            �5�  jI_ ?�K  Uj�B @�  T T2p 	�\	  P�C           �b�  U��  	�,�7  � � U�1  	�,=  A 5 U�Z 	�,GJ  � � Xbdf 	��7  c W Vֳ  	��    � V�U 	�\	  _ I Xp 	��  Y K V/� 	�&	  � � V�n 	��  : 4 VhV 	�{	  � � e�  	�^�C     W�Z 	�:��  g�  V� 	�&	  � � V.� 	�&	  � �  :�  ��  Vb 	�&	   � >@�  VE- 	��   } V<v 	��  � � ;��C     . ��  9Uv  8'�C     . 9U��9T0   hb�  {�C       p�  	�M�  3�    3s�  j d >p�  5��  � � K��  ��5��  � � \��  6��  ��C     7��  ��C     �       ��  5��  a S 5��    � 5��  < 8 5��  z x 5��  � � 5��  � � ]�  `�C             5�  � �   ;��C     ?�  �  9U} 9T FDB9Q��9R�� ;��C     	- /�  9U��9Q~  8��C     - 9U��9T~    8��C     (. 9Uv   _"g 	>\	  �  `��  	>&�7  `^�  	?&e  bbdf 	A�7  a��  	BC	  a�U 	C\	  W�  	�W�c 	�Fbp 	T�  a��  	U&	  acC  	V&	  a�y 	WC	  a/� 	X&	  a�n 	Y�  Fa� 	o&	     kr 	)J�  `��  	)$�7  bbdf 	+�7  Fa^�  	0e    _d ^\	  ��  `^�  ^e  `��  _�7  aڰ  a�  a�U b\	  a�a dA  a�R  ezA  aZL  f��  arP hC	  a�i  j�  asj  ke  afP m�  a�] nC	  bnn p	  af qC	  &UV s"��  	�	G     E�  �[U�  a�f �&	  aU �&	  a�X �,&	  bx �8&	   [g�  a�B �zA   [z�  C�B zA   FC�B UzA  FCo oC	     	zA  T4l GG   p�C            �*�  pa G!U  Upb H!U  TVXP JzA  � � V_P KzA  � � V�\ MC	  � � V�\ NC	   
  cUX 9 D     )       �~�  U^�  9!e  9 3 Vڰ  ;�  � � <0D     J-  S*q C D     �      ���  -��  C�7  � � 0ڰ  E�  + ' 0�i  F�F  e a :��  �  0^�  re  � � 8	D     - 9Ts�  M�  �D      p�  c��  3#�  � � >p�  5/�    � ];�  �
D     H       5<�  W U 8�
D     - 9Ts�
    MĚ  �D      ��  g��  3њ  ~ | >��  5ݚ  � � 8�D     - 9Ts�
   YRD     ��  9Us  YdD     ��  9Us  YvD     �  9Us  Y�D     %�  9Us  ;�D     J- =�  9Uv  ;�D     J- U�  9Uv  ;Y	D     J- m�  9Uv  Yz	D     ��  9Us  ;�	D     J- ��  9Uv  ;�	D     J- ��  9Uv  ;�	D     J- ��  9Uv  ;�	D     J- ��  9Uv  ;�	D     J- ��  9Uv  ; 
D     J- �  9Uv  ;
D     J- )�  9Uv  ;4
D     J- A�  9Uv  ;N
D     J- Y�  9Uv  ;h
D     J- q�  9Uv  ;�
D     J- ��  9Uv  8�
D     J- 9Uv   ,�e �\	   0D     g      ���  -^�  �"e  � � -��  �"�7  �  �  -�' �"	  )" !" -�[  �"	  �" �" -\  �"�  �" �" '�U �\	  ��02Y �\	  q# _# 0xf ��  D$ <$ 0�a ��  �$ �$ 0�a ��  ?% 9% 0�` ��  �% �% 0^ ��  �% �% 0�V ��  J& B& 0ua ��  �& �& 0�i  ��F  ' �& I�  61D     :��  &�  Hi �	  �' �'  :��  �  0ah �  �' �' 0�1  �7	  �( �( :��  J�  Hm M	  �) �) 0�^ O�  ;* 5* :��  ��  0�� U�  �* �* =� w6D       0�  X3	 �* �* 3� �* �* >0�  5�	 + 	+ 5�	 P+ L+    4~:D     O       'a�  e�  ��8�:D     �- 9U	@G     9T09Q| 9R0   :`�  ��  0/� �&	  �+ �+ >��  0ڰ  ��  �+ �+ 0Mp  �		  F, :, 04` ��  �, �, '�e �[  ��0:W  �o?  B- 6- 0�P �&	  �- �- 0Ue �!&	  #. . :��  7�  0�d  �w  r. p. N�7D     9Uv 9T~ 9Q|   ;B7D     V- n�  9U��~9T 9Q09R~ 9X09Y�� ;n7D     V- ��  9U��~9T49Q09R~ 9X09Y�� 8�8D     V- 9U��~9T49Q��~9R��~9X��~9Y��   MY�  �3D       P�  C�  3j�  �. �. 3j�  �. �. 3v�  �. �. >P�  5��  V/ R/ 5��  �/ �/   qY�  �3D            ��  Jj�  Jj�  Jv�  4�3D            5��  �/ �/ ?��    MY�  �3D      ��  ��  3j�  0  0 3j�  0  0 3v�  '0 %0 >��  5��  S0 O0 5��  �0 �0   8H6D     s�  9U   MY�  �4D        �  o�  3j�  �0 �0 3j�  �0 �0 3v�  1 1 > �  5��  t1 p1 5��  �1 �1   qY�  (5D     (       ��  Jj�  Jj�  Jv�  4(5D     (       5��  G2 C2 ?��    qY�  Z5D     #       �  Jj�  Jj�  Jv�  4Z5D     #       5��  2 }2 ?��    Y�0D     9�  9U 9Txibs9Qv 9R0 Y�0D     S�  9U 9Tv  Y�0D     {�  9U 9TCLBC9Qv 9R0 Y1D     ��  9U 9TTDBC9Qv 9R0 Y?1D     ��  9U 9Tv  YL1D     ��  9U 9Tv  YY1D     ��  9U 9Tv  Yf1D     �  9U 9Tv  Y�1D     *�  9U 9Tv 9Q0 Y�1D     I�  9U 9Tv 9Q0 Y�1D     h�  9U 9Tv 9Q1 Y�1D     ��  9U 9Tv 9Q1 Y�1D     ��  9U 9Tv  Y$2D     ��  9U 9Tv  Y<2D     ��  9U 9Tv  YL2D     ��  9U 9Tv  Y\2D     	�  9U 9Tv  Yi2D     #�  9U 9Tv  Yz2D     >�  9U 9T�U ;�2D     �	 a�  9U 9T19Qv  Y4D     {�  9U 9Tv  ;P4D     �	 ��  9U 9TE9Qv  ;�4D     �	 ��  9U 9TF9Qv  ;�4D     �	 ��  9U 9T2 Y�8D     �  9U 9Txibs9Qv 9R0 ;�:D     �	 )�  9U 9T@9Qv  ;g;D     �	 L�  9U 9TA9Qv  ;�;D     �	 o�  9U 9T19Qv  ;�;D     �	 ��  9U 9TA9Q0 8B<D     �	 9U 9T@9Qv   ,@Y �\	  `_D     K      �[ -^�  �"e  �2 �2 -��  �"�7  44  4 -�' �"	  5 5 -�[  �"	  ~5 v5 -\  �"�  �5 �5 0�U �\	  N6 J6 0�-  �   �6 �6 0�i  ��F  
7 �6 0�  �	  h8 \8 :` ��  0ϖ ��  �8 �8 06e  �n	  %9 !9 8�_D     4. 9T	׷F     9Q1  1@gD     @       V�  05a ��  ]9 [9 ;MgD     A. 5�  9Us 9T	��F      8\gD     4. 9T	��F     9Q0  1gD     (       ��  05a ��  �9 �9 ;%gD     A. ��  9Us 9T	��F      84gD     4. 9T	��F     9Q0  :�	 � 0ڰ  (�  �9 �9 '�q *C	  ��~0��  ,C	  : : 0�  -C	  K: E: 0�  /		  �: �: 0)�  0		  �: �: 0��  1		  H; 4; 0ga 2		   < < 0�' 4	  }< m< 0nZ 6�  A= += 0Q 7�  >> *> : 
 ��  0(o qC	  ? ? 0�[ rC	  Z? T? 04Q r)C	  �? �? Hp t�  �? �? Hi u&	  u@ m@ ;hD     =- 8�  9Us  ;�hD     �- a�  9Us 9T| 9Q} 9R4 ;-iD     �- ��  9Us 9T| 9Q~ 9Rv  8?iD     N. 9U 9T~ 9Qv   Y#fD     ��  9U} 9Travf9Qs 9R��~ ;dfD     J- ��  9U| 9T  ;ofD     J-   9U| 9T~  Y�fD     :  9U} 9Tfylg9Qs 9R0 Y�fD     b  9U} 9T2FFC9Qs 9R0 Y�fD     �  9U} 9T FFC9Qs 9R0 ;�gD     �- �  9U| 9T��~9Q��~ ;�gD     �- �  9U| 9T��~9Q��~ ;]jD     �- �  9Us 9T��~ ;{jD     |-  9Us 9T��~ ;�jD     �- 7 9Us 9T2 ;�jD     |- W 9Us 9T��~ ;�jD     |- w 9Us 9T��~ ;kD     |- � 9Us 9T��~ 8AkD     |- 9Us 9T��~  M[ �_D      �  3z �@ �@ 3m �A �A >� 5� �B �B K� ��~5� �C �C 5� �C �C 6�  `D     MJ�  K`D      @ {� 3g�  yD mD 3g�  yD mD 3[�  E �D >@ 5s�  �E �E K�  ��~K��  ��~5��  aF MF 5��  MG 7G 5��  JH 8H 5��  6I I 5��  kJ WJ 5��  lK <K 5��  zM lM 5��  )N N 5��  &O O 6�  WaD     Lz�  � � 5{�  �O �O L��   _ K��  ��~8�oD     Y. 9Us 9Q��~  ;PoD     �, w 9U  ;ioD     �, � 9U  ;�oD     �, � 9U  <wpD     �-  L!�  P � ?&�  52�  BP 8P 5>�  �P �P 5J�  �P �P  LU�  � � 5Z�  �Q xQ ;�cD     �, ! 9U  ;�cD     �, 9 9U  ;dD     �, Q 9U  ;dD     �, i 9U  ;dD     �, � 9U  8AdD     �, 9U   Lg�  	 � 5l�  R R  ;i`D     �- � 9U 9T	�	G     9Q��~ ;:aD     �- � 9Us 9Q��~ ;baD     J-  9Us  ;naD     J- 3 9Us 9Tw  ;BbD     �- X 9Us 9TP9Q��~ ;cD     V- � 9Us 9T09Q09X09Y��~ ;JcD     V- � 9Us 9T89Qw 9Xw 9Y��~ ;ycD     �, � 9U  ;cdD     J- � 9Us 9Tv  ;kdD     e.  9U~  ;vdD     J- % 9Us 9T~  ;QlD     �, = 9U  ;llD     r. h 9Uw 9Q89R	p�C      ;EnD     V- � 9Us 9T19Q��~4$#9R��~9Xv 9Y��~ ;,pD     ~. � 9U~ 9Tv  <SpD     �.   L� @	 � 5� BR >R ;�aD     �-  9U 9T	�	G     9Q}� ;�iD     V- I 9U��~9T89Q09X09Y��~ ;�iD     �, a 9U  ;�iD     �, y 9U  8�iD     �, 9U   ;`D     =- � 9U  ;`D     �- � 9U 9T��~ ;?`D     �, � 9U 9Ts  8UeD     �- 9U��~9T89Q��~   ;�dD     �. , 9Us 9T	��F      ;�eD     �, D 9Us  N�eD     9U} 9Ts   @�` W\	  � A^�  We  A��  X�7  Cڰ  Z�  C�U [\	  Dtag \C	  C�  \C	  '
i ^"�  	�	G     E)f nFDn �	    @T "�  �	 A�!  "G   A"  #G   Y %N	 �!  'G    "  (G   T )�   �] +	 N	 [	 p	 @   
 `	 'Tb .p	 	 
G     Dcur @�	 	[	 C��  @�	  TUo �\	  �D     �      �� U��  �"�7  �R yR Uhq �"		  3S %S U}W �"�B  �S �S Vڰ  ��  <T 8T &�U �\	  ��V�Y  �q  ~T rT Xn �		  U U Xrec ��2  �U �U V^ �	  �V �V V�\ �	  �W �W VVc �	  �W �W V�Y �	  �X �X VV �	  KY ;Y V�d ��  �Y �Y Va �U  �Z oZ I�  +D     1�D     �       � 0^�  
e  k[ i[ ;�D     V- _ 9U| 9T 9Q09X09Y�� ;D     �, w 9U~  ;D     J- � 9U|  8ED     b- 9U~   ND     9Us 9T|   TBd \q   �C     �       �� U�, \(�2  �[ �[ Uڰ  ](�  �[ �[ V�: _q  #\ \ Xlen `&	  s\ m\ V�* `&	  �\ �\ Xn `&	   ] �\ V�K a�  �] �] &�U b\	  �\8K�C     V- 9U�T9T19Q09Rs����9X09Y�\  T<X 9q  ��C     �       �� U�, 9(�2  �] �] Uڰ  :(�  ^ ^ V�: <q  e^ _^ Xlen =&	  �^ �^ V�* =&	  _ �^ Xn =&	  B_ 8_ V�K >�  �_ �_ &�U ?\	  �\8�C     V- 9U�T9T19Q09R|����9X09Y�\  ,)e ��  `�C     
       � -ϖ �$�  ` ` -2*  �$=  S` O` Rj�C     �. 9U	�G     9T�T  ,Hp V\	  p�C     t       �� -��  V&�7  �` �` -�7 W&J  ,a  a -n/ X&J  �a �a 'T Z�I  �@':�  Z �I  �P0�U [\	  Pb Hb ;��C     5�  � 9Us 9T	��F     9Q�P 8��C     5�  9Us 9T	��F     9Qw   @jc =  M A��  �7  C�  	  Dwin 	  C^ 	  C�Y  =   @�V =  � A��  "�7  C�U \	  Cڰ  �  Dmm �P  C�  &	  CԚ  �  C;�  �N  C�  	  Dwin 	  C^ 	  Di &	  Dj &	  C�Y  �   Dp �   Eek �E�q �[3 Dlen $&	   [� C�i  z�F  C��  |7	  C�}  }&	  CO�  �   FCcy  �&	  C�U ��   Ds ��     [� C�~  ��0  FDt ��     FC��  ��  C��  �� Dh �'$  FDv �     �  � @    @\ ��   n A#�  �	  Bbuf ��   Dp ��   Dq ��   Dtmp �n C�q �	  C�i �	  Di �	   �   ~ @    ,/P _�  ��C     �       � -��  _ �7  �b �b Pid ` 		  T.win a PD  �b �b /^ b PD  RHn d	  Bc <c >��  0}W l�2  �c �c   @xd $�   � Aڰ  $%�  A^�  %%e  A�, &%�2  A�P '%�P  A�W (%�  C�U *\	  C�Y  ,�   Dr -q  Dp .e6  Dlen /&	  E�U S @�Q ��   K Aڰ  �#�  A^�  �#e  A�, �#�2  A�P �#�P  A�W �#�  C�U �\	  C�Y  ��   Dr �q  Dp �e6  Dlen �&	  E�b  Q�f )� Bkey )*U  Blen **Z   A��  +*�  Bout ,*_   CKl  .�  C�] /N   Dh1 1�  Dh2 2�  Dh3 3�  Dh4 4�  Dc1 6�  Dc2 7�  Dc3 8�  Dc4 9�  C� ;� Di =
G   [U Dk1 B�  Dk2 C�  Dk3 D�  Dk4 E�   FC�
 n�  Dk1 p�  Dk2 q�  Dk3 r�  Dk4 s�    	�  @r �  � Bh �   ,�W G   ��C            �� .c G   d 	d  T�c �G   p�C     "       �2 pc �G   UXcc �S   Gd Ed  T
m �&	  �XD     �       �� U��  �*  rd jd U{ �*�  �d �d V�H  ��7  @e 8e Xi �&	  �e �e VV �&	  �e �e 4 YD     /       &��  �q  �HV�U �\	  /f -f ru   YD       YD            �� 3<u  Xf Rf 3/u  �f �f 3"u  �f �f 4 YD            ?Iu  ?Vu  ?cu  ?pu  \}u  8YD     r 9Uv 9Ts 9Q�H   8+YD     �. 9U}    _bg �\	  � `��  �$  `x �$&	  `_| �$n	  `�H  �$&	  a��  �q  a�U �\	   _�X }\	  A `��  }�7  iidx ~&	  itag J1  `�  �J1  `��  �J1   TgX P_   ��C     �       �� j��  P �7  Ugtag Q �.  �f �f V�B S_   4g ,g  s� 0PD     V       �6 t U3 �g �g t Qt( Rt4 X]� TPD     ,       34 �g �g 3( 	h h 3 .h ,h 3 Uh Qh 3 �h �h   s��  �PD     U       �L 3��  �h �h 3��  mi _i K��  P1�PD            � 5�  j j R�PD     ��  9U�U9T�T9Q1  7��  �PD            8 3��  �j �j 3��  �j �j 4�PD            5��  k k ]r �PD            ?�  8�PD     m�  9Us     R�PD     �  9Q1  s��  �PD     ?       �� 3��  /k )k 3��  �k {k 5��   l �k K�  PL��  0 � 3��  Pl Ll 3��  �l �l >0 ?��  5�  �l �l 8QD     ��  9Uu    RQD     ��  9Q1  s��  0QD     ?       �� 3��  �l �l 3ȿ  /m %m 5տ  �m �m K�  PL��  ` � 3ȿ  �m �m 3��  5n 3n >` ?տ  5�  Zn Xn 8ZQD     ��  9Uu    RHQD     ^�  9Q1  s!�  pQD     \       �r 33�  �n }n 3@�  o �n 5M�  �o �o L!�  � K 3@�  �o �o 33�   p p >� 5M�  [p Yp \Z�  8�QD     	- 9Uv 9Qs�   N�QD     9Us 9Tpamc9Qv 9Rs�  uu  @WD     Q      �� 3"u  �p ~p 3/u  }q iq 3<u  hr Tr 5Iu  Cs ?s 5Vu  �s ys 5cu  vt jt 5pu  u �t \}u  L�u  � C 5�u  �u �u 7�u  �WD     /       . 5�u  �u �u  8XXD     �v  9Us   L�u    r 5�u  �u �u 8�XD     �v  9Us   YjWD     � 9U0 N�WD     9U}   su  �XD     &       � 3"u  3v -v 3/u  �v v 3<u  �v �v ?Iu  ?Vu  ?cu  ?pu  R�XD     r 9U�U9T�T9Q�Q  s� �YD     r       �� 3� )w #w 3� {w uw 3� �w �w 3� gx [x ?� ?� hu  �YD      ` �� 3<u  �x �x 3/u  y y 3"u  qy ky >` ?Iu  ?Vu  ?cu  ?pu  \}u    ^� � 3� �y �y 3� z z 3� az [z 3� �z �z >� K� �X5� { { vu  �YD            �� J<u  J/u  J"u  4�YD            ?Iu  ?Vu  ?cu  ?pu  \}u  8�YD     r 9U�U9T�T9Q�X   8�YD     �. 9Uv 9Qs ����    s��  �]D     B       �� 3��  ^{ T{ 3��  �{ �{ 3Ő  m| g| 5Ґ  �| �| ?ߐ  L��  � � 3Ő  �| �| 3��  } } 3��  ^} X} >� KҐ  P5ߐ  �} �} \�  R2^D     �- 9U�T9T	@G     9Q�U#�   N
^D     9Us 9T�Q9Qv 9R0  s(�  `^D     �       �! 3:�  ~ ~ 3G�  �~ �~ 5T�  � � ?a�  L(�   �  3G�  � � 3:�  \� R� > 5T�  ހ Ԁ 5a�  U� M� \ʈ  ;�^D     �- q  9U| 9T	�G     9Q}  ;_D     �- �  9U| 9T	�G     9Q}  ;(_D     �- �  9U| 9T	`G     9Q}  RT_D     �- 9U�T9T	PG     9Q�U#�   N�^D     9Us 9T2/SO9Q| 9R0  s��  �pD     �       �A" 3��  Ł �� 3��  l� `� 5��  �� � 5��  |� x� 7��  �pD     :       
" 3��  �� �� 3��  � � 4�pD     :       5��  "�  � ?��  ]��  �pD     :       5��  K� E� 5��  �� �� 8/qD     . 9Uv 9T@    ;MqD     . '" 9Uv 9T8 8\qD     . 9Uv 9T8  u �uD           ��# 3) � �� 36 m� c� 3C � �� 3P O� G� Kj ��5w �� �� 5� D� >� 5� �� �� 5� �� � 6� IvD     3] L� J� ;�uD     �- # 9Uw 9Q�� ;�uD     �, # 9U  ;�uD     �, 7# 9U  ;IvD     �, Q# 9U�� ;[vD     J- i# 9U~  ;uvD     J- �# 9U~  8�vD     �, 9U��  u� �vD     1      ��$ 3� |� t� 3� � ܈ 3� a� Y� 3� ȉ �� K ��5 3� '� 5 �� �� 5) � � 54 p� l� 6A �wD     3� �� �� ;�vD     �- ^$ 9Uw 9Q�� ;wD     �, v$ 9U  ;!wD     �, �$ 9U  ;�wD     �, �$ 9U�� ;�wD     J- �$ 9U~  ;�wD     J- �$ 9U~  8�wD     �, 9U��  s� �wD     G
      ��, 3 �� Ћ ? ?% ?2 w?  7� ExD     �       & 3 �� �� 4ExD     �       5 ܌ ڌ K% ��K2 ��5? � � ;\xD     ~ �% 9Uv 9Tt 9Q��9Rr  ;�xD     A" �% 9R	p�C     x] 1 8�xD     �# 9R	p�C     x� 1   yM �xD      �xD     O	      #3_ F� >� 4�xD     O	      Kl ��5y �� �� 5� ύ Ǎ K� ��K� ��K� ��5� 3� +� K� ��K� ��5� �� �� 5� 4� 2� 5� r� X� 5 �� |� 6 �|D     6 PzD     L3 �
 �' 58 �� � ?E 5R C� =� K_ ��Ll  �' 5m �� �� Kz ��5� �� �� Y�yD     p' 9Uv 9Q�� <�yD     (. ;�yD     �- �' 9U~ 9Q�� ;�yD     �. �' 9U|  8HzD     J- 9U~   Y~D     �' 9Uv 9Q�� 86~D     (. 9U   L� @ �( 5� � ؓ L� � �( 5� ]� Q� =� �zD         �3 � ߔ 3 S� I� >  5% �  50 {� i� K; ��5H >� 6� 5U �� �� 5b �� r�    ;tzD     �- �( 9U~ 9Q�� <�zD     �.  L� � `+ 5� X� R� K� ��5� �� �� MK �|D      � �<+ 3s !� � 3� �� �� 3f � � 3Y �� z� >� 5� � ޜ 5� 9� -� 5� 
� �� 5� �  � 5� � �� 5� Ӡ �� 5� �� �� 5� � � 5� r� l� 5� Т ʢ 5 0� (� 5 �� �� 7 �|D     �       K* 5$ У ƣ 50 ~� r� 5< 7� 3� 5H {� o�  LU @ �* 5V 6� 0� 5c �� � 5o S� C� 5{ � � 5� ި ʨ  M� D      � �
�* 3� �� ��  M� aD      P �
�* 3� �� ��  M� iD       �
+ 3� 3� 1�  =� }D      ` �
3� Z� V�    ]� �D     '       5� �� ��   L  � \, 5% �� �� ;׀D     ~ �+ 9Uv 9Tt 9Q��9Rr  ;�D     �# �+ 9R	��C     x� 0 ;�D     (. �+ 9U|  ;��D     A" 	, 9R	��C     x] 0 ;ׁD     ~ 4, 9Uv 9Tt 9Q��9Rr  8��D     ~ 9Uv 9Tt 9Q��9Rr   NyD     9Uv 9T��9Q��9R09X��    zM  M  �{�X �X 1N{�i �i 1�z�O �O 1>z[l  [l  �z@G  @G  �z�]  �]  �z�a  �a  �zKS  KS  �z�<  �<  �z]>  ]>  �z!`  !`  �ze  e  �zva  va  �z�Z  �Z  �{�s  �s  2�{�I  �I  2�z�D  �D  �z�k  �k  �zHg  Hg  �zw  w  �zd  d  z�^  �^  �z�[  �[  �{�`  �`  2v|BY  8Y  3 |D  D  3 z2n  2n  {�k  �k  (k{�p �p '{�r  �r  (z{��  ��  4{��  ��  4"{Ne  Ne  42z�b  �b  8z$i  $i  -|/�  %�  3 {=\ =\ 5�z~l  ~l  |{�  �  6Xz)p  )p  vzO  O  qz�?  �?  4zF>  F>  k{�  �  4zu  u  2y{j�  j�  4 �  +[  m&  �� �:  @�D     ��      �� K�  (\  �@   K,  i   �S   K�  nint o.�   @�   
�  �    
p   	G   
�  #	G   
X  &	G   
�  )	G    
�  ,	G   (
�  -	G   0
/  2Z   8
�  5Z   < �   K�  #�   �  8"c   	+  K  �   	%  L  	�  M  K'  K;  K�  s&  Z   �  -   )  A"i  o  .�   ��  
�  �a    
��  ��  
<h ��  
�I  ��   �  X�  �  $a   �  ]  @    �   m�  �  0�  ]  a    f  �    $a   )  ]  @   @   a    J   �"5  ;  �  PH�  Ǟ  J8   ֳ  KS   ?pos LS     N�  /[  O�   �K P  (�R QE  0ڰ  S]  8O�  T8  @��  U8  H p�  ��  c<v �@   c��  �a    �  ��  ""  �    $S   8  )  S   8  S    >  K�  �   R  X  0c  )   v  :@   .�  L�  1x Nc   1y Oc   �  Qo  #�  .~   w�  

  yc   
�!  yc  
�   zc  
H  zc   "  |�  �  (q  M} -    5�  -   `�  	Z   _| 
8  
!  <  ?   >  2   >  B  a     �  �  #q  �  (Q�     S5   0�  T5  N5  V�  �   W�   H� X�  �1  ZZ     �  5  �  \�  �  J�  -   �C  �!   /�   pmoc/�  stib/u!  ltuo/�  tolp :  �  �8  5"]  c  ^�$  �4  S�  ?x U5   ?len V<  e� W>   �#  Yh  #�  �%  {�  �  0�  Z   Z   �  a    �  �#  ��  �  $Z     Z   Z   a    �.  �  #  08  Z   Z   a    �8  `��  .   �   �; �  �1  Z   �5  �  �+  �   `(  �  (�/    0�  a   8*  �  @ ~  �  qu(  
8  #�  �2  (�  �  $Z     a      P  �3  ;  $  0/  P   v)  ]<  B  0W  P  8  S    �3  yd  j  $Z   �  P  S   a    H7  ��  �  $Z   �  P  �   �  51  0�  y2  �C   � ��   �/  *
 �W  / ��   $ �  ( 2$  ��  -4  l>  +  �8  K�  $8  �>  #?  K    ��   #V  {"  �5  !  �<  \   �Z   �  �-   }  �@   )$  �S   �   @   c,  +Z   C*  6a   +D  CG   �]  P4    :   �3	  ?xx ��   ?xy ��  ?yx ��  ?yy ��   5  ��  #3	  8  �p	  ��  �P   ��  �   $  �E	  c   ��	  �	  0�	  a    �  ��	  Kl  �a    �  �}	   s  ��	  �"  $�	  �	  �   +
  �� -�	   �W .�	  Kl  /a    %  DJ
  uR F�	   �
 G�	   }  I
  d-   (��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<  5�  >c   ��  ?c  �"  Ac  �"  Bc  i!  Cc   %!  Ec  (2!  Fc  0�  Gc  8   I�  �"   s{  ��  ug   5�  vg  ֳ  xc  !  zc  m  {c   v  }&  J  �#�  �  Z�!  �}Y  ڰ  ]   {3  �  S0  �  �/  �  �1  ��  �1  �#  6Y/  �J
  6�*  ��  (6�)  �Y  06+:  � #  86<8  �0#  X6�*  �  � �3  �"f  l  �(  ��  Oe ��"   �-  ��  ڰ  �]   U  �"�  �  �  8�  ah !�"   Oe "�  U1  #J
   ;+  $�  0 i(  �$    l;  ���  ah ��"   Oe �
#  y2  �C   {:  �0  (�� �P  h/ ��  p�� ��  x T   � �  �  _  �W  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"    8�  �  @`  !  Hd  "�  P�@  $�	  X�;  )�  h�   +s  ��  ,g  �
  -g  ���  .g  �?!  0g  ��  1g  ��  3g  ��  4g  �ȩ  6�  �ֳ  7W  ��� 8  �K <�  �ڰ  =]  �^�  >)  �U  @J
  �t  B�	  �k  Ca   ��L  E:  � "   d  j  1  Xm�  ��  o�   �@  p�	  �e q�  �L  r�  P @  $%�  �  Z  0\  �-  ^�   ��  _�  �W `�  x a�  �@  b�	   �e d  0�"  e�  pi"  f�  x� g�  ���  iC  �.a kq  ��  l  �J  m  �Mj  o�  ��  q�  ��  r�  �6M  ta    6Z  u@   6_"  wc  6(   xc  6Ud za    6�L  |  ( �!  F#  !  Z!  Ah  ��  C�   T D-  �!  Es  "  Fs   JS  -   �-  Y   /�  bmys/�  cinu/�
  sijs/    bg/�  5gib/F  snaw/  ahoj/�    bg/�  sijs/=    bg/�  5gib/�
  snaw/k  ahoj/�  BODA/t  EBDA/�  CBDA/  1tal/�  2tal/�   nmra �  h  0  `)G  M  �"  �e�  �1  g3	   H+  h�   x+  i  0��  km!  8�)  n#�"  h�'  q,  p��  rC  t�*  y  x V  {    �  �)�  �  �!  H�*  $  �a    7:  ��  s4  ��   b  8H�  !  Js   m  Ks  A� M�  �� N�  �  Pc  
  Qc   ��  Rc  (�  Sc  0 �  U*  x   �$�  �  .�!  0'  
ad  )   
�1  *s  
&D  +  
2B  ,  
x� -3	     �)%  +  �"  P��  ��  ��   �1  ��  �&  �   �3  �3	  ]7  ��  0�7  �a   @�1  �C  H P6  �  ?tag �   Kl  �   �6  	�  �  J�5  -   
  i7   �&  9  F9  8%  �*   �,  
�  ./   6
t  b 8
   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�    J�8  -   ��  �:   4,  �6  $  �/  l9   �2  ��  J�[  -   �   Y   zS  �e   ti  �M   �#  ��  �'  �    $�  +  Y   �2  �7  =  0H  Y   l/  �T  Z  $�  n  Y  n   �   .;)  H��  
�#  ��   
:  ��  
�5  ��  
F1  ��  
,8  ��   
2*  ��  (
�*  �
  0
`1  �+  8
��  �H  @ b  �-  �t  #�  d)  s  !  $�  0  a    9  F#A  #0  .�$  @J�  
�#  L�   
y2  MC  
W� O  
�� P7  
�,  Q�   
M4  RT  (
�;  S�  0
�*  T�  8 c/  X!�  �  .�-  (q  
�-  s�   
Oe t  
��  uC  
� v�   <  �/  )  #  $�  7  �  �   g%  .C  I  0T  �   �.  1`  f  0{  �  {  �   @	  73  6�  �  0�  �  �   �  �8  :�  �  $�  �  �  �   "3  >  $)  Y�  �  $�    �  �  �  �   �6  _    $�  ;  �  �  {  �   �3  fG  M  0b  �  �  �   ;0  ln  t  $�  �  �  �  �   .�&  x��  
ah � �   
y2  � C  H
�8  � �  P
�8  �   X
�'  � ;  `
� � b  h
�9  � �  p   �.  ��  ."9  H2W  
Mj  4�   
H5  5�  (
�)  6�  0
�  7�  8
�  8�  @ �0  :  .T%  �=�  
ڰ  ?]   
�0  @�  
q5  A�  
L)  B�  
)  C   
Ǟ  EW  
�  FW  `
Ud Ha   � X+  J�  c  1  �  �  $�     )  �      �   �&  &,  2  0=  �   �1  *I  O  $�  ^  W   �6  -j  p  0{  W   w-  1�  �  $�  �  �   �;  4�  �  0�  �   =;  8�  �  $�  �  W  t   B$  <�  �  $�    W  �   2  @    $�  5  �  W  �  C   7  GA  G  $�  e  �  �  �  �   q8  Nq  w  $�  �  �  )   )2  S�  �  $�  �  �  �  �  C  �   �  .k.  ���  
ah ��   
#,  ��  H
�4  ��  P
,;  ��  X
EY ��  `
/q �   h
Z)  �=  p
�#  �^  x
'0  �{  �
.  ��  �
��  �  �
� �5  �
`9  �e  �
��  ��  �
5  ��  �
U#  ��  � �2  ��  �  0t  P&�  �  ^�h  �V  m�  �  0�  �  �  �  �   a   @   EU  �      0'   �  a    j]  �3   9   0I   �  �   �l  �U   [   $�  ~   �  �  W  �  C   .t>   ��   
�=  �$'    
[I  �$�  
�d  �$   
��  �$I    � �~   #�   .8S  ��   
�d  �n   
�W  ��   C  ��   #�   �&  0�m!  y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  �
!  *  V'�!  �!  ^�0  .�*   u�!  
|#  w�   
�#  x�  
� y�  
C4  z�   �&  |�!  �'  ��!  �!  $�  
"  z!  �  
"   p	  �9  �"  ""  02"  z!  
"   A2  �>"  D"  $�  b"  z!  �     b"   �!  8(  �"  ��  )�!   $�  )"  �-  )2"   )  h"  #�"  3  <�"  �� >%�"   ��  ?%z!   �"  #  A�"  �"  �  �(  �l  �  %Y   #  +S    %  0#  +S    %�  @#  +S    H'  �%  _�� -   N�(  ��  ۻ ޫ (�y A�x i	� {�� �4� �(� �T� ��� �"� �v� c� � .Y� 8�� X�� x�� �>� ��� �� �ԕ �� ��  � 4�� T�� t�� �e� �E� �� �!� i� 4� M{� ��� �#� ��� �Μ �e� 0� >Q� ^(� ~}� ��� �� ��� ��� ��  � )�� BЎ [�� t� ��� �� �&� �jv �ߐ ˂ 5�� U�u un� ��� �	� �Z� �2� �� 5> U?� u�� �C� ��� ��� � x �� 5[� ]�� q-� �$� �)� ��� �Ջ ��y ��� 	'� L	�� m	�x �	� �	� �	̾ �	�� 
[� 
� -
Z� ?
�� N
φ z
!� �
1� �
W� �
;� �
�� �
�� �
�� ͨ /}� O�� qk� ��z �1y �(w �$� �� (�� 4�� L� \m� l� z4� �Y� ��� ��z ��� ��� �"t ù �� 7ɲ TɊ n�� �7� �ܬ ��� ��� �!� �� J�t N� n� �\x ��� ��� �ф �ͺ ��� �{ �� -m� A�� i9� �D� �� �� �O� �	� � 61� ^�� ~�� ��� ��� �Y} ��� �� �Hy �� 1�� ]	� u�� �o� ��t ��� ��v �ۛ �[� �� 5e� MX� i� u�� �� ��� �� �߽ �_� ��� ;� w� �� ��� �� ��t � f� M#  %�   �(  P #�(  M� "�(  J� -   C;*  ��  A� �| 		� �� � �~ ̓  ʝ $5� +�� .ȇ 5t� :�� ?+� Es� K
� P�� Sd� Z�� a� f�� i� p� v�� |M� ��� ��� ��� �ј ��� �j� ��� �ر �g� �u� ��� �I� ��{ ��| �.� �� ��� �� �f� �u� ��z �� ��� �S� �fu �f| �ʥ ��� ��� �� �)� ��� �أ � �� ��(  	� �s*  �: ��(   �  �s   �� �H*  #s*  %�*  �*  P #�*  N~ ��*  .:� M�*  1org Oc   1cur Pc  1fit Qc   "� S�*  W� S�*  �*  O� �&+  +  Z�� x2 T,  ڰ   V]   A�  X�  �  Yc  ��  [�  q	  \c   �0   ^  (��   _  ,N5   `q=  0q5   b  8D�  c  <H�  dBA  @�~   fHA  H6"�  hP  6�  iP  6�e  k�,   6+�  mc  (6�  nc  06
�  v�@  8 .� 0��,  
��  ��   
A� ��  
�� ��  
� �c  
q	 �c   
�L  ��  (
�1  �P  , 2� �,  �� ��,  ,  �� �(�,  �,  "� H��,  ހ �4   $� ��,  �� �   80� �(4  @ 5� �-  -  $�  -  �,  �   �� �+-  1-  0A-  �,  �,   r� �M-  S-  0^-  �,   ɸ �j-  p-  0�-  �,  �-  �-   c  � ��-  �-  $�  �-  �*  �,   � ��-  �-  $�  �-  �  �*  �-  �,   �  J�� -   
.  �  �y B� C� �  s� �-  Bw @�.  *� .   zt (�  � (�,  } (-  � (A-   ]� (^-  (՟  (�-  0�� !(�-  8 8� #&.  #�.  �� %,�.  #�.  �.  J6� -   >E0  ��  E� �� z� � �~ @� *� �� ݌ 	9� 
?� ̻ �� ~� ��  ũ �� � L� (� �� =� +� �v � !� 	� Q� 5� � D�  D� !	� "�� #� $;� %� &�� '[� (�� )�| *�w +J� ,� -[� .� /�� 0x� 1� 2�� 3� 4�� 5� 6>� 7K� 8m� 9֖ : �� E�.  x� H}0  ��  JP   ��  KP   �� MR0  #}0  `� Q)�0  �0  �� (T�0  � VE0   ;� Y�0  ~ Z�0  � \   0� ^n    �� `�0  #�0  u b%1  #	1  1  Jͷ -   �w1  �y  �{ et �| H� L� S� V� ä �� 	*� 
 h� �!1  J�� -   ��3  ��  s� x� �� $� 5� ߼ � �� +� 	m� 
�� �� |� H� � 6� ā �� �~ �� �� �� �� �� }| �� ]�  � x� �� s� ��  �� !*� "�� #�� $�� %H� &�� ' � (;� )&� *޴ +ڳ ,e� -R� .�� /�v 0~� 1�� 2�� 3P� 4�� 5� 6� 7̼ 8�� 9�u :�� ;X� <� =�� >K� ?P� @e� Au� B�| CU� D՚ E� FȢ Gt� Hy I�� J�� K̐ LK� MQ� N�w O`� P� Q�� R
� S`� T�� U !� ��1  (� ��3  l�  ��3   *� �.  � �E0  �� �;*  e� �w1   �� ��3  #�3  �� �$"4  #4  4  � �'54  ;4  U1�  !i�4  
��  !k�   
�� !l�  
�� !m�<  
�� !u�  
�e !w�<   2�� !{s  �2�� !~c  �2�� !�c  �2�� !�c  �2�� !�c  �2�� !��  �2ϖ !��5  � �~ ��,  Q�(  "	�PG     `�*  "�	�HG     .a� H##y5  
ah #%�"   
� #'�  
�� #(�  
� #*    
�'  #,   !
iO  #-y5  $ %  �5  +S    � #/�5  5  	�-  #2	  %�.  �5  P #�5  	\� !!�5  	v� $!1  	�� $'1  	 � $-1  	T� $31  	ޭ $91  	�� $@1  	� $F1  	п $L1  	� $R1  	�� $X1  	e� $^1  	*� $d1  	 � $j1  	�� $p1  	�� $v1  	�� $|1  	� $�1  	G� $�1  	�� $�1  	k� $�1  	Lz $�1  	�� $�1  	�� $�1  	G� $�1  	]� $�1  	� $�1  	_� $�1  	ҵ $�1  	� $�1  	(u $�1  	�� $�1  	x� $�1  	� $�1  	�� $�1  	� $�1  	�� $�1  	�� $�1  Gx $1  �u $1  t� $1  ˃ $1  8� $1  �� $ 1  ș $&1  r� $,1  !� $21  ۔ $91  /� $@1  � $F1  6� $M1  $� $S1  ؠ $Y1  /� $_1  \w $g1  ڷ $m1  O� $s1  �� $y1  n� $�1  %1  �8  P #�8  	� !+�8  	�� %V4  	� %]4  	�� %d4  	2{ %k4  	G� %r4  	�� %y4  	m� %�4  	e� %�4  	t~ %�4  	�� %�4  	ۤ %�4  	� %�4  	� %�4  	�� %�4  	�� %�4  	� %�4  	5~ %�4  	~� %�4  	:� %�4  	� %�4  	�� %�4  	�� %�4  	�� %�4  	�} %�4  	 %�4  	�� %�4  	x� %�4  	�� %�4  	�� %�4  	\� %�4  	T� %�4  	р %�4  	� %�4  	3� %�4  	+� %�4  	�� %�4  	� %�4  	�u %�4  	�� %�4  	�� %�4  	qw %�4  	�� %�4  	|� %�4  	�� %�4  � %4  2� %	4  ƽ %4  �� %4  Mu %4  �� %4  � %4  �� %4  �� %4  c� %4  � %4  �} %4  	t %4  .� %4  �� % 4  5� %'4  �� %74  u� %>4  �� %E4  �� %L4  fy %S4  �� %Z4  %� %a4  �� %h4  �v %o4  M� %v4  �� %}4  �� %�4  6� %�4  ]{ %�4  � %�4  �� %�4  Lt %�4  % %�4  �� %�4  9� %�4  G� %�4  h� %�4  �� %�4  � %�4  s� %�4  %4  �<  P #�<  	�� !5�<  s  %�,  =  +S   T _� -    !(=  D�  )� &�  X�  *=  _J� Z    /e=  �� �� e�� � ec� ~ 3�  74=  �  �#}=  �=  .~� P �.>  
�1   �s   
'�  �,  
�  �,  1ox  �c  1oy  �c  1fx  �g  1fy  �g  1x  �c   1y  �c  (1u  �c  01v  �c  8
�W  �q=  @
��  �q=  H Ű  �#:>  @>  3� P !?  �1   
?   ?dir  ,  ?pos  g  ��  g  5z  g  ܁  g  ��   g  
{�  !?  +�  .>  ��  .>   Q�  .>  (�  c  0?len  c  8��   q=  @��   q=  H ��  �#-?  3?  8� X  �?  �  "g   ^�  #c  ?pos  $c  �1   &?  ?dir  ',  1�  (�   \�  *�*  (��  +!?  0Q�  ,!?  8�  -  @��   /.>  H��   0.>  P 7�  �=  �  @>  կ  23?  f�	 G:@  X�  I:@   6V�  JJ@  � %�?  J@  +S    %@  Z@  +S    Z u �	 7�@  `�  9     :  X�  ;.>  ��  @  @�  A  V�  B!?  ��  De=   
�  K@  ( c�  NZ@  ?z  N�@  Z@  f@ r"A  H�  t"A   N5   u2A  @ %q=  2A  +S    %�?  BA  +S   _ q=  %�@  XA  +S    ��  x+  	ۢ &�.  .�� H&M�A  1ref &O�*   
�� &P�*  
�  &Qc  0

  &Rc  8
�1  &S�  @ �� &UqA  � &U�A  qA  UX� 0I&X�B  
1� &Z�   
�� &[c  
�� &]�  
Չ &^�B  2�� &_c  �2M�  &`c  �2!� &a   �2y� &d�  �2��  &e�B  �2� &g�   I2l� &hc  (I %�*  �B  +S    %�A  �B  +S   �  � &j�A  �� &j�B  �A  U� ��&m�B  
ah &o�4   
��  &p�  H
�~  &q�B  P %�B  C  +S    �� &s�B  �� &sC  �B  	Nv '�.  .ƍ 8'@fC  1ref 'B�*   
�� 'C�*  
�1  'D�  0 7� 'F1C  J� 'F~C  1C  U P9'I7D  
1� 'K�   
�� 'Lc  
�� 'N�  
Չ 'O�B  2�� 'Pc  �2M�  'Qc  �2!� 'R   �2�� 'U   �2y� 'V�  �2��  'W7D  �2� 'Y�  @92l� 'Zc  H9 %fC  GD  +S   � � '\�C  � '\_D  �C  U&� �r'_�D  
ah 'a�4   
��  'b�  H
�~  'c�D  P %GD  �D  +S    � 'eeD  �t 'e�D  eD  d-   (�G  �v  i� �x L� ߇ �� 8� �� �� ԩ 	� 
O� `� а | �� (� � �� �� � ��  � ![� "=� #9| $$� %8� &�� '�� (x� 0� 17� @N� A�� Q� R� S?� T]� Up� V�� W�� X$v `�u a�| b�x cD� p�� ��� ��� �)� �y� �� ��w ��� ��� ��� �x� ��� �� �Ս ��� ��� �� ��� �� �� ��� ��� �t� ��� �o� ��� �� ��� �f� �� �%� �3� �� �\� ��� ��� ��� �̒ ��w ��� �1� �� ��� �a~ �E� �w �I� � s� ) C  #G  .j� p)"�G  1x1 )$c   1x2 )$c  1t1 )%c  1t2 )%c  
�� )&c   
� )&c  (
i� )'c  0
	� )'c  81w0 )(c  @
� )(c  H
�� )(c  P
!� )*�  X
� )+c  `
�� ),G  h
{ )-G  l �� )/G  S{ )/H  G  `%C  @		�HG     	� *�.  QH  <	@HG     %�0  AH  P #6H  	�� $!AH  	H� $'AH  	�� $-AH  	m� $3AH  	�{ $9AH  	{ $@AH  	q� $FAH  	�� $LAH  	k� $RAH  	�w $XAH  	&� $^AH  	� $dAH  	u� $jAH  	!� $pAH  	B� $vAH  	�w $|AH  	T| $�AH  	K� $�AH  	�} $�AH  	Ѕ $�AH  	S� $�AH  	9� $�AH  	az $�AH  	ݙ $�AH  	֑ $�AH  	�v $�AH  	� $�AH  	Y� $�AH  	� $�AH  	Ѧ $�AH  	K� $�AH  	�� $�AH  	� $�AH  	�� $�AH  	�� $�AH  	�} $�AH  	�� $�AH  � $AH  �� $AH  S� $AH  �� $AH  N� $AH  �� $ AH  8� $&AH  i $,AH  ܏ $2AH  !� $9AH  ɛ $@AH  �� $FAH  � $MAH  T� $SAH  x $YAH  r� $_AH  �� $gAH  �� $mAH  � $sAH  �� $yAH  �� $�AH  	�� $!AH  	�� $'AH  	�� $-AH  	�} $3AH  	5� $9AH  	~ $@AH  	Z� $FAH  	� $LAH  	=� $RAH  	�� $XAH  	q� $^AH  	X� $dAH  	۪ $jAH  	� $pAH  	� $vAH  		� $|AH  	�� $�AH  	{� $�AH  	�� $�AH  	�� $�AH  	� $�AH  	� $�AH  	>� $�AH  	�z $�AH  	d� $�AH  	x� $�AH  	�� $�AH  	t� $�AH  	߶ $�AH  	g� $�AH  	9� $�AH  	o� $�AH  	� $�AH  	� $�AH  	V� $�AH  	�� $�AH  	�� $�AH  P� $AH  �� $AH  �� $AH  � $AH  �~ $AH  מ $ AH  v� $&AH  �� $,AH  g� $2AH  S� $9AH  �� $@AH  � $FAH  j� $MAH  �� $SAH  � $YAH  -� $_AH  �� $gAH  �� $mAH  � $sAH  � $yAH  �� $�AH  	Z� +�.  �5  	 HG     �5  	�GG     �5  	�GG     �5  	@GG     �5  	 GG     �5  	�FG     6  	�FG     6  	@FG     #6  	 FG     /6  	�EG     ;6  	�EG     G6  	@EG     S6  	 EG     _6  	�DG     k6  	�DG     w6  	@DG     �6  	 DG     �6  	�CG     �6  	�CG     �6  	@CG     �6  	 CG     �6  	�BG     �6  	�BG     �6  	@BG     �6  	 BG     �6  	�AG     �6  	�AG     7  	@AG     7  	 AG     7  	�@G     +7  	�@G     77  	@@G     C7  	 @G     O7  	�?G     [7  	�?G     g7  	@?G     s7  	 ?G     7  	�>G     �7  	�>G     �7  	@>G     �7  	 >G     �7  	�=G     �7  	�=G     �7  	@=G     �7  	 =G     �7  	�<G     �7  	�<G     8  	@<G     8  	 <G     8  	�;G     (8  	�;G     58  	@;G     B8  	 ;G     O8  	�:G     \8  	�:G     i8  	@:G     v8  	 :G     �8  	�9G     �8  	�9G     �8  	p9G     �8  	P9G     �8  	09G     �8  	9G     �8  	�8G     �8  	�8G      9  	�8G     9  	�8G     9  	p8G     $9  	P8G     09  	08G     <9  	8G     H9  	�7G     T9  	�7G     `9  	�7G     l9  	�7G     x9  	p7G     �9  	P7G     �9  	07G     �9  	7G     �9  	�6G     �9  	�6G     �9  	�6G     �9  	�6G     �9  	p6G     �9  	P6G     �9  	06G     �9  	6G     :  	�5G     :  	�5G      :  	�5G     ,:  	�5G     8:  	p5G     D:  	P5G     P:  	05G     \:  	5G     h:  	�4G     t:  	�4G     �:  	�4G     �:  	�4G     �:  	p4G     �:  	P4G     �:  	04G     �:  	4G     �:  	�3G     �:  	�3G     �:  	�3G     �:  	�3G     �:  	p3G     
;  	P3G     ;  	03G     $;  	3G     1;  	�2G     >;  	�2G     K;  	�2G     X;  	�2G     e;  	p2G     r;  	P2G     ;  	02G     �;  	2G     �;  	�1G     �;  	�1G     �;  	�1G     �;  	�1G     �;  	p1G     �;  	P1G     �;  	01G     �;  	1G     <  	�0G     <  	�0G     <  	�0G     (<  	�0G     5<  	p0G     B<  	P0G     O<  	00G     \<  	0G     i<  	�/G     v<  	�/G     �<  	�/G     �<  	�/G     �<  	p/G     �<  	P/G     �<  	0/G     �<  	/G     Q�5  
J	�.G     Q�8  
X	 -G     Q�<  
f	@*G     Q�M  u	 *G     `eA  '	�)G     .}� x,%&W  
��  ,(�   
0� ,)(4  
�7  ,,�*  
�e ,-�,  
�&  ,.    
^� ,/3	  (
� ,0�  H1pp1 ,1�  X1pp2 ,2�  h d� ,5�V  �� ,5>W  �V  � -�oW  ��  -��   ?map -��<   @} -�DW  � -��W  ��  -��   ��  -��   &� -�|W  �<  .�W  �W  $�  �W  Y  n  �      s=  .$�W  �W  $�  X  Y  n  a    �  .) X  #X  .#P  .)HX  
R  .+�W   
bD .,�W   7�� �X  	�)G     %!  oX  +S    #_X  7�� �oX  	�)G     r�� #�   	`)G     �5  ,	 )G     ,FH  /; 	�(G     ,K  /A 	�(G     ,RH  /H 	�(G     ,K  /S 	 (G     ,^H  /l 	�'G     ,+K  /s 	�'G     ,jH  /z 	�'G     ,7K  /� 	�'G     ,vH  /� 	�'G     ,CK  /� 	�'G     ,�H  /� 	�'G     ,OK  /� 	@'G     ,�H  /� 	 'G     ,[K  /� 	'G     ,�H  /� 	 'G     ,gK  /� 	�&G     ,�H  /� 	�&G     ,sK  /� 	�&G     ,�H  /� 	�&G     ,K  /� 	�&G     ,�H  /� 	�&G     ,�K  /� 	p&G     ,�H  /� 	`&G     ,�K  /� 	P&G     ,�H  /� 	@&G     �K  /  	0&G     �H  / 	 &G     �K  / 	�%G     �H  / 	�%G     �K  /, 	 %G     �H  /: 	%G     �K  /@ 	%G     I  /F 	�$G     �K  /O 	�$G     I  /V 	�$G     �K  /] 	�$G     I  /c 	�$G     �K  /k 	x$G     *I  /q 	`$G     �K  /x 	P$G     6I  / 	@$G     L  /� 	8$G     BI  /� 	 $G     L  /� 	�#G     NI  /� 	�#G     L  /� 	�#G     ZI  /� 	p#G     'L  /� 	@#G     fI  /� 	#G     3L  /� 	�"G     rI  /� 	�"G     ?L  /� 	�"G     �I  /� 	�"G     cL  /� 	`"G     ~I  /� 	P"G     KL  /� 	 "G     �I  / 	 "G     WL  /	 	�!G     �I  / 	�!G     oL  / 	�!G     �I  / 	� G     {L  /C 	  G     �I  /Y 	�G     �L  /a 	�G     �I  /g 	`G     �L  /y 	@G     �I  / 	0G     �L  /� 	 G     �I  /� 	G     �L  /� 	�G     �I  /� 	�G     �L  /� 	�G     �I  /� 	�G     �L  /� 	 G     J  /� 	�G     �L  /� 	�G     J  /� 	�G     �L  /� 	�G     J  /� 	�G     �L  /� 	�G     )J  /� 	�G     �L  /� 	pG     6J  /� 	`G     M  /� 	PG     CJ  / 	@G     M  / 	0G     PJ  / 	 G     M  / 	 G     ]J  / 	�G     *M  /! 	�G     jJ  /' 	�G     7M  /- 	�G     wJ  /5 	�G     DM  /< 	pG     �J  /D 	`G     QM  /J 	@G     �J  /S 	0G     ^M  /Y 	 G     �J  /d 	�G     kM  /j 	�G     �J  /u 	�G     �M  /{ 	�G     �J  /� 	`G     xM  /� 	PG     �J  /� 	@G     �M  /� 	0G     �J  /� 	 G     �M  /� 	 G     �J  /� 	�G     �M  /� 	�G     �J  /� 	�G     �M  /� 	`G     �J  /� 	PG     �M  /� 	 G     K  /� 	�G     �M  / 	�G     %G  Ha  +S   ? #8a  @�� 	-Ha  	�G     [�s 	��b   �� 	�%�G   �7  	�%�*  adim 	�%(=   /� 	�%�   �� 	�%�-  �~  	��@  N5  	�q=  � 	��  l� 	�c  )nn 	�  ��  	�  `� 	�#  )X1 	�  )X2 	�  )w 	�  � 	�G  X� 	�.>  "Gb  )X 	�   "Zb  �� 	Z    "�b  �� 	.�  +� 	/c  xx1 	0c  xx2 	0c   !� 	`�  � 	ac    V� 	HP�D     �      ��d  L�� 	H.�G  UL1� 	I.�  T-�� 	J.c  L� F� bxx1 	K.c  �� �� bxx2 	L.c  ٫ ի -� 	M.G  � � LX� 	N..>  � L`� 	O.  ��� 	Q  l� d� � 	Q  � � �� 	Q%  E� 9� :nn 	R  �� �� @^� 	S�d  ��}!� �c  �� 	]c  T� J� � 	^c  6� *� :w 	_c  (� "�  38�D     h       �d  :len 	yc  �� ~� :y0 	zc  �� � :y 	{c  � � :idx 	|  o� i� s��  8�D      � 	z��  �� �� ��  � ߳ � ��  � � ��  U� Q�    0 :idx 	�  �� �� ` � 	�G   � �� 
� 	�G  �� ��    %G  	e  +S   @ g(� ��  we  �e �(�,  � �(a   4idx �(-   � �(we  y�  �(we  ��  ��  x ��   �  h�� bn  0�D     �      ��f  Hp b+n  � ҵ �e c+�,  � � � d+a   t� h� /� e+�f  � �� ��  g�  Ѹ ϸ ch h�  	� �� ��  h�  � չ buf i�f  R� F� !�9 df  �  o�  � ڻ  !: �f  �  t�  V� J�  W��D     �  -   �  t�� Y�f  ��  Y#�  4buf Z#a    h� Pa   �D            ��f  B��  P"�  U g� A�  @g  0� A+(4  ހ B+4  p� C+�<  �� D+    <X� ��  0�D     p      ��r  ϖ �+�5  �� � �  �+�  ս ѽ ֳ  �+W  � � x �+�  O� K� �1  �+C  �� �� �U ��  �� �� ڰ  �]  � � 7�7  �r  �Ț7��  �r  �Й��  ]�D      �& Ph  Ǹ  G� E� ��  n� j�  �}  ��D       ' �h  �}  �� �� �}  �� ��  uz  ��D      p' �r  �z  � �� �z  0� ,� �z  v� l� �z  �� �� �z  �� �� p' �z  (�  � �z  �� �� �z  � � �z  s� i� �z  �� �� �z  �� �� 
{  5� #� '{  ���"{  � 
� i.{  A:{  �� �� F{  �� �� CR{  ��D     C[{  ��D     ^}  F�D      �' +j  �}  � � {}  P� L� o}  �� �� �' �}  �� �� e�D     ��  Us T�ؙQ���   C�  _�D      �' ;.k  o�  ;� 5� |�  �� �� b�  �� �� U�  B� @� �' ��  �� h� ��  �� �� ��  �� �� ��  =� 5� '��  ���Cʻ  }�D     \ӻ  *ܻ  @( ݻ  �� �� X�D     �j  Uv  X+�D     �j  Uv  6�D     � k  U~ Tv  ��D     � U~ Q���    ('|  �( [m  '(|  ���'5|  ����  ��D      �( 
�k  ��  �� �� ��  %� #� �( ��  W� S� ��  �� ��   ��  �D       ) �k  ��  �� �� ��   ) ��  �� �� ��  B� >�   �  ��D       0) -6l  (�  �� }� (�  �� }� 5�  �� ��  ��  !�D      `) @#�l  ��  � � ��  7� 5� `) ��  `� \� ��  �� ��   ��  X�D      �) 1�l  ��  �� �� ��  � � �) ��  /� +� ��  r� n�   N�D     � m  Us T��� ��D     �  m  Us Q0 ��D     � >m  Us T|  ��D     
 U��T|   D|  �D      �) �ap  m|  �� �� a|  �� �� U|  %� !� �) y|  g� c� �|  �� �� �|  �� �� �|  3� 1� �|  t� n� '�|  ��'�|  ���|  �� �� �|  � � �|  \� V� '�|  ���C�|  ��D     5}   �D     �       �n  
}  �� �� }  �� �� M��   �D      * ��n  ��  � �� ��  .� *� * ��  l� h� ��  �� ��    �D     ��  �n  9�x  �Й9�x  s  M�D      T���  5#}  ��D     �       �o  $}  �� �� 0}  � � M��  ��D      P* ��o  ��  >� <� ��  d� b� P* ��  �� �� ��  �� ��   ��D     ��  �o  9�x  �Й9�x  s  ��D      �o  T��� 5�D      U�Șs T�Ș  k�D      p  U�B$T�Ș X��D     +p  U T��Q�� h�D     $ Cp  Us  ��D     � Us T���   (d{  �* �p  'i{  ����D     1 �p  U��� R�D     
 U���T���  ��  ��D      �* �	q  ��  � 	� ��  3� 1� �* ��  \� X� ��  �� ��   (w{   + �q  |{  �� �� 5�{  q�D     �       �q  �{   � � �{  _� Y� �{  �� �� �{  � � �{  A� ?� �{  f� d� �{  �� ��  I�{  ��D     2       �{  �� �� �{  �� ��   (|  P+ �q  |  �� �� |  "�  �  X8�D     r  U T��� XN�D     )r  U�ȚT  r�D     > \r  Us T����Q����	�
(! ��D     � ur  Uv� u4�D     U����T�ȚQs R    D}  ��D      �+ �r  Q}  J� H�  ��D     ��  U�Ț  %XA  �r  +S     %&W  �r  +S     A"� �@�D            �.s  B̖ �"Y  U <>� ��  ��D     H       �vs  B̖ �"Y  Uϖ ��5  s� q�  <c� ��  ��D     
       ��s  ϖ �"Y  �� �� 2*  �"n  �� �� O��D     K U	�)G     T�T  <܉ =�  �D     �      �pv  ̖ =!Y   � � �1  >!n  �� �� <v ?!a   � �� �U A�  �� �� ϖ B�5  +� � � C�  �� �� �� D�  �� �� � F   �� �� 3 �D     !       u  Cp L"pv  d� ^� 70� M"(4  �h0�D     2x  T�hQ�U  3 �D            Gu  val Xvv  �� �� ހ Z4  �� ��  3T�D            ru  val cvv  (� $�  3p�D     (       �u  Cp l!|v  e� a� 70� m!(4  �h��D     2x  T�hQ�U  3e�D            �u  val y�v  �� ��  3��D     @       3v  iO  ��v  �� �� val ��v  �� ��  &��D            �'  �   #� !� val ��v  H� F�   oW  �  �W       N�� k�  2x   ̖ k!Y   �1  l!n   <v m!�   �h  n!   �U p�  ϖ q�5  "w  � zvv  )ss {�  ހ �4    "$w  �� �vv   "Bw  Cp �!|v  0� �!(4   "\w  )s �n  )w �@    "nw  � ��v   "x  iO  ��v  )x1 �  )y1 �  )x2 �  )y2 �  )x3 �   )y3 �$  )x4 �(  )y4 �,  )dp �y5  )s �n  )ep ��   )i �Z     ""x  s !n  nsd "@    �'  -�v    R� I�  ��D     f       ��x  -��  I2�  u� k� -�� J2�x  �� �� -ϖ K2�5  �� x� �U M�  �� �� @0� N(4  �X��D     ��  T�X  (4  EA� VC  uz  ��  V+2W  ��  W+�  M�  X+c  ϖ Z�5  �   \s  � ]�  � ]�  `� ^�  Z� ^�  M� ^1�  �� ^>�  %� _  x1 `  y1 `  x2 `  y2 `  x3 `   y3 `$  x4 `(  y4 `,  D-� �D4� �DP� �""z  � �  m� �  x �   "Mz  � �  m� �  x �   � �  m� �  x �    N(� ��  D|   ��  �$2W   ϖ �$�5   ��  �$�   x �$�   �1  �$C  �U ��  ֳ  �W  
� ��  �  ��  �� �  �m  ��  �7  ��*  $� ��,  '} ��,  �� ��  ހ �4  c� ��.  D�  ID4� "w{  �} �3	   "|  �~  ��@  "�{  �� �!?  Ɩ �!?  c� �c  �� �c  V� �c  �u �c  �� �c   �� �c  �� �c    "'|  �� �c  �� �c   �;  �  � �    NL� Y�  >}   ��  Y62W   ��  Z6�   '} [6�,  �U ]�  �  _�  0� `(4  c� a�.  I�  c>}  ,� ec  N� fc  E� h   Mp  k�  � l�  � n3	  ]�  �"#}  	� ��  �� �)�   �� ��  �� �)�    �  [t� H^}   ��  H2W   N� +�  �}   ��  +2W   ϖ ,�5   ��  -�  �U /�   [z} �}   ��  "2W   �7   "�*   E� ��  n~  x �*�  �7  �*�*  Mj  �*�-  �e �*C  �U ��  dim �Z   �~  ��B  F�  ��D     ��  �G  1� �  �� c    8�� ���  �7  �'�*  4dim �'(=  �~  ��@  V� �!?  �� �!?  � ��  {� �!?  �`  �!?  � �  ހ �4  � �	1  � �   "a  �� ��*  �� �!?  Ɩ �!?  	� �?  Ԍ �?    "h�  Ɩ #!?  "�  K{ Ec  � Ec  �� E&c  n� Fc  P  Fc  P  F#c  �� F+c  �� F2c   � �c  K{ �c  � �#c  �� �/c  n� �c  w� �c  ��  �%c  P�  �-c  �� �c  �� �c     "ɀ  �� !?  Ɩ !?  �� !?  �� c  a� c  & c  �� $c   �� Jc  �j  l!?  R  l!?     8]� �+�  �7  �-�*  Ǟ  �-!?  Q� �-!?   A�� pP�D     I       ���  �7  p.�*  b� ^� Hdim q.(=  �� �� � r.!?  �� �� �� s.!?  0� *� �  uc  �� |� b� uc  �� �� N� vc  � � ��D     9�  Q�T9�  �U  E�� �
c  ��  �7  �
/�*  4dim �
/(=  5�  �
/c  b� �
/c  �� �
/�  �� �
/�  �e �
C  �~  �
�B  �  �
c  �} �
  <  �
  D�� e"ׂ  �� �
c  �� 	c  � �     ��  #c  �� Oc     v�� z
c  {�  Չ z
"�*  /� {
"�  5�  |
"c  n ~
�  �� 
c  D� �
c  ��  �
c  w �
c  �  �
c    <�� !
�   �D     �       �P�  B�7  !
)�*  UB�e "
)C  Tt $
�  @� :� "� %
P  �� �� � %
#P  �� �� ��  &
�  2� 0� ;y�  (�D      p )
��  W� U� ��  W� U� ��  |� z�   8&� �	C�  �7  �	7�*  �e �	7C  �~  �	�@  {� �	!?  �� �	!?  �� �	�B  1� �	�  bb �	�  �� �	�*  �� �	   �� �	c  �� �	�A  i� �	   �� �	$   �� �	5   �  �	c  ~� �	        E�� �	�  ��  �7  �	2�*  �� �	2�  Չ �	2��  4dim �	2(=  �U �	�   �*  <J� 8�  �D     5      �G�  �7  80�*  �� �� Hdim 90(=  :� 0� �~  ;�@  �� �� �U <�  1� )� ڰ  =]  �� �� C� >�B  @� :� ހ @4  � A	1  �� �� � C    � �� X� E.>  f� `� T� F.>  �� �� seg G.>  � �� 1� L�  �� �� �� Mc  >� 0� 2� Nc  �� �� `� Oc  (� "� F�  �	��D     !@ 7�  �  �!?  y� u� ee �  �� �� 3��D     )       ��  {� �!?  �� �� �  �c  .� (�  � 7{� �!?  ��G��  <�D      <�D            ��  ��  ��  �� �� &<�D            ��  �� �� ��  0� ,�   �D     %�  U��R���X��Y��   3��D     i       ��  �  �!?  q� k� ee �  �� �� � {� �!?  �� �� �  �c  :� 4�   !  ��  V� 	!?  �� �� �� 	!?  �� �� {� 	!?  � � 0 ��  	  �� {� �� !	  �� �� p N� ,	   !� � � Ɩ E	!?  �� � #� F	.>  �� �� &کD     :       �� T	c  `� ^� �{ U	c  �� ��      ��  ��D      � ���  ��  �� �� ��  �� �� � ��  � � ��  N� J�   ��D      �  U@ ��D      2�  U Ts  �D      Ts   A�� �p�D     �      �G�  �7  �0�*  �� �� �� �0�  �� �� Չ �0��  � � Hdim �0(=  D� @� �~  ��@  �� }� X� �.>  � � T� �.>  )� '� � �c  R� L� 
� �"c  �� �� w5} �-c  �Sd  �9c   � � ˿ �.>  I� C� #� �.>  �� �� � r� �c  �� �� {� �c  � � � min �c  �� �� max �c  �� �� len �c  ]� [�  �  �c  �� �� y� �c  �� �� � �#c  � � @ �� c  *� &�      <>� �  ��D     �	      �  �7  3�*  ~� v� Hdim 3(=  �� �� �e C  1� /� �~  �@  ^� V� ڰ  ]       �U �    g  ��  	.>  � � 7� 
�?  ��~2 BA  � � ǟ BA  � � �� e=  � � m� !e=  d J j� c  } w F�  �КD     3U�D     &       ȍ  c q=  � � ��  q=      3T�D     ,       �  c *q=   w ��  +q=  � �  !� ݐ  c 8q=  '  ��  9q=  � � �� :Z   � q �x ?c  
 �	 ͋ @c  �
 �
 5z Ac  � � ܁ Bc  � r ٮ Cs  � � �� Ds  V > t� Ec  p Z �� Fc  u ] �� H   � u y� J.>  x j }x Lc    ȋ Mc  � � 0z Nc  A ' ׁ Oc  | b Ԯ Ps  � � �� Qs  � � o� Rc  S 9 � Sc  � t   u nc  � � v nc  N B ;��  ЗD      � >��  � � ��  � � ��  '  � 'ɺ  ��~պ  /  C�  �D     *�    �      ��  �  �  �  Q! I! C�D     X ��  U��~TPY��~ �D     X U��~TPQ0X0      &��D     �       X� x.>  �! �! �� y.>  �! �! � ��  ~q=  " " ��  q=  �" �" D� �c  �" �" 9� �c  j# d# 3��D     &       ��  p �q=  �# �#  &,�D     &       p �q=  �# �#     A�� �P�D            ��  B�e �2C  UBN� �2�-  TB,� �2�-  Q Ax� ���D     <       ���  �e �,C  >$ 6$ $� �,�,  �$ �$ ֯D     ��  {�  Us Tv Q0 O�D     ��  U�UT�TQ1  A0� �P�D     U      �"�  �e �0C  % % $� �0�,  �% �% Hdim �0(=  =& -& 1� ��  �& �& �� �c  h' d' �~  ��B  �' �' nn ��  i) W) !  �  � ��B  5* +* �� ��A  �* �* ` ��  �c  + + �  �c  X+ T+ k� �c  �+ �+ ��  ��  �+ �+ � ��  
, , 3 �D     �       ��  � �c  w, q, �  �c  �, �, �� ��  - - ��  Q�D      � ���  ��  8- 2- ��  �- �- � ��  �- �- ��  . .   �D     d U   ;��  ��D     	 � ���  @. >. ��  e. c. � ��  �. �. ��  �. �.     !  ��  5�  2�*  / / Y��  8�D      8�D            5��  ��  D/ B/ &8�D            ��  l/ h/ ��  �/ �/    !� ��  �� V�A  �  Wc  !� ŕ  P�  gc  �/ �/  ��  խD         Z�  ��  ��  0 0   ��  c0 _0 ��  �0 �0   ��  U�D      ` aI�  ��  ��  ` ��  ��    ;��  2�D      � \��  ��  � ��  �0 �0 ��  &1 $1    3��D     K       ז  �� ��A  i ��  &ɮD     '       b ��A    ;��  a�D      P B��  ��  K1 I1 P ��  �1 �1 ��  �1 �1    <R� x�  PE     O      ���  �e x+C  2 2 ��  y+�  r2 j2 �U {�  �2 �2 �� }  ?3 73 F�  ��E     ��  �E      �B �A�  ՙ  �3 �3 ș  �3 �3 �B �  �3 �3 �  W4 O4 '��  ��	�  �4 �4 '�  ��#�  %5 5 '0�  ��=�  z5 t5 *H�   C I�  �5 �5 'V�  ��G	e  =E      =E            X�  Oe  �5 �5 Be  )6 #6 5e  �5 �5 (e  z6 x6 e  �6 �6 &=E            \e  �6 �6 ie  �6 �6 [E     q T Q
R��   3E     }e  U~ Tv Q��R��    �E     } b�  Us Tcinu �E     � ��  Us Tw  �E     ��  ��  Uv Ts  �E     z�  Uv Ts   8�� 3e�  �e 33C  ��  43�  � 6   �� 6   � 7�  �� 7�  � >�  �t ?a   *� Cu�  p Dn  x O�  T� P-     %�   u�  +S    #e�  <I� @Z   �E     �      �!�  �e @1C  7 7 ��  A1�  R7 N7 7�� C!�  ��y7� D!�  ��|}� F�  �7 �7 � G�  O8 ?8 �� I�A  9 	9 �U J�  �9 �9 �~  K�B  �9 �9 Mj  L�  J: 6: sc N4  bss P;*  bs Q1�  <= 4= j� Sc  �= �= 7� Z�  ��x�t [a   �= �= !�> �  p ln  C> -> �� m�-  6? .? �� n�-  �? �? �  oc  �@ �@ 
  pc  �A �A ! ? �  x ��  �B �B y�  ��  �B �B *� �  iC OC � �!  �D tD b� �5  FE 4E N5  ��  5� �c  F F k� �   �F �F i �-   kG [G 7T� �-   ��x!�? �  �� �c  0H H �  �   RI BI ! @ ��  nn �  J  J ��  �  DJ <J ��     �J �J P@ &�   �J �J pp   AK -K   !�@ B�  � =c  +L L �� >  �L �L �W >  4N  N �� ?  TO BO O� ?)  /P P z� @  ^Q <Q � @*  �R �R �  Ac  rT FT A :� �c  <Y 0Y `A <u �c  ��  �  �Y �Y ��  �  �Z �Z hit �   �[ �[ 0� �  p\ h\ }u �  �\ �\ ^� �   K] I] �A l2r �   v] p] d �c  �] �]     G	e  �E      �E            �ן  Oe  �^ �^ Be  _ _ 5e  9_ 7_ (e  ^_ \_ e  �_ �_ &�E            \e  �_ �_ ie  �_ �_   �E     > U~ Q1  GE     }e  T��wQ��xR��x  3^E     =       k�  ref �c  �_ �_ �� �c  5` 3` � �   m` k`  jb�  %E     l       �Ġ  {�  o�  &%E     l       ��  �` �` ��  ��  �` �`   kb�  �E     {       �{�  o�  &�E     {       ��  'a !a ��  ��  ua sa    !�A ѡ  i ��  7W� �7�  ��x!�B o�  a ��-  �a �a b ��-   b �a  xG�  0B �b�  U�  0B o�  @b 8b z�  �b �b ��  *��  `B ��  �b �b ��  c �b     &�
E     G       0� (4  <c 8c p� �<  {c wc i �  �c �c   %c  1�  +S   2 �*  %�A  G�  +S   	 8�� ��  /� &�  �B &��  i �  j �  uL  �A  a "c  b "c    �A  V¶ <`E            �Ԧ  -�e <2C  �c �c -��  =2�  Ld Fd @�7  @�r  ���|]�  �!p= ��  �U O�  �d �d x P�  �d �d :dim QZ   2e "e @��  RԦ  ���}$� S�,  �e �e ހ U4  f 
f � V	1  If Ef @� ]�  ���|�t ^a   �f �f :p an  g g 3�E     :       ��  @T� w-   ���}l	e  �E      �E            ���  Oe  ?g =g Be  ?g =g 5e  ?g =g (e  eg cg e  �g �g &�E            \e  �g �g ie  �g �g   �E     }e  Ts Q���|R���}  ! > ��  �~  ��B  h �g  u ��@  ^h Zh :seg �.>  �h �h ��  �.>  �h �h �� �#.>  �i �i @I� ��  ���|!0> T�  �  �c  �i �i  �E     G�  r�  Uv T|  �E     G�  ��  Uv T0Q0R|  _E     ��  U���|Tt   !p> �  �~  ��B  +j !j n� �c  �j �j  My�  �E      �= �+�  ��  0k ,k ��  0k ,k ��  hk fk  E     > H�  U| Q1 EE     � n�  U���}T0Q
�� �E     �  Uv T}�  M��  �E        = I��  Ǹ  �k �k ��  �k �k  E     ��  Uv   %C  �  +S     y�� `�   �e `0�D   N� a0�-   ,� b0�-   RR� R�  ��D            ���  -x R(�  �k �k -�7  S(�*  /l +l -Mj  T(�-  ll hl -�e U(�D  �l �l O��D     ��  U�UT�TQ�QR�R  R@� I�  0�D            ��  L�7  I'�*  U-�e J'�D  �l �l O5�D     B�  Uu T�T  VO� @ �D            �u�  -�e @*�D  #m m -$� A*�,  `m \m O�D     r�  U�UT�T  R]� $�  �E     e       �M�  -�e $)�D  �m �m -��  %)�  n  n �� (  kn gn E     } ��  Us Tcinu 2E     � �  Us T|  KE     f�  0�  Uv Ts  SE     �	 Uv 9��  s   85� ���  �7  �,�*  4dim �,(=  1� �,�  �� �,c  N5  �q=  #z �q=  c �q=   A��  ��D     P      �[�  �7   4�*  �n �n Hdim !4(=  *o  o N5  #q=  �o �o �� $q=  p p 2 %BA  Zp Pp ǟ &BA  �p �p x� '�  q q c (q=  �q �q t�  )q=  t t �>  *q=  at Ut F�� �`�D     Fr� y��D     �% ��  Fq=  sz F q=  �t �t [�  @�D      0& u	{�  ��  bu ^u ��  �u �u u�  �u �u i�  0& ��  ��  ��  ��  ɭ  խ  �  �  c�D     ��  Rv    G[�  ��D      ��D     ;       �+�  ��  v v ��  ;v 7v u�  uv sv i�  &��D     ;       ��  ��  ��  ��  ɭ  խ  �  �  ��D     ��  T| Q��Rs    G[�  ��D       ��D     5       ��  ��  �v �v ��  �v �v u�  �v �v i�  !w w &��D     5       ��  ��  ��  ��  ɭ  խ  �  �  �D     ��  U~ Ts�Rs    Y	�  ��D      ��D     T       |	/�  Hw Dw #�  �w �w �  �w �w &��D     T       <�  �w �w G�  cx _x     8�� �	�  4p1 �q=  4p2 �q=  ~�  �q=  �|  �q=  p �q=  u �c  v1 �c  v2 �c  u1 �c  u2 �c  d1 �"c  d2 �&c  1� �    8�t �U�  4p1 �q=  4p2 �q=  4ref �q=  p �q=  �� �c   A��  �D     �      ���  �7  6�*  �x �x Hdim 6(=  �x �x N5  q=  Ey Cy �� q=  ky iy �~  �@  �y �y V� !?  Oz Kz �� !?  �z �z x� �  �z �z F�� �U�D     P c  q=  { { {� !!?  Z{ H{ � u &c  9| %| ou &c  } } fu &c  �} �} �� 'c  �} �} � min _�  �~ |~ max _�  �~ �~ mid _!�  � � � `c  � � !� (�  nn k�  �� |�    �j  �!?  Ӏ ̀ R  �!?  ��  3�D      P ���  ��   � � ��  E� C� P ��  w� s� ��  �� ��   Wx�D           8,� ���  �7  �4�*  4dim �4(=  �~  ��@  X� �.>  T� �.>  seg �.>  "M�  {� �!?  c �q=  ��  �q=  ��  �!q=   {� �!?  c �q=  ��  �q=  ��  �!q=    8� ��  �7  �'�*  Mj  �'�-  c �q=  ��  �q=  vec ��  tag ��    <ۗ ��   �D     m      �y�  �7  �)�*  � �� Mj  �)�-  ˂ �� 7�U ��  ��N5  �q=  �� �� -Q  ��  � � �N  ��  Ԅ �� A�  �  )� !� �� �  �� �� � c  �� � q	 c  �� �� ڰ  ]  I� C� F�  ���D     Fz nY�D     !� �  c bq=  �� �� �� cq=  ؉ ̉ ��  f�  d� ^� L� g  � ي !� ��  vec l�  ^� X� tag m�   �� �� �� ng   � �� end oq=  �� � �� pq=  +� � � q  �� � ` �o  vc  \� Z� �o  vc  �� �� ��  V�D      � ~"b�  ��  ��  � ��  ގ ڎ ��  !� �   ;��  ~�D      � "��  ��  � ��  `� \� ��  �� ��     ! �  2 �BA  � ޏ ǟ �BA  R� D� end ��  � � idx �5  U� M�  &P�D     �      W� �  �� �� 2 �BA  � � ǟ �BA  W� Q� !@ N�  ��  �q=  �� �� �W �q=  
� � �� �q=  _� S� '� �!q=  � � �o  �c  o� G� �o  �c  � Ė � � e=  ;ո  ��D        �  � �� �  m� a�   ��  �� �� �  3� /� �  p� l�     !@ ֶ  �j  Fc  �� �� C  Fc  D� @� �o  Gc  �� �� �o  Gc  L� H� t� Iq=  �� �� ϑ Jq=  ߜ ݜ  � t� {q=  � � ϑ |q=  )� '� W�D     �    �D     � -�  U~  �D     X W�  Uv T8R Y�� s�D     X Uv TPY��  8{� ���  �7  �,�*  �e �,�,   A�~ ��D     "      ���  �7  �'�*  R� L� ڰ  �]  dim �Z   �� �� 3�D     �       �  �~  ��@  �� � "�D     � :�  Uv  J�D     � R�  Uv  x�D     � j�  Uv  ��D     � Uv   ̰D     � ��  Uv  ��D     � Uv   8C� �ո  �7  �'�*  ڰ  �']   E�� �e=  %�  4dx �!c  4dy �!c  ll �c  ss �c  dir �e=   RV� c�  ��D     x      ���  -�~  c)�@  X� H� -� d)  � � bdir e)e=  z� j� -� f)   5� %� -ڰ  g)]  �� � -� h)��  � Ρ @�U j�  ��{� k!?  �� �� V� l!?  3� 1� z�  ���D     � -Q  y  a� W� �N  z  � ң �� {  �� }� &�D     X g�  TXY�� ��D     X TXQ0X0Y��   !?  N�x &�  �   �~  &,�@   ڰ  ',]   ˕ (,�  �U *�  ��  +.>  ]�  Y-Q  8  �N  9  �� :    .>  E,� 
�   C�  0� 
�-(4  J�  
�-�   E�� 
��  �  0� 
�2(4  J�  
�2�  Ũ 
�2�  �� 
�2�  �e 
��,  l�  
��3  c� 
��.  ހ 
�4  �U 
��  D�  
�D]�  
�ڰ  
�]    �,  {t� 
~ �D     }       ���  0� 
~)(4  ˤ �� 0  ڰ  
�]  A� =� nn 
��  3J�D     :       ��  ހ 
�"4  y� w� c� 
�"�.  �� �� w�D     � U|   O��D     � T�U   <�u 
K�  ��D     ?      �˿  ��  
K)�  �� � �� 
L)�x  ]� U� ϖ 
M)�5  Ǧ �� |�U 
O�   ڰ  
P]  >� <� 0� 
Q(4  m� c� F�  
w0�D     ˿  ��D      �& 
n��  ܿ  � ާ �& �  � � ��  B� >�  �  � y� �  Ш ̨ �  � 	� #�  b� \� -�  �� �� C9�  ��D     5B�  M�D     4      �  G�  ש թ S�  �� �� _�  <� 4� 5k�  `�D     k       ��  p�  �� �� '|�  ��p�D     � ��  Uv T�� ��D     � Uv Q��  I��  ��D     }       ��  6� *� '��  �� �D     � �  Uv T~  ]�D     � Uv T~ Q��   5��  ��D     !       O�  ��  �� �� ��D     � Uv T|   5��  ��D     :       v�  ��  ߫ ݫ  ��D     } ��  Uv Tcinu  �D     � Uv T��   %�D     � Q��  NG� 
��  ��   0� 
�;(4  �U 
��  ��  
��  �� 
�  p� 
��<  )ss 
��  )i 
��  �� 
��  D�  

"��  ހ 
�4  � 
�	1  x  
��0  "��  �_ 
��  J�  
��   �_ 
��  J�  
��    "��  ހ 
�4   "��  J�  
�   nn 
�    N�� )�  &�   x )*�   �7  **�*   Mj  +*�-   �e ,*�,  �U .�   R�� �  ��D     3       ���  L�7  )�*  UL�e )�,  T}y�  ��D      ��D            ��  � � ��  � � ��  *� (�   E�� ��  J�  x �&�  �7  �&�*  Mj  �&�-  �e �&�D  �U ��  dim �Z   F�  2	z�D     �� 	�G  1� 	�  �� 	c    8� ���  �7  �,�*  4dim �,(=  �~  ��@  V� �!?  �� �!?  {� �!?  g� �   seg �.>  "��  c �q=   �� �c  c �q=      8� X�  �7  %�*  4dim %(=  �~  �@  V� !?  �� !?  � �  {� !?  �`  !?  �� c  ��    @v !   � "c  D�  �"��  �� 3�*  �� 4!?  Ɩ 4!?   "��  Ɩ j!?   ";�  �� !?  Ɩ !?  �� !?  �� c  a� c  & c   �j  a!?  R  a!?    <� �c  ��D     \      ��  �7  �'�*  U� M� {� �'!?  Ŭ �� Ɩ �'!?  l� `� �`  �'c  � �� Hdim �'(=  �� �� K{ �c  � � �� �c  �� �� � �c  � � n� �c  �� �� w� �c  ױ ű � �c  � � ҧ �c  6� $� � �c  =� 5� ٧ �%c  �� �� �� �-c  K� ;� �  �c  �� �� �  �c  Y� O� F�  ��D     ��D     ��  Q�XR| v 9��  �U  8W� {O�  �7  {+�*  Ǟ  |+!?  Q� }+!?   8g� a��  �7  a,�*  4dim b,(=  � c,!?  �� d,!?  �  fc  N� hc   EQ� �c  Y�  �7  �-�*  4dim �-(=  5�  �-c  �� �-�  �� �-�  �e ��D  �~  �SD  �  �c  �} �  <  �   D�� V�� c    <�� �c  p�D     w       �B�  Չ � �*  Է ̷ /� � �  >� 6� B5�  � c  Qn ��  �� �� �� �c  � ܸ D� �c  7� /� ��  �c  �� �� &��D     "       w �c  �� �� �  �c  &�  �   <v{ h�  ��D     �       ��  B�7  h%�*  U�e i%�D  �� �� t k�  � غ "� lP  L� B� � l#P  ɻ �� ;y�  ��D      ` o��  B� @� ��  B� @� ��  g� e�   A��  �D     �      �n�  �7  3�*  �� �� �e 3�D  ˼ Ǽ Hdim 3(=  � � �~  �@  G� A� {� !?  Ƚ ƽ �� !?  � � cjk SD  +� '� 1� �  �� �� f� c  � � 3��D           �  bb *�  6� 4� �� +�*  ^� Z� �� ,c  �� �� 0 �� 1rC  � � �v 2   &� "� �� 2(   r� p� &�D     ~       �  Gc  �� �� �F  H�*  � � Y��  d�D      d�D            V��  ��  7� 5� &d�D            ��  ^� Z� ��  �� ��      ;��  n�D      � ��  �� �� ��  � � � ��  K� G� ��  �� ��    Ey ��  ��  �7  �0�*  4dim �0(=  �U ��   EA� ��  }�  �7  �.�*  4dim �.(=  �~  ��@  �U ��  ڰ  �]  C� �SD  X� �.>  T� �.>  seg �.>  1� ��  �� �c  D�  �D�� �"��  �  !?  �� c  ee   "��  {� $!?  �  %c  �� 1.>  ˿ 8.>  a� 9c  �� >.>      {� U!?    V� �!?  �� �!?  {� �!?  �� �  �� �  N� �   Ɩ �!?  #� �.>  �� �c  �{ �c        8{ P��  �7  P.�*  4dim Q.(=  �~  S�@  X� T.>  T� U.>  �� Ve=  ˿ W.>  #� W.>  � Xc  �� Yc  "I�  �  kc  min rc  max sc  len tc    �� �.>  �� �.>  seg �.>  �� �.>      EC� $�  %�  �7  $1�*  4dim %1(=  �~  '�@  X� (.>  T� ).>  �U *�  seg +.>  pt 6q=  ��  7q=  f0 8�  f1 9�    Aq�  �D            �r�  B�e .�D  UBN� .�-  TB,� .�-  Q A�� ���D     X       � �  �e �(�D  �� �� $� �(�,  8� 0� �D      �  ��  Us Tv Q0 O��D      �  U�UT�TQ1  A�{ ���D     �      �v�  �e �,�D  �� �� $� �,�,  	� � Hdim �,(=  o� k� 1� ��  �� �� �� �c  �� �� �~  �SD  &� � nn ��  �� �� � �� �rC  H� @� �  �c  (� $� !� ~�  ��  �c  �� �� P�  �c  �� �� ��  ��D      � �i�  ��  � � ��  Y� U� � ��  �� �� ��  � 
�   �D      T   ��  X�D       � ���  ��  z� x� ��  �� �� � ��  �� �� ��  	� �   ��  ��D      � �*�  ��  F� D� ��  k� i� � ��  �� �� ��  �� ��   ;��  ��D      0 ���  � � ��  0 ��  9� 5� ��  |� x�     <ʭ ��  �E     `       �p�  �e �'�D  �� �� ��  �'�  &� � �� �  �� �� �E     } ��  Us Tcinu �E     � �  Us T|  �E     f�  5�  Uv Ts  �E     �  S�  Uv Ts  �E     �	 Uv 9��  s   8� @�  �e @/�D  ��  A/�  � C   �� C   � D�  �� D�  � K�  �t La   *� Pu�  p Qn  x \�  T� ]-     A��  �D     �      �f�  �e -�D  �� �� ��  -�  *� &� 7�� !�  ��y7�� !�  ��|�� !�  p� b� }� "�  � � |# $   �� �� �� &rC  <� 4� �U '�  �� �� �~  (SD  � � Mj  )�  v� h� sc +4  ,� *� bss -;*  T� P� bs .1�  �� �� 7� 5�  ��y�t 6a   �� �� �; p Hn  *� � �� I�-  �� �� �� J�-  p� h� !< a�  x l�  &� $� �� mc  Q� I� *� n  �� �� N5  o�  7T� q-   ��y!`< ��  nn �  o� k� ��  �  �� �� ��  �  � � �< pp �  �� u�   G	e  ��D      ��D            ��  Oe  	� � Be  	� � 5e  	� � (e  /� -� e  W� U� &��D            \e  |� z� ie  �� ��   ��D     }e  G�  Us T} Q��yR��y ��D     > U~ Q1  3�E     ?       ��  ref c  �� �� �� c   � �� ��    7� 5�  jb�  z E     g       ��  {�  o�  &z E     g       ��  e� _� ��  ��  �� ��   kb�  � E     {       �{�  o�  &� E     {       ��  �� �� ��  ��  ?� =�     Vd� E��D            ���  -�e E.�D  � w� -��  F.�  �� �� @�7  I�r  ��}]�  �!�: ?�  �U X�  6� 0� x Y�  �� � :dim ZZ   �� �� @��  [��  ���~$� \�,  {� y� ހ ^4  �� �� � _	1  �� �� @� f�  ��}�t ga   J� D� :p jn  �� �� 3K�D     :       m�  @T� {-   ���~l	e  {�D      {�D            �H�  Oe  �� �� Be  �� �� 5e  �� �� (e  �� �� e  &� $� &{�D            \e  K� I� ie  s� q�   q�D     }e  Ts Q��}R���~  !0; l�  �~  �SD  �� ��  u ��@  �� �� :seg �.>  V� R� ��  �.>  �� �� �� �#.>  "� � @I� ��  �ܴ}!`; 	�  �  �c  �� ��  >�D     G�  '�  Uv T|  U�D     G�  O�  Uv T0Q0R|  ��D     ��  U�ܴ}Tt   !�; ��  �~  �SD  �� �� n� �c  P� F�  My�  �D       ; ���  ��  �� �� ��  �� �� ��  �� ��  ��D     > ��  U| Q1 ��D     � #�  U���~T0Q
�r �D     �  Uv T}�  M��  �D       P: Rt�  Ǹ  $� "� ��  K� G�  ��D     ��  Uv   %�D  ��  +S     V7� �@�D     �      �b�  -/� �*vv  �� �� L�B �*�*  T-�  �*c  � � :i ��  �� �� :j ��  � � e� ��  ]� M� �� �c  � � :sum �c  H� B� uL  ��*  �� ��  [�� ���   /� ��   �B ��-  )i ��  )j ��  uL  �c   NVJ  �C  ��  aa �C  ab �C  )ret �.  )tmp �.   =��  ��D     �      ���  ��  	� �� ��  �� �� ��  n� l� ��  �� �� ��  ��  ��  �� �� �  h� R� �  G� � &�  �� �� 3�  U� E� C@�  ��D     (I�  �  ��  J�  O� I�  �D     Y�  ��  Qq  3�D     Y�  Qq   =��  �D     Q       �9�  ��  ��  ��  ��  ��  �� �� ��  �� �� Ʊ  �� �� ӱ  � 	�  =��  @�D           ���  �  B� .� (�  =� � 5�  �� �� B�  � �� SO�  � �  �  \�  �� �� i�  _� G� v�  N� &� ��  �� �� ��  w� c� C��  (�D     (��  �  1�  ��  �� �� *��  �  ��  � �� *Ƃ  ! ǂ  �� ��    *ׂ  @! ؂  5�  �D     8       f�  �  W� Q�  X�D     ��  ~�  Qq  ϷD     ��  Qq    =��  ��D     K       ���  ��  �� �� ��  �� �� �  p� f� �  �� �� �  &� "� 5��  ȹD            s�  ��  _� ]� �  �� �� �  �� �� ��  �� �� &ȹD            �  �D     ��  9��  s 9��  v    ��D     �  Us Tv   =n�  �D     �      ���  ��  /  '  ��  �  �  ��  �  �  ��  ��D       �! ��  ��  5 1 ��  o k �! ��  � � ��  � � ��    ��  ` ^ ��  � � 5��  @�D     L       ��  ��  � � ��  � � �  "  �  d `  $�D     G�  U T|    *n�  �! ��  � � ��  % ! �! ��  }�  ��D      �! H�  ��  c [ ��  � � �! ��  - # ��  � � ��  Q M ��  � � ��  I ? ��  � � ��  5	 1	  �  �	 �	 5�  .�D     �       ��  �  
 
 *�  @"  �  U
 Q
 -�  �
 �
 :�      (I�  p" 2�  J�  B 8 W�  � � *d�  �" e�     *r�  �" s�  @ :    ׺D      U�   ;��  s�D       # ��  � � ��  � �  # ��  H B ��  � � ��   � ��  � { �   � �  A 9 "�  � � /�  r n <�  � � \I�  CR�  ؼD     (��  `# ��  ��     ��  ) % �  g _ *�  �# �  � � &�  1 ) *3�  �# 4�  � � *A�  $ B�  � � O�    *\�  `$ ]�  Y U j�  � �      ��  ֽD       �$ �  ��  � � ��  � � �$ ��   � ��  E A   ([�  �$ ��  `�  � � m�  � � z�  $ " (��  �$ ��  ��  L H ��  � � *��  0% ��  � � I��  ��D     ^       ��  � � ��  6 0 *��  `% ��  � �     I��  ��D     �       '��  ��G��  �D      �D            gQ�  ��  ��  � � &�D            ��  #  ��  y u   ��D     %�  U��Q} 8$8&R0X��Y��   ��D      U@      =[�  ��D           ���  i�  � � u�  = 3 ��  � � ��  � � ��  Y M ��  � � ��  � � ��  � � ɭ   � խ  = 7 �  � � �  � � I��  h�D     t       ��    ��  ��D      �% ��  ��  ��  ; 7 �% ��  z v ��  � �   {�D      T} v    =�x  0�D     �      �C�  �x   � �x  �x  �x  y   w y  !y  � � .y  g a ;y  � � Hy    � Uy  V  N  by  �  �  oy  1! +! |y  �! �! �y  " �! �y  �" �" �y  # # �y  x# p# �y  �# �# �y  J$ @$ �y  �$ �$ C�y  ��D     C�y  2�D     C�y  X�D     ��  �D      p& �j�  ��  '% %% ��  P% J% p& ��  �% �% ��   & �%   5Mz  2�D     F       �  Nz  U& S& [z  hz  z& x& =�D      ��  Ts  ^�D     d ��  U|  $ &Tv  $ &Q  $ & l�D      U~ ����Ts   5"z  ��D     h       ��  'z  �& �& 4z  Az  �& �& ��D      a�  Ts  �D     d ��  U|  $ &T~  $ &Q��� $ & �D      U ����Ts   G��  0�D      0�D            �)�  ��  
' ' ��  /' -' &0�D            ��  V' R' ��  �' �'   5�y  p�D     �       ��  �y  �' �' 	z  z  ( ( ��D      y�  Ts  ��D     d ��  U|  $ &T  $ &Q��� $ & ��D      U���@$����Ts   Y�D      ��  U�B$ ��D      
�  Ts  ��D      "�  T}  e�D      Uv ����Ts   =�v  ��D     4      �|�  �v  F( :( �v  �( �( �v  ) �( �v  �) �) i�v   �v  �) �) 3 �D     @       ��  �v  �v  �* �* �+ w  �* �*   !�+ ��  w  �* �*  *�v  , �v  D+ 8+ �v  �+ �+ �v  I, -, �v  |- x- , �v  �- �- �v  (nw  P, L�  sw  �- �- w  *. (. �w  Q. M. �w  �. �. �w  �. �. �w  �. �. �w  '/ #/ �w  b/ ^/ �w  �/ �/ '�w  ��I�w  q�D     n       �w  �/ �/ '�w  ���w  ��D     � *�  U| T��Q: ��D     � U| T��Q:   5\w  ��D            s�  aw  �/ �/  5$w   �D     @       ��  )w  0 	0 '5w  ���D     2x  T��Qv   5"x  ��D            ��  #x  00 .0  (Bw  �, +�  Gw  W0 S0 Qw  �0 �0 ��D     � U| T0Q:  Ix  	�D            	x  �0 �0 x  �0 �0 �D     � U| T0Q:     =ca  0�D     �      �2�  pa  1 1 |a  �1 �1 �a  .2 "2 �a  �2 �2 �a  ,3 "3 �a  �3 �3 �a  4 4 �a  ?4 =4 �a  d4 b4 �a  �4 �4 �a  �4 �4 �a  45 *5 
b  �5 �5 b  ?6 96 b  �6 �6 +b  �6 �6 ~�a   57b  ��D            ��  <b  t7 p7  M��  ��D      �, 	���  ��  �7 �7 ��  �7 �7 �, ��  	8 �7 ��  �8 �8   M��   �D      - 	�.�  ��  /9 -9 ��  T9 R9 - ��  ��    (Gb  �- I�  Lb  9 w9  (Zb  �- Y�  _b  �9 �9 lb  : : yb   ; �: �b  �; �; ��  ��D      . 	X��  ��  *< (< ��  O< M< . ��  x< t< ��  �< �<   u�D      ��  T�� ��D     �b  Uu Tt Q'v t  $ &��t  $ &��?&"#��@&Rv X} Y	~ 2$~ "1$  I�b   �D     g       �b  �< �< �b  = = ��  �D      `. 	d��  ��  F= @= ��  �= �= `. ��  �= �= ��  > �=   ;��  ?�D      �. 	f��  ?> => ��  d> b> �. ��  �> �> ��  �> �>     =��  ��D     �      �Q�  ��  ? ? ��  V? H? ��  �? �? ��  4@ 0@ ��  v@ l@ �  (��  �. ��  ��  �@ �@ ��  GA AA ��  �A �A ��  �A �A �. ��  rB jB �  �B �B \�  ��  ��D      @/ )		%�  �  �C �C �  XD 8D @/ �  �E �E )�  ,F F 6�  G �F C�  H �G P�  EH )H ]�  yI cI j�  wJ eJ w�  UK =K ��  lL VL ��  vM TM C��  #�D     (��  �/ ��  ��  �N �N ��  -O %O ��  �O �O ;O�  4�D      00 Zw�  P P w�  P P ��  @P >P ��  @P >P j�  eP cP ]�  �P �P 00 ��  �P �P ��  �P �P T�D     ��  Q��~�9��  ~     (��  `0 g�  ��  Q Q O�   �D      �0 �	^�  w�  {Q yQ w�  {Q yQ ��  �Q �Q ��  �Q �Q j�  �Q �Q ]�  �Q �Q �0 ��  R R ��  RR PR C�D     ��  Q��~�9��      O�  x�D       1 �	�  w�  wR uR w�  wR uR ��  �R �R ��  �R �R j�  �R �R ]�  �R �R  1 ��  S S ��  NS LS ��D     ��  Q��~�9��      ��D     X�  5�  U Ts Q} R0X0 p�D     X�  U Ts Q} R��~X��~�  (��  `1 ��  ��  wS qS ��  �S �S �  ,T &T �  }T uT  �  �T �T -�  .U &U  �  r�D      �1 V	 �  '�  �U �U 4�  �U �U 4�  �U �U A�  �U �U A�  �U �U  *;�   2 <�  %V V I�  �V �V G�  ��D      ��D            v��  '�  �V �V 4�  W W 4�  W W A�  DW BW A�  DW BW  G�  )�D      )�D            t�  '�  iW gW 4�  �W �W 4�  �W �W A�  �W �W A�  �W �W  W �D     d    J�  #�D      P2 *		�  e�  �W �W X�  YX OX P2 r�  �X �X �  xY pY ��  �Y �Y ��  �Z �Z ��  [ [ *��  �2 ��  5[ 1[ 5��  ��D     L        �  ��  m[ k[ I��  ��D     >       ��  �[ �[   *��  �2 ��  �[ �[     5 �  ��D     �       N�  '!�  ��~'.�  ��~';�  ��~M�  ��D       3 #	"�  h�  �[ �[ [�  \ \ [�  \ \ ��  <\ :\ u�  a\ _\ 3 ��  �\ �\ ��  �\ �\ ��  �\ �\ ;��  ��D      @3 ���  ��  <] 8] @3 ��  �] �] ��  �] �]     ��D     |�  U��~T��~Q��~R��~  ��D     n�  k�  U T1 ��D     �  ��  U T��}Q1 �D     U�  ��  U��~T|  �D     ��  ��  U��~T|  F�D     ��  9��  { 9��  ��}   �D     �  �  U T��} r�D     n�  /�  U T0 ��D     �  U T��}Q0  =�}  ��D     =      �-	 �}  ^ ^ �}  x^ Z^ �}  �_ �_ �}  �` �` ~  va ja ~  &~  (�}  p3 � �}  
b b �}  vb nb �}  �b �b �}  d �c p3 ~  �d �d ~  &e e &~  *f "f \3~  P�  +�D      �3 �	N  k�  �f �f ^�  �f �f �3 x�  g g ��  ^g Zg ��  �g �g ��  �g �g ��  5h 1h *��   4 ��  th rh Ƅ  �h �h ӄ  �h �h ��  ji bi (�  @4   �  �i �i ��  2j 0j �  Wj Uj �  |j zj *"�  p4 #�  �j �j (0�  �4 ��  1�  l l Y��  ��D      ��D            
��  ��  dl ^l &��D            ��  �l �l ��  <m 8m    Y��  0�D      0�D            �	��  ��  }m wm &0�D            ��  �m �m ��  6n 2n     ;��  ��D      �4 �	��  ��  �4 ��  ��       n~  i�D       5 	 �~  }n qn |~  %o o 5 �~  qp ep �~  q q �~  lq Tq �~  zr lr �~  ds <s �~  1u u �~  w �v �~  2x 0x �~  Zx Xx   �x �x (a  �5 � f  
y �x (�   6 � �  �y �y �  �y �y �  Bz >z 	�  �  �z �z #�  &{ "{ 0�  u{ i{ =�  | | IJ�  {�D     �       K�  �| �| X�  } }   (s  p6 Y x  Z} T} �  �} �} �  �  �} �} �  7~ 1~ �  �~ �~ �  �~ �~ �  "  M�D     +�  U} T��}�Qs Rv   R�D     +�  U} T��}�Qv Rs   (  �6 �   y m *  � � 7  ـ π (D   7 � E  P� H� R  Ɓ ��  ��D     +�  U T1Rv   (h�  @7 h m�  8� 4� z�  v� p� ��  ł �� ��  � � ��  p� j� ��  ȃ �� ��  e� a�  *ɀ  �7 ʀ  �� �� G��  n�D      n�D            [� �  � � �  � � �  � � �  >� <� �  >� <�  *׀  �7 ؀  g� a� �  �� �� W��D     d     ��  ��D      08 	# Ұ  �� � Ű  `� X� 08 ߰  Ć �� �  g� _� ��  ˇ Ç �  +� '� 5M�  �D     9       � N�  g� a� [�  �� �� h�  ۈ ׈ u�  � �  I�  �D     9       �  >� 8� %�  �� �� 2�  �� �� ?�  � �    C�  ��D       �8 �: |�  � � o�  O� K� b�  �� �� U�  ъ ˊ �8 ��   � � (C�  �8  |�  k� i� o�  �� �� b�  �� �� U�  � ߋ �8 ��  � � �D     G�   U Tv Q��}#hR0 �D     ��  U T0   ��D     G�  U T0   C�  ��D       �8 �O |�  +� )� o�  Q� O� b�  ~� |� U�  �� �� �8 ��  ߌ ی (C�  09 4 |�  � � o�  =� ;� b�  j� h� U�  �� �� 09 ��  �� �� �D     G�   U Tv Q~��R1 �D     ��  U T1   ��D     G�  U T1   5D~  0�D     q       � 'E~  ��~'R~  ��~'_~  ��~M�  T�D       p9 	W h�  ٍ ׍ [�  �� �� [�  �� �� ��  $� "� u�  I� G� p9 ��  r� n� ��  �� �� ��  Ԏ Ύ ;��  p�D      �9 ���  ��  $�  � �9 ��  r� n� ��  �� ��     G�D     |�  U��~T Q��~R��~  `�D     U�  � U Ts  j�D     ��  � U Ts  ��D     ��  9��   9��  ��~   ��D     �  � U T��~ �D     9�  Q��}�R��~X0Y| �  =�f   �D            �k	 Sg  USg  TS%g  Q2g  � ��  =�f   �D            ��	 S�f  US�f  T =p�  �E     �       �& ~�  7� -� ��  �� �� ��  �� ֐ ��  [� Q� '��  ����  ב ͑ '��  ����  M� G� '��  ����  �� �� *��  �< ��  �  � '�  ��G	e  $E      $E            e�
 Oe  <� :� Be  f� `� 5e  <� :� (e  �� �� e  ߓ ݓ &$E            \e  � � ie  ,� *� BE     q T| Q
R��   E     }e  Us Tv Q��R��   =	e  �E     :       �� e  S� O� (e  �� �� 5e  ͔ ɔ Be  
� � Oe  I� C� \e  �� �� ie  �� �� �E     q Tv Q
R�R  >�Q  �Q  �T�s  �s  0�T�`  �`  0vT@  @  �>�a  �a  >CA  CA  E>�C  �C  w>\P  \P  >%O  %O  �>zE  zE  �>�J  �J  �
>F>  F>  kT�I  �I  0�>e  e  �T>m  >m  1y>@R  @R  8>�E  �E  WD  D  3 >Q  Q  ^>�_  �_  A>�n  �n  �T$  $  2. ˛   �b  &  �� �:  �E     �=      '= ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  s&  G   �  N   )  	A"]  c  �   	��  �  	�U    ��  	��  <h 	��  �I  	��   �  	X�  �  U   �  Q  -    �   	m�  �  �  Q  U    f  	��  �  U     Q  -   -   U    J   	�")  /  �  P	H�  Ǟ  	J,   ֳ  	K@   pos 	L@     	N�  /[  	O�   �K 	P�  (�R 	Q9  0ڰ  	SQ  8O�  	T,  @��  	U,  H �  	��  <v 	�-   ��  	�U    �  	��  ""  	�    @   ,    @   ,  @    2  �  �   	F  L  W     v  
:-   �  
L�  x 
NW   y 
OW   �  
Qc  	�  ~   
w�  
  
yW   �!  
yW  �   
zW  H  
zW   "  
|�  �  (
e  M} 
N    5�  
N   `�  
	G   _| 

,  
!  
0  ?   
2  2   
2  B  
U     �  
�  	e  �  (
Q�     
S)   0�  
T)  N5  
V�  �   
W�   H� 
X�  �1  
ZG     �  )  �  
\w  �  �  N   
�7  �!   �   pmoc�  stibu!  ltuo�  tolp :  
��  �8  
5"Q  W  �$  �4  
S�  x 
U)   len 
V0  e� 
W2   �#  
Y\  	�  �%  
{�  �  �  G   G   �  U    �  �#  
��  �  G     G   G   U    �.  
�    ,  G   G   U    �8  `
��  .  
 �   �; 
�  �1  
G   �5  
�  �+  
�   `(  
�  (�/  
  0�  
U   8*  
�  @ r  �  u(  

,  	�  �2  
(�  �  G   �  U   �   D  �3  
;    #  D   v)  
]0  6  K  D  ,  @    �3  
yX  ^  G   w  D  @   U    H7  
��  �  G   �  D  �   �  51  0
�  y2  
�7   � 
��   
�#  *
 
�K  / 
�w   $ 
�  ( 2$  
��  -4  l2  +  �,  �  $8  �2  	3  ?    ��   	J  {"  �)  	[  !  �0  \   �G   �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U   +D  C4    :   �	  xx ��   xy ��  yx ��  yy ��   5  ��  		  8  �\	  ��  �D   ��  �x   $  �1	  c   �v	  |	  �	  U    �  ��	  Kl  �U    �  �i	   s  ��	  �"  $�	  �	  �   +
  �� -�	   �W .�	  Kl  /U    %  D6
  uR F�	   �
 G�	   }  I
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<  5�  >W   ��  ?W  �"  AW  �"  BW  i!  CW   %!  EW  (2!  FW  0�  GW  8   I�  �"   sg  ��  u[   5�  v[  ֳ  xW  !  zW  m  {W   v  }  J  �#�  �  �!  �}E  ڰ  Q   {3  �x  S0  �x  �/  �x  �1  ��  �1  �|!  Y/  �6
  �*  ��  (�)  �E  0+:  ��!  8<8  ��!  X�*  �x  � �3  �"R  X  �(  ��  Oe �c!   �-  �t  ڰ  �Q   U  �"�  �  �  8�  ah !i!   Oe "d  U1  #6
   ;+  $�  0 i(  �$�  �  l;  ��o  ah �i!   Oe �v!  y2  �7   {:  ��  (�� �D  h/ �w  p�� ��  x T   � |  �  _  �C  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"  x  8�  �  @`  !x  Hd  "�  P�@  $�	  X�;  )�  h�   +l  ��  ,[  �
  -[  ���  .[  �?!  0[  ��  1[  ��  3[  ��  4[  �ȩ  6�  �ֳ  7C  ��� 8�  �K <�  �ڰ  =Q  �^�  >  �U  @6
  �t  B�	  �k  CU   ��L  E&  � "   P  V  1  Xm�  ��  oo   �@  p�	  �e q�  �L  r�  P @  $%�  �    0\�  �-  ^t   ��  _o  �W `�  x a�  �@  b�	   �e d  0�"  e�  pi"  f�  x� g�  ���  i7  �.a ke  ��  lx  �J  mx  �Mj  o�  ��  q�  ��  r�  �M  tU    Z  u-   _"  wW  (   xW  Ud zU    �L  |  ( �!  F#    Z!  AT  ��  Co   T D  �!  El  "  Fl   S  N   �  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  T  0  `)3  9  �"  �e�  �1  g	   H+  h�   x+  ix  0��  k�  8�)  n#]!  h�'  q   p��  r7  t�*  yx  x J  g  �  �  �)�  �  �!  H�  $  �U    7:  ��  s4  ��   b  8H�  !  Jl   m  Kl  A� M�  �� N�  �  PW  
  QW   ��  RW  (�  SW  0 �  U  x   �$�  �  �!  0'  ad  )x   �1  *l  &D  +x  2B  ,x  x� -	     �)    �"  P��  ��  ��   �1  ��  �&  �  �3  �	  ]7  ��  0�7  �U   @�1  �7  H P6  �  tag �   Kl  �   �6  	�  �  �5  N   
�  i7   �&  9  F9  8%  �*   �,  
�  ./   6
`  b 8
�   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(m    �8  N   ��  �:   4,  �6  $  �/  l9   �2  �s  3  �#  ��  �'  ��  �  �  �  E   �2  ��  �    E   l/  �    �  .  E  .   �   ;)  H��  �#  ��   :  ��  �5  ��  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  ��  8��  �  @ V  �-  �4  	�  d)  s�  �  �  �  U    9  F#  	�  �$  @Jw  �#  L�   y2  M7  W� O�  �� P�  �,  Qi   M4  R  (�;  SA  0�*  T�  8 c/  X!�  �  �-  (q�  �-  st   Oe t�  ��  u7  � v�   �  �/  )�  �  �  �  w  �   g%  .  	    w   �.  1   &  ;  w  ;  �   ,	  73  6M  S  c  w  c   �  �8  :u  {  �  �  w  w   "3  >�  $)  Y�  �  �  �  �  �  �  �   �6  _�  �  �  �  �  �  ;  �   �3  f    "  �  �  c   ;0  l.  4  �  M  �  �  �   �&  x��  ah � �   y2  � 7  H�8  � �  P�8  � �  X�'  � �  `� � "  h�9  � �  p   �.  �M  "9  H2  Mj  4�   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :�  T%  �=�  ڰ  ?Q   �0  @�  q5  A�  L)  B�  )  C  Ǟ  E  �  F  `Ud HU   � X+  J�  #  1  �  �  �  �    o  x  x  �   �&  &�  �  �  o   �1  *	    �    C   �6  -*  0  ;  C   w-  1G  M  �  \  �   �;  4h  n  y  �   =;  8�  �  �  �  C  `   B$  <�  �  �  �  C  �   2  @�  �  �  �  �  C  �  7   7  G    �  %  o  �  �  �   q8  N1  7  �  K  o     )2  SW  ]  �  �  o  �  �  7  �   �  k.  ��d  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q ��  hZ)  ��  p�#  �  x'0  �;  �.  �\  ���  ��  �� ��  �`9  �%  ���  �K  �5  �y  �U#  ��  � �2  �p  �  �&  0��  y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  �v  *  V'�  �  �0  �*   u?   |#  w�   �#  x�  � y�  C4  z�   �&  |�  �'  �W   ]   �  v   �  �  v    \	  �9  ��   �   �   �  v    A2  ��   �   �  �   �  �    �    ?   8(  !  ��  )K    $�  )|   �-  )�    )  �   	!  3  <J!  �� >%J!   ��  ?%�   !  #  A!  P!  �  �(  �X  �  E  �!  @    �  �!  @    �  �!  @    H'  �%  ��  ��#  ��  �x   ��  �x  *�  �3  ��  �3  	��  �3  
�  �3  .�  �#  ��  �#  (��  �#  <�  �#  X0�  ��  pY�  �x  xA�  �x  |M�  �,#  ���  �,#  ���  �3  �W�  �3  ���  �  ��  �  ���  �<#  �[�  �<#  ���  ��  ���  ��  ���  ��  ��  �L#  � [  #  @    [  ,#  @   	 l  <#  @     [  L#  @    [  \#  @    c�  ��!  8�  �\#  �  $�  )$�#  �#   P�  p��#  ڰ  �Q   _� ��*  !��  ��*  8 a�  ,�#  �#  �  �#  Q  �#  �#   h#  z#  ;�  1$  $  +$  z#  �  �  �  �   w�  87$  =$  H$  z#   *�  ;}$  � =�#   �� >�#  �� ?+$   � AH$  M�  A�$  H$  ��  h!�$  �$  ��  ��  u-�$  5%  ��  8V5%  �7  X�$   ��  Y:%  �R Z�%  �� [W%  �� \~%   �� ]�%  (a� ^�%  0 	�$  t�  �F%  L%  W%  �$   S�  �c%  i%  ~%  �$  �  �   !�  �c%  ��  ��%  �%  �%  �$  �   e�  
�%  �%  �  �%  �$  �   |�  1�%  �%  �  &  �$  &  z#  �   �  l� `�$  �  �!$&  *&  ì  ��  �-<&  �&  �  8��&  �7  �&   ��  ��&  �R �X'  O� ��&  �  �'   y� �0'  (a� �'  0 	B&  ��  ��&  �&  �&  &   ��  ��&  �&  '  &  �  x  �   i�  �'  '  0'  &  �  �  D   p�  &='  C'  X'  &  �  D   !�  De'  k'  �  '  &  �   %�  j�'  �'  �  �'  &  &  z#  �   �� �B&  ��  ��'  ��  �(   �� �(  � �/(   �$  (  E   �'  �$  (  E   (  /&  /(  E    (  ��  ��'  	5(  0� @|(  org Bx   cur CW  fit DW   M� FG(  � F�(  G(   �� �J�(  /� L�   Չ M�(   |(  �(  @    �� O�(  �� O�(  �(   ]� �R))  n� T�(   !W� U�  �!J� V�  � @� X�(  �� XA)  �(  l� 0\�)  0� ^x   l� _x  � `x  r� ax  �� cW  z�  dW  )� eW   �� fW  ( h� hG)  n� h�)  G)   �� k*  /� m�   �� n*   �)  *  @    [� p�)  �� p,*  �)   �� 8t�*  � v*   !v� w*  !J� x*  !� y*  	!0�  {�   !Y�  |x  (!� }x  ,!A�  ~x  0!��   4 �� �2*  � ��*  2*  ))  �*  @    �� �!+  � �G    g� �W  0� �W   }� ��*  #� �9+  �*  �� 4 K+  Q+  O� E�+  pos Gx   len Hx  �1  I�   "�� N   7�+  � ��  � <�+  � T�+  ��  V�   �� W�  �7  X?+   5� Z�+  L� Z�+  �+  � ^F,  $� `�   �� a�  Vu  b�  t�  c�   �� e,  �� e^,  ,  U� i�,  |� k�   T� l�  �� mR,   � od,  Z� o�,  d,  �� 0s�,  �7  u�+   �� v�,  �� w�,    	� y�,  3� y-  �,  ?� xY-  ڰ  �Q   �U ��  �  �D  I� ��+  _� �Y-   �,  i-  @    �� �
-  �� ��-  
-  4� !�-  �-  �� 03.  � 5x   K{ 6x  �� 7W  �� 8W  �1  9�  �  :�-   � ;x  ( i�  CD.  1� E�   �� F�  min GW  max HW   z� J.  _� J\.  .  �� HM�.  �� O�   ��  P�  �7  Q�-  �  R�.  Q� S�.  � T�   �� U�.  (�y  VP.  0�� W�,  8�� X�,  @ �-  D.  i� Zb.  �� Z/  b.  b� ]$(/  ./  �� H��/  �� �/   �W �/  2 ��/  �1  ��  �� ��  �� �    d� �   !�� ��-  (G� �W  0�� �W  8.� �W  @ 5� ^$�/  �/  j� �0  �k �/   /� ��   G   a20  p� #�� �� #�� ~C�  4� ��1  ��  ��   D� ��  N5  �/  H� ��/  ڰ  �Q  Mj  �&   0� �z#  (N� �1  0<  �  ��� �x  ��� �x  �z� �  �9� �  �]� �  �>� �  �L� �  � �.   1  @    � �20  �� �81  20  N   ��3  ;�  �� "� � ?� Q� �� � '� � 	m� 
�� �� �� �� � .� }� �� {� �� :�  �� !�� "�� #�� $� %�� &�� '� (F� 0V� 10� @�� AU� Qo� R� Sa� T�� U�� V�� W0� X1� `�� a�� b~� c� p�� ��� �|� �q� ��� ��� ��� ��� ��� �-� �O� ��� ��� �v� �� ��� ��� ��� ��� ��� �y� ��� �x� �5� ��� ��� ��� �	� �� �� ��� ��� ��� �^� ��� �N� ��� �o� ��� �� ��� ��� ��� ��� �� ��� �B� �  �� �3  ah i!   �� i-  ��  }$  ���  
&  �� !�'  � �� #�3  �3  $^� _B(  	�eG     %]4  h�  	`eG     &I� �+4  '�� �,+4   �'  (F� �p(E     �       ��5  )�7  �&  �� �� )_� ��  M� I� )/� �x  �� �� )Ԛ  ��  ږ Ԗ *O� ��5  ��}+y �W  ,� &� ,X$ �x  z� v� +n �x  �� �� -�:  )E      )E            ��5  .(;  � � .;  p� n� .;  �� �� .;  �� �� /)E            05;  1/)E     S}  2Uw 2T��}�2Q~ 2R��}   1�(E     ]�  2U   W  �5  @    (h� ��E     9       ��6  3�7  �&  U4_;  �E      �E     8       �.z;  � �� .m;  � � -�C  �E      �E            BS6  .�C  -� +�  4�C  �E      �E            C.�C  T� R�    &� u�6  '�� u,�6   
&  (A� f(E     V       ��7  )�7  f�$  �� z� )_� g�  ҙ ̙ )Ԛ  h�  $� � *O� j�7  �P-�:  C(E      C(E            p�7  .(;  r� p� .;  �� �� .;  �� �� .;  � �� /C(E            05;  1](E     S}  2Uv 2T| 2Q12Rw    5)(E     ]�  5:(E     ]�   W  �7  @    (1� `PE     9       ��8  3�7  `�$  U4_;  PE      PE     8       b.z;  � � .m;  -� +� -�C  ^E      ^E            By8  .�C  R� P�  4�C  sE      sE            C.�C  y� w�    6�� ;�  9  '�7  ;u-  't�  <�  7�U >�  87ڰ  DQ  9dim E�,    &n� �9  '�7  'u-  '�� '�  'Vu  'D  7�U �  :WD  489dim �,  7ڰ  Q  7�� �  7�Q �    &�� �:  '�7  �$u-  't�  �$�  '�� �$�  'Vu  �$D  7�U ��  :WD  89dim ��,  7ڰ  �Q  7�� ��  7�Q ��    &�� �a:  '�7  �u-  't�  ��  7�U ��  :WD  �87ڰ  �Q    &�� y�:  '�7  y u-  '_� z �  'O� { �  7�U }�  :WD  �89dim ��,  7ڰ  �Q  7/� �x  9idx ��:    x  �:  @    &�� I_;  '�7  Iu-  '_� J�  '/� Kx  'O� Lt#  9dim N�,  87�U b�  7ڰ  cQ    &O� <�;  '�7  < u-  'I� = �+   &Z� 2�;  '�7  2u-  'ڰ  3Q   &;� $�;  '�7  $u-  7ڰ  &Q   6S� �  <  ;dim #�,  't�  #�  'ڰ  #Q   6�� ��  �<  ;dim �+�,  '�� �+x  '�� �+x  '�� �+x  'ڰ  �+Q  7�U ��  7/� ��  7y� �R,  :�   <�� ��  �%E     �      ��?  =dim �*�,  �� �� =pos �*x  �� r� =len �*x  #� � )ڰ  �*Q  ̝ �� )�� �*�?  �� �� ,�U ��  � u� ,�1  ��  � � >�  ��&E     ?�J ,�� �R,  ޠ ڠ +idx ��  � � +max ��  �� z� ,�� �?+  D� 8� @I  U&E      �J �T>  .3I  ݢ ٢ .&I  #� � .I  r� n� ?�J A@I  �� �� AMI  � �� BZI  ��CgI  �&E     1�&E     wI  2U}2T��2Q��   @�M  �&E      0K ��?  .�M  ;� 7� .�M  �� {� .�M  � � ?0K A�M  L� H� A�M  �� �� A�M  ٥ ӥ D�M  E�M  'E      'E     `       `.N  (� $� .N  (� $� . N  b� ^� .N  �� �� /'E     `       A,N  �� �� A8N  � � BDN  ��1B'E     j�  2U��2T<2R	�����2Y��     1t&E     �K  2Ts    x  <4� r�   QE     4      �C  =dim r/�,  I� 5� )�; s/D  4� &� )�� t/�  � Ҩ )\� u/�  �� ~� )t�  v/�  .� *� )ڰ  w/Q  u� g� ,�U y�  � � >�  �kQE     @C  'QE       0_ }mA  ./C  Q� M� ."C  �� �� .C  ȫ ī ?0_ B<C  ��-JC  ?QE       ?QE            iJA  .XC  � �� .XC  � � .eC  � � /?QE            ArC  	� � FC  CQE            A�C  D� @�    1gQE     wI  2U 2T~ 2Q��   GMH  �QE      `_ �.�H  �� �� .�H  � � .yH  �� �� .lH  �� � ._H  `� X� ?`_ A�H  ̰ ư A�H  � � D�H  @I  �QE      �_ @�B  .3I  k� g� .&I  �� �� .I  � � ?�_ A@I  %� � AMI  x� p� BZI  ��CgI  8RE     18RE     wI  2U 2T~ 2Q��   H�H  �_ �B  A�H  ز ֲ A�H  � �� A�H  N� L� A�H  }� q� A�H  � �  1�QE     �|  2Uv2Tv2Qs 2R~ I M  v     6�� a�  JC  ;dim a*�,  't�  b*�  'ڰ  c*Q  7�� eR,   &� N�C  ;dim N(�,  't�  O(�  7/� Q�  87�� VR,    &Z� +�C  '_� +$�,   &��  �C  '_�  $�,  'ڰ  !$Q   <}� ��  �)E     �      ��F  )�B �+�,  �� �� )ڰ  �+Q  � � ,v�  �x  {� i� ,}�  �x  B� :� J�U ��   >�  �*E     @�G  *E      �K  E  .�G  �� �� .�G  �� � .�G  .� *� ?�K A�G  h� d� A H  �� �� AH  � � AH  E� A� A%H  � {� A2H  Ÿ �� A?H  � ��   G�F  �*E      �K .�F  g� c� .�F  g� c� .G  �� �� .�F  � ۹ .�F  .� *� ?�K AG  j� d� CG  �*E     K:G  0L A;G  �� �� AHG  � � AUG  :� 8� AbG  o� i� AoG  �� �� H|G  �L }F  A�G   � �� A�G  �� �� A�G  � � @�L   ,E      �L �IF  L�L  L�L  .�L  r� p� ?�L A�L  �� ��   1�+E     �|  2U��#2T��#2Q���2R��  F�G  4+E     [       A�G  Ž �� 1_+E     v�  2Q ����1$ ����"3$      6F� ��  �G  '�B �'�,  'v�  �'�  '}�  �'�  'ڰ  �'Q  7�U ��  :�  �M:G  7�S  ��   87*� �R,  7=� �R,  7�� ��  7�Q ��  7�� �x  M�G  9pos ��  7�K ��  7�  ��   87��  �F,     6� sx  MH  '�B s0�,  'v�  t0�  '}�  u0�  7*� wR,  7=� xR,  9p1 y�  9p2 z�  7�� {�  7�Q |�  7/� }�   6&� 6�  I  '�B 6+�,  '�; 7+D  '&� 8+�  '�� 9+�  'ڰ  :+Q  7�U <�  7�� =R,  :�  l87�K L�  7�� Mx  7�  N�  7�� Ox  9val Px    6l� �  qI  '�B &�,  'ڰ  &Q  '� &qI  7�U �  7/�  �  7�� !R,  :�  . R,  N0� ��  �#E     �       ��J  O�B �'�,  2� *� Oڰ  �'Q  �� �� O� �'qI  � � P/� ��  }� w� ,�U  �  ̿ ƿ ,�� R,  � � >�  $E     G�J  '$E      �I 	.�J  j� h� .�J  j� h� .�J  �� �� .�J  �� �� ?�I A�J  �� �� AK  � � BK  �L1E$E     j�  2U�T2TH2R| ����2Y�L    Q�� ��  K  R�B �(�,  R/� �(�  Rڰ  �(Q  S-Q  ��  S�N  ��  S�U ��   T�� �0E     �       ��K  O�B �&�,  T� N� Oڰ  �&Q  �� �� P/� ��  �� �� P�� �R,  3� -� UiM  `E      G ��K  .�M  �� ~� .vM  �� �� 1pE     ��  2Uv   1�E     ��  2Uv 2Ts   N�� ��  �%E     Q       ��L  O�� �R,  �� �� Vidx ��  c� [� Oڰ  �Q  �� �� P�U ��  G� A� Wp ��  �� �� X�  ��%E     1�%E     �|  2Uv2Tv2Q| 2R�QI M  v   Y�� ��L  R�� �R,  Zidx ��  [p ��   Q�� �x  M  R�� �R,  Zidx �x   Q,� ��  iM  R�� �R,  R/� ��  Rڰ  �Q  S-Q  ��  S�N  ��  S�U ��   Y�� |�M  R�� |R,  Rڰ  }Q   Q�� R�  �M  R�B R'�+  Rڰ  S'Q  R�� T'�M  S�U V�  S/� W�  S�� X?+  \�  l ?+  Q7� =�  QN  R�B =(�+  R/� >(�  Rڰ  ?(Q  S-Q  A�  S�N  B�  S�U C�   Yp� 2wN  R�B 2&�+  Rڰ  3&Q   N�� Y/&  @E            ��N  ]ϖ Y%E  U N�� Q�$  0E            ��N  ]ϖ Q%E  U NZ� I�$   E            �
O  ]ϖ I*E  U N>� 3�  �E     �       �5P  Oϖ 3%�3  �� �� Pڰ  5Q  �� �� Wph 6U   � � U�;  �E      �F 9�O  .�;  =� ;� .�;  b� `�  ^R  E      E     !       ;�O  .R  �� ��  ^�6  -E      -E     B       =P  .�6  �� ��  E4  vE      vE     B       @.4  �� ��   T� (pPE     �       �R  Oϖ (%�3  � �� _�;  �PE      P^ -L�;  ?P^ A�;  Q� O� @�C  �PE      �^ )>Q  .�C  v� t� L�C  @QN  �PE      �^ %Q  .jN  �� �� L^N  1�PE     ��  2Uv   `�PE     K  "Q  2Us� 2Tv  1�PE     K  2Us� 2Tv   G�C  �PE       _ *.�C  �� �� .�C  �� �� -QN  �PE      �PE            %�Q  .jN  � � .^N  2� 0� 1�PE     ��  2Uv   `�PE     K  �Q  2Us�2Tv  1�PE     K  2Us� 2Tv      &$� R  '�� 2R   }$  (u� �PE     �      ��U  )0� �'z#  \� X� )A� �'�  �� �� )�� �'�  �� �� )� �'�  i� e� )q	 �'�  �� �� +dim �5)  '� !� @A[  �E       0D �U  .i[  }� w� .\[  �� �� .O[  #� � ?0D Av[  �� �� A�[  �� �� A�[  Y� Q� a�[  �E     d       �S  A�[  �� �� Gat  E       `D � .|t  @� <� .rt  z� v� ?`D A�t  �� �� A�t  '� �    H�[  �D  U  A�[  �� �� @at  �E      �D �T  .|t  � � .rt  4� 0� ?�D A�t  p� l� A�t  �� ��   @at  �E       E �gT  .|t  �� �� Lrt  ? E A�t  � � A�t  Z� V�   @at  �E      0E ��T  .|t  �� �� Lrt  ?0E A�t  �� �� A�t  � ��   Gat  E      �E �.|t  >� <� Lrt  ?�E A�t  e� a� A�t  �� ��    K�[  �E A�[  �� �� A�[  M� I� A�[  �� �� A�[  �� �� A�[  �� �� A\  )� %� K\  F A\  m� _� Gat  0E      pF  .|t  6� 2� .rt  z� r� ?pF A�t  �� �� A�t  j� b�       `�E     W_  �U  2U{ 2T0 1�E     W_  2U{ 2T1  <�� ��  0E     �      �0Z  )ڰ  �"Q  �� �� )��  �"�#  >� 8� )�� �"�#  �� �� ,0� �z#  �� �� *�U ��  ��bE0E     A      Z  ,/� ��  G� C� ,�K �0Z  �� }� c`N �V  +dim �5)  � � ,�  ��(  ?� 7�  c�N )W  +dim �5)  �� �� ,�  ��(  �� ��  bS1E     �       �Y  ,Z� ��  1� /� ,� �[  ^� T� -�Z  X1E       X1E     4       ��W  .[  �� �� .[  � 	� .�Z  G� E� /X1E     4       A[  n� j� F+[  p1E            A,[  �� ��    -�Z  �1E       �1E     +       ��X  .[  ,� *� .[  Q� O� .�Z  v� t� /�1E     +       A[  �� �� F+[  �1E            A,[  �� ��    -�Z  �1E       �1E     +       �Y  .[  U� S� .[  z� x� .�Z  �� �� /�1E     +       A[  �� �� F+[  �1E            A,[  � ��    -�Z  �1E       �1E     ,       ��Y  .[  ~� |� .[  �� �� .�Z  �� �� /�1E     ,       A[  �� �� F+[   2E            A,[  ,� &�    1+2E     ��  2U
�  `-1E     #\  �Y  2U��2Q��2X  1S1E     #\  2U��2Q~ 2X}   160E     ��  2U} 2T
p2Q��  [  &� laZ  '0� l%z#  87ڰ  pQ    &�� %�Z  '��  %'�*  'Q� &'x  '�� ''x  'J� ('-+  7�B * *  7/� +�  7�� ,W  7�y  -�)  7n� .x   6� [  ;[  ;num )�  '
Q );[  '�� )[  7/� �  87J� [    g  &�� o#\  '��  o%�*  '1� p%�  '�� q%W  7/� s�  9num t�  7�B u *  M�[  7�  �x   M�[  7�y  ��)   87�� ��)  7�� ��)  7�� ��  7�Q ��  7  � *  7�V � *  87
�  �W     T�� �0.E     �      �}^  O.  �#�*  �� �� O/� �#�  +� � O��  �#0Z  X� P� OF� �#�  �� �� O��  �#0Z  @� 6� OF�  �#x  �� �� O�V �#x  � � P�� � *  n� j� P~� �  *  �� �� P�� ��  �� �� P�� � �  �� �� b�.E     J       o]  ,�y  �)  6� .� /�.E     @       ,�� x  �� ��   c�M �]  ,�y  *�)  �� �� /�.E     :       ,�� /x  >� <�   c N (^  +dim @x  k� a� +top @x  �� �� +bot @ x  %� � ,�� @%x  �� �� ,�y  A�)  �� ��  `w.E     �  T^  2U02Rr 2Xv I�^  �U 1�.E     �  2U12T} 2Q~ I�^  �U  Y�� �W_  R.  �*�*  R�� �*  R*� �*�  R�K �*0Z  R�� �* *  R~� �* *  S�� ��  S�� ��  S��  �  \w  �8SD� �x  S�� �!x  S/� ��  S�� ��)  S�y  ��)  [top �  8S� �x     Tr� *�E     �       ��`  O0� **z#  �� ~� Oh� +*�  �� �� Wdim -5)  �� �� Pn� .�(  �� }� P/� /�  � � P5�  0�(  F� >� P�� 1�(  �� �� P1� 2�  � � c�C �`  Ww ?W  R� L� P�  ?W  �� �� _at  �E       D BL|t  .rt  �� �� ? D A�t  � � A�t  ^� Z�    Eat  �E      �E     !       7L|t  .rt  �� �� /�E     !       A�t  �� �� A�t  � �    d�� �  �a  '�� #u-  'Mj  #&  '0� #z#  ';:  #�  7q�  1  7ȩ  ,1  7�U �  7_� !x  :�  �87� A5)  7� B5)  7A� D�  7�� E�  7=� G�  7~� H�  7��  J�  7k� K�  7�� M    &�� �c  'ȩ  �2,1  '_� �2x  9dim �5)  71� ��  7�� ��  72 ��/  7D� ��  :=� 87�k �/  7��  �/  7�W �/  7c �/  7U� ��  87� �W  70� �W  7�� �$W  7.� �+W  7[� �W  7�� �W  7�� �$W  7A� ��     &�� �d  'ȩ  �3,1  '_� �3x  9dim �5)  71� ��  7ڰ  �Q  71� �d  7T� �
d  7-� ��  7N5  �/  7� �/  7c �/  M�c  7�U �   M�c  7�>  d   87�j  ?/  7R  ?/  9nn @�  89u aW     /  /  d  @    &D� ��d  'ȩ  �3,1  '_� �3x  9dim �5)  71� ��  7/� ��  7c �/  87�� ��-  87�� �W     &�� l.e  '��  l*�*  'ȩ  m*,1  7�B o *  7�y  p�)  7�� q�  7y� r�  7c s/  89y xW  Me  7�� �W   87�� �W     &�� *f  'ȩ  ,,1  '_� ,x  7�B #
/  7�� $R,  7|� %�  7��  &�  7�� 'x  9dim )5)  71� *�  7�  +x  M�e  7�W <�  87/� A�  7c B/    Mf  7/� Q�  7c R/   87/� ^�  7c _/    &�� �{g  '�B �6
/  'c �6/  '/� �6�  '�  �6x  '�� �6x  7�  ��.  7��  ��  87�� �x  7G� �W  M�f  9nn ��  87�� ��-  9d �W    Mg  9nn ��  87�� ��-  9d �W    89nn ��  7K� ��  7�� � �  MKg  7�� ��-  9d �W   Mig  7�� ��-  9d �W   87�� �-      &�� 	 h  'ȩ  	),1  9n �  :w  y:h� L:'� =M�g  7��  /  7c /  7�j  /  7R  !/   87c T/  7�j  T/  7R  T!/    6S� ��  oi  'ȩ  � ,1  'Mj  � &  '�� � u-  '0� � z#  7�U ��  7ڰ  �Q  :�  M�h  7��  ��  7�W ��  9n �%�  7N5  �/  72 ��/  87/� ��  7c �/    87N5  �/  7c �/  9vec ��  9n ��  87�� �x  7h� �x  9dxi �W  9dyi �W  9dxo �W  9dyo � W     &�� [�i  'ȩ  [%,1  '_� \%x  9n ^�  7c _/  9vec `�  7�   a�    &z� 9j  'ȩ  9%,1  '_� :%x  9vec <�  7c =/  7/� >�   6�� G   jj  ;dx W  ;dy W  9ax !W  9ay !W  7�Y  "G    &�� �j  'ȩ  ,1  7ڰ  Q   &�� �ak  'ȩ  �-,1  9n ��  :w  87��  �/  7�k �/  9end � /  7�j  �%/  7R  �-/  7�j  �W  7C  �W  7�o  �W  7�o  �%W  7�� �x  7�� �x  7�� �x    &�� N�k  '�B N/
/  '0� O/z#  '_� P/x  'ȩ  Q/,1  7�� S�-  7/� T�   (� ��2E     z      �9p  )�� � �-  Q� A� )0� � z#  � �� )_� � x  �� �� )ȩ  � ,1  C� -� +dim �5)  R� *� ,1� ��  S� O� ,�� ��  �� �� ?O +pos �W  )� � +len �W  �� �� ,d� �x  � �� ,b� �W  �� �� ,� �!+  �� N� c0P �n  ,�  ��-  �� y� c�P �m  ,� �W  �� �� ,�� �%W  � � ,M�  W  �� �� ,z�   %W  �� �� @at  3E      �P �m  L|t  .rt  �� �� ?�P A�t  3� /� A�t  v� r�   1�7E     �k  2U} 2T| 2Rw   b�8E     @       3n  ,�� @W  �� �� ,8� AW  �� �� ,&� BW  C� ?� ,�� CW  �� ~�  @�p  �3E      Q W�n  .�p  �� �� .�p  "� � .�p  �� �� K�p   Q A�p  c� Y�   G9p  P4E      PQ ]!.Xp  �� �� .Kp  �� �� ?PQ Aep  )� #� Arp  �� ��    @at  �2E       �O �6o  .|t  �� �� .rt  L  J  ?�O A�t  s  o  A�t  �  �    -at  3E       3E            ��o  .|t  �  �  .rt  - ) /3E            A�t  i e A�t  � �   GaZ  g5E       �O �	.�Z  � � .�Z  g _ .|Z  � � .oZ  q i ?�O A�Z  � � A�Z  � y A�Z   � A�Z  7 - A�Z  � �     6�� ��  �p  ;pos �,�  ;len �,�  7��  ��  7P�  ��   6�� XW  �p  ;dim X.5)  ;len Y.W  'd� Z.  87�� `W    Y]� ��q  R�B �1
/  R�� �1R,  S�� �x  [val �x  SO�  ��  [idx ��  S��  ��  S/� ��  MXq  7�� �-  87�Q �    89i1 5x  9i2 5x  7�� 6�-  7�� 6�-  7�  7�.    Q�� ��  Fr  R�B �(
/  R�7  �(�+  R�� �(�,  R�� �(�,  Rڰ  �(Q  S/� ��  S�U ��  \�  �M%r  S�  ��-  S�K �?+   M7r  S�� �R,   8[idx ��    Y$� ��r  R�B �/
/  R�� �/R,  S�� �x  [val �x  SO�  ��  [idx ��  S��  ��   Th� `�E     �       �zs  ]�B `*
/  UVidx a*�  + ' P�� c�-  j d ?@C P\� u�.  � � P/� v�  , * P�� w�-  S O _7t  6E       �C LHt  LHt  .Tt  � � .Tt  � �    Y�� P�s  R�B P.
/  S/� R�  S�� S�-   T�� ?�E     m       �7t  O�B ?(
/  � � Oڰ  @(Q  	 	 `�E     ��  
t  2Uv  `�E     ��  "t  2Uv  1E     ��  2Uv   Q�� 5x  at  R�� 5�-  R�� 6�-   QVJ  �7  �t  Za �7  Zb �7  [ret �"  [tmp �"   e�p  �E     C      �"v  .�p  m	 g	 L�p  L�p  A�p  �	 �	 A�p  T
 L
 Aq  �
 �
 Aq  #  Aq  _ [ A*q  � � ^zs  �E       �E     -       ��u  .�s  1 + .�s  � } /�E     -       A�s  � � A�s  � �   a6q  *E     .       �u  A;q  \ Z FHq  ;E            AIq  �    KXq  @G AYq  � � Aeq    Aqq  6 4 A~q  [ Y A�q  � ~   e*f  E     �      ��w  .Ef  � � .Rf  > : f_f  Xflf  YL8f  L8f  Ayf  v t A�f  � � K�f  pG A�f  � � A�f  � � Hg  �G Tw  Ag  v p Ag  � � A g  2 * H-g  H w  A2g  � � A?g  � �  aig  } E     #       /w  Ajg  $    KKg  @H APg  ^ Z A]g  � �   H�f  pH �w  A�f  � � K�f  �H A�f    A�f  N H   F�f  � E     X       A�f  � � F�f  !E     ;       A�f  � � A�f   �     e�q  �!E     #      �z  .�q  \ P .�q  � � .�q  � x .�q    L�q  L�q  A�q  H 6 B�q  ��C�q  t#E     Hr  �H �x  Ar    Ar  s k  H%r  I Fy  A*r  � � _Fr  �"E       PI �	._r  &   ._r  &   .Sr  u s ?PI Akr  � � Awr  0 * A�r  � � A�r  � � A�r  P N 1>#E     �r  2Uu 2T|    H7r  �I {y  A8r  } s 1o#E     �r  2Uu 2T|  `�!E     j�  �y  2U| 2T82Q02R} 2X02Y�� `"E     j�  �y  2U| 2T02Q02Rw 2X02Y�� 1?"E     j�  2U| 2T 2Q02R}����2X02Y��  e:  `$E     �       ��|  .!:  � � ..:  � � g;:   K:  �I ..:  8 , .!:  � � ?�I A;:  E ? CH:  �$E     KQ:  0J AR:  � � @C  �$E      pJ ��{  ./C  � � ."C  � � .C  , * ?pJ B<C  �X-JC  �$E      �$E            i�{  .XC  W Q .XC  � � .eC      /�$E            ArC  ,  (  FC  �$E            A�C  g  c     1�$E     wI  2Us(2T| 2Q�X   4C  �$E      �$E     '       �L/C  ."C  �  �  .C  �  �  /�$E     '       B<C  �X-JC  �$E       �$E            i�|  .XC  ! ! .XC  R! N! .eC  �! �! /�$E            ArC  �! �! FC  �$E            A�C  �! �!    1�$E     wI  2Us� 2T| 2Q�X       eM  %E     t       �S}  .,M  V" P" .8M  �" �" L M  L M  ADM  )# ## APM  ~# r# B\M  �\1i%E     j�  2U�R2T12Rs ����2Y�\  e�:  �'E     �       ��}  .;  $ $ .;  �$ �$ .;  % % .(;  ?% 9% A5;  �% �% KB;  `K AC;  0& .& AP;  U& S& 1�'E     �<  2U} 2X0   e6Z  P)E     Q       �q~  .DZ  �& y& F6Z  X)E     H       .DZ  �& �& FQZ  X)E     H       ARZ  4' 2' h�)E     ��  2T�U    e�8  @,E     u       ��  .�8  c' W' .�8  �' �' A�8  o( m( K�8   M .�8  �( �( .�8  ) ) ? M A�8  �) �) K�8   M A�8  �) �) A�8  =* 1* @�;  Z,E      @M H�  .<  �* �* .�;  �* �* .�;  5+ 1+ -JC  Z,E      Z,E            �  .XC  }+ o+ .XC  5, ', .eC  �, �, /Z,E            ArC  - - FC  ^,E            A�C  C- ?-    1~,E     �C  2Us82T|   G�;  �,E      pM K.<  �- �- .�;  �- �- .�;  . . -JC  �,E       �,E            Ȁ  .XC  q. k. .XC  �. �. .eC  / / /�,E            ArC  F/ B/ FC  �,E            A�C  �/ ~/    h�,E     �C  2U�U#h      e}^  �,E     f      ��  .�^  �/ �/ .�^  J0 D0 .�^  �0 �0 f�^  Rf�^  XA�^  �0 �0 A�^  1 1 A�^  �1 �1 C�^  �-E     .�^  �1 �1 K�^  �M A�^  
2 2 A_  �2 �2 A_  �2 �2 A#_  s3 m3 A/_  �3 �3 A;_   4 �3 FG_   .E            AH_  v4 t4    e�`   9E           ��  .a  �4 �4 .a  6 6 .a  �6 �6 .)a  :7 7 B6a  ��}0Ca  APa  �8 �8 A]a  9 9 Cja  �9E     @ h  A9E      �Q 9Z�  .Yh  : : .Lh  �: �: .?h  A; 3; .2h  �; �; ?�Q Bfh  ��|Ash  �< �< C�h  h?E     H�h  0R _�  A�h  ]= U= A�h  �= �= A�h  > 	> A�h  ;> /> A�h  �> �> K�h  pR A�h  ? �> A�h  ~? v?   H�h  �R ̄  A�h  �? �? A�h  ]@ W@ Ai  �@ �@ Ai  (A  A Ki  �R Ai  �A �A A+i  bB TB A8i  ?C 7C AEi  �C �C ARi  D �C A_i  kD cD @j  S;E       S �"Z�  .8j  �D �D .,j  E E ? S ADj  CE ;E APj  �E �E A\j  �E �E   @j  �;E      PS �#��  .8j  ;F 1F .,j  �F �F ?PS ADj  /G #G APj  �G �G A\j  XH TH   5�<E     ��    @�i  (=E      �S �/�  .�i  �H �H .�i  I �H ?�S A�i  �I �I A�i  J �I Aj  iJ eJ   i�j  �S �e�  L�j  L�j  ?�S A�j  �J �J C�j  �=E     K�j   T A�j  $K  K A�j  jK ZK A�j  ,L L A�j  M �L A�j  WM KM Ak  �M �M Ak  qN iN Ak  �N �N A+k  �O �O A8k  IP CP AEk  �P �P ARk  �P �P `1>E     ��  :�  2U��{2T~ 2Q} 2R  1�>E     ��  2U} 2T��|2Q 2Rs     `�9E     j�  ��  2Us 2TH2Q02X02Y��| `:E     j�    2Us 2T@2Q02X02Y��| `2?E     �w  �  2U��~2Q��|# 2R��|#(2X��|I�q  ��|#I�q  ��|#8 1d?E     �w  2U��~2Q��|#P2R��|#X2X��|I�q  ��|#HI�q  ��|#h   -jj  �9E      �9E     T       ��  .xj  JQ HQ /�9E     T       A�j  rQ pQ `�9E     �s  ˇ  2U��~2Ts  `�9E     �s  �  2U��~2Ts  `�9E     ��  �  2Us  1�9E     ��  2Us    Ksa  `T Ata  �Q �Q A�a  S �R A�a  sT gT A�a  U �T A�a  �U �U A�a  �V �V A�a  PW JW A�a  �W �W A�a  @X ,X @at  �?E      �T P�  .|t   Y Y .rt  EY CY ?�T A�t  rY nY A�t  �Y �Y   i�d  U {��  L�d  L�d  L�d  ?U 0�d  A�d  �Y �Y 0�d  A�d  4Z *Z A�d  �Z �Z K�d  PU A�d  �Z �Z a
e  SLE     |       �  Ae  �Z �Z  Fe  �LE            Ae  /[ +[     -�i  q@E      q@E     �       m	 �  .�i  u[ e[ .�i  ;\ +\ /q@E     �       A�i  ] �\ A�i  �] �] Aj  7^ 3^   i{g  �U p	܊  L�g  ?�U A�g  }^ m^ C�g  PAE     C�g   AE     D�g  H�g  �U ��  A�g  -_ '_ A�g  �_ x_ A�g  �_ �_ A�g  ` `  K�g   V A�g  C` ;` Ah  �` �` Ah  a a    -ak  gAE       gAE     @       s	��  .ok  �a |a .ok  �a |a .�k  1b +b .�k  �b �b .|k  �b �b /gAE     @       A�k  �b �b A�k  `c \c 1�AE     �k  2UsP2T| 2Q��|�2R��}   @.e  �AE      pV y	��  .Ie  �c �c .<e  �c �c ?pV AVe  Jd Dd Ace  �d �d Ape  �d �d A}e  .e "e A�e  �e �e A�e  g g A�e  zg vg A�e  �g �g H�e  �V �  A�e  lh fh F�e  aBE     O       A�e  �h �h A�e  �h �h `�BE     �t  ��  2U I�p  v  1�BE     "v  2Uu 2Tt 2Qs 2R~ 2X��|�2Yy I8f      af  �CE     @       �  Af  i �h Af  *i &i  a�e  �JE     K       ��  A�e  di bi A�e  �i �i `�JE     �t  d�  2U  1�JE     "v  2Uu 2Tt 2Qs 2R~ 2X��|�2Yy I8f     1�AE     ��  2U    id  �V |	�  L5d  L(d  ?�V 0Bd  0Od  0\d  Aid  �i �i Kvd  0W Awd  	j �i K�d  �W A�d  �j yj @at  yDE      �W �n�  L|t  .rt  Qk Mk ?�W A�t  �k �k A�t  �k �k   -at   JE       JE            �,Ԏ  L|t  .rt  l l / JE            A�t  7l 3l A�t  zl vl   5KE     ��      @c  �DE      X }	�  .&c  �l �l .c  )m !m ?X A3c  �m �m A@c  $n n AMc  �n �n AZc  �n �n Bgc  ��|Atc  �o uo A�c  3p /p A�c  qp ip A�c  �p �p H�c  `X ��  A�c  �q �q  H�c  �X ��  A�c  �q �q A�c  _r ]r A�c  �r �r H�c  �X �  A�c  Zs Rs 5�ME     ��   @at  IJE      0Y LU�  L|t  .rt  �s �s ?0Y A�t  �s �s A�t  =t 9t   Gat  �KE      `Y \L|t  .rt  |t xt ?`Y A�t  �t �t A�t  �t �t    a�c  �KE     )       �  B�c  ��|1�KE     j�  2U 2T82Q02X02Yv   1�FE     ��  2U 2Tv    @�a  �FE      �Y ~	!�  .b  ?u 9u .�a  �u �u ?�Y Ab  �u �u A b  #v !v A-b  bv \v A:b  �v �v AGb  �v �v CTb  wGE     K]b  �Y A^b  %w w Akb  yw ow Axb  �w �w A�b  �x �x A�b  y y H�b  Z n�  A�b  ]y Uy A�b  �y �y A�b  iz cz A�b  �z �z A�b  5{ /{ A�b  �{ �{ A�b  %| !| A�b  c| [| @at  �HE      `Z �(��  L|t  .rt  �| �| ?`Z A�t  } } A�t  N} J}   @at   IE      �Z ��  L|t  .rt  �} �} ?�Z A�t  �} �} A�t  �} �}   -at  �HE      �HE            �Q�  L|t  .rt  4~ 0~ /�HE            A�t  s~ q~ A�t  �~ �~   1mHE     ��  2U��|2T~   @at  RIE      �Z �"��  L|t  .rt  �~ �~ ?�Z A�t  �~ �~ A�t  - )   4at  �IE      �IE            �L|t  .rt  j h /�IE            A�t  � � A�t  � �      -oi  �GE      �GE     �       �	��  .�i  � � .}i  N� L� /�GE     �       A�i  x� t� A�i  �� �� A�i  ր Ԁ A�i  �� ��   `�?E     ��  ϔ  2U��|2Tv 2Qs  `�?E     %R  �  2R02X0 1�JE     %R  2T��|2Q��|2R02X0   e�`  0NE            ���  .a  "� � .a  _� [� .a  �� �� .)a  ف Ձ 06a  0Ca  0Pa  0]a  jENE     �   ea:  PNE           �͘  .o:  � � .|:  �� �� .�:  1� %� g�:   Ka:  [ .�:   �� .|:  � � .o:  � � ?[ A�:  �� {� C�:  PE     K�:  P[ A�:  ؅ ʅ A�:  �� }� 0�:  B�:  ��@<  �NE       �[ ���  LZ<  .M<  �� �� .@<  � � .3<  ]� W� .&<  �� �� ?�[ Ag<  |� j� At<  @� <� B�<  ��C�<  APE     @�L  jOE       �[ �;�  .�L  �� ~� .�L  �� ~� .M  �� �� K�L  @\ L�L  L�L  .M  � �   @�L  �OE       �\ ���  .�L  � � .�L  � � .M  /� -� K�L  0] L�L  L�L  .M  T� R�   @�L  �OE       �] ��  .�L  y� w� .�L  y� w� .M  �� �� K�L   ^ L�L  L�L  .M  ŋ Ë   `�OE     wI  /�  2U	s ��"#82T} 2Q�� `�OE     �K  M�  2Tv 2Q}  `APE     �K  k�  2T~ 2Q}  1`PE     �K  2T| 2Q}    5�NE     ]�  5�NE     ]�  1�NE     �<  2U~ 2Q| @&2R} 2Xv      e9  `RE     �       �
�  .9  � � .9  o� g� .*9  ی ь 079  K9  �_ .*9  Z� P� .9  ׍ ύ .9  C� 9� ?�_ A79  �� �� CD9  �RE     KM9  0` AN9  �� � A[9  }� {� Ah9  �� �� Au9  ߏ ۏ `�RE     �?  ԙ  2Us2Tv 2Q02R| 2X02Y~  1�RE     �?  2Us� 2Tv 2Q| 2R} 2X02Y~      e�9  �RE     �       �]�  .�9  � � .�9  �� �� .�9  � � .�9  �� }� 0�9  K�9  p` .�9  � �� .�9  �� {� .�9  � � .�9  n� d� ?p` A�9  � � C�9  iSE     K�9  �` A�9  '� � A�9  �� �� A�9  Д ̔ A:  
� � `JSE     �?  '�  2Us2T} 2Q| 2Xv 2Y~  1eSE     �?  2Us� 2T} 2Q02R| 2Xv 2Y~      k�s  �s  7l�I  �I  �ln  n  l�s  �s  �k\P  \P  l�`  �`  vkQ  Q  ^k�l  �l  Rke  e  � S   !i  &  �� �:  �SE     S)      �x ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  s&  G   �  N   v  :-   �  L�  x NQ   y OQ   �  Q]  	�  ~   w�  
  yQ   �!  yQ  �   zQ  H  zQ   "  |�  �  (_  M} N    5�  N   `�  	G   _| 
_  
!  0  ?   e  2   e  B  U     e  �  �  �  	l  �  (Q�     S)   0�  T)  N5  V�  �   W�   H� X�  �1  ZG     �  )  �  \~  	�  �  �  N   �C  �!   �   pmoc�  stibu!  ltuo�  tolp :  �  �8  5"]  c  �$  �4  S�  x U)   len V0  e� We   �#  Yh  	�  �%  {�  �  �  G   G   �  U    �  �#  ��  �  G     G   G   U    �.  �  #  8  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(  �  (�/    0�  U   8*  �  @ y  �  u(  
8  	�  �2  (�  �  G     U      P  �3  ;  $  /  P   v)  ]<  B  W  P  _  @    �3  yd  j  G   �  P  @   U    H7  ��  �  G   �  P  �   �  51  0�  y2  �C   � ��   �/  *
 �W  / ��   $ �  ( 2$  ��  	  
�� &+   )  A"=  C  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  1  -    �   m�  �  �  1  U    f  ��  �  U   �  1  -   -   U    J   �"	    �  PH�  Ǟ  J_   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q  0ڰ  S1  8O�  T_  @��  U_  H �  ��  <v �-   ��  �U    �  ��  ""  ��  �  @     �  @   _  @    �       *  �   -4  	le  +  	�B  �  $8  	�e  	I  U    	��   	`  {"  	�)  !  	�0  \   	�G   �  	�N   }  	�-   )$  	�@   _]  	-   �   	-   c,  	+G   C*  	6U   +D  	C4    :   	�=	  xx 	��   xy 	��  yx 	��  yy 	��   5  	��  	=	  8  	�z	  ��  	�Z   ��  	��   $  	�O	  c   	��	  �	  �	  U    �  	��	  Kl  	�U    �  	��	   s  	��	  �"  	$�	  �	  �   	+)
  �� 	-�	   �W 	.�	  Kl  	/U    %  	DT
  uR 	F�	   �
 	G�	   }  	I)
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @
<#  5�  
>Q   ��  
?Q  �"  
AQ  �"  
BQ  i!  
CQ   %!  
EQ  (2!  
FQ  0�  
GQ  8   
I�  �"   
s�  ��  
uq   5�  
vq  ֳ  
xQ  !  
zQ  m  
{Q   v  
}0  J  
�#�  �  �!  �}c  ڰ  1   {3  ��  S0  ��  �/  ��  �1  ��  �1  ��!  Y/  �T
  �*  �	  (�)  �c  0+:  ��!  8<8  ��!  X�*  ��  � �3  
�"p  v  �(  ��  Oe ��!   �-  ��  ڰ  �1   U  
�"�  �  �  8	  ah !�!   Oe "|  U1  #T
   ;+  $�  0 i(  
�$    l;  ���  ah ��!   Oe ��!  y2  �C   {:  �  (�� �P  h/ ��  p�� ��  x T   
� �  �  _  �
a  �!  
�   �  
�  �  
�    
�  �  
�   �U 
�  (�  
�  03"  
�  8�  
�  @`  
!�  Hd  
"�  P�@  
$�	  X�;  
)�  h�   
+}  ��  
,q  �
  
-q  ���  
.q  �?!  
0q  ��  
1q  ��  
3q  ��  
4q  �ȩ  
6�  �ֳ  
7a  ��� 
8  �K 
<�  �ڰ  
=1  �^�  
>�  �U  
@T
  �t  
B�	  �k  
CU   ��L  
ED  � "  
 n  t  1  X
m�  ��  
o�   �@  
p�	  �e 
q�  �L  
r�  P @  
$%�  �    0
\  �-  
^�   ��  
_�  �W 
`�  x 
a�  �@  
b�	   �e 
d#  0�"  
e�  pi"  
f�  x� 
g�  ���  
iC  �.a 
kl  ��  
l�  �J  
m�  �Mj  
o�  ��  
q�  ��  
r�  �M  
tU    Z  
u-   _"  
wQ  (   
xQ  Ud 
zU    �L  
|"  ( �!  
F#%  +  Z!  
Ar  ��  
C�   T 
D7  �!  
E}  "  
F}   S  N   
�7  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  
r  0  
`)Q  W  �"  �e�  �1  g=	   H+  h�   x+  i�  0��  k�  8�)  n#{!  h�'  q6  p��  r7  t�*  y�  x `  �    �  
�)�  �  �!  H�4  $  �U    7:  ��  s4  ��   b  8
H�  !  
J}   m  
K}  A� 
M�  �� 
N�  �  
PQ  
  
QQ   ��  
RQ  (�  
SQ  0 �  
U4  x   
�$�  �  �!  0'"  ad  )�   �1  *}  &D  +�  2B  ,�  x� -=	     
�)/  5  �"  P��  ��  ��   �1  ��  �&  �*  �3  �=	  ]7  ��  0�7  �U   @�1  �7  H P6  
�  tag 
�   Kl  
�   �6  
	�  �  �5  N   

  i7   �&  9  F9  8%  �*   �,  

�  ./   
6
~  b 
8
   5�  
9
�  ��  
:
�  5  
;
�  Q(  
<
�    -  
I
(�  )  �8  N   
��  �:   4,  �6  $  �/  l9   �2  
��  �#  ��  �'  ��  �  �    c   �2  �       c   l/  �,  2  �  F  c  F   �   ;)  H��  �#  ��   :  ��  �5  ��  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  �  8��  �   @ l  �-  �L  d)  s�  �  �    U    9  F#  	  �$  @J�  �#  L�   y2  MC  W� O�  �� P
  �,  Q|   M4  R'  (�;  ST  0�*  T�  8 c/  X!�  �  �-  (q�  �-  s�   Oe t�  ��  uC  � v�     �/  )�  �  �  
  �  �   g%  .    '  �   �.  13  9  N  �  N  �   J	  73  6`  f  v  �  v   �  �8  :�  �  �  �  �  �   "3  >�  $)  Y�  �  �  �  	  �  �  �   �6  _�  �  �    	  �  N  �   �3  f     5  	  �  v   ;0  lA  G  �  `  	  �  �   �&  x��  ah � �   y2  � C  H�8  � �  P�8  � �  X�'  �   `� � 5  h�9  � �  p   �.  �`  	�  "9  H2/  Mj  4�   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :�  T%  �=�  ڰ  ?1   �0  @�  q5  A�  L)  B�  )  C*  Ǟ  E/  �  F/  `Ud HU   � X+  J�  ;  1  �  �  �  �  �  �  �  �  �   �&  &  
    �   �1  *!  '  �  6  a   �6  -B  H  S  a   w-  1_  e  �  t  �   �;  4�  �  �  �   =;  8�  �  �  �  a  ~   B$  <�  �  �  �  a  �   2  @�  �  �    �  a  �  7   7  G    �  =  �  �  �  �   q8  NI  O  �  c  �  �   )2  So  u  �  �  �  �  �  7  �   �  k.  ��|  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q ��  hZ)  �  p�#  �6  x'0  �S  �.  �t  ���  ��  �� �  �`9  �=  ���  �c  �5  ��  �U#  ��  � �2  ��  �  -   �&  0��  y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��  *  V'      �0  �*   u]   |#  w�   �#  x�  � y�  C4  z�   �&  |   �'  �u   {   �  �      �  �    z	  �9  ��   �   �      �    A2  ��   �   �  �      �  *  �    ]   8(  +!  ��  )i    $�  )�   �-  )�    )  �   	+!  3  <h!  �� >%h!   ��  ?%    8!  #  A=!  n!  �  �(  �v  �  c  �!  @    �  �!  @    �  �!  @    H'  �%  N   �$  ��  �� � �� � �� m� /� � `� 	/� 
w  �� w� m� W  �� � �� � R� ��  �  !�� "z #&� $� %� &�� '�� (�� 0�� 1� @P� A� Q�� R�� S�� TU� U� V6� W�� X�� `z� a�� b�  c�� p�� �T� ��� ��� �/ �p� �S� ��� ��� ��� �E� �p� �~� ��  ��� �M� ��� ��� ��� �.� �� ��� �Y� �� ��� �.� �K� �L ��� �=  �� �� ��� �@� ��� ��� ��� �A� ��� ��� �6� ��� �p� �  �1� �_� ��� �  Int 4G   �  5N   !  6)  !  70  �� 8-   �� 8"�  ,$  9@   �� ;e  �� ;"_  04  <�   � H�$  x JN$   y KN$   p� M�$  �  N   W�$  ��  �� L� �  � ^�$  �� a%  � @d�%  X f�   �� g�%  �  h[$  �1  iA$  ��  mN$   �k nN$  (�� p$  0�W s�%  8 � b�%  	%  6� w�%  �� x�%  �%  {� }�%  �Z 4$   G�  �4$   �� ��%  � �"&  �� ��F(  �� �$   �� �$  �� �$  �� �$  �� �$  � �$  � �[$  q� �[$   z� �[$  (top �[$  0�U ��  8� �$  <arc ��(  @C� �A$  H�� ��$  P�� �N$  X�� �N$  `�  �N$  h�� �N$  p9� �A$  x(� ��$  z�� ��$  {�� ��%  ��� ��%  �
� ��%  ���  ��$  �.  l  �Mj  �  �8� N$  �C� 4$  �<� 	�(   P� 
�(  
� �(  j �(  �� u$   �� �$  !4� �(  (�� �(  8�� $  x �� �2S(  &  � �f(  {(  F(  {(  {(   4$  j� ��(  �(  F(  4$  �  �  �%  �%    ��(  �(  F(   �$  Y(  �(  �(  �$  �(  @   ` �%  )  @    �� )  ڰ  U     !� !,)  )  J� �?)  E)  P)  �(   !%  �	`fG     
!+  �  "c)  �	�eG     #�� ^�  PzE     %      �b+  $�� ^(	  R� @� $�  _(�   � � $t `(�  �� �� $�t  a(�  @� ,� %�U c�  ��~&Mj  db+   � � &.a eh+  y� o� &ڰ  f1  �� �� &yW  gQ  I� 3� &�b  hQ  L� 8� %\  j�  ��~'�  ��{E     (�zE     �R  �*  )Us )T2)Q|  (&{E     �R  �*  )U~ )T��~)Q}  (O{E     �R  �*  )U )Q0)X0)Y��~ *�{E     +  )T��~ (|E     �R  '+  )U  (?|E     �R  ?+  )U  +p|E     �R  )U~ )T��~)Q}   �  l  ,�� QzE     ?       ��+  $�� Q&	  5� 1� $�  R&�  t� n� $�'  S&v  Ǜ Û -OzE     �R  )U�T#�)T�Q  .m� 6�  F,  /�� 6+	  /�  7+�  /�3  8+N  /�� 9+�  0�U ;�  '�  J�|E      #�� )�   dE            ��,  $�� )%	  �  � $y� *%�  V� R� $Kl  +%�  �� �� 12dE     )T�T)Q�Q  #�� �  �cE     !       �-  $�� !	  Ҝ ̜ 2
dE     )T0)Q0  3]� �G   �vE     :      �H.  4�� �-P  &� � 4\  �-�  �� �� 5Mj  �H.  �� � 5� ��  j� ^� 6�  �N.  ���~6_| �^.  ���~7 0  �wE       g �820  �� �� 9 g :?0  {� u� ;{Q  �wE       0g .  8�Q  ȟ ğ 8�Q  � 
�  (�xE     M0  ,.  )Uw )T0 +=yE     M0  )Uw )T1    �  �%  ^.  @     N$  o.  <@   � 3^� �G   �cE            ��.  =�� �!P  U=t �!h$  T=E�  �!U   Q >�� ��cE            �/  =�� �P  U=%� ��$  T=�  �h$  Q >3� �@dE            �l/  4�� �!)  J� D� 5ڰ  �1  �� �� -KdE     �R  )T�U  3�� �G   �yE     9       ��/  4ڰ  �!1  נ Ѡ 4�� �!�/  )� #� 6�U ��  �\5�� �)  y� u� +�yE     �R  )Uv )T8)Q�\  )  ?�� W 0  @�� W!)   A`e  �  M0  @�  F(  B�U �   3m� �G    iE     l      �:  4�  �F(  ̡ �� 4�� �&�$  � � Ci �4$  1� +� Dj �4$  XCk �4$  �� z� ;-B  �iE      �a �5  8LB  � � 8?B  Ȥ �� 9�a :YB  �� �� :dB  }� u� EqB  �b {4  :rB  ަ ڦ :B  � � ;�B  	jE      �b �f4  8�B  \� R� 8�B  
� � F�B  8�B  �� x� 9`c :�B  �� �� :�B  d� F� :�B  �� ث :�B  �� �� :C  � 
� :C  Ю ® : C  �� e� :-C  �� �� G:C  �mE     HCC  HLC  HUC  I^C  WjE            72  JcC   IqC  `jE            V2  JvC   I�C  kE     ;       �2  :�C  V� P� :�C  �� �� I�C  (kE            �2  J�C   +6kE     �H  )U~   E�C  �c }3  :�C  Բ Ĳ :D  �� |� :D  �� s� :D  ?� +� :+D  � � :7D  b� \� IVD  �kE            73  J[D   ECD   d J3  JHD   (�kE     zD  b3  )U~  +)vE     zD  )U~ )Yv   I�C  XlE            �3  J�C   E�C  Pd 4  J�C  :�C  �� �� :�C  A� 9� I�C  �lE            �3  J�C   (�lE     �F  �3  )U~  +mE     �F  )U~ )Xs   ( lE     �H  >4  )U~ )Tv )Q|  +1nE     �F  )U~ )Qs )Rv )X|    +�nE     �P  )Uu   7�O  �nE      �d 
8�O  �� �� 9�d :�O  }� m� :P  3� '� KP  �d :P  �� �� :P  � � (7oE     ,P  �4  )Uu  +HoE     ,P  )T}      7:  �oE      �d �8:  �� �� 9�d :+:  9� !� :6:  ;� 5� :C:  �� �� :P:  4� � :[:  +� � :f:  \� X� :s:  �� �� L�:  ��L�:  ��:�:  �� �� :�:  #� � :�:  �� � :�:  � �� :�:  a� ]� J�:  :�:  �� �� :�:  � � L�:  ��L
;  ��L;  ��G$;  �rE     G-;  �tE     G6;  isE     ;B  �oE     	  e �
s6  8B  �� ��  MB  �oE      �oE     	       �
�6  8B  �� ��  ;B  �oE      Pe �
�6  8B  � �  ;�A  XpE      �e �
47  8�A  :� 6� 8�A  v� p� 9�e :�A  �� �� :�A  d� \� :B  �� ��   ;|A  tE      �e 9�7  8�A  � � 8�A  A� ;� 9�e :�A  �� �� :�A  7� +�   ;|A  �qE      �e �
�7  8�A  �� �� 8�A  � 	� 9�e :�A  �� v� :�A  6� (�   ;�A  �qE      0f �
C8  8�A  �� �� 8�A  � � 90f :�A  g� [� :�A  �� �� :B  0� ,�   ;�A  @tE      `f �
�8  8�A  j� f� 8�A  �� �� 9`f :�A  � �� :�A  �� �� :B  �� ��   E?;  �f �8  :@;  � �  ;|A  �sE      �f 09  8�A  5� 1� 8�A  q� k� 9�f :�A  �� �� :�A  g� [�   *qE     99  )U~ )T��)Q�� (/rE     A  Q9  )Uu  (9rE     A  i9  )Uu  *�rE     �9  )U~ )T )Xs )Y}  *vsE     �9  )U~  (�tE     A  �9  )Uu  (�tE     A  �9  )Uu  *�tE     �9  )U~ )T )Xs )Y}  2EuE     )U~     A�  t
�$  O;  @�  t
F(  Ny v
4$  B�� v
4$  Bq�  v
 4$  NP x
�%  NQ x
�%  B� x
�%  Bb� x
!�%  B�� z
4$  B� z
4$  Ntop z
!4$  Bv� z
&4$  B�� z
.4$  Nx1 |
N$  Nx2 |
N$  Nxs |
N$  Ne1 |
N$  Ne2 |
#N$  B�� ~
�%  B�� 
�%  B� 
�%  O`� 	O�� GOA� PB�� �
$    >�� f
�cE            �~;  =�  f
F(  U > � �	�aE     �      ��<  =�  �	F(  UQy �	/4$  �� �� Qx1 �	/�  _� Q� Qx2 �	/�  � �� 4�  �	/�%  �� �� 4c� �	/�%  }� m� Ce1 �	N$  A� 1� Ce2 �	N$  �� �� Cpxl �	N$  n� b� 5c� �	�$  �� �� Cf1 �	u$  {� y� R�  `
=bE     SPbE     l      5�� 
$  �� ��   >�� �	`aE     p       ��=  =�  �	F(  UQy �	/4$  �� �� Qx1 �	/�  �� �� Qx2 �	/�  0� (� 4�  �	/�%  �� �� 4c� �	/�%  �� �� 9�a Ce1 �	N$  � � Ce2 �	N$  }� u� S�aE     *       Nf1 �	u$  5c� �	�$  �� ��    >C� �	PaE            ��=  =�  �	F(  UTmin �	+{(  TTmax �	+{(  Q >�� �	@aE            �!>  =�  �	F(  U >/� 	�_E     �      �L?  =�  	F(  UQy 	-4$   � � Qx1 	-�  �� �� Qx2 	-�  �� �� 4�  	-�%  <� ,� =c� 		-�%  YCe1 	N$  � �� Ce2 	N$  �� �� Cpxl 	N$  �� �� Cc1 	4$  Q� E� Cf1 	4$  �� �� R�  �	�_E     S�_E     O      5�� 1	$  P� B�   >�� �p^E     	      ��@  4�  �F(  6� 0� Qy �-4$  �� �� Qx1 �-�  �� �� Qx2 �-�   � �� 4�  �-�%  =� 9� 4c� �-�%  z� v� Ce1 �N$  �� �� Ce2 �N$  z� v� 5.  ��@  �� �� 5�� �
$  � �� S�^E     �       Cc1 �$  t� r� Cc2 �$  �� �� Cf1 �u$  � �� Cf2 �u$  9� 7�   u$  >L� �@^E     %       �A  =�  �F(  UTmin �){(  TQmax �){(  `� \� 5`�  �N$  �� ��  >�� j�]E     �       �|A  4�q  j�%  �� �� Cold l�%  � � 5�  l�%  � y� 5�W l�%  �� ��  ?�� G�A  @�q  G�%  @@  H�%  Nold J�%  B�  J�%   ?�� (B  @�q  (�%  @@  )�%  Nold +�%  B�  +�%  Nx ,N$   ?a� 'B  Ul 'B   �%  A�� ��$  �B  @�  �F(  @�� � $  Ni �$  B�k �'$  PB�� ��%  No ��$    As� ��$  zD  @�  �F(  @��  �%A$  @��  �%A$  @�� �%$  Bw  ��  BnX  ��  BJ  ��  BN5  ��  Bc ��  B��  ��  B�   ��   Ntag �'$  OM�  �OWD  �O?j  MO�l  �VqC  BuL   N$   V�C  BuL  N$   V�C  Nx 9N$  Ny 9N$  PBuL  ?N$    V�C  BuL  KN$   V�C  B�R  P�  Nx QN$  Ny QN$  PBuL  \N$    PNx1 }N$  Ny1 }N$  Nx2 }N$  Ny2 }N$  Nx3 }!N$  Ny3 }%N$  VVD  BuL  �N$   ViD  BuL  �N$   PBuL  �N$     3�� V�$  p[E           ��F  4�  VF(  � � Qcx1 VN$  �� �� Qcy1 WN$  �� �� Qcx2 XN$  /� +� Qcy2 YN$  l� h� Qx ZN$  �� �� Ty [N$  � Cy1 ]N$  �� �� Cy2 ]N$  b� Z� Cy3 ]N$  �� �� Cy4 ]N$  R� J� Cx4 ]N$  �� �� 5� ]"N$  8� 2� 5� ])N$  �� �� 5�� ]0N$  �� �� 5"� ]7N$  %� � 5�� ^�$  r� n� OWD  �W�a XF  Co ��$  �� �� (_\E     �P  7F  )Uu )Ty  +u\E     *Q  )Uu )Tt )Qq   (�\E     TJ  �F  )Us )T3)Q	`VE      X�\E     O  +j]E     DK  )Us )T3)Q	`VE       3J� ��$  �YE     �      ��H  4�  �F(  �� �� Qcx �N$  �� �� Qcy �N$  �� �� Qx �N$  � � Qy �N$  N� J� Cy1 �N$  �� �� Cy2 �N$  � �� Cy3 �N$  � w� Cx3 �N$  �� �� 5�� �N$  e� _� 5� �$N$  �� �� 5�� ��$  � � OWD  /WPa /H  Co �$  [� W� (eZE     �P  H  )Uu )Ty  +{ZE     *Q  )Uu )Tt )Qq   (�ZE     TJ  YH  )Us )T2)Q	�UE      X�ZE     �O  +J[E     DK  )Us )T2)Q	�UE       3�  q�$   gE           �TJ  4�  qF(  �� �� Qx qN$  =� %� Qy rN$  N� 8� M�L  8gE      8gE     H       ��I  8�L  :� 6� 8�L  y� u� 8�L  �� �� 8�L  �� �� 8�L   � �� 8�L  )� %� 8�L  e� a� S8gE     H       :�L  �� �� :�L  �� �� +hgE     M  )Us )R| )Xv    (�gE     �P  �I  )Us  (hE     *Q  �I  )Uu )Tt )Qq  (IhE     M  J  )Us )R| )Xv  (�hE     �P  3J  )Us  +�hE     *Q  )Uu )Tt )Qq   3�� @�$   YE     [       �DK  4�  @F(  �� �� 4N  @$$  ;� 7� 4�� A$2)  x� t� 4G B$N$  �� �� 4Y� C$N$  !� � Carc E�(  r� p� 5�Y  F�$  �� �� 5(� F�$  �� �� +\YE     DK  )Uv )R�X)X�R  Y�� ��$  WE           ��L  4�  �F(  �� �� 4N  �"$  w� s� 4�� �"2)  �� �� 4G �"N$  P� D� 4Y� �"N$  �� �� Cy1 �N$  L� B� Cy2 �N$  �� �� Ce �N$  �� x� Ce2 �N$  �� �� Ce0 �N$  J� @� Nf1 �4$  Carc ��(  �� �� B�� ��(  Ctop �[$  �� �� ZFin FXE      A�� ��$  M  @�  �F(  Ux1 �N$  Uy1 �N$  Ux2 �N$  Uy2 �N$  @G �N$  @Y� �N$  B�Y  ��$  B(� ��$   3�� ��$  PdE     �      �O  4�  �F(  �� �� Qx1 �N$  U� E� Qy1 �N$  � �� Qx2 �N$  �� �� Qy2 �N$  w  k  4G �N$  	 �  =Y� �N$  � CDx �N$  � ~ CDy �N$  � � Ce1 �$  '  Ce2 �$  � � Cf1 �$  , & Cf2 �$  | v 5ֳ  �$  � � CIx �N$  a Y CRx �N$  � � CAx �N$  � � Ctop �[$  d ` (eE     �R  �N  )U��)Q  (�eE     �R  �N  )T��)Q  (pfE     �R   O  )U��)T} s )Q  +�fE     �R  )T��)Q   >	� �`VE     �       ��O  =Ǟ  ��(  UCa �N$  � � Cb �N$  S K Cc �N$  � �  >�� ��UE     d       ��O  =Ǟ  ��(  UCa �N$  � � Cb �N$  >	 .	  A)� L�$  ,P  @�  LF(  Nn NA$  Np O�%  PBv� Y$  Ntop Y$    3�� �$  UE     �       ��P  =�  F(  UQy  $  
 
 5k� [$  �
 ~
 Cn $  �
 �
 9 a Cy2 )$  � �   3'� ��$  pTE     �       �*Q  =�  �F(  U4�� ��$  � � Ch �N$  "  9�` 5�� ��%  � �   3� ��$  �SE     �       �{Q  =�  �F(  U=�� �"�$  T=�� �"�$  Q ?*  E�Q  @�  EF(  @
� E%$   [�+  �|E     S       ��R  8�+  � � 8,  � � 8,  N J 8,  � � \),   I�+  �|E            �R  8�+  � � 8,    8,  + ) 8,  P N S�|E            :),  u s G5,  �|E     +�|E     �R  )Us�   +�|E     	S  )Us�)T�Q  ]�_  �_  �]�a  �a  ^�I  �I  �^�s  �s  �^@  @  �^�`  �`  v]e  e  
�]-R  -R  ]CA  CA  E �A   �n  &  � �:  �|E     #      �� �  �  �  v  :N   ,  �  Ly   x NB    y OB    �  QU   y   ~   w�   
  yB    �!  yB   �   zB   H  zB    "  |�   N`  -   �!  	�T   	jt  	�C  	�H  	�H  	�K  	RR  	Zs  	WO   
�  (�  M} -    5�  -   `�  	�  _| 
�  
!  �  ?   �  2   �  B  �    int �  �  �  �  !  �  
�  (Q2     S2   0�  T2  N5  V9  �   W?  H� XQ  �1  Z�    ;  y   E  �  E  2  �  \�  W  �P  �v  |  �  �  �  �   �   m\  v  �N  4�  �  �  �  �  �  �   �s  X�  �  �     �  �  �  �   
K[  0�c   �i   - ��  �
 ��  Q ��  m�  ��   �� �B   ( �l  �   c  �  -   ��  	�!   �   pmoc�  stibu!  ltuo�  tolp :  �u  �8  5"�  �  �$  
�4  S  x U2   len V�  e� W�   �#  Y�    �%  {.  4  N  �  �  N  �     �#  �a  g  �  �  �  �  �   �.  ��  �  �  �  �  �   
�8  `�5  .   5   �; ;  �1  �  �5  !  �+  !   `(  T  (�/  �  0�  �  8*  �   @ �  A  u(  
�  B  �2  (a  g  �  {  �  {   �  �3  ;�  �  �  �   v)  ]�  �  �  �  �  ;    �3  y�  �  �  �  �  ;   �   H7  �     �    �     O  
51  0��  y2  ��   � �T   ��  *
 ��  / ��   $ ��  ( 2$  �   �  | /+�  (\  �N   i   �;   �   @<  �  ?   p   	�  �  #	�  X  &	�  �  )	�   �  ,	�  (�  -	�  0/  2�  8�  5�  < �  8"�  +  KT  <  %  LT  �  MT  '  �M  �  N   �  ;    s&  �  �  -   )  	A"�  �  �   	�  �  	��   ��  	�  <h 	�)  �I  	�K   �  	X    �  )  �  N    �   	m5  ;  K  �  �   f  	�W  ]  �  {  �  N   N   �   J   	�"�  �  
�  P	H(	  Ǟ  	J�   ֳ  	K;   pos 	L;     	NN	  /[  	ON	   �K 	PZ	  (�R 	Q�	  0ڰ  	S�  8O�  	T�  @��  	U�  H �  	�N	  <v 	�N   ��  	��   �  	�(	  ""  	�f	  l	  ;   �	  {  ;   �  ;    �   	�	  �	  �	  {   -4  
l�  +  
��	  �  $8  
��  �	  �	    
�E  �	  {"  
�2  !  
��  \   
��  �  
�-   }  
�N   )$  
�;   �   
N   c,  
+�  C*  
6�  +D  
C�  �]  
P�  
 :   
��
  xx 
�7
   xy 
�7
  yx 
�7
  yy 
�7
   5  
�x
  �
  
8  
��
  ��  
��	   ��  
�
   $  
��
  c   
�    #  �   
�  
�N  Kl  
��   �  
�   s  
�#  �"  
$h  n  
�   
+�  �� 
-[   �W 
.[  Kl  
/�   
%  
D�  uR 
F[   �
 
G[   }  
I�  -   �"  	10   	�(  	Q;  	�4  	�(  	�0  	*  	/  	d2  	�+  		a0  
	~5  	�0  	k*  	�,  	U5  	l1  	�.  	�)  	�/  	l,  	a-   	.  !	�5  "	-5  #	�%  $	�*  %	�-  &	_:  '	N*  (	�8  0	a#  1	(  @	�$  A	I,  Q	.  R	6  S	^6  T	�9  U	L3  V	�(  W	�:  X	�7  `	Z'  a	�,  b	�7  c	�%  p	U.  �	I8  �	�,  �	�5  �	+  �	r'  �	�9  �	U$  �	-  �	�4  �	�4  �	�1  �	i$  �	@-  �	#(  �	�0  �	/7  �	�+  �	�+  �	E:  �	x0  �	+'  �	'  �	�'  �	�)  �	�%  �	,  �	
8  �	9.  �	0  �	|;  �	�:  �	54  �	�5  �	+-  �	�2  �	�-  �	�2  �	+6  �	�3  �	�9  �	�6  �	�%  �	39  �	�$  �	8#  �	�:  � 
�  @<�  5�  >B    ��  ?B   �"  AB   �"  BB   i!  CB    %!  EB   (2!  FB   0�  GB   8   I"  
�"   s  ��  u�	   5�  v�	  ֳ  xB   !  zB   m  {B    v  }�  J  �#  #  �!  �}�  ڰ  �   {3  �
  S0  �
  �/  �
  �1  �
  �1  �#  Y/  ��  �*  ��  (�)  ��  0+:  �(#  8<8  �8#  X�*  �
  � �3  �"�  �  
�(  �-  Oe ��"   �-  �  ڰ  ��   U  �":  @  
�  8�  ah !#   Oe " !  U1  #�   ;+  $5  0 i(  �$�  �  
l;  ��  ah �#   Oe �#  y2  ��   {:  ��  (�� ��  h/ ��  p�� �2  x T   �     
_  ��  �!  
   �  
  �  
    
  �  
   �U T  (�  T  03"  
  8�  Z  @`  !
  Hd  "`  P�@  $N  X�;  )�   h�   +�	  ��  ,�	  �
  -�	  ���  .�	  �?!  0�	  ��  1�	  ��  3�	  ��  4�	  �ȩ  69  �ֳ  7�  ��� 8�  �K <-  �ڰ  =�  �^�  >{  �U  @�  �t  BN  �k  C�  ��L  E�  � "   �  �  
1  Xm9  ��  o   �@  pN  �e q1  �L  rf  P @  $%F  L    0\�  �-  ^   ��  _  �W `9  x a
  �@  bN   �e d�  0�"  e7
  pi"  f7
  x� gy   ���  i�  �.a k�  ��  l
  �J  m
  �Mj  oW  ��  q
  ��  r>  �M  t�   Z  uN   _"  wB   (   xB   Ud z�   �L  |�  ( �!  F#�  �  
Z!  A�  ��  C   T D�  �!  E�	  "  F�	   S  -   ��  	Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  0  `)�  �  
�"  �eT  �1  g�
   H+  hy    x+  i
  0��  ku!  8�)  n#�"  h�'  q�	  p��  r�  t�*  y
  x �	    �  �  �)s  y  
�!  H��  $  ��   7:  �G  s4  �1   
b  8H1  !  J�	   m  K�	  A� M7
  �� N7
  �  PB   
  QB    ��  RB   (�  SB   0 �  U�  x   �$K  Q  �!  0'�  ad  )
   �1  *�	  &D  +
  2B  ,
  x� -�
     �)�  �  
�"  P�$  ��  �5   �1  �
  �&  ��	  �3  ��
  ]7  �y   0�7  ��  @�1  ��  H 
P6  O  tag +
   Kl  Q
   �6  	$  O  �5  -   
�  	i7   	�&  	9  	F9  	8%  	�*   �,  
b  
./   6
�  b 8
�   5�  9

  ��  :

  5  ;

  Q(  <

    -  I
(	  �  �8  -   �G  	�:   	4,  	�6  	$  	�/  	l9   �2  �  �	  �#  �Q
  �'  �r  x  D
  �  �   �2  ��  �  �  �   l/  ��  �  Z  �  �  �   L  ;)  H�S  �#  �+
   :  �
  �5  �S  F1  �7
  ,8  �7
   2*  �;  (�*  �f  0`1  ��  8��  ��  @ �	  �-  ��  d)  sr  x  D
  �  �   9  F#�  �  �$  @J  �#  L
   y2  M�  W� Oh  �� P�  �,  Q    M4  R�  (�;  S�  0�*  T&  8 c/  X!     �-  (qb  �-  s   Oe tb  ��  u�  � vy    �  �/  )t  z  D
  �    9   g%  .�  �  �     �.  1�  �  �    �  �   �
  73  6�  �  �    �   �   �8  :    D
  &       "3  >t  $)  Y>  D  D
  b  �  9  G  �   �6  _n  t  D
  �  �  9  �  �   �3  f�  �  �  �  9  �   ;0  l�  �  D
  �  �  +
  Q
   �&  x�M  ah � Y   y2  � �  H�8  � 2  P�8  � b  X�'  � �  `� � �  h�9  � M  p �  �.  ��  S  "9  H2�  Mj  4W   H5  59  (�)  69  0�  7
  8�  8>  @ �0  :d  T%  �=5  ڰ  ?�   �0  @
  q5  A
  L)  B
  )  C�	  Ǟ  E�  �  F�  `Ud H�  � X+  JA  �  1  S  Y  D
  |  {    
  
  \   �&  &�  �  �     �1  *�  �  D
  �  �   �6  -�  �  �  �   w-  1�  �  D
  �  9   �;  4  
    9   =;  8!  '  D
  ;  �  �   B$  <G  M  D
  a  �  +
   2  @m  s  D
  �  9  �  
  �   7  G�  �  D
  �    
  
  9   q8  N�  �  D
  �    {   )2  S�  �  D
       
  
  �      7
  k.  �� !  ah �Y   #,  �
  H�4  �
  P,;  �
  XEY �G  `/q �|  hZ)  ��  p�#  ��  x'0  ��  �.  ��  ���  �a  �� ��  �`9  ��  ���  ��  �5  �  �U#  �;  � �2  �!  "   
�&  0�u!  y%  �Q
   �/  �Q
  �'  �Q
  �6  �Q
  �+  �Q
   �6  �Q
  ( �7  �!  *  V'�!  �!  �0  �*   u�!  |#  w
   �#  x
  � y
  C4  z
   �&  |�!  �'  ��!  �!  D
  "  �!  
  "   �
  �9  �$"  *"  :"  �!  "   A2  �F"  L"  D
  j"  �!  
  �	  j"   �!  
8(  �"  ��  )�!   $�  )"  �-  ):"   )  p"  �"  
3  <�"  �� >%�"   ��  ?%�!   �"  #  A�"  �"  Y  �(  ��  S  �  (#  ;    e  8#  ;    y   H#  ;     H'  �%�  -   ��%  	�  	� 	g 	� 	+ 	 	� 	� 	� 	J 		� 
	� 	� 	�
 	� 	� 	
 	 	_ 	S 	� 	]  	�	 !	� "	� #	0 $	 %	1	 &	e '	� (	^ 0	P 1	� @	� A	> Q	f R	� S	4 T	r U	� V	� W	�	 X	 `	" a	� b	< c	� p	� �	� �	� �	� �	� �	:
 �	z �	Z �	F �	]	 �	_ �	� �	� �	� �	z	 �	� �	� �	 �	� �	2 �	� �	d �	�
 �	� �	4 �	�	 �	) �	" �	T
 �	� �	t
 �	y �	�
 �	� �	 �	e �	 �	� �	/ �	� �	 �	� �	�
 �	O �	F �	� �	� � � �N    ��  �%  Y ��   ��%  �%  
X �&  x ��%    ��%  �r  ��%  �W ��%   � ��%  
w �T&  �t  ��   `�  ��   � �)&  �  ��'  �Y  �y   ex ��%  @ey ��%  D� ��%  H� ��%  L
 ��%  P� ��%  T�r  ��%  X ��%  \m  ��  `� ��'  h
 ��%  pS	 �k
  x
 �k
  �x ��%  �y ��%  �Mj  �W  �.  �T&  � �!  �1 ��  ��+  ��'  �� ��   �%    �'  ;   	 � �a&  � ��'  a&  
�
 ��'  ڰ  ��    | � (  �'  !ei  Up  	�hG     "�  �	`hG     �$  _  �#   _  �.  "_  #0(  �	�gG     #<(  �	`gG     #H(  �	�fG     $� �D
  ��E            �1)  %�� �-�  � � %�  �-9  � � %t �-G    %�t  �-�  T P &��E     �*  'U�U'T�T'Q�Q'R�R'X4  $	 �D
  ��E            ��)  %�� �+�  � � %�  �+9  � � %t �+G    %�t  �+�  H D &��E     �*  'U�U'T�T'Q�Q'R�R'X3  $� �D
  ��E            ��*  %�� �'�  � � %�  �'9  � � %t �'G   � %�t  �'�  a ] &��E     �*  'U�U'T�T'Q�Q0�Q $@L$.( 'R�R'X0  (@ qD
  �E     j      ��.  )�� q/�  � � )�  r/9  � � )t s/G  � � )�t  t/�   � )k u/G  � � *�U wD
  ��~+Mj  x�.  � � +.a y/  � � +ڰ  z�  � � +yW  {B   ` L +�b  |B   J 4 +� }
  M 1 +/ ~
  1  *\  �B  ��~,�  l\�E     -�h h-  +� �T  � � +�S  �T  (  .i �
  � � .j �
      /��  -   D  <  /5�  -   �  �  /`�  �  ,! &! 0sub 9  }! y! 1O�E     CA  �,  'U~  2[�E     �,  'T��~ 1��E     CA  �,  'U~  2ƍE     �,  'T��~ 12�E     CA  �,  'U~  2>�E     -  'T��~ 1H�E     PA  +-  'U��~'T��~'Q��~ 1(�E     \A  K-  'Tv 'Q��~ 3g�E     gA  'U��}'Tv   4x�E     �      +.  /`�  =�  �! �! 0sub ?9  �! �! 1ЎE     CA  �-  'U~  2܎E     �-  'T��~ 11�E     CA  �-  'U~  2=�E     .  'T��~ 1��E     CA  .  'U~  5��E     'T��~  6��E     gA  1�E     CA  ^.  'U~ 'T| 'Q}  1#�E     sA  �.  'Us 'T 'Q��} 1��E     �A  �.  'U��}'Q0'X0'Y��~ 2N�E     �.  'T��~ 1��E     gA  �.  'U��} 3،E     CA  'U~ 'T| 'Q}   W  �  7 dЉE     ?       ��/  )�� d%�  !" " )�  e%9  `" Z" )�'  f%�  �" �" &�E     �A  'U�T#�'T�Q  8z ID
  �/  9�� I*�  9�  J*9  9�3  K*�  9�� L*�  :�U ND
  ;�  ]ߖE      (� =D
  p}E            �Z0  )�� =$�  �" �" )y� >$+
  B# ># )Kl  ?$Q
  # {# <�}E     'T�T'Q�Q  (\ D
   }E     g       ��0  )��  �  �# �# .sub $9  $ 
$ 5`}E     'T0'Q0  $%
 }�  �|E            �
1  =�� }(�  U=t ~(;   T=E�  (�  Q > r�|E            �W1  =�� r&�  U=%� s&�  T=�  t&;   Q > f�}E            ��1  %�� f �  q$ k$ /ڰ  h�  �$ �$ &�}E     gA  'T�U  $� S�  ��E     9       �H2  %ڰ  S �  �$ �$ %�� T {  P% J% !�U VD
  �\/�� W�'  �% �% 3��E     PA  'Uv 'T8'Q�\  $* ��  ��E     �      ��2  %�� �0�  �% �% %\  �0  �& �& /Mj  ��2  ' ' /� �5  �' �' !�  ��2  ��}3��E     �2  'Uw   d  �'  �2  ;     $� ��  �E     �      �J5  %�  ��'  P( F( /�!  ��%  �( �( /H  ��%  �( �( !_| �J5  ���~/��  ��  k) i) 0n ��  �) �) 0y ��%  1* )* ! �[5  ���~/N �k5  �* �* /< �
�  �* �* ?�g /5�  ��%  ~+ r+ /�U ��  , , @L6  ��E      h �5  AZ6  \, Z, ?h Bg6  �, , Cr6  Ph Bs6  �, �, B�6  �, �, B�6  5- /- B�6  �- - 1�E     �6  �4  'U~ 'Q| 'R  1*�E     �6  �4  'U~ 'Q| 'R  2I�E     �4  'U| 'Q}  3��E     �6  'U~ 'Q| 'X1    1`�E     �A  .5  'T0'Qw  3��E     q5  'U~ 'T    &  [5  D;   � �%  k5  ;    �%  $� c�  �E     �       �L6  %�  c�'  �- �- %< d"�  V. R. /�U f
�  �. �. 1�E     �A  �5  'Uw  6�E     �A  1�E     �A  )6  'Uw #�'T	�hG     'Qw  6�E     �A  3�E     �=  'Uw   E� �6  F�  �'  Gy 
�  HI/ �%  Gx �%  I �%  I�r  �%    >� ��}E     C      ��7  %�  ��'  / / Jx � �%  �/ �/ Jy � �%  o0 a0 %e� � �%  1 1 %u � �%  �1 �1 -`g g7  /& ��7  `2 \2 5-~E     'U�Q'T:'Qs�  Kh~E     {       0q ��  �2 �2 0c ��  �3 �3 &�~E     �A  'Q	�X $ &     $L ��  p�E     *       �h8  %� �$�  �3 �3 %� �$�  64 24 Jto �$�  s4 o4 %�  �$�'  �4 �4 3��E     v>  'U�RL:  �UL:  �TL:  �Q  $�
 ��  ��E     $       ��8  %��  �$�  5 �4 Jto �$�  ?5 ;5 %�  �$�'  ~5 x5 3��E     F?  'U�QL�:  �UL�:  �T  $m ��  �E     )       �S9  Jto �#�  �5 �5 %�  �#�'  6 6 32�E     _;  'U�T  $= ��  @�E     G       ��9  Jto �#�  ]6 Y6 %�  �#�'  �6 �6 0x ��%  7 �6 0y ��%  Y7 S7 3p�E     v=  'U| 'Tv 8&'Qs 8&  E MO:  F�  M�'  F� M1�  F� N1�  Mto O1�  IB QO:  Garc R9  Nt	 � y   _:  ;   0 ET -�:  FǞ  -!9  Ga /�%  Gb /�%  Gc /�%   E� �;  F�  ��'  F��  �1�  Mto �1�  IB �;  Garc �9  Gdx ��%  Gdy ��%  IS ��  IC ��   y   -;  ;     E� �_;  FǞ  �!9  Ga ��%  Gb ��%   >� QP�E     �      �v=  %�  Q�'  �7 �7 %� Q$�%  8 8 %� R$�%  ^8 L8 0dx T�%  09 "9 0dy T�%  �9 �9 0fx1 U�%  �: k: 0fy1 U�%  �; ~; 0fx2 U�%  = �< 0fy2 U�%  �= �= 0ex1 V�%  G> 3> 0ey1 V�%  =? ? 0ex2 V�%  �@ �@ 0ey2 V�%  �A qA OEnd �@�E     -�h =  / ��%  �B rB /X �N   C C / �N   WC SC 3ӆE     v=  'U~ 'T| 'Q}   1��E     v=  +=  'U~ 'Tv 'Q|  1ƈE     v=  U=  'U~ 'T���'Q��� 3��E     v=  'U~ 'Tv 'Q}   >�	 ;ЄE            ��=  %�  ;�'  �C �C Jex ;#�%  -D %D Jey <#�%  �D �D 6E�E     �=   ># �~E     �       �v>  %�  �'  �D �D / �'  :E 2E // �%  �E �E 0x �%  �E �E ,cs /`E     3yE     �A  'T1  P�9  ��E     �      �F?  A�9  @F 8F Q:  Q:  Q:  Q:  Q:  Q:  R+:  ��yB8:  �F �F SE:  ��E     @_:  ��E       i �%?  Am:  JG FG ? i Tz:  T�:  B�:  �G �G   3T�E     _;  'U} 'T| 'Qv   P�:  ��E     �      �B@  A�:  �G �G Q�:  Q�:  Q�:  Q�:  R�:  ��{B�:  7H #H B�:  I I B�:  tI rI B;  �I �I B;  kJ _J @-;  ÕE      0i !	@  A;;  K K ?0i BH;  *K &K BS;  hK `K   1)�E     _;  -@  'Uv  3S�E     _;  'Uv   P�/  ��E     S       �CA  A�/  �K �K A�/  L L A�/  WL SL A�/  �L �L U�/   V�/  �E            &A  A�/  �L �L A�/  M 
M A�/  4M 2M A�/  YM WM K�E            B�/  ~M |M S�/  ��E     3��E     CA  'Us�   3ߖE     �A  'Us�'T�Q  W�a  �a  X�`  �`  vYBY  8Y   X�s  �s  �W�_  �_  �X�I  �I  �X@  @  �YD  D   X�p �p 'X
 
 �X�c  �c  |Xo o �XD  D  0XbU  bU  #WCA  CA  E =;   �s  &  % �:  �E     �0      <� ,  i   	�@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  �  
N   )  A"P  V  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  D  -    �   m�  �  �  D  U    f  ��  �  U     D  -   -   U    J   �"  "  �  PH�  Ǟ  J   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q,  0ڰ  SD  8O�  T  @��  U  H �  ��  <v �-   ��  �U    �  ��  ""  ��    @       @     @    %  �  �   9  ?  J     v  :-   ~   w�  
  yJ   �!  yJ  �   zJ  H  zJ   "  |V  �  (#  M} N    5�  N   `�  	G   _| 
  
!  0  ?   %  2   %  B  U     �  �  	#  �  N   �s  �!   �   pmoc�  stibu!  ltuo�  tolp :  �5  �8  5"�  �  �$  �4  S�  x U)   len V0  e� W%   �#  Y�  	�  �%  {�  �    G   G     U    �  �#  �!  '  G   @  G   G   U    �.  �M  S  h  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(    (�/  @  0�  U   8*  �  @ 0    u(  
h  	  �2  (!  '  G   ;  U   ;   �  �3  ;N  T  _  �   v)  ]l  r  �  �    @    �3  y�  �  G   �  �  @   U    H7  ��  �  G   �  �  �     51  0�C  y2  �s   � �   �_  *
 ��  / ��   $ �A  ( 2$  ��  �  $8  �%  	W  c  !  �0  �  �N   }  �-   )$  �@   c,  +G   C*  6U   +D  C4   N   �
  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � W  �   H'  �%C  N   �d  m  H  � � � { | �   	� 
� � �    k � & � i    !� "< #� $� %� &* 'Z (� 0C 1F @� A� Q R  Sl Tm UH V W X] `� a� b4 c� p, �( �[ �c � �! �  �� �� �� �� �� �T �� �� �� �� �; �� �� �� �a �� �� �� �� �� �� �� �U �� �B � �t �| � �> �Q �� �H �� �� �8 �l  �� �D �2 � �� �%  g �N   	p  z �@    �d  	�  6 �p  	�  � ��  � �U   
�  ��  �   
9  ��   
�	  �G   
�  �G   
Z  �G   - ?    �  4  �  p  p   8 @@  F  V  �  �   � pD  � E   s Fp  H G�   I  � Jp   � K�  (msg M�   0��  N o  8� P	  @W Q4  H R�  P] TG   X� U�  `Y  V�  h �  � (o  t !   sub +2  � .G   �  /p  � 1`       ? WV  � Y�  u  
 G   
 �   
� �   � ��  �  �  �  �  �  p   �  e #�  	�  � !  ��  E   Ǟ  p   E  � d    d   g    !  pad 
p    )s  � p  t �   sub /[  ��  0p  (� 3p  ,� 4	�  0f  58  8y 6
  @end 7
  H�K 8
  P�  9
  X$ :�  `� ;	�  h 3  ()  � 0�  t !�   len $p  sub /F  � 2d  9 3d  g 48   r 58  ( N   �  3Y     �   � H DRY [ BAD 	 N �   $2  �B %p   ad  &p    '2  bb (p  tb )8   �  �  +U  = -U       "�  �  #
p  * *�  u .>    |  �  !@    	�  "� +�  	`G     ",  /�  	�~G      |  �  !@    	�  "/ 2�  	`~G     "� 6�  	�}G     #� 
|  	#� |   �  6  $@   � 	%  "� 6  	�mG      �  a  !@    	Q  " �a  	�lG      |  �  !@    	|  "� �  	�lG     N   �  o  LEN ` � � � LIT � END � 	 � �  &"  s '8   C (p   +F  get ,p   �  -p   %t  �* )�  lit *
p  �,  ."    |  �  !@    	t  "� �  	 lG     N     �  ^y  � � � � � 0 � � 	� 
# S �  � �  &2  was '�   C (�   $`  - %
p  � )  # *
p   g  %� � ��  �; �   ^�  �  ڰ  �D  * �u  �k ��  �� ��  �&_| ��  �'pos ��  � &O�  �
  � &��  �
  �   W    $@   � ! �  f  (=\ ��  ��E     �       �8  )ڰ  �'D  �M �M )� �'
  ,N "N )o �'8  �N �N )� �'h  �O �O )� �'�   P �O *^�  �u  ��~+err �G   tP bP ,A�E     7  �  -Uw -T/ ,R�E     1#    -Uw -T4 ,a�E     ?-  #  -Uw  .��E     ?-  -Uw   �  (w< k�  ��E           ��  )^�  k"  9Q /Q )�; l"  �Q �Q /�U n�  S S /ڰ  oD  BS >S +zip p  �S xS 0�  �X�E     1 q �  /� ��  ST IT 1�q 0  /� �
  �T �T 1�q   //� ��  \U TU 2.  *�E      �q ��  3<  �U �U 4�q 5I  �U �U .3�E     ?-  -U}   ,��E     �  �  -U} -T0-Qv -R  ,�E     �  �  -U} -T0-Q0-R0 ,�E     �:  �  -U| -Tv  .��E     �:  -U| -T}   .��E     �:  -U| -T -Q��  6�  �E      pq �3  <V 0V 4pq 7  ��5   �V �V 5-  XW LW ,�E     �:  �  -Uv  ,m�E     �:  �  -Uv -T�� ,��E     �:  �  -Uv -T~  8��E     �:     2W  [�E      �p ��  3�  �W �W 3v  4X ,X 3i  �X �X 4�p 5�   Y �X 5�  �Y �Y 9�  ��E     ,��E     �  g  -Uv  ,��E     �:    -Uv  .��E     7  -U}-T	�   ,�E     �  �  -Uv  ,L�E     �:  �  -U| -T
� -Q�� .��E     �:  -U| -T}   :� S�  ;  ;^�  S-  <�U U�  <� V�  <�Y  W�   =6 F@   ��E     	       ��  )^�  F&  Z Z )�  G&@   IZ EZ )_| H&  �Z �Z )/� I&@   �Z �Z +zip K   [ �Z >��E     �  -T�T-Q�Q-R�R  ?� 0��E     �       ��  )^�  0$  A[ 7[ +zip 2  �[ �[ /ڰ  3D  �[ �[ 2.  ��E      pi 9�  3<  -\ +\ 4pi 5I  V\ P\ .��E     ?-  -Us   ,��E     �:  �  -U| -Ts  .�E     �:  -U|   :Y ��  M  @zip �!  @pos �!�  ;_| �!
  ;/� �!�  <�Y  ��  <�U ��  0�  "V�E     A<�� �    :� ��  �  @zip �*  ;/� �*�  <�U ��  <�� ��   =� ��  `�E     �      ��  Bzip �*  �\ �\ /* ��  �] �] /�U ��  "^ ^ 4@o +err �G   �^ �^ 2�  ��E      �o ��  3�  �^ �^ 4�o 5�  U_ K_ 5�  �_ �_ 5�  W` G` C��E     -Uv -Q| -R
    .��E     1#  -U} -T0   :� x�  �  @zip x)  <* z�  <^�  {  <ֳ  |�   :� \�  .  @zip \$  <^�  ^  <�U _�  A<* d�    Dx EW  @zip E#  <* G�   :� �  �  @zip #  ;^�  #  ;�; #  <* �  <�U �  E�  ? F� ��  ��E     .      �v   G^�  �$  (a  a H�U ��  �a �a "uR �v   �\0�  �E     Io�E     =       z  Jlen �z  �a �a ,�E     �:  e  -Us -Tv  .��E     ;  -Us   I�E            �  Jc �z  �a �a .�E     ;  -Us -Tv   I@�E     "       �  +c z  b b .K�E     ;  -Us -Tv   ,��E     �:     -Us -T0 ,¡E     ;  ?   -Us -T�\-Q4 ,��E     ;  \   -Us -T6 .��E     ;  -Us -T2   W  �   !@    K? �@�E            �&!  G ��  cb _b Lptr ��  �b �b M"  @�E      @�E            �36"  �b �b 3*"  c c >E�E     �:  -U�U-T�T   F� ��  p�E            �"  G ��  Wc Sc G. �N   �c �c Gֳ  �N   �c �c NC"  p�E      �i �3l"  d 
d 3`"  Kd Gd 3T"  �d �d 4�i 5x"  �d �d 7�"  �l5�"  8e 4e .��E     �:  -U�U-T�Q�����T����-Q�l    O� �C"  Pڰ  �D  P�& ��   Q� }�  �"  Pڰ  }D  P. ~p  Pֳ  p  Rsz ��  S�U ��  Rp ��   F� �  @�E     2      �1#  G� �  se oe Lbuf �  �e �e Llen 
p  _f Qf Js1 @    g �f Js2 @   �h �h Jk 	G   Hj @j  T� �G   �E     b      �-  Lz ��  �j �j Lf �G   Lm Dm Jr �G   �m �m Jb �p  zo po U\.  ��E       0j ��,  3�.  �p p 3w.  �u �u 3m.  �v �v 40j 5�.  gw -w 5�.  z �y 5�.  �| =| 5�.  �� =� 5�.  ń �� 5�.  g� +� 5�.  ˈ �� 2�0   �E      �j WU&  3�0  � �� 3�0  k� g� 3�0  �� �� 4�j 5�0  �� ۍ 5�0  -� � 5�0  � Տ 5�0  s� K� 5�0  ;� �� 5�0  �� �� 5�0  � Ǘ 51  �� Q� 51  �� �� 51  � ѝ 5$1  � �� ,�E     �1  6%  -U| -Ts -Q	� ,��E     �1  X%  -U��~-T��~ ,��E     �1  z%  -U��~-T��~ ,8�E     �1  �%  -U| -Ts -Q1 ,s�E     �1  �%  -U| -Ts  ,g�E     �1  �%  -U| -Ts  ,ۺE     �1  �%  -U| -Ts -Q	� ,��E     �1  &  -U| -Ts  ,r�E     �1  9&  -U| -Ts  .��E     �1  -U| -Ts    Vo0  (�E      (�E            Z�&  3�0  Y� U� 3�0  Y� U� 3|0  �� ��  W/  0l �&  5/  á �� 5/  �� �� 5/  G� C� 5)/  �� ��  Ui3  ��E       �l ��'  3�3  � � 3�3  n� f� 3�3  ޤ Ф 3�3  �� �� 3{3  F� >� 4�l 5�3  �� �� 7�3  ��5�3  D� <� X��E     �'  -TC-Q4 ,�E     �3  �'  -U��~-TC-QC-R0-X0 X9�E     �'  -T��~ X2�E     �'  -T��~ C4�E     -T��~   W5/  �l r*  76/  ��7B/  ��7N/  ��7Z/  ��5f/  �� �� 2�2  �E      `m =�)  353  � � 3)3  8� 0� 33  �� �� 33  +� !� 33  �� �� 3�2  5� +� 3�2  �� �� 3�2  � � 3�2  k� i� 4`m 5@3  �� �� 7K3  ��5W3  ì �� ,�E     �3  >)  -U��~�����2$��"-T���#-Q0-R	`~G     -X	�}G     -Y�� X3�E     T)  -T��~ X,�E     n)  -T
 -Q4 ,s�E     �3  �)  -U��-T��~�-Q
-R	`G     -X	�~G     -Y�� X��E     �)  -T��~ C`�E     -T��~   6/1  d�E        n K3l1  '� %� 3l1  '� %� 3a1  L� J� 3V1  u� q� 3K1  �� �� 3@1  � � 4 n 5v1  '� %� Cl�E     -T1-Q0    W�.  �n �+  5�.  N� J� 5�.  �� �� 5�.  Ʈ ® 5�.  � � U/1  U�E      �n �#D+  3l1  ^� Z� 3l1  ^� Z� 3a1  �� �� 3V1  � � 3K1  0� ,� 3@1  l� h� 4�n 5v1  �� �� C]�E     -T1-Q0   Yj2  U�E      U�E             ��+  3�2  � ް 3�2  � � 3�2  D� B� 3�2  n� l� 3|2  �� ��  .5�E     �1  -Ts -Q	�  ,��E     �1  �+  -Ts -Q	� ,��E     �1  ,  -Ts -Q1 XɰE     +,  -T O 
�?5%O"#�-Q4 ,>�E     �1  I,  -U| -Ts  ,��E     +;  i,  -Tv -Q��~ ,��E     �1  �,  -Uw -Ts  ,�E     �1  �,  -Ts  ,k�E     �1  �,  -Ts -Q	� ,(�E     �1  �,  -Ts  .��E     �1  -Ts    .`�E     �/  -Ts   Q' RG   ?-  Zz S�  Zw TG   P��  U
  Py VG    T7 DG   ��E     ~       ��-  Lz E�  ȱ �� M3.  �E      �E     5       J3P.  +� '� 3E.  c� a� ,��E     �/  �-  -Uv -Ts -Q0 C�E     -Tv    F� 6G   `�E     R       �3.  Lz 7�  �� �� .��E     �/  -T�U-Q0  :� |G   \.  @s }`  @z ~�   Q� wG   s/  Zs x`  Zz y�  Zr zG   Rt |p  Rb }	�  Rk ~p  Rp 
  Rn �p  Rq �
  Rm �p  [/  Rbl �p  Rbd �p  Rtl �8  Rtd � 8   [5/  \h 8  \i p  \j p  \c p   A\bl 6p  \bd 6p  \tl 78  \td 78  \c 8U    Qm X`  �/  Zz Y�  Zc Z�  Zw [p  Rs ]`   ]` C��E     �       �i0  Ls D`  � � Lz E�  E� ?� Lc F	i0  �� �� Yo0  �E      �E            MO0  3�0  г γ 3�0  г γ 3|0  �� �  CQ�E     -U0-T0-Q0  �  O� ��0  Zc �U  Zz ��   Q5 PG   /1  Zs Q`  Zz R�  Zr SG   Rj Up  Rt V8  Re Wp  Rb X	�  Rk Yp  Rp Z
  Rn [p  Rq \
  Rm ]p  Rf ^
  Rc _U   Q� :U  �1  Zbl ;p  Zbd ;p  Ztl <8  Ztd =8  Zz >�  Rc @U   F� G   ��E     A      �j2  Ls `  !� � Lz �  �� �� Lr G   � �� Jn p  � u� Jp 
  �� � Jq 
  N� >� X �E     )2  -T -Q~  ,9�E     +;  G2  -T -Q~  X��E     \2  -Tw  8�E     +;   :� �G   �2  @bl �2  @bd �2  @tl ��2  @td ��2  @z ��   �2  �  :i GG   c3  @nl Hp  @nd Ip  @c J2  @bl K2  @bd L2  @tl Mc3  @td Nc3  @hp O8  @z P�  \r SG   \hn Tp  \v U
2   8  :B +G   �3  @c ,2  @bb -2  @tb .c3  @hp /8  @z 0�  \r 3G   \hn 4p  \v 5
2   F� _G   �E     �      ��5  Lb `2  � �� Ln ap  �� z� Ls bp  !� � Ld c�5  ]� Y� Le d�5  �� �� Lt ec3  ո Ѹ ^m f2  � ^hp g8  �^hn h�5  �Lv i2  � � Ja qp  k� _� _c r�5  ��}Jf sp  � 	� Jg tG   � غ Jh uG   �� m� Ji vp  u� S� Jj wp  �� Խ Jk xG   �� �� Jl yG   (� � H�� zp  �� �� Jp {
2  J� � Jq |8  f� \� Jr }�  �� �� _u ~6  ��~Jw G   � �� _x ��5  ��~Jxp �
2  �� �� Jy �G   � �� Jz �p  .� �  �  p   p  6  !@     8  6  !@    `"  0�E            �m6  3*"  U� Q� 36"  �� �� >5�E     �:  -U�U-T�T  `C"  P�E            �7  3T"  �� �� 3`"  � � 3l"  I� E� 5x"  �� �� 7�"  �l5�"  �� �� .f�E     �:  -U�U-T�Q�����T����-Q�l  a-  �E     �      ��8  3-  <� 0� 3-  �� �� b2-  pc&-  �7  Us/  ��E       �i }38  3�/  j� d� 3�/  �� �� 3�/  � � 4�i 5�/  Y� Q� X��E     �7  -T1-Qp XݤE     �7  -T8-Q
� X��E     �7  -T1-Q}  ,%�E     �/  8  -Uv -Ts -Q0 X��E     !8  -Tv  C��E     -Tv    XV�E     L8  -T1-Q( ,2�E     �-  d8  -Us  ,��E     ?-  |8  -Us  .ȥE     ?-  -Us   `�   �E     �      ��:  3�  �� �� 3�  �� v� 3�  Z� L� 3  � �� d   d   W�  0p �9  e�  3  �� �� e�  e�  40p 5  � � 5  �� �� f,  g=  pp 5>  �� �� ,d�E     +;  m9  -U} -Q|  ,��E     +;  �9  -Qv  .��E     �  -Us     2�  ��E      �p �-:  3�  	� � 4�p 5  A� ?� 5  i� e� h  `�E     O       :  5  �� �� .i�E     �-  -Us  8��E     �:    iM  ��E       ��E     m       3l  �� �� 3_  s� q� j��E     m       5y  �� �� 5�  �� �� .R�E     �  -Us     k�s  �s  �k�`  �`  vlM  M  �l�f  �f  �l�Z  �Z  �k�U  �U  {l�G  �G  �lw  w  �l�k  �k  �l�D  �D  �mBY  8Y   n�1.1.4  �   z  &  �" �:  ��E     �      �� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  �  8"W   	+  K�   �   	%  L�   	�  M�   '  ;  �  
s&  G   )  A"K  Q  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  ?  -    �   m�  �  �  ?  U    f  ��  �  U     ?  -   -   U    J   �"    �  PH�  Ǟ  J   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q'  0ڰ  S?  8O�  T  @��  U  H �  ��  <v �-   ��  �U    �  ��  ""  ��  �  @       @     @       �  
�   4  :  E     v  :-   ~   w�  
  yE   �!  yE  �   zE  H  zE   "  |Q  �  (  M} N    5�  N   `�  	G   _| 
  
!  +  ?      2      B  U     
�  �    �  N   �n  �!   �   pmoc�  stibu!  ltuo�  tolp 
:  �0  
�8  5"�  �  �$  �4  S�  x U$   len V+  e� W    
�#  Y�  �  
�%  {�  �  	  G   G   	  U    �  
�#  �  "  G   ;  G   G   U    
�.  �H  N  c  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(    (�/  ;  0�  U   8*  �  @ +  �  
u(  
c  �  
�2  (  "  G   6  U   6   {  
�3  ;I  O  Z  {   
v)  ]g  m  �  {    @    
�3  y�  �  G   �  {  @   U    
H7  ��  �  G   �  {  �   
  51  0�>  y2  �n   � �   �Z  *
 ��  / ��   $ �<  ( 
2$  ��  -4  l   �  $8  �   !  �+  \   �G   �  �N   }  �-   )$  �@   
c,  +G   
+D  C4   N   
�
  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � ^  H'  	�%>  N   
�Y  �*  Q" G, ' �, �' �$ �& �& g% 	<$ 
W# r( �  b+ M( �$ �+ �# �& �' �'  ! !9& "�! #�* $�) %0% &�, '^$ (", 0�( 1�  @�, Ar' QF+ R5" S�" T�# U�+ Vc, W-! X!+ `�' a	+ b�( c�+ p�! �n" �g! ��( ��* ��( ��% �B# ��* �.# ��) ��) �S' ��% ��) ��# �" �8' �' �e* ��$ ��! �H! �~% �# ��  �$ ��, ��% ��" � " �* �O% �s& �s) ��+ �( ��  �) �& ��+ �F* �~! �_& ��) �U) ��# � .( N   2�  |$  �$ �' )  ;, 9Y  �& �q�  ^�  s�   
- tv  W& v�  �, w�  �@ x�  �% yK   T$ z�  (�� |�  0V }v  4- ~�  8$� ��  <- ��  @% ��  D�* ��  H�# ��  L- ��  P��  ��  X�( �
  `0$ ��  h�� �
  p#! ��  x4J ��  �j( ��  ��; �  �ڰ  �?  � ^  �  @    j  ^  	  @   ? �# ��  �( �!  �  �) B�  �; D   ^�  E  ڰ  F?  lzw G	  _| I�  � pos J�  �!O�  K
  �!��  L
    ^  �  "@   � �' N�  '  #,  �  ��E     �      �A  $��      (�  � $_|  
  �� �� $%  �  � � %�Y  �  �� � %�# �  �� f� %�* �  �� �� %- �  � �� &�  ���E     'Eof �K�E     &�! A��E     (�s   )�� ^  ��*c 2  +��E     (  �  ,T2 +��E     5    ,T��,Q1 -W�E     T  ,Us   (Ps �  .c =2  D� 8� %�* >�  �� �� +G�E     T  e  ,Us  +]�E     �  }  ,Us  +L�E     �  �  ,Us  -��E     �  ,Us   /e  x�E     �s �0v  �� �� 1�s 2�  -� '� 2�  ~� x� 2�  �� �� 3�  ��+��E     B  (  ,T3,Q��,Y�� -��E     N  ,Q��    45* ���E     �       ��  5��  �"  	� � 6ڰ  �?  W� U� 7K  ��E     �r ��  0X  |� z�  +�E     Z  �  ,Uv  -%�E     Z  ,Uv   4, ���E     �       �K  5��  �"  �� �� 8�; �"  T9K  P�E     P�E     )       �0X  �� ��   :;( �e  ;��  �#   <=) �G   �  ;��  �)  =^% ��  =v  ��  =ڰ  �?  =�U ��   >�* wG   ��E     �       �T  5��  w(  � �� 1Pr 6ڰ  {?  �� }� ?�U |�  �\6^% }�  �� �� 6v  ~�  � � -M�E     B  ,T1,Y�\   >�& <2  P�E     �      �#  5��  <&  �� �� 6$� >�  � � 6�  ?�  �� �� @p @
  [� U� 6�Y  Av  �� �� A#  ��E      r Z04  �� �� 1 r 2@  	� � -��E     5  ,Ts    <n# G   M  ;��  $  =/� �   #�- W�  ��E     4      ��  $^�  W!  I� ?� $�; X!  �� �� B�U Z�   %ڰ  [?  ;� 7� .zip \�  � q� &�  �8�E     C�  @�E     �r w|  0"  � � 0  U� Q� 0
  �� �� 1�r 2.  �� �� 2:  � �� DF  +|�E     O  `  ,Uv  -��E     �  ,U~ ,Tt    +��E     O  �  ,Uv  +��E     f  �  ,U| ,T
,Q�L -��E     Z  ,U| ,T}   E�# J@   ��E     ,      ��  $^�  J%  T� P� $�  K%@   �� �� $_| L%  � � $/� M%@   � s� .zip O�  � � /�  ��E     t R0�  K� A� 0�  �� �� 0�  ,� "� 0�  �� �� 1t 2�  �� �� 2�  �� �� F�  C�E     G�  @t �  2�  �� �� Cg  ��E     �t $f  0x  �� �� 1�t 2�  !� � 2�  p� n� 2�  �� �� -��E     �  ,Us,T~ ,Q
    +N�E     r  ~  ,Q|  -��E     r  ,Qv   C�  p�E     �t    0�  �� �� 1�t 2�  �� �� 2�  � � 7K  ��E     �t �   0X  +� )�  -z�E     (  ,T0   /  ��E      u 	0"  ^� P� 0   � �� 1u 2.  :� 6� G:  Pu r  2?  t� r�  HL  �u 2M  �� �� 2Y  � � +?�E     �  �  ,U ,T0,Q
  -q�E     �  ,U ,T0,Q~        I�! 7`�E     L       ��  $^�  7#  V� P� .zip 9�  �� �� %ڰ  :?  �� �� C�  q�E     s @x  0�  � � -}�E     A  ,Us  -��E     Z  ,U| ,Ts   <�% ��    Jzip ��  Jpos ��  ;_| �
  ;/� ��  =�Y  ��  =�U ��  K�  )LM�� �    <�% ��  g  Jzip �(�  ;/� �(�  =�U ��  NL  =�� ��   L=�� ��  =>+ ��    <% ��  �  Jzip �(�  Olzw �  =/� ��  =�U ��   <�" ��  �  Jzip �"�  =^�  �  =�U ��   P�  ��  Jzip �!�   <�* h�  O  Jzip h!�  ;^�  i!  ;�; j!  Olzw l  =�U m�  Q�  � >�$ S�  ��E     c       ��  5^�  S#  K� =� 6�U U�  �� �� ?uR V�  �nR�  b��E     +��E     (  �  ,Us ,T0 -�E     }  ,Us ,T�n,Q2  ^    @    SK  ��E     *       �(  TX  U UM  M  �U�h  �h  �V�I  �I  �Vn  n  V�s  �s  �V�`  �`  vWBY  8Y   U�D  �D  � ބ  W  s&  -H �:  ��E     ��      �� (\  �9   S,  i   �L   S�  tint S�  u�   @�   �  �    p   	@   �  #	@   X  &	@   �  )	@    �  ,	@   (�  -	@   0/  2S   8�  5S   < �   S�  "�   �  8"c   A+  K  �   A%  L  A�  M  S'  S;  S�  "<  s&  S   �  Z   T4 S   �F Z   )  A"�  �  �   ��  �  �a    ��  ��  <h ��  �I  �   �  X�  �  a   �  |  9    �   m    %  |  a    f  �$  *  a   H  |  9   9   a    J   �"T  Z  �  PH�  Ǟ  JW   ֳ  KL   Dpos LL     N  /[  O   �K P'  (�R Qd  0ڰ  S|  8O�  TW  @��  UW  H j�  �  k<v �9   k��  �a    �  ��  ""  �3  9  L   W  H  L   W  L    ]  S�  �   q  w  %�  H   v  :9   �  L�  +x N�   +y O�   �  Q�  "�  ~   w  
  y�   �!  y�  �   z�  H  z�   "  |�  �  (�  M} Z    5�  Z   `�  	S   _| 
W  
!  <  ?   ]  2   ]  B  a     �    "�  �  (Q     S5   0�  T5  N5  V  �   W�   H� X  �1  ZS     �  5  �  \�  �  Z�  Z   �b  �!   3�   pmoc3�  stib3u!  ltuo3�  tolp :  �$  �8  5"|  �  V�$  �4  S�  Dx U5   Dlen V<  e� W]   �#  Y�  "�  �%  {�  �  %�  S   S   �  a    �  �#  �    S   /  S   S   a    �.  �<  B  %W  S   S   a    �8  `��  .   �   �; �  �1  S   �5  �  �+  �   `(    (�/  /  0�  a   8*    @ �  �  vu(  
W  "�  �2  (    S   *  a   *   o  �3  ;=  C  %N  o   v)  ][  a  %v  o  W  L    �3  y�  �  S   �  o  L   a    H7  ��  �  S   �  o  �   �  51  0�2  y2  �b   � �   �N  *
 �v  / ��   $ �0  ( 2$  ��  -4  l]  "?  +  �a  "P  S�  $8  �]  "h  t    ��   "  {"  �5  !  �<  "�  \   �S   "�  �  �Z   }  �9   )$  �L   �   9   c,  +S   C*  6a   +D  C@   �]  P-    :   �f	  Dxx ��   Dxy ��  Dyx ��  Dyy ��   5  �#	  "f	  8  ��	  ��  �y   ��  ��   $  �x	  c   ��	  �	  %�	  a    �  ��	  Kl  �a    �  ��	   s  ��	  �"  $
  
  �   +R
  �� -
   �W .
  Kl  /a    %  D}
  uR F
   �
 G
   }  IR
  OZ   -��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<L  5�  >�   ��  ?�  �"  A�  �"  B�  i!  C�   %!  E�  (2!  F�  0�  G�  8   I�  �"   s�  ��  u�   5�  v�  ֳ  x�  !  z�  m  {�   v  }Y  J  �#�  �  P�!  �}�  ڰ  |   {3  ��  S0  ��  �/  ��  �1  ��  �1  �Z$  	Y/  �}
  	�*  �2  (	�)  ��  0	+:  �j$  8	<8  �z$  X	�*  ��  � �3  �"�  �  �(  ��  Oe �4$   �-  ��  ڰ  �|   U  �"�  �  �  82  ah !:$   Oe "�  U1  #}
   ;+  $  0 i(  �$?  E  l;  ���  ah �:$   Oe �G$  y2  �b   {:  �p  (�� �o  h/ ��  p�� �  x T   � �  �  _  ��  �!  �   �  �  �  �    �  �  �   �U   (�    03"  �  8�    @`  !�  Hd  "  P�@  $�	  X�;  )  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7�  ��� 8A  �K <�  �ڰ  =|  �^�  >H  �U  @}
  �t  B�	  �k  Ca   ��L  Ez  � "   �  �  1  Xm�  ��  o�   �@  p�	  �e q�  �L  r+  P @  $%�  �  P  0\A  �-  ^�   ��  _�  �W `�  x a�  �@  b�	   �e dL  0�"  e�  pi"  f�  x� g�  ���  ib  �.a k�  ��  l�  �J  m�  �Mj  o  ��  q�  ��  r  �	M  ta    	Z  u9   	_"  w�  	(   x�  	Ud za    	�L  |r  ( �!  F#N  T  Z!  A�  ��  C�   T D`  �!  E�  "  F�   ZS  Z   �`  Y   3�  bmys3�  cinu3�
  sijs3    bg3�  5gib3F  snaw3  ahoj3�    bg3�  sijs3=    bg3�  5gib3�
  snaw3k  ahoj3�  BODA3t  EBDA3�  CBDA3  1tal3�  2tal3�   nmra �  �  �C  HT  0  `)�  �  �"  �e  �1  gf	   H+  h�   x+  i�  0��  k_   8�)  n#�!  h�'  qP  p��  rH  t�*  y�  x   �  A  �S  I�  �  �)8  >  �!  H�w  $  �a    7:  �&  s4  ��   b  8H�  !  J�   m  K�  A� M�  �� N�  �  P�  
  Q�   ��  R�  (�  S�  0 �  Uw   x  t�  x   �$  #  �!  0'r  ad  )�   �1  *�  &D  +�  2B  ,�  x� -f	     �)  �  �"  P��  ��  �   �1  ��  �&  �?  �3  �f	  ]7  ��  0�7  �a   @�1  �H  H �  ~�  P6  .  Dtag �   Kl  �   �6  	  .  Z�5  Z   
y  i7   �&  9  F9  8%  �*   �,  
A  ./   6
�  b 8
y   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  �  Z�8  Z   �&  �:   4,  �6  $  �/  l9   �2  ��  h  �#  ��  �'  �Q  W  �  f  �   �2  �r  x  %�  �   l/  ��  �  9  �  �  �   �   "�  ;)  H�7  �#  ��   :  ��  �5  �7  F1  ��  ,8  ��   2*  ��  (�*  �E  0`1  �f  8��  ��  @ �  �-  ��  "=  d)  s[  a  �  p  a    9  F#�  "p  �$  @J�  �#  L�   y2  Mb  W� OQ  �� Pw  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!  	  �-  (qK  �-  s�   Oe tK  ��  ub  � v�   |  �/  )]  c  �  w  �  �   g%  .�  �  %�  �   �.  1�  �  %�  �  �     s	  73  6�  �  %�  �  �     �8  :�  �  �    �  �   "3  >]  $)  Y'  -  �  K  2  �  &     �6  _W  ]  �  {  2  �  �     �3  f�  �  %�  2  �  �   ;0  l�  �  �  �  2  �  �   �&  x�6  ah � =   y2  � b  H�8  �   P�8  � K  X�'  � {  `� � �  h�9  � 6  p 2  �.  ��  "9  H2�  Mj  4   H5  5  (�)  6  0�  7�  8�  8  @ �0  :H  T%  �=  ڰ  ?|   �0  @�  q5  A�  L)  B�  )  C?  Ǟ  E�  �  F�  `Ud Ha   � X+  J%  �  1  7  =  �  `  H  �  �  �  ;   �&  &l  r  %}  �   �1  *�  �  �  �  �   �6  -�  �  %�  �   w-  1�  �  �  �  �   �;  4�  �  %�  �   =;  8    �    �  �   B$  <+  1  �  E  �  �   2  @Q  W  �  u  �  �  �  H   7  G�  �  �  �  �  �  �     q8  N�  �  �  �  �  H   )2  S�  �  �     �  �  �  H      �  k.  ���  ah �=   #,  ��  H�4  ��  P,;  ��  XEY �+  `/q �`  hZ)  �}  p�#  ��  x'0  ��  �.  ��  ���  �E  �� �u  �`9  ��  ���  ��  �5  ��  �U#  �  � �2  ��    a   �&  0�_   y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��  *  V'x   ~   V�0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |�   �'  ��   �   �  �   l   �  �    �	  �9  �!  !  %$!  l   �    A2  �0!  6!  �  T!  l   �  ?  T!   �   8(  �!  ��  )�    $�  )!  �-  )$!   )  Z!  "�!  3  <�!  �� >%�!   ��  ?%l    �!  #  A�!  �!  �U  �,�!  �!  �B  �#"  �� �m   Oe �#"   fP  �,/"  �"  4I  P��"  ֳ  ��   �� ��"  �q ��"  R` �#  �W �?#   P �#k#  (�U  �#�#  0�v  �#�#  8�v  �#�#  @�J  �#$  H "5"  ��  ��!  wq  ��"  �"  �  �"  �!  �   �J  �#  #  %#  �!   �\  �%#  +#  �  ?#  �!  U   \  �K#  Q#  �  e#  �!  e#   U  U  �w#  }#  �  �#  �!  �!  U  U   �O  ��#  �#  �  �#  �!  U  U   �n  ��#  �#  e#  �#  �!  |   ;O  ��#  �#  e#  $  �!  |  U   -k  ��#  *�  �5"  "#$  =  �(  ��  <  �D  &�  �  j$   L    N  z$   L    �  �$   L    wH'  �%2  ��  8 Y%  ��   [   ��   \  п   ]  �U  ^  ��   _   �   `�  (W�   a?  0�   b�  2�   c�  4 ��   e�$  �   p$2%  �$  ��  � ��&  ��   ��   ��   ��  *�   �h  ��   �h  	��   �h  
�   �h  .�   ��&  ��   ��&  (��   ��&  <�   ��&  X0�   ��  pY�   ��  xA�   ��  |M�   ��&  ���   ��&  ���   �h  �W�   �h  ���   �?  ��   �?  ���   ��&  �[�   ��&  ���   ��  ���   ��  ���   ��  ��   ��&  � �  �&   L    �  �&   L   	 �  �&   L     �  �&   L    �  �&   L    c�   �8%  �   �#�&  8%  8�   ��&  ��   >'  ��   h   +�   >'  r�        �  [�   "'  P0�    ((  ��   *�   �~   +�  U�   -(  ª   ./(  (��   /?(  �	|�   1   	P�   2   	��   4O(  	��   5_(  �	n�   7�  (	��   9o(  0	��   A(  �	��   B�  �   /(   L       ?(   L    D'  O(   L    &%  _(   L    �&  o(   L    �  (   L    �  �(   L    ��   D�(  Q'  Z�  Z    4�(  �   5�  B�  �  ��   �   <�(  $�  !)$�(  �(  VP�  a�  !,)  
)  �  #)  |  #)  ))   �&  �(  ;�  !1;)  A)  %`)  �(  �  �  �  �   w�  !8l)  r)  %})  �(   *�  !;�)  � !=�(   �� !>/)  �� !?`)   M�  !A�)  })  ��  !h!�)  �)  V��  ��  !u-�)  ^*  ��  8!V^*  �7  !X�)   ��  !Yc*  �R !Z�*  �� ![�*  �� !\�*   �� !]�*  (a� !^�*  0 "�)  t�  !�o*  u*  %�*  �)   S�  !��*  �*  %�*  �)  �      !�  !��*  ��  !��*  �*  %�*  �)  �   e�  !
�*  �*  �  �*  �)  �   |�  !1	+  +  �  -+  �)  -+  �(  &     �  !�!@+  F+  Vì  ��  !�-X+  �+  �  8!��+  �7  !�3+   ��  !��+  �R !�t,  O� !��+  �  !�,   y� !�L,  (a� !��,  0 "^+  ��  !��+  �+  %�+  3+   ��  !��+  ,  %,  3+  �  �      i�  !�,,  2,  %L,  3+  �  �  y   p�  !&Y,  _,  %t,  3+  �  y   !�  !D�,  �,  �  �,  3+  �   %�  !j�,  �,  �  �,  3+  -+  �(  &   ��  !�-  ��  !�-   �� !�)-  � !�>-   �)  -  �   -  �)  )-  �   -  K+  >-  �   /-  ��  !��,  �  !� ^-  D-  jhG  "5�-  Qnum "7�  Qstr "8�   *f  ":d-  �_  "=�-  +key "?�-   Kl  "@@    �K  "D$�-  �-  �d  "H�-  �-  �  �-  �-   �-  �r  "K.  	.  ?  .  �-  �-   Uj  ("Oy.  ��  "Q�   ֳ  "R�  [M "S�  �V  "U�-  �F  "V�-  �B "Xy.    �-  �@  "\ �.  .  N�  ##�.  �.  U  �.  �   :�  #)�.  �.  �  �.  �   8�  #/�.  �  #5/  V #7U   x #8�   ��  #:�.  ��  #=$/  %/  ��  (#?Z/  I_ #A�"   J�  #B�  �m #CZ/    /  f�  #Ml/  r/  �  �/  �  �   �  #U�/  �/  %�/  �  �   ��  #Y�/  �/  �  �/  |  /  �  `/  �/  �   r�  #a�/  �/  �  0  /  U   ��  #e0  0  U  .0  /  e#   ��  @#i�0  4v #k �.   �y #m �/  v #n �/  Ty #o 0  hn #q �.   S�  #r �.  (��  #s �0  0��  #t �0  8 ".0  q�  #i�0  �0  C  �   $I1  ��  $K�   ��  $L�  ��  $M�  R` $O1  K�  $P1   �  7  ��  $R�0  ��  $R41  �0  I�  $ZU1  ��  $\�    A�  $^:1  MĿ  $a�2  ��  $c%   ת  $dU1  8�  $e�&  @*�  $f   ��  $h�(  (T $i1  0��  $k3  P�  $l3  X��  $m3  `��  $o�  h+ $p�2  p��  $q�2  x��  $r.  ��  $t�  ��o $u�2  ��" $v�2  �C�  $w�2  ���  $yh  ���  $zh  �}�  ${f	  �	�  $|�  �j�  $}  �[ $~�   �  $��   3  �    ��  $�a1  ��  $��2  a1  ��  ($�<3  N  $��   ��  $��  �  $��  ��  $��  A�  $��    \�  $�H3  �2  �  $��3  v�  $��   }�  $��  +x $��  +y $��   \�  $��3  N3  I�  X$�4  ��  $�?   o�  $�  )r  $��  (dS  $��  0"�  $�<3  81�  $��  @��  $��3  H'�  $��  P �  $� 4  �3  ��  $�!24  84  M��  x$��4  ah $�   �O  $��2  �Q  $��  g  $��  �  $��  �  $��4   d  $�5  @E�  $��(  P��  $��  X��  $��  \��  $��  `f�  $�>'  h�  $��  p m  5   L    A  5   L    �I  `%U6  Q  %W�   �g  %X�  �;  %Z�  �U  %[�  �B %]�   �o  %^�  "Y  %`6  (+I  %a6  8
  %c�  H�!  %d�  J�   %e�  LH  %f�  N�`  %h�  P�X  %i�  RO  %k�  T,G  %l�  V�t  %m�  X �  6   L    I  %o5  �g  8%� 7  ��  %��   )r  %��  dS  %��  
�B  %��  �P  %��  �p  %��  �K  %��  =  %��  me  %��  +^  %��  �]  %��  �u  %� 7  
h  %��  $^K  %��  &tR  %�a   (%?  %�a   0 �  7   L    �]  %�"6  �S  8%?8  ��  %A�   )r  %B�  dS  %C�  
�B  %D�  �A  %F�  �n  %H�  �n  %I�  �W  %J�  me  %K�  +^  %L�  �]  %M�  �u  %O 7  
h  %Q�  $�V  %R�  &tR  %Xa   (%?  %Ya   0 �u  %[7  JW  �%xI:  ��  %z�   =  %{�  �<  %|�  tB  %}�  �k  %~�  �m  %�  
�D  %��  gJ  %��  !X  %��  �S  %��  5f  %��  ?X  %��  �a  %��  �_  %��  �a  %��  Gf  %��  �=  %�I:   �E  %��  0F  %��  8�A  %��  @F  %��  H�E  %�Y:  P5D  %��  TH  %��  V#l  %��  X$r  %��  Z_S  %��  \'N  %��  ^?_  %��  `L  %��  b�O  %��  h�O  %��  p~e  %��  x [  %��  z0m  %��  |�M  %��  ~rM  %��  �]  %��  ��g  %��  � h  Y:   L   	 P  i:   L    �X  %�8  kE  @%�;  �^  %��   zp  %��  dv  %��  �i  %��  �<  %��  �F  %��   �D  %��  (�p  %��  03X  %��  8 �b  %�v:  K_  @%��;  ��  %��   �J  %��  �<  %��  e  %��  $� %��  dk  %��  ![  %��  L^  %��  �`  %��;  yN  %�<  ,ma  %�<  4�Z  %�P  :�q  %�P  ;r  %�h  <�u  %�h  = P  <   L    P  <   L    P  !<   L    	l  %�;  �M  (%8=  ��  %:�   �T  %;�  �P  %<�  
�K  %=�  B  %>�  ^  %?�  �g  %@�  /o  %A�  %B  %B�  �O  %C�  �<  %D�  �]  %E�  *w  %F�  dW  %G�   �F  %H�  " e=  %J.<  |[  &O^=  �� &Qh   �\  &Rh  +red &Sh  q  &Th   �[  &V=  �?  (&��=  `a  &��   �L  &��=  r  &��=  &W  &��  �F  &��=    �  Ik  &�j=  ��  'L >  }W 'N   ��  'O�  ��  'P�   ��  'R�=  8y  h'lA>  �~  'n�   ��  'o�  �~  'pA>    >  Q>   L    `�  'r>  ,�  0'��>  }W '�   ��  '��  +def '��  ��  '��  +tag '��   cy  '��  ( ˣ  '�]>  ��  '��>  Ԛ  '�    cy  '��  �}  '��   	�  '��>  U�   '�U?  �~  '��   ��  '��  ˧  '��  �~  '�U?  i{  '�[?   �>  �>  �  '�?  >i   (J�?  +tag (L�   ��  (M�  /� (N�  �f  (O�?   �  2\  (Qm?  G   (�@  +Tag (��   g  (��  �=  (��  Ja  (��   mn  (�@  �?  �v   (�~@  �T  (��   �Y  (��  D  (��  S  (��  E]  (��  ;C  (��  �: (�3   �[  (�@  DQ  (�@  E]  (�   ;C  (�  �: (3   �i  (�@  >M  0(.AA  ��  (0�   �Z  (1�  vv  (2�  �r (3AA  =P  (4�  �Q  (5GA   ^�  (6H  ( ~@  �@  �p  (8�@  CE  (Y�A  �B  ([�   b  (\�   Pq  (^�A  ZA  �m  (x�A  ��  (z�   �R  ({�  Up  (|�A   �=  (~�A  �U  (�B  �  (P   
  ( P  Sd  (!h  �Q  ("P  �G  (#P  �v  ($P  �=  (%P  sD  (&P  �\  ('P  �X  ((P  	`N  ()�B  
 P  �B   L    �T  (+�A  >t  (�C  �>  (��B   � (��B  !  (�h  m  (�h  �[  (�h  SX  (�h   �<  (�C  �B  x@  ("aC  �  ($�   �`  (%�  TL  (&1  �o ('aC   gC  P  �h  ()C  �Z  (<�C  �  (>�   �f  (?gC   fR  (AzC  x(Z�C  lj (\mC  l�Y (]�C   ms   (VD  �  (X?   �r (_�C   J  (a�C  �t  (r!D  "D  VU<  �c  ((��D  �B (�3   �c  (�3  �y (�3  �Y  (��  cC  (��   �  (�?  $ 	\  (�'D   L  (� �D  �D  P�i  �(�gI  ah (�   �u  (��?  �	�v  (��  	�R  (��   	o  (�@  (	�& (�6  0	�Q  (�7  �	@  (�=  �	5�  (�?  �	<  (�8  �	�`  (��  0	�a  (�MA  8Jos2 (�i:  h	F�  (�;  �	j  (�3  0	 M  (��  8	w_ (�8K  @	�>  (�iK  H	�A  (��K  P	^Z  (��K  X	�f  (��K  `	KT  (��K  h	�i  (�a   p	Q  (�a   xJmm (�a   �Jvar (�a   �	g  (�a   �	�Y (��A  �	Fq (�!<  �	jQ  (��  �	nQ  (�C  �	m  (D  �	�P  (�=  	@  (�  @	B  (L  H	�u  (?  P	�u  (^=  Q	�;  (�  X	zQ  (3  `	FN  (�  h	T  (3  p	!u  (�  xJcvt (L  �	2i  (gI  �	)  ()�	  �	�  (+�  �	�j  (-�  �	:>  (.�  �	�_  (0?  �	S?  (3?  �	E�  (4D  �	�W  (6U  �	XA  (8�  �		K  (9�  �	�c  (?�  �	][  (@�  �	�J  (B�  �	'<  (C3  �		Z  (E3   	�q  (F�  	�G  (G�  	�T  (H�  	�a  (I3   	�\  (K3  (	�u  (L�  0	o  (ML  8	^C  (N�  <	:W  (O�2  @	_  (Q3  H	�@  (R�  P	>  (S�  X	}?  (TU  \	m?  (UU  `Jbdf (X�D  h	�k  (\�  �	�Z  (]�  �	Pl  (h�  �	(a  (i�  �	i (ma   �	�d (na   � �Q  (�[  �g  (�"�I  �I  P�t  x(�8K  ��  (��D   ֳ  (��L  ȩ  (��  �m  (�  �1  (��   x (��  (^�  (�H  0��  (��  8   (��  <�;  (�  @�C  (��  `� (��  d"f (��  h�I  (�?  lDpp1 (��  pDpp2 (��  �Ǟ  (��L  ��y  (��L  �	BJ  (��L  	�<  (�3  	bL  (��   	Ud (�a   (	�W  (��  0	r�  (��  4Jpp3 (��  8Jpp4 (��  H	O�  (�3  X	��  (�3  `	�k  (�}
  h �^  (EK  KK  �  iK  �D  �  H  �?   �D  (*vK  |K  �  �K  tI  �  �  �   �b  (A�K  �K  �  �K  tI   SQ  (Q�K  �K  %�K  tI   Z�=  Z   (TL  �G   �v  k_  <L  ok   �`  (_�K  ^=  H  �j  @(��L  ڰ  (�|   �0  (��  q5  (��  
0�  (��     (��  Dorg (�  Dcur (�  " (�   �   (�3  (H� (�1  0�>  (��  8 ,L  (�%L  @\  (�'�L  �L  V�r  �d  (�  M  M  V�a  
�  @)E�M  ^�  )GH   �k )H�  ��  )I�  /� )J�  T�  )Kh  z�  )L�   ��  )M�  (�f  )O�?  0Vu  )P3  8 �  )RM  M��  )U�M  ��  )W�   �  )X�  /� )Z�  c�  )[�M  = )\�M   �  �M   L   � ��  )^�M  Y�  ()acN  ��  )d�   �  )e�  c�  )g1  ��  )h1  "�  )j�   �  )k�  $ ��  )mN  -�  )r�N  ��  )y�   ��  )z�2   8�  )|oN  9�  )��N  z  )��   �  )��  �  )��   �  )��N  �  )��N  ّ  )��N    �N  ��  )��N  J�   )�`O  ��  )��   ��  )�`O  �  )��  ��  )��  ��  )�fO   �N  O  ��  )�O  ��  )��O  O  ��  )�!�O  �O  PU�  �)R�Q  �-  )T�   ^�  )UH  ڰ  )V|  ��  )W�  �!  )X�   �  )Y�  ${3  )[h  (S0  )\h  )G�  )]h  *��  )_�  ,�_  )a?  0�  )c�M  8Y�  )d�M  x�  )e�M  �T )g�M  �	�  )hcN  	��  )j�M  8	9�  )k�M  x	��  )l�M  �	x�  )m�M  �	*�  )o  8	1�  )r�2  @	��  )u�  H	�y )v�2  P	v�  )w3  X	x�  )x�  `	Ω  )zX  h	��  ){�  0	��  )| X  8	9�  )~�W  8	�  )�Q-  X	Q  )��0  `	��  )��  h	��  )�0X  p	:�  )�  x	%�  )�  �	��  )��	  �	��  )�lO  �	ת  )�6X  � ��  0)�[R  ��  )�?   ��  )�?  �  )��O  ��  )��  3�  )��  L�  )�   ��  )��   +BV )�L  ( 4�  )��Q  ;�  )�xR  "gR  �Q  Ma�  H)��T  ��  )��   ��  )��  ��  )��  п  )��  �U )��  ��  )��  W�  )�?  �  )��   �  )��  (�  )��  0��  )��  8[@ )��  <}�  )�f	  @�  )�?  `��  )��  h	�  )��  p��  )��  �j�  )�  ��  )��  �	�  )��  ���  )��  ��  )��  ���  )��  ���  )��  �ɼ  )��  �=�  )��  �6�  )��  �!�  )��  �"�  )��  �6�  )��  ���  )��   ��  )��  �  )��  $�  )��  n�  )��   ��  )��  (&�  )��  0��  )��  4�  )��  6ɰ  )��  85�  )��  @ Z�  )�~R  [�  )�$�T  �T  P��  �)/�U  �  )1�T   	�  )2bW  H	E�  )5[R   	3�  )6�  PJNDV )7   X	��  )A3  `	!�  )B3  h	��  )C�  p	��  )D�  t	x�  )F�M  x	)�  )G�2  �	.�  )JU  � M׬  �)�2W  *�  )�h   ��  )�h  ��  )�h  �  )�h  .�  )�2W  ��  )�BW  x��  )�2W  ��  )�BW  8	0�  )�  �	Y�  )�  �	A�  )�  �	M�  )�  �	��  )�  �	��  )h  �	W�  )h  �	��  )	RW  �	[�  )
RW   	��  )?  �	�  )�  �	��  )�  �	��  )�  �	��  )�  �	��  )�  �	�  )�  �	��  )�  �	��  )�  �	y�  )�  �	��  )�T  � �  BW   L    �  RW   L   	 �  bW   L    ��  )�U  ��  )|W  �U  7�   )�W  ��  )h   �  )�  Kl  )"3  ��  )#�  M�  )&�  ��  )'�  �  )(h   ׵  )*�W  ��  )*X  �W  ��  )L�T  �T  0X   L   � %  U1  ��  `*,dX  ah *.   m */�  X ��  *1pX  <X  M��  H*<�X  ah *>�   �� *@?  0��  *A?  1A� *C�  8�� *D�  @ ��  *F�X  vX  M�  *QY  �  *S�(   ��  *TY   �(  Y   L   � ;�  *V!Y  �X  xX  h+*vY  ah +,M$   �q  +.�  8�'  +/?  <iO  +0vY  @��  +1H  ` �  �Y   L    Y  +3�Y  'Y  ��  +?-�Y  �Y  �  `+�:Z  *�  +�3   O�  +�		  z�  +�		  �� +��  6�  +��   ��  +��  $�K +��2  (h�  +��2  0ڰ  +�|  8�� +��Z  @ ��   +X|Z  �� +[�Z   �q +`�Z  +add +c�Z  U1 +i�Z   �  �Z  �Y  �  |   |Z  %�Z  �Y   �Z  �  �Z  �Y  �  �  �   �Z  H�  +k:Z  "�Z  ��  +�"�Z  �Z  ;�  �+�V[  O�  +�3   Ǟ  +�3  ��  +�3  �U +��  ڰ  +�|   �� +��_  ( ��  +�"b[  h[  Q�  +��[  �k +�3   ��  +�3  b +�w\   K�  +�"�[  "�[  �[  �  0+�@\  �  +�   ��  +K]  b +�\  ��  +W]  �  +�  ֳ  +h  C�  +�   ��  +	�  $��  +�  ( W��  Z   +�w\  ��   }�  ��  ��  �  ��   I�  +�@\  ��  +�h[  W"�  Z   +��\  :�   G�  ��  Z�  z�  !�  ��  d�   �  \�  	��  
��  Ѻ   ��  +��\  W��  Z   +�K]  ��   ��  F�  r�  ػ  ��  ��  _�  j�  ��  	 e�  +��\  [�  +�c]  i]  %y]  �  �   1�  +�[  ��  h+uK^  �� +xe^   �q +~v^  �Y +�v^  �L +�v^  ; +��^   �> +��^  (nD +��^  0�M +��^  8�: +�_  @�[ +�-_  H�l +�S_  P` +�|_  X�9 +�|_  ` %e^  �Z  3  3  |   K^  %v^  �Z   k^  �  �^  �Z   |^  �  �^  �Z  �   �^  �  �^  �Z  3  		  �?  ?   �^  �  �^  �Z  �  �^   �  �^  �  _  �Z  �     �   �^  %-_  �Z  V[   _  %M_  �Z  V[  �  M_   �  3_  �  |_  �Z  �[  �  �  �?   Y_  :�  +��]  "�_  ��  +��_  ;�  p+4�`  ڰ  +6|   ��  +7�  ȩ  +8�X  ��  +9  Ǟ  +:-+   �  +;-+  (��  +=a  0��  +>a  8�C  +@  @� +A  H�;  +C�  P.�  +D?  X�� +E?  Y8�  +F?  Z��  +H?  [�  +I?  \�� +K�`  ` ��  +��`  �� +��`   �q +��`   %�`  �`  a   ?   �_  �`  %�`  �`   �`  ��  +��`  "�`  �  ��  +bLa  Ǟ  +d3   ��  +e3  O�  +f3   Q�  +ha  (�  +lfa  la  �  �a  �D  �  �2  �?   ;�  +r�a  �a  %�a  �D  �2  �   Pw�  �+w�c  �I +y�_   �� +{�c  pJtop +|   �	�� +~�c   	�y  +�c  �	a�  +��  �	�  +��  �	�  +��c  �Jcff +��O  	��  +��T   	��  +�d  (	��  +�a  0	׹  +�?  8	��  +��  <	P�  +��  @	"�  +��  D	c�  +��  H	��  +��  L	T�  +��2  P	0� +��2  X	�o +��2  `	�  +��  h	;:  +�&  l	zd +�?  p	��  +�&Ya  x	��  +�&�a  �	Q  +��0  �	��  +��  �	Z�  +��2  �	��  +�.  �	}�  +�f	  �		�  +��  �	E�  +��(  �	f�  +�>'  �	��  +��  � �  �c   L   0 La  �c   L    La  �  d   L    �	  ��  +��a  �  +�##d  )d  ��  �+<4e  ڰ  +>|   ��  +?�  ȩ  +@�  ��  +A  Ǟ  +B-+   �  +C-+  (��  +E�  0��  +F�  8�C  +H�  @� +I�  P�;  +K  `˹  +L�f  ��� +M?  �8�  +N?  ���  +P?  �b�  +Ra   ��  +Sa   ��� +U�f  � ^�  +�Ae  Ge  �  [e  d  �   G�  +�he  ne  %�e  d  �  �  h   r�  +��e  �e  �  �e  d  �  �   h�  +��e  �e  �  �e  d    �  +��e  ��  +��e  �e  %f  d   ؽ  @+��f  �� +��f   �q +��e  VY +�$4e  c +�$[e  f +�$�e   2 +�$�e  (�J +�$�e  0� +�$�e  8 %�f  d  �  �  �  ?   �f  ��  +�f  "�f  Z��  Z   +��f  >�    �  /�  i�   v�  +��f  f�  +W)d  ��  +v6g  O�  +x3   Ǟ  +y3  ��  +z3   ��  +|�f  ��  +|Pg  �f  �  +/cg  ig  P��  �+��h  �I +��f   �� +�j  �Jtop +�>'  �	�� +�j  �	�y  +�Cg  x
	Q  +��0  �
	�  +��  �
	�o +��2  �
	��  +��  �
	��  +��  �
	+ +��2  �
	��  +��2  �
	��  +�.  �
	}�  +�f	  �
		�  +��  �
	a�  +��  �
	�  +��  �
	�  +��c  �
	E�  +��(  `	;:  +�&  h	��  +�Di  p	�� +��i  x	f�  +�>'  �	��  +��  �	zd +�?  �	��  +��	  � �   +�Di  �� +��i   �q +��i  ;U +��i  �" +��i   õ  +�Qi  Wi  �  ki  Vg  �   �  �i  Vg  �  �  �  �2  �(  ?  &  Di   ki  %�i  Vg   �i  �  �i  Vg  3  �   �i  �  �i  �i  3  �   	d  �i  '�  +��h  "�i  �  j   L   � 6g  /j   L    D�  +� <j  ��  �+TGk  ڰ  +V|   ��  +W�D  ȩ  +X�X  ��  +Y  Ǟ  +Z-+   �  +[-+  (��  +]�  0��  +^�  8�C  +`�  @� +a�  P�;  +c  `.�  +e?  ��� +f?  �8�  +g?  ���  +i?  �b�  +ka   ��  +la   ��� +n�l  � 9�  +�Tk  Zk  �  nk  nk  �   /j  ��  +��k  �k  %�k  nk  �  �  h   �  +��k  �k  �  �k  nk  �  �   ��  +��k  >�  +��k  �k  %�k  nk   ש  +�l  l  �  l  nk   ��  @+��l  �� +�l   �q +�k  VY +
%Gk  c +%tk  f +%�k   2 +%�k  (�J +%�k  0� +%�k  8 %�l  nk  �D  dX  �X  ?   �l  �  +l  "�l  ^�  +�	m  Ǟ  +�3   ��  +�3  O�  +�3   ��  +��l  P��  �+��n  �I +�/j   Dcff +��O  ��� +��c  �Jtop +�   h	�� +��n  p	�y  +��n  	a�  +��  	�  +��  	�  +��c  	��  +��  �	��  +��  �	0�  +�?  �	׹  +�?  �	��  +��  �	f�  +��n  �	P�  +��  �	"�  +��  �	c�  +��  �	��  +��  �	T�  +��2  �	0� +��2  �	�o +��2  �	�  +��  �	;:  +�&  �	zd +�?  �	��  +��T  �	��  +�&Ya  �	��  +�&�a  � 	m  �n   L    	m  �  �n   L    �  +�m  +�  +�3o  �� +�go   �*  +��o  �" +��i   %ao  ao  �D  dX  �X  ?  &  Ya  �a   �n  3o  �  �o  ao  dX  �   mo  �  +��n  "�o  �  +�#�o  �o  ��  (+p  ڰ  +|   ^�  +�p   +4  F�  +	q  w�  + a     ӫ  +�?p  �� +�]p   �q +�np  �i +��p   �  ]p  �o  |  3  3   ?p  %np  �o   cp  �  �p  �o   tp  ��  +�p  "�p  ��  +�#�p  �p  ��   0�p  O�  23   Ǟ  33  ��  43  V 6�   �  	q  �  		  a    �p  R�  +-.q  iq  ��   +/iq  f�  +1#"   ]J +2#"  ��  +3#"  V +4#"   ""q  �I +6"q  "nq  ��  X+A)r  8�  +D!)r   ��  +E!/r  �  +F!5r  ��  +G!;r  կ  +JVr   *�  +Okr  (��  +R�r  0��  +W�r  8�  +[q  @��  +^!�r  H�  +`"�r  P �Z  �_  �f  
j  %Vr  3  		  �   Ar  U  kr  U   \r  %�r  �i  a   ?   qr  %�r  �  �&  �T   �r  �p  �o  a +b�q  �4 +e�r  "�r  W!c Z   ,-		s  �-  eQ A5 }4 �C c^  m,;Es  Qs ,=�   Qf ,>�  Qi ,?�  Qu ,@�  Qb ,A?   �] ,8ks  b ,:�r   +u ,C	s   "P ,EEs  e_ ,E�s  Es  OZ   -��u  /P  4 �/ �X :L #6 �7 �j �K �c 	�S 
�3 �Q a/ 4K oX '8 b �b �G �A ZU  ~H !)R "(e #3G $V5 %^ &�M '�V (�G 0XT 1�P @$W ApI Q< RhO SFe T�D U�k V�E W�` X�[ `Z3 aQ< b�C c!A p�\ ��B ��\ �?^ ��/ ��^ �]1 ��= ��5 �i ��E �9 �vb ��1 �/ ��V ��l �p0 �{V �}l ��] ��d �>` ��0 ��f ��@ ��. �= �L? �43 �i- �0= ��R ��\ �(7 ��\ ��M �d ��> ��2 ��- ��a �8 ��d ��1 ��U ��N � OZ   (�u  f  c �? G]  W)K Z   ��w  �_  �[ 5 �Z �W ?@ �K �< �6 �6 	W. 
P @ QX �] �@ �> �K �= �L R 9B B �[ �T rc �X E8 �O 9D �j �A Q  �< !GS "�K #	L $L %�< &�e '�= (= )�8 *[f +S= ,�c -�4 .e /�D 0M0 18i 2I 3�5 4tf 5 X 6+Z 7�P 8�O 9\ :�_ ;�1 <�f =�l >�_ ?�4 @�4 A�_ BR2 C\j D�` E�` F'l GLC H�. I�N JWZ K @7 �u  �  �w   L   I "�w  !4/ �w  	��G     A1 .!�l  A? .$a  A,C .'+I  A8�  /)�Z  A��  /,�_  A�  //�f  A��  0 
j  B/ 1&#gx  mx  }g 81(�x  I_ 1*�"   �F 1,�=  W 1-�.   �  1/�  (�o 10�x  0 �  A�a 16/$  AeW 19/$  �` 1D&�x  �x  J (1F.y  I_ 1H�"   ��  1I�  /� 1J�  ZL  1K1    A�E 1Q/$  A[g 1_/$  �_ 2EH  "Fy  OZ   -��{  }h  K; cC *_ 0 k �_ F �g jj 	9X 
�9 �R �B dJ ;T 'V �G Y E  h %4  C !x^ "O6 #�Z $LO %sL &HQ '�? (aS 03 1�Y @wY A�_ Q;Z R�f S�6 TQi UU V�H W�E X�F `�S aT b]] c�i p4; �[ �TL �[7 �M �6I �ri ��5 ��j ��V ��F �o_ �F_ �k. ��H �5Y �vG �.M �?J ��Q ��< ��@ �`2 ��k ��i ��M �ZA ��c ��W ��R �cK �4? ��k �|] ��7 ��< �.: ��H �-a ��9 �@- ��L �<P �t5 �&2 ��1 �Ff � �_ 31H  W�9 Z   3O�{  �f  �: 6<  �F 3U�{  k@ @43M|  ڰ  45|   �U 46M|  �4 48@   8T 49@   8 4:@    /� 4;@   (�k 4<@   0+ptr 4>a   8 �  �Z 4@�{   H 4@p|  "_|  �{  |A  5.�|  �U 50M|   �k 51y  +end 52y  +ptr 53y   D2 55v|  l 55�|  v|  �B 6=b  WG Z   6A}  �Q �d �/ VV  . 6L_}  +a 6NFy   +b 6OFy  +c 6PFy  +d 6QFy  +tx 6RFy  +ty 6SFy   �U 6U}  "_}  M#\ �7?  ڰ  7A|   �U 7B�  _ 7D?  �D 7E?  �2 7F�|  �h 7L_}  C 7M_}  ,@ 7N_}  D� 7OFy  \E�  7R[R  `y�  7So  �3�  7To  �+NDV 7U   ��j 7Wb  �O 7YFy  �0O 7ZFy  �Mj  7]ۀ  �LM 7^�i  ��d 7_�T  �Mk 7c?   �j 7d?   [ 7f?  �g 7hvY  ,� 7kFy  $N� 7lFy  ($/ 7mFy  ,,/ 7nFy  0�A 7p?  4��  7sÅ  8��  7uT�  � �G 6Z.!  "  p}  �3 6[ 3  �W  8v�  �1  8xo   ad  8y@   m 8{Fy  u4 8|Fy  1� 8}Fy   �d 6[.�  "�  3  �T H6f�  +pt0 6h�   +pt1 6i�  +pt2 6j�   +pt3 6k�  0+op 6mb  @ yQ 6o�  �] 6o�  "�  �  -[ 6s,�  4E 86|�  �I 6~��   _F 6��   W 6���  �; 6���  B 6�b   ڰ  6�|  (�U 6�M|  0 �J 6t-��  �  |: 6x��  ��  %��  �  �   �N @9�ۀ  ah 9�
�   LM 9��i  8 �N 9���  5 9��  ��  h+x  :!	��G     h7x  :+	 �G     hx  :A	 �G     aCx  :I	��G     aOx  :X	��G     d��  :g�p  	��G     d�  :q{q  	`�G     ax  :{	 �G     d�  :��o  	 �G     bVP :��r  	��G     d�(  :�I  	@�G     \  ��   L    "Ё  bO +��  	��G     a�x  �	`�G     a�x  �	 �G     n.y  	��G     n:y  e	@�G     WfR Z   ,��  cb  �- \4 wd }N Jl �0 P Ng �S 	sH 
D< B6 �P Ec �B �8 �L >] _ u: �A �R �J _ �C k �j  W^ LA�  �  �   L    "�  �Z P�  ��  ;!5�  ;�  �  J�  �   m�  ;$V�  \�  �  z�  �O  �T  �      �  ;*��  ��  h  ��   X  �   �  ;.��  ��  ?  Ѓ  gR  �  �      d�  ;4܃  �  �   �  gR  �  �      B�  (;:O�  ��  ;<$)�   �  ;=$J�  Y�  ;>$z�  ��  ;?$��  ��  ;@$Ѓ    " �  ��  ;:`�  O�  OZ   8V��  {k �8 : ok �? Pc   OS   8h��  3�F   pyEd ���| �j 8�	�  �H 8�Fy   sR 8�Fy  0 8�Fy  `d 8�Fy  �f 8�?   IW 8���  M�a P8���  1� 8�Fy   /� 8�o  ,] 8�?  h; 8�?  	Ah 8�Fy  m 8�Fy  �5 8�Fy  A 8�Fy  �b 8�'   �2 8�'  @�y  8���  ` 	�  Å   L    00 8��  "Å  �< 8��  "ԅ  �  OZ   <. �  �0 ` �; 0<F\�  �U <HM|   �d <J?  Z <K?  	`- <M@   1T <N@   �� <P\�    h  l�   L    �` <R �  > <R��  "x�   �  �h <Uކ  [M <W?   +min <YFy  +max <ZFy  QG <\Fy  �d <]Fy   �T <_��  "ކ  �U <_��  ��  OZ   <y�  �N � M�S (<~��  �  <�   �/ <���  �[ <�_|  �d <�?  Mk <�?  1� <�Fy  /� <�o   �^ <�o  ${� <���  ( �  '  ��   L   � �] <��  �U <���  "��  M|< �I<���  �  <�   �K <��  Q <���  �a <���  8�/ <���  `0�[ <�S|  �H�8 <�Fy  �H�S <�Fy  �H�8 <�Fy  �H,N <��  �H^ <�?  �H%9 <�?  �H�^ <�?  �HV <�?  �H�7 <�_|  �H1. <�_|  �HEg <�x�   I�A <�Fy  I��  <���  IC"  <�Fy  I�  <�Fy  IS <�Fy   I�8 <�Fy  $Id <��  (I�k <��  8I/ <��  HIB1 <��  XI�k <��  hI�> <�?  xI�L <�b  |IfF <��  �IzS <��  �I�a <��  �IqF <��  �I υ  &b <�͇  �A <�Ӊ  ͇  ��  ='�  �  �  ��  �  ��   Q>  �z  =+�  �  �  +�  �  +�   1�  a?  9~  =/C�  I�  �  b�  �  �  >'   "�  =6n�  t�  �  ��  �  �      ��  ==C�  �  =Bn�  ��  =G��  ��  �  ˊ  �  �   Ӏ  =KC�  ݓ  =P�  �  �  �  �  �2  �  �  +�      `�  =Wl  ��  =Zn�  3�  =_6�  <�  �  U�  �  �2      y  `=d��  �~  =f"ى   -�  =g"7�  g�  =h"��  ��  =i"ˊ  7�  =j"�   Y�  =k"b�  (�  =l"��  0&�  =m"��  8U�  =n"�  @A�  =o"*�  HY�  =r׊  P��  =s�  X "U�  g�  =d�  ��  QN :<�  +j <@    �- =Fy   < ?�  �; ?T�  �  m>1��  Qr >3Fy  Qf >4�{  Qi >5b   �0 >/��  +u >6Z�   b >8�{   7 >:��  �D (>=�  ڰ  >?|   �U >@M|  _| >A�  +top >B�  �  >C�    ��  fI >E�  ��  OZ   ��  �h  K ya H fP . �? �N �e eG 	uP 
�Q if �A {\ �5 u3 �2 �S �? <4 IR �5 q7 Sa N �F k< K �/ �: �Z  OZ   ��  5S  (I J �^ �Z �8 �e c\ �= �g 	rl 
�T �l �Q kb �e 2j �Q |F �h �9 y1 oh I. �8 T �R �8 :f TS �g CV 0\  => !�^ "�T #Z $M3 %�P & /6 E��  �� E	�   4d �n�  �� �	�  /� �b  m�  �b  ��  ���  �K �b  8idx �b  8i �b  2tmp -��    4CA ���  �� �	�  :num �o   4] �Ə  �� �!	�  :idx �!o  :val �!Fy   0�J �Fy  ��  �� �!	�  :idx �!o   0:k �Fy  �  �� �"	�   0d4 �b  ,�  �� � 	�   4. {R�  �� {#	�  :val |#Fy   4�U kx�  �� k!	�  :val l!b   0)D do  ��  �� d	�   42h T��  �� T	�  2ڰ  X|    0�S 5	�  
�  ڰ  5|  :e 6M|  �  7�  �U 9�  �� ;	�   0�1 j?  (�  :buf j�|   0�U Pb  F�  :buf P!�|   ,�N ��BF     c/      ���  �  �1  `� 8� 7buf �1�|  ;� )� �K �1�  � � gV �1  �� �� ND �1?  @� <� W: �1Fy  {� y� \: �1Fy  �� �� 5�  �1��  �� �� 
�g ��  T� B� 
LM ��i  (� � 
�U �M|  "� � 
ڰ  �|  �� �� 
�8 �Fy  _� S� 
j �Fy  �� �� 
u8 ��  �� e� 
�i �?  � �� 
MI �?  �� �� !�s ���  ���~
�8 ��  P    
�A �Fy  � � 
�G �	�  �  
�  ��  n b op1 �h  T  !�y  ���  �غ~!�P ���  ���~
u;  U  � s !E[ S|  ���~!�- ?  ���~
9� �|  F ( 
=0 b  � � !�7 S|  �ع~!1. S|  ���~!Eg l�  ���~!Kh ��  ���~;�  ��PF     T�> N#�PF     *       m�  
�S  ��  � � �PF     �  Uu   $�� ��  
��  ��  � � ��  W^F      � ��  ��  i a ��  i a �  � � �  S C � %�   � 2�  � � ?�  � � J�     U�  @ < x�  y^F       � �V�  ��  � v ��  � v  Kb�  p� ��  c�  6 . p�  � � �g �^F       �� �ӕ  �g � � �g   �� �g 7 3 �g z v   ��  _F      � �g�  ��  ��  � � ��  � � <x�  
_F       
_F            �N�  ��  D > ��  D >  Bh_F     Uu 5��  {   �^F     Ə  ��  Uu T{  �^F     Ə  Uu Tz  I_F     n�  Uu T} s    ]3PF     Ӗ  Us  ]\PF     �  Us  lPF     �  Uu   #�RF     p       ʗ  idx ao  � � 
/� bo  � � x�  �RF       �RF            b}�  ��  0 . ��  0 .  �RF     Ə  ��  Uu Tv  �RF     Ə  ��  Tv �RF     �  U���~  $� ؘ  idx xo  [ S 
/� yo  � � isX {?  � � $P� c�  v �Fy    uRF     �  H�  U���~ �RF     Ə  Uu T|   x�  ,RF        � y��  ��  [ S ��  [ S  @�  SF      SF     	       ��  � � �  � �   $Щ �  
/� �o  � � idx �o  N @ #RWF     �       Q�  x1 �Fy  � � y1 �Fy  ' # x2 � Fy  _ ] y2 �$Fy  � � x3 �(Fy  � � y3 �,Fy  � � ]WF     Ə  ��  Uu Tvz lWF     Ə  Ι  Tv{ ~WF     Ə  �  Tv| �WF     Ə  ��  Tv} �WF     Ə  �  Tv~ �WF     Ə  .�  Tv �WF     ��  U���~R~ Y|   x�  (WF      � ���  ��  !    ��  !     �  *^F      *^F            �ɚ  �  l  j  �  l  j   �]F     Ə  �  Uu Tv  	^F     Ə  ��  Tv *^F     �  U���~  $�� ��  
ug �b  �  �  #RVF            l�  val ���  �  �  YVF     ��  c �UF       � ��  � ! ! t w! u! � � �! �! L� �UF        � � �! �!  �! �!    ��  �VF      P� <�  ��  " " ��  i" g" ��  �" �" P� �  # �"   S�  ZF      ZF     7       ���  �  _# ]# r�  �# �# e�  �# �# &ZF     7       ��  �# �#   6VF     �  Uu   $� ��  op2 (h  #]\F     &       �  !R 1%��  	 �G      #2\F     &       k�  !R I%��  	�G     X\F     ��  U T���~Q� R���~X	�G     Y0  $� ��  !R a%��  	 �G     \F     ��  U T���~Q� R���~  #�[F            �  !R y%��  	��G      $ � ��  v0 �%Fy  $ $ v1 �)Fy  a$ [$ v2 �-Fy  �$ �$ isV � ?  �$ �$ ��  �bF       @� �Ҟ  ��  E% A% ��  �% �% ��  �% �% <x�  �bF       �bF            ���  ��  & & ��  & &  B�cF     5��  2  ��  cF       �� �g�  ��  ~& z& ��  �& �& ��  '  ' <x�  cF       cF            �U�  ��  @' :' ��  @' :'  B�cF     5��  4  �SF      r ��  5��  s  �bF     Ə  ��  Uu T0 �bF     Ə  ��  T2 �bF     Ə  ̟  T4 �bF     Ə  �  T1 cF     Ə  Uu T3  #�pF     %       v�  
&D  �#Fy  �' �' 
2B  �#Fy  �' �' �pF     ��  T�  Uu  �pF     ��  qF     R�  Tt   #�pF            �  
&D  �#Fy  �' �' 
2B  �#Fy  ( ( �pF     ��  ͠  Uu  �pF     ��  �pF     R�  Tt   #�pF            I�  arg #Fy  I( G( �pF     ��  1�  Uu  �pF     R�  Tt �  $� E�  
P   �  x( l( 
�?  b  ) �( 
kd -b  d) ^) 
�C   �  �) �) 
� .�  3* /* 
��  &4  �* |* !Wl $�|  �ػ~!2> $Fy  ���~
�T b  �* �* 
}[ b  7+ /+ ady  �  �+ �+ adx !�  , , asb "�  �, �, $� ��  
ȩ  g'�  �, �, 
��  h'  ;- 7- 
7B  i'  z- t- �kF     � Ţ  U���~T2 6lF     � ݢ  Us  QlF     � U���~� $ &  �  �mF       P� �n�  '�  �- �- 4�  @. 6. 4�  @. 6. P� A�  �. �. 6N�  ��~B�mF     T��~   �  �nF       �� ��  '�  �. �. 4�   / / 4�   / / �� A�  K/ G/ 6N�  ��~B�nF     T��~   2kF     �  ��  Uu  :kF     �  AkF     ��  JkF     ��  RkF     ��  �lF     $ J�  U} Tv  mF     $ h�  U} T|  EmF      � ]mF     �s ��  Tv Q�ػ~5n�  }  �mF     F�  ٤  U~ T�ػ~Q�з~R�ط~X1Y0 8nF     �s �  T| Q�ػ~5n�  ���~ qnF     F�  U~ T�ػ~Q�з~R�ط~X1Y	s ���~�  #�jF     �       ٥  
; �"Fy  �/ �/ 
#; �)Fy  �/ �/ 
�I �"�`  �/ �/ �jF     ��  ��  Uu  �jF     ��  �jF     ��  �jF     ��   #RpF            �  arg �#Fy  0 0 ZpF     ��  Uu   #pF            }�  
@. 	#Fy  50 30 
�T 
#Fy  \0 X0 &pF     ��  o�  Uu  -pF     ��   #�oF            �  
�[ #Fy  �0 �0 
); #Fy  �0 �0 �oF     ��  Ԧ  Uu  �oF     ��   $� b�  
fX *#Fy  �0 �0 
9�  +#Fy  31 +1 pF     ��  pF     ��  :�  Uu  pF     ,� CpF     �  KpF     �   $�� ��  arg E#Fy  �1 �1 �oF     ��  Uu   #GoF            �  
&D  U#Fy  �1 �1 
2B  V#Fy  �1 �1 OoF     ��  �  Uu  VoF     ��  eoF     R�  Tt   $�� �  
�` gb  E2 +2 
&i hb  j3 L3 
/� io  �4 �4 
�D jo  �7 �7 #�gF     �       ,�  idx �!�  �: �: 
�` �!�  �: �: H0 hF      hF            � �  Z0 �: �: g0 6; 4; hF     ~v U���~#T15Z0 ���~  �hF     ��  U���~  $�� 
�  
E�  #�(  ^; Z; 
��  #�  �; �; nn /�  �; �; mm 3�  *<  < 
�� #o  �< �< 

Q #o  j= `= $ � �  tmp D&Fy  �= �= �g (gF       0� I#%�  �g )> '> �g N> L> 0� �g u> q> �g �> �>   ��  OgF      `� O��  ��  ��  �> �> ��  3? -? <x�  SgF       SgF            ���  ��  �? |? ��  �? |?  B�lF     Uu 5��  z   gF     Ə  ת  Uu Tz  (gF     Ə  Uu   �gF     n�  Uu Tx y   #LfF     `       d�  idx ^#�  �? �? 
E�  _#�(  @ @ pfF     �  �fF     9�  #/fF            ��  
@. w'Fy  ,@ *@ 
�T x'Fy  S@ O@ >fF     ��  EfF     ��   #fF            �  
�[ �'Fy  �@ �@ 
); �'Fy  �@ �@ fF     ��  &fF     ��   #�eF     0       �  
�O �'Fy  �@ �@ 
$5 �'Fy  A A �g �eF      �eF            �Ŭ  �g 4A 2A �g YA WA &�eF            �g �A |A �g �A �A   �eF     ��  �eF     ��   #�eF     .       G�  
fX �'Fy   B �A 
9�  �'Fy  %B #B �eF     ��  �eF     ��  �eF     ,�  #3eF     P       ��  idx �#b  JB HB 
E�  �#�(  oB mB UeF     �  qeF     ��   #�dF     M       �  idx �#b  �B �B 
E�  �#�(  �B �B eF     �   #�dF     0       ��  
&D  'Fy  �B �B 
2B  	'Fy  C C 
�Y 
'Fy  MC IC 
= 'Fy  �C �C �dF     ��  �dF     ��  �dF     ��  �dF     ��   $@� �  r !'Fy  �C �C �+ ^dF      p� -Ѯ  �+ D 
D  �dF     ,�  Uu   #�lF     <       #�  i 7!�  dD ^D �lF     ��  Uu   x�  /dF       � ~Y�  ��  �D �D ��  �D �D  �  �gF      �gF     	       ��  �  G 
G �  G 
G  H0 �hF      �hF            ��  Z0 1G /G g0 YG WG �hF     ~v U���~#T65Z0 ���~  � %iF      �� �/�  � �G }G  ��  LiF      �� e�  ��  �G �G ��  �G �G  � @iF      @iF            ���  � H H   dF     �  ��  Uu  (dF     �  �iF     ,�  ݰ  Uu Tt  �iF     ,�  Tt   #ejF     %       W�  val {#Fy  ;H 9H idx |#b  `H ^H mjF     �  I�  Uu  ujF     ��   #FjF            ��  idx �b  �H �H NjF     �  Uu   #jF     ,       ?�  
&D  �#Fy  �H �H 
2B  �#Fy  �H �H 
�Y �#Fy  I I 
= �#Fy  EI AI "jF     ��  �  Uu  *jF     ��  2jF     ��  9jF     ��   #�iF     8       ��  r �#Fy  I {I U�+ �iF      �� ��+ �I �I   #oF     )       `�  
�O �#Fy  J J 
$5 �#Fy  CJ AJ �g .oF      .oF            �:�  �g hJ fJ �g �J �J &.oF            �g �J �J �g �J �J   &oF     ��  R�  Uu  .oF     ��   #woF     F       ��  arg �#Fy  :K 2K #�oF     /       �  
ah �!�  �K �K 
]h �!�  �K �K �oF     ,� Uv Ts   oF     ��  Uu   #mpF            P�  arg �#Fy  �K �K upF     ��  ;�  Uu  |pF     ,�  Tt   #�pF            ´  
&D  �#Fy  3L /L 
2B   	#Fy  mL iL �pF     ��  ��  Uu  �pF     ��  �pF     ,�   $@� �  idx 	b  �L �L 
ֳ  	o  �L �L $p� (�  
}R 	!o  nM jM E`F     Ə  Uu   x�  `F      `F            	j�  ��  �M �M ��  �M �M  `F     �  Uu   #qF     �       �  idx /	b  �M �M 
/� 0	b  �N �N ��  !qF      !qF     �       8	�  $�  �N �N �  wO sO �  �O �O &!qF     �       0�  �O �O <�  �P �P H�  Q �P T�  �Q �Q <x�  3qF       3qF            ���  ��  ZR VR ��  ZR VR  K^�  � ��  _�  �R �R  @� �qF       �qF     )        �R �R  �R �R    qF     �  �  Uu  qF     �   (�   XF      � (#H�  9�  <XF     l Ur   �cF     ��  `�  Uu  �cF     ��  roF     ��  Uu   #`ZF     �       �  
; s	Fy  7S 5S 
�I t	�`  \S ZS hZF     ��  ٷ  Uu  �ZF     ��   #�`F     6      �  
�T �	b  �S �S 
}[ �	b  �S �S !Wl �	�|  �ػ~!2> �	Fy  ��~
P  �	�  �S �S ��  daF      �� �	��  �  \T ZT �  \T ZT �  �T �T B�aF     Ts   ��  �aF      �aF     "       
�  �  �T �T �  �T �T �  �T �T B�aF     Ts   �`F     �  )�  U  �`F     �  �`F     ��  �`F     ��  aF     �  s�  U���~Q�ػ~ daF     F�  ��  U~ T�ػ~Q�з~R�ط~X1 �aF     �  ӹ  U���~Tv Q�ػ~ �aF     F�  U~ T�ػ~Q�з~R�ط~X1Y0  $О %�  !BN 6
��  �ػ~!�P 7
l�  ��~��  �NF       � :
��  0�  �T �T #�  (U $U �  gU aU 	�  �U �U ��  �U �U  ��  yOF      P� ?
̺  ��  7V 5V ��  _V ]V  �OF     ��  �  U��~T~  �OF     1�  U�ػ~T�ع~Q���~R��~X0Y0  $�� o�  
/� �
o  �V �V idx �
o  �V �V #MF     �       ��  x1 �
Fy  gW cW y1 �
Fy  �W �W x2 �
 Fy  �W �W y2 �
$Fy  �W �W x3 �
(Fy  #X !X y3 �
,Fy  HX FX MF     Ə  �  Uu Ts  !MF     Ə  �  Ts 3MF     Ə  3�  Ts ?MF     Ə  K�  Ts KMF     Ə  c�  Ts ZMF     Ə  {�  Ts |MF     ��  U���~R~ Y}   x�  �LF      �LF            �
�  ��  oX kX ��  oX kX  �  �WF      �WF            �
"�  �  �X �X �  �X �X  �LF     Ə  @�  Uu T}  �LF     Ə  X�  T} �LF     �  U���~  #�KF     �       *�  
/� �
o  �X �X 
�� �
o  �X �X idx �
o  [Y OY $`� �  x1 �
Fy  �Y �Y y1 �
Fy  7Z 3Z x2 �
 Fy  oZ mZ y2 �
$Fy  �Z �Z x3 �
(Fy  �Z �Z y3 �
,Fy  �Z �Z �KF     Ə  b�  Uu Tv  LF     Ə  z�  Ty  LF     Ə  ��  Tv LF     Ə  ��  Tv ALF     ��  о  U���~R| Y|  wLF     Ə  Uu Tv   @x�  �KF       �KF            �
%��  [ [ ��  [ [   $@� ��  
/� �
o  *[ &[ 
�� �
o  d[ `[ idx �
o  �[ �[ $p� ��  x1 �
Fy  c\ _\ y1 �
Fy  �\ �\ x2 �
 Fy  )] '] y2 �
$Fy  N] L] x3 �
(Fy  s] q] y3 �
,Fy  �] �] �JF     Ə  �  Uu Tv  KF     Ə  /�  Uu Tv  )KF     Ə  G�  Ty  5KF     Ə  _�  Tv CKF     Ə  w�  Tv iKF     ��  U���~Q~ X| Y}   @x�  �JF       �JF            �
%��  �] �] ��  �] �]   $�� Q�  
/� o  �] �] 
�� o  N^ J^ idx o  �^ �^ 
;c 	?  #_ _ $ � ��  x1 Fy  a_ Y_ x2 Fy  �_ �_ x3 Fy  Z` T` y1 #Fy  �` �` y2 'Fy  a a y3 +Fy  �a �a �TF     Ə  ��  Uu Tz  �TF     Ə  ��  Tv  �TF     Ə  �  Tx  �TF     Ə  #�  Ts  &UF     ��  I�  U���~Q} Yv  {UF     Ə  g�  Uu Tz  �UF     Ə  �  Tv  �UF     Ə  ��  Tx  �UF     Ə  ��  Ts  �UF     Ə  ��  T|   [F     Ə  T|   �  �JF      � H�  �  �a �a �  �a �a  @x�  �TF       �TF            %��  b 	b ��  b 	b   $�� �  v Nb  �b �b 
�` Pb  �b �b 
�^ Qb  c c (�  pJF      �� P��  9�  �YF     l Ur   (�  �JF      � Q�  9�  �YF     l Uu   �JF     R�  Uu Tt   #�ZF            _�  v bb  ,c (c �ZF     R�  Uu Tt   $@� ��  v ob  oc ec (�  �XF      p� u��  9�  �XF     l Ut   �XF     R�  Uu Tt   $Ъ 7�  v �b  �c �c (�  b[F       � ��  9�  t_F     l Uu   �[F     R�  Uu Tt   $0� ��  v �Fy  td rd 
�` �U  �d �d 
�^ �U  �d �d 
�_ �U  e e 
$_ �U  Ge Ee (�  �\F      p� �+��  9�  `F     l Uu   (�  �\F      �� �+�  9�  �_F     l Us   (�  �\F      Ы �+F�  9�  �_F     l Us   (�  �\F       � �+{�  9�  �_F     l Uu   4]F     R�  ��  Uu Tt  O`F     ,�  Uu   ��  �DF      �� -��  #�  te je �  �e �e 	�  Hf Ff ��  qf kf ��  �f �f ��  g g ��  ng jg ��  �g �g ��  �g �g ��  �g �g ��  }EF      � N��  0�  Jh Hh #�  oh mh �  �h �h 	�  �h �h ��  �h �h  ��  �EF      p� S�  0�  �h �h #�  i i �  0i .i 	�  Wi Ui ��  |i zi  ��  �EF      �� Xb�  0�  �i �i #�  �i �i �  �i �i 	�  j j ��  >j <j  h EF      � I��  � gj ej � �j �j � �j �j u �j �j  �DF     D� U���~T0Q
�I  ��  (CF      @� � ��  ��   h kCF      �� F�  � �j �j � (k $k � `k ^k u �k �k  h �CF      � ��  � �k �k � �k �k � �k �k u l l  h %DF       �  ��  � Gl El � ml kl � �l �l u �l �l  ��  uDF      P� &�  ��  �l �l ��  m m  ��  �FF      �� LE�  ��  @m ,m  �  �FF       �FF            V z�  �  (n &n  ��  �FF      К XI�  �  On Kn ې  �n �n ϐ  �n �n К 6�  �ػ~��  &o o �FF     O� ��  U| T(Q�ػ~ GF     [� 3�  U| T8Q0R} X0Y�ػ~ D[F     g� U|    � 0GF       � d��   �o �o � �o �o �XF      U���~TA  
�  �GF      `� v��  �  fp Vp �  fp Vp  �  }HF      }HF            ��  �  ,q *q �  ,q *q  (�  �HF      �HF            �?�  9�   � �PF      �� �u�   Sq Oq  �q �q  ��  �HF      �� ���  ��  �q �q UB �HF      Л �O �q �q Л [ r r IF     g�    B 0IF       � �,�  O Cr Ar  � [ lr jr YIF     g�   B uIF      @� �u�  O �r �r @� [ �r �r �IF     g�   B �IF      �� ���  O �r �r �� [ s s �IF     g�   ��  �IF      �IF     '       �H�  ��  -s +s =��  �IF     "       ��  Rs Ps JF     g� ,�  Us  JF     g� Us T    �  QJF      QJF            ���  �  ws us �  ws us  x�  �MF      �MF            n
��  ��  �s �s ��  �s �s  x�  �MF      �MF            U
�  ��  �s �s ��  �s �s  x�  lNF       lNF            
P�  ��  t t ��  t t  � QF      P� �	y�  � Lt Ht  ��  9QF      �� �	��  ��  �t �t ��  �t �t  � -QF      -QF            �	��  � �t �t  c �QF      �� �	b�  � u u t +u )u �� 1� C� �QF      �QF            � Tu Ru  {u yu    x�  0SF      0SF            N��  ��  �u �u ��  �u �u  ��  �VF      �� ���  ��  v v <^F     �t U���~  c 	YF       	YF     U       !u�  � {v uv t �v �v &	YF     U       � �v �v L� YF       �� �  w w  Gw Ew    x�  e`F      0� �	��  ��  pw jw ��  pw jw  ��  �`F      `� �		��  ��  �w �w hbF     �t U���~  x�  �`F       �`F            �	.,�  ��  +x )x ��  +x )x  NF     ��  D�  Uu  *NF     ��  \�  Uu  �NF      r ��  U| T���~#�Q R���~X�Y���~5��  ���~ QF     L�  ��  U���~ qSF     ��  ��  Uu  �SF     L�  ��  U���~ �YF     Ə  �  Uu T0 $[F     L�  +�  U���~ �[F     Ə  H�  Uu T0 �[F     Ə  e�  Uu T0 �]F     ��  ��  U���~Ts  �bF     Ə  Uu T0  Fy  Fy  ��   L    Fy  ��   L    Fy  ��   L    @   K  ��   L    "��  /XD ��  E�  �!sR  �G �!	�  ��  �!o  �� �o  Ǟ  �o  i �o  j �o  ��  �o  2��  ��  sum �Fy    Ry  ,U O /F     �      ���  �G O	�  Vx Nx W: P��  �x �x \: Q��  $y y Kh Rǉ  �y �y R S��  �y �y y9 T?  Iz =z !$g V��  ��idx Wo  �z �z sV X?  top Yb  i Yb  �{ �{ j Yb  �{ �{ $P� ��  
�g o?   | | 
kL rFy  \| X| �/F     Ə  ��  Us  m0F     Ə   �  B0F      B0F            �#�  �  �| �| �  �| �|  �/F     Ə  A�  Uu T~ !0F     ��  [�  U��~ B0F     ��  ��  U��~R X} Y��~� �0F     Ə  ��  Uu Ty �0F     Ə  Uu   K  Fy  ��   L    /Td z�  �     �G  	�  �I  _|  5�   ��  �-  z�  �3  Fy  i  o  /� !o  �` "?  �  %Fy  T�  H2nY 5ކ    ?  4^c ���  �  �&x�  `- �&@   8i �@   �� �o   4xK ���  �  �$x�  9� �$�|  `- �$@   8i �@    0�. l@   "�  �  l)x�  `- m)@    09F e3  @�  �  e*x�   4de Zf�  �  Z&x�  :val [&?   0�Y S?  ��  �  S+��   0�d L?  ��  �  L-��   4�6 B��  �  B$x�  �U C$M|   /�= p��  �@ p/ǉ   ,7 �,F     F      ��  �@ )ǉ  } } 7x1 )Fy  }} s} 7y1 )Fy  �} �} 7x2 )Fy  ^~ V~ 7y2 )Fy  �~ �~ 7x3 )Fy    cy3 )Fy  � !i> Fy  ��!Rf Fy  ��!r> $Fy  ��!�@ .Fy  ��XP0 �  ��P1 �  � y P2 �  *� $� P3 �  �� �� �  C-F       �� 4k�  4�  �� �� )�  #� !� �  H� F� �  m� k�  -F     ��  ��  Uu R} X Yy  1-F     ��  ��  T| Qv R~ X� �Yy  t.F     `�  �.F     $�  ��  Us TsQ��Y0 /F     1�  UsY0  ,QF � +F     �      �L�  �@ �(ǉ  �� �� 7x �(Fy  � � 7y �(Fy  {� s� !C"  �Fy  ��!�  �Fy  ��XP0 ��  ��P1 ��  �� ڂ 
�R �?  9� 7� �+F     ��  ��  Us R| Xv Yy  x,F     1�  �  UsY0 �,F     $�  >�  Us TsQ��Y0 �,F     `�   ,�I ��)F     �       ���  �@ �(ǉ  e� ]� 7x �(Fy  ΃ ă 7y �(Fy  N� @� ��  �)F      �� ���  ��  � � e*F     �t  I*F     1�  Uv Y0  ,�e ���E     �      �`�  9�@ �/ǉ  U7x1 �/Fy  +� #� 7y1 �/Fy  �� �� 7x2 �/Fy  �� �� 7y2 �/Fy  i� a� cx �/��  Y7y �/��  φ ˆ dx �Fy  � � dy  Fy  � ܇ �  �E       �z �  4�  �� �� )�  ܈ ڈ �  � � �   �g @�E      @�E            +r�  �g )� '� �g Q� O� &@�E            �g y� w� �g �� ��   �g I�E      �z D��  �g ȉ Ɖ �g �� � �z �g � � �g ^� Z�   �g X�E      X�E            F6�  �g �� �� �g Ê �� &X�E            �g � � �g 0� ,�   �g ��E      ��E            `��  �g m� k� �g �� �� &��E            �g �� �� �g � ��   �g p�E       { y��  �g � 
� z�g Ι} { �g 6� 2� �g y� u�   @�g ��E      ��E            {�g �� �� �g ތ ܌ &��E            �g 
� � �g M� I�    ,	X �p*F     �       �$�  �@ �*ǉ  �� �� �k �*�  �� � !\  ��  ���*F     �i ��  Us TsQ��R��X| Yv 5T�  �� ]�*F     �  Tw  +F     L�  Us   o_` &`#F     �      ���  �@ &.ǉ  Y� M� ;A '.��  � � �W (.  )� � Tk ).�  �� �� �R *.?  ߏ ۏ !\  ,�  ��~
Q> .  "� � 
�N /  �� �� 
�3 1�  � �� 
�O 2?  ;� /� ��  �#F      p� J	�  ��  ɒ Ò ��  ɒ Ò ��  � � ��  � � ��  R� L� ��  R� L� ��  �� �� ��  �� �� ��  � � ��  � � ��  N� H� ��  N� H� p� 1��  1��  1�  �  �� ��  �  �� �� �g $F      �� �L�  �g !� � �g F� D� �� �g m� i� �g �� ��   �g  $F       � ���  �g � � �g  � �g � � �g W� S�   �g �%F      �� ���  �g �� �� �g �� �� �� �g � � �g ,� (�   �g $&F      �� �6�  �g �g �� �g k� g� �g �� ��   �g Q&F       P� ���  �g � � �g D� B� P� �g m� g� �g Ø ��   �g �&F      �&F            ���  �g � �� �g ?� =� &�&F            �g h� b� �g �� ��   J&F     ,�   �$F     �i E�  Us Ts�0Q��R��Yy 5T�  �� ^%F     �i ��  Us T~ Q��R��Yy 5T�  �� �%F     �i ��  Us T~ Q��R��Yy 5T�  �� �%F     �i ��  Us T~ Q��R��Yy 5T�  �� ]�%F     �  T��~ (F     �i H�  Us T��~Q��R��Yy 5T�  �� m(F     �i q�  Us T��~5T�  �� �(F     �i Us Ts�05T�  ��  '�3 �?  ,�  �@ �8ǉ  )u1 �8  )u2 �8  )v1 �8  )v2 �8  �3 �8  u ��  v ��  w ��  �G  �Fy  s �Fy   /�I ���  �@ �+ǉ  ;A �+��  )ppt �+  )x �+Fy  )y �+Fy  pt ��   /~W ��  �@ *ǉ   /sU 81�  �@ 8-ǉ  �  9-  �K :-�  �8 ;-Fy  �7 =-_|  1. >-_|  Eg ?-x�  �A @-Fy  ��  A-��  ,N B-   ,�7 % F     �
      �?�  ;A %$��  � � �7 &$_|  �� z� 1. '$_|  {� g� Eg ($x�  y� U� �W )$Fy  � �� bN *$?  #� � 
�C ,3  �� �� 
�  .  �� �� !�k /l�  ��
`- 1@   !� � i 1@   y� _� 
QA 2h  �� �� #�F     X       ��  !��  g'  ��~.�  �F      �� j��  ;�  ɣ ţ  �F     ?�  ��  Us T�Q��~ �F     ?�  Us T��~Q�  $Ѕ 0�  !j9 }'  ��~!�/ }&'  ��~z�  fF       fF             �>�  ��  � �  z�  zF       zF             �s�  ��  �� ��  $ pF       � ���  P &� � C �� �� 6 � �  � ] G� ;� j զ ͦ w ?� 1� � � ا � �� �� ��  �F      `� �$�  ��  � �  ��  F      �� *M�  ��  m� i�  >�  _F      _F            >	��  L�  �� ��  U>�  �F      �� 8	L�  թ ѩ    ?F     H�  ��  Uu T��~Qv R~ X��~� aF     H�  �  Uu T��~R~ X��~� �F     ?�  Us T��~Q��~  #�F     k       ��  !{� �'  ��~!m  �'  ��~.�  �F      �� �	��  ;�  � �  .�  /F      /F     $       �	��  ;�  P� N�  XF     ?�  Us T��~Q��~  $�� ��  !j9 �'  ��~!�/ �('  ��~F     H�  G�  Uu T��~Qv R��~X  �F     H�  u�  Uu T��~R��~X  �F     ?�  Us T��~Q��~  $ � z�  
nY  �  w� s� c GF       GF     2       !H�  � �� �� t �� �� &GF     2       � $� "� L� QF       P� � I� G�  p� n�    @��  yF      yF             %��  �� ��   "�  �F      �F             [��  3�  ϫ ͫ  ��  wF       @� F��  ��  �� �� ��  3� /� @� ��  q� i� ��  � � L��  wF      p� �
�  Z� V� 	�  �� �� =��  �F            �  έ ʭ 	�  � � C� �F       �F            r 4� 2�  Z� X�      B�  �F      �� q�  P�  �� }� �� ]�  � �� h�  �� � � �F      `� ��  � 6� .�  Ks�  �� ��  x�  �� �� K��  �� (�  ��  �� }� ��  7� )� ��   � � ��  ֳ ȳ ��  ȴ �� ��  � ֵ ��  �� �� ��  U� K� ��  ̹ ʹ ��  �� � �  M� G� �  �� �� K"�  P� �  6#�  ��~�F     � T��~  Uz�  UF       �� ��  �� �   ��  �F       �F             �]�  �  E� 9�  z�  �F     	 �F             ���  ��  � ��  �F     ,� �F     ,�  =3�  �F     �       14�  c F       �� 9E�  � �� �� t � ޼ �� 1� C�  F        F             � � �  ,� *�    @��  tF      tF             J�      @�  �F      �F            3��  Y�  Q� O� M�  w� u�  Z�  =F       =F             ��  l�  �� ��  ��  �F       �� :�  ��  � � ��  -� )�  UF     1�  Qv R��Y1  ,�Y W��E     �      �B�  ;A W(��  r� f� j9 X(�  � �� �/ Y(�  ο �� 
�^ [o  �� �� i�- ^?  
O[ _�  (� $� 
�? `�  t� ^� #��E     V       ��  
 X �Fy  g� c� 
�f �Fy  �� �� �g ��E      @z ��  �g �� �� �g �� �� @z �g �� �� �g 4� 0�   ��E     C�   $ z ��  
4B �o  w� o� 
gE �o  �� �� 
/� �o  � ��  z�  )�E       �y ���  ��  �� ��  ��  ��E      ��E             �4�  ��  �� ��  k�E     C�   /z` �C�  ;A �)��  i �@   j �@   ^3�  �- �?  2�j �Fy  9 �Fy  ;Q �Fy  3 �Fy  uB �Fy  �] �Fy  �- �Fy  �d �Fy  ��  �Fy  �i �Fy  ?C �Fy  �b �?  2�X <�     2fh 8H�    .�h KFy  ��E           ���  9;A K!��  Um L!Fy  �� �� $`y G�  i Vo  a� M� �g 7�E      �y t��  �g �g �y �g 5� 1� �g x� t�   @�g ��E      ��E            i�g �� �� �g �� �� &��E            1�g 1�g    @�g `�E      `�E            Q�g  � � �g H� D� &`�E            �g �� �� �g �� ��    /J7 ,��  ;A ,"��   'A %?  ��  ;A %+ȇ   /�B >�  ;A #��  �  #  bN #��  �[ #_|  1� #Fy   /I: Z�  �� �   'uE ?  z�  �� )�   0�P �?  ��  �� �&�   0 D �?  ��  �� �&�   0�g �?  ��  �� �#�   0�0 �?  ��  �� �'�   0�- �?  �  �� �$�   0k6 �?  .�  �� �%�   4�e �H�  �� � �   Yk ZPF     �      ���  ?�� Z&�  U-�I [&k|  :� 2� ?WG \&@   Q-�  ]&  �� �� -�W ^&Fy  )� � -1� _&Fy  �� �� ?v� `&?  � (5�  bFy  5� � (lE c��  �� |� Nc wF      � h(��  � �� �� t 3� /� � � k� i� L� �F       P� � �� ��  �� ��    N>�  F      �� ���  L�  � �  L�g .F      Ѐ ��g -� +� �g R� P� Ѐ �g y� u� �g �� ��    �  0�X Eb  @�  :x1 E&Fy  :y1 F&Fy  :x2 G&Fy  :y2 H&Fy   /�R 
ti�  Mj  
t#�  LM 
v�i   /�i 
f��  Mj  
f#�  LM 
h�i   ',5 
\Fy  ��  LM 
\&�i   '�V 
RFy  ��  LM 
R&�i   '�J 
b  �  LM 
+�i  ug 
+b  )buf 
 +�|  idx 
"o   /�G 
�\�  LM 
�)�i  )buf 
 )�|  ��  
&4  Kl  
�	   '�5 
��  ��  LM 
�(�i  x 
�(�  )buf 
�(�|  )�  
��	  �U 
��  ��  
�&4  �O  
��2  inc 
�#�!  2�. 
�3  ��  
��    /a 
��  LM 
�'�i  )buf 
�'�|   .Gj 
��  `F     �       �S�  LM 
�&�i  �� �� �* 
�&b  f� ^� 7buf 
�&�|  �� �� gid 
�b  F� D� !9� 
�3  �PXlen 
��  �X
�U 
��  k� i� +  �F       � 
�<�  J  �� �� =  �� �� � W  #� � b  q� m� o  �� �� B�F     U�T   B�F     Qw R�X  'E 
xb  ��  LM 
x,�i  ug 
y,b  )buf 
z,�|  idx 
|o   '7b 
mb  ��  LM 
m&�i   /�M 
`��  LM 
`)�i  /� 
a)��  Kl  
b)��   a  /�M 
S,�  LM 
S$�i  /� 
T$��  Kl  
U$��   /�6 
Fb�  LM 
F#�i  /� 
G#��  Kl  
H#��   /�; 
9��  LM 
9#�i  /� 
:#��  Kl  
;#��   /�C 
%��  LM 
%$�i  Ah 
&$��  m 
'$��  �5 
($��   'TM 
Fy  ��  LM 
�i   'n\ 
Fy    LM 
�i   '�D 
�Fy  ;  LM 
��i   '�i 
��  �  LM 
�)�i  )len 
�*�  )vec 
�*�  ��  
��D  mm 
��   o  '%S 
��  �  LM 
�!�i   'H 
�xO  �  LM 
��i   '�c 
��T  �  LM 
� �i   .�c 
4�  rF     Z      �� LM 
4/�i  �� �� �. 
5/3  I� +� ��  
6/�  �� �� 
ڰ  
8|  �� �� !�U 
9�  ��~
�  
:  I� ?� 
�  
<?  �� �� $�� � 
�I 
k�`  L� 2� 
K 
l�Y  p� j� 
�J 
n?  �� �� 
Lb 
pP  %� � 
P  
t�  �� �� Xbuf 
u�|  ��!x� 
v_}  ��
39 
wFy  1� +� 
Mk 
y?  �� }� 
��  
z?  (�  � 
 �rF      �� 
��  �� �� L �� �� ? �  � 2 H� D� % �� ��  � lsF      lsF             
�# � �� ��  � psF      Э 
�w � �� �� � �� ��  � � Э  f� d� �sF     ,� U�C$   * �sF      � 
�- c �� �� V y� i� I M� 9� < F� 6� � p �� �� 6} ��~6� ��~� �� �� _� fzF     � �sF       � �
 � �� �� � �� ��  � � t� p� � �� �� � �� �� � &�  �  �� ��  �  �  �� �� ( � � 65 ��~6B ��~  ?tF      ?tF            F� -   Kb � ; c �� �� p � 
� } N� D� ��  !uF      �� �:    � huF       huF     +       �	 � �� �� � �� �� � � � � 6� 4� � ^� \� � �� �� � &huF     +       1� 1� 1 E E E' �uF     B| U| Tv Rs�X0   ��  �uF      а �, ��   � �uF        � �� � �� �� � �� �� � �� �� � � � � B� @� � i� g� �  � 1� 1� 1 E E E' vF     B| U| Tv Rs�X}    � gvF      0� ��
 � �� �� � &� � 0� � �� �� � �� �� � �� �� � D� >� � �� �� � �� �� 
 N� B�  �� �� " f� ^� . �� �� : F� >� F �� �� R .� � \ �� �� h �� �� N��  �vF      � dH ��  (� &� ��  M� K� ��  u� s� ��  �� �� �vF     ,� T�B$  Nb�  �vF      � i� p�  ��  �� �� }�  �� ��  <,�  �vF      �vF            j� :�  T�  � � G�  C� A�  <��  �vF      �vF            k	 �  �  m� k� �  �� ��  <��  �vF      �vF            lT	 ��  ��  �� �� ��  �� ��  <��  �vF      �vF             �
�	 ��   Kt @� �	 u � � � �� �� � k� e� � �� �� � � �  N�g YF      �� �($
 �g i� g� �g �� �� �� �g �� �� �g �� ��   N�g �F      � �%y
 �g :� 8� �g a� ]� � �g �� �� �g �� ��   �xF     ,� �
 U@<$ `}F     ,� �
 U@<$T|  �}F     s� �
 U
��Qv  $ & �~F     ,� U@<$T|    � �|F       � �	� � !� � � v� r� � �� �� � �� �� � A� =� � {� w� � � 1� 1� 1 E E E' �|F     B| U| Tv Y0   �uF     ,� � U�?$ �|F     ,� � U��~T��~ �~F     ,�  U��~T��~ (�F     ,� $ U�?$Tw  J�F     ,� U�?$  =O �}F     �       T �� �� ;  �}F      `�  � M  �� �� g  � �� Z  X� R� `� t  �� �� �  �� �� B�}F     T��~Q0R��~X0   ]~F     � U~� B%~F     T~     i�  �yF       �yF            x w�  �� �� w�  �� �� &�yF            ��  8� 6� zF     ��   @�  TzF       TzF            *� N�  ]� [� &TzF            [�  �� �� ]zF     Ci � Uu 5�. v  fzF     ��   -zF     F�  Us T��Q} R��~X0Y0   @� |zF       |zF            
�� �� �� � �� �� &|zF            �        Z �{F      �� 
`�  I  G  s g p  n   �{F     O� Uw T
�Q��~  'wD 
)�  
 LM 
)#�i   /�: 

Z LM 

)�i  A� 
)��  �� 
)��  Mk 
)z�  ��  
)z�   4�> 
�� Mj  
�"�  ڰ  
�"|  �U 
�"M|   Y�; 
�`3F     F      �D -�K 
�1�  �  �  -\  
�1�  6 * (�U 
��  � � (Mj  
��    �I 
��`  < / t3F      t3F            
� J/ � � ?/ � � 2/ &t3F            U/   �3F     �w Us    <H0 �3F      �3F            
�� Z0 g0 V T �3F     ~v UsT3  N�/ �3F      `� 
�[ 0 ~ z 0 � � �/ � � �/ `� 0 2 . =+0 �3F     )       ,0 j h 90 � �    N�/ �3F      �� 
�� 0 � � 0 
  �/ \ V �/ �� 10 F+0  � ,0 � � 90 � �    L�/ �3F      0� 
�0 � � 0 2 . �/ n j �/ 0� 10 F+0 p� ,0 � � 90 � �     Y"- 
��AF     x       �� -�K 
�1�  � � -\  
�1�  u o (�U 
��  � � (Mj  
��   � (�I 
��`  � z < / �AF      �AF            
�G J/ � � ?/ 	 	 2/ A	 ?	 &�AF            U/ h	 d	 �AF     �w Us    L�/ �AF        � 
��/ �	 �	 �/ �	 �	 �/ C
 =
  � �/ �
 �
 H0 �AF      P� �� Z0 �
 �
 g0   BF     ~v UsT15Z0 s   {8BF     �v    Y�D 
��F            �� -�K 
�1�  ? ; -\  
�1�  | x (Mj  
��  � � (�I 
��`  � � �F     Ci Uu 5�. s   4 > 
k� :ptr 
ka   �  
m  2ڰ  
r|    4�^ 
\� Mj  
\#�  5�  
]#Fy  LM 
_�i   0
Z 
A�  $ x� 
A*$ �j 
B*b  �[ 
DFy   k}  '[k ��  � �  �+  9� �+�|  x� �+$ 39 �+��  �g ��  gV ��  �Z �Fy  �- �?  T�  , 4g �� �  �&  x� �&$ LM ��i  �Z �?  ��  �� �W �?  �W �Fy  Uh �Fy  P�  �T  � Fy  �\ o  2    ^b ��  T�   2L4 �Fy  N� �Fy  �j �b    lO  4`B 4� L4 4%Fy  � 5%Fy  	m 6%Fy  �8 7%��  �Z 8%Fy   [ 9%?  �g :%M_  �? nFy  �P n"Fy  �1 o�  e-� �e4� �eP� �28x1 }�  8y1 ~�  8x2 �  8y2 ��  8x3 ��  8y3 ��  8x4 ��  8y4 ��  ^� � ��  m� ��  8x ��   ^� � ��  m� ��  8x ��   2� ��  m� ��  8x ��     42@ 	,$ �U 	,M|  <v 	-�   '8l �?  � ��  �'��  j9 �'�  �/ �'�  _I �Fy  �f �Fy  �; �Fy  91 �?  i �o   4�B B� ��  Bԅ  �  C  LM F�i  �X HFy  �h IFy  �I JFy  �a L@   UK M@   �^ N@   V O@   .F Qa  e0 Ra  1 Sa  l Ta  8i V@   �9 WFy  �2 WFy  2j @    e Fy  �0 Fy    "Fy  |6  Fy    Yg= ���E     Y       �c -J= �$_|    |ptr �$�  � ~ #��E            N (�  �@   � � (S �a   = 9 ��E     9� Tv   ��E      Us   0�I �a   � J= �0k|  :idx �0@   S �a    0f[ �a   � J= �/k|   0-J �@   � J= �*k|   4�l �� J= �%_|   4�T � J= �(_|  !G �(@    G)g _?  ��E     �       �B -J= _._|  � | -!G `.@    � p�  ��E     $`{  b�U e�  �\(ڰ  f|   { (3Q h@   � � <� w�E       w�E            y�  3 1  Z X  T�E     [� T1Rv Y�\  L� �E       �{ �  }  � �   4�; Lh J= L(_|  ڰ  N|   4�/ 8� J= 8$_|  ڰ  9$|  �U :$M|  �4 ;$@    .M ;	�  �F     	      �� LM ;	&ao  � � ֳ  <	&dX  M E x =	&�  � � 
�I ?	nk     cff @	�O  � � sub A	�T  � � i�U B	�   
��  D	T�  : 6 ;�  o	�F     #�F     a       � 
��  J	h  z t #�F            � 
�  [	�  � � 
�L  \	Y  � �  B�F     Us�&T�Q  U}  AF      �� f	�    �  7 5 �� �  ^ \ =}  CF            �  � � �  � � &CF            1�       ,X> 	`@F     �       �+  LM 	6ao  � � ��  	6�D  #  ֳ  	6dX  ` \ �  	6�X  � � n�  	6?  � � ;:  	6&  . ( �6 	6Ya  ~ | �S 	6�a  � � cff  	�O  � � }  �@F      p� -	� �  	  �  . , p� �  U S =}  �@F            �  z x �  � � &�@F            1�      �@F     �3 Us T�TQ�QR�RX�X�  'C\ ��  }  )cff �.�O  �_ �.�  n ��  ��  ��  ��  �T�   'IU ��  �  X@ ��  ��  ��  �Y  ��   o�l ���E     �       �Q! LM � Vg  � � 
ڰ  �|    .8 ��E      0{ �<! <8 = ; 0{ I8 b `   c�E     g� Uv   .mN ��  `F           ��" LM �)Vg  � � ��  �)�    ֳ  �)�  � � �  �)�  � � �o �)�2  ` V E�  �)�(  � � n�  �)?  Z X ;:  �)&  � ~ ��  �)Di  � � $@� �" 
Q  ��0  � � �� 
ϖ ��    
6e  ��  D @ �F     �� T	׷F     Q1   �F     W8 Us T} Q��R~ X �  .0U ��  ��E     �      �$ 9LM �)Vg  U�. �)3  ~ z ��  �)�  � � 
�y  �Cg  � � ip �3  J 0 
��  �3  m a 
�I �d  � � ;<d ��E     ;��  ��E     T��  ��x top �>'  (  op ���  � � 
<v �H  � �  y 
A�  F�  �  �     }�4 ��  �F     �       ��$ -LM �3�i  ^! V! -�_ �3�  �! �! Rn ��  " " ({ �7  |" v" (Q  ��0  �" �"  � (}W �  # # 'F     �� T}    .%m YU  ��E            �O% Aq Y+/  ?# ;# ��  Z+e#  |# x# 
��  \&4  �# �# 
Q  ]�0  �# �# f��E     U�UT�T  .y= M�  ��E            ��% Aq M,/  	$ $ ��  N,U  F$ B$ 
��  P&4  �$ $ 
Q  Q�0  �$ �$ f��E     U�UT�T  ,�F A��E     (       �K& Aq A&/  �$ �$ 
��  C�  #% !% 
ڰ  D|  I% G% ��E     g�  .)` *�  @�E     6       ��& Aq *&/  y% q% ��  +&�  �% �% 
��  -&4  & & 
ڰ  .|  S& O& 
Q  /�0  �& �& fn�E     T�UR	0�E     X0  .�2 "�  0�E            �=' 9��  ""&4  Ucidx #"�  T G�R �U  ��E     d       ��' -I_ �,�x  �& �& ?��  �,e#  T(�Y  ��  @' .' (��  �U  ( �' ;�  �E      GaM ��  ��E            �( ?I_ �-�x  U-��  �-U  �( �( (�Y  ��  :) 8)  Yea ���E            �A( ?I_ �'�x  U GM/ ��  P�E     %       ��( ?I_ �'�x  U?��  �'�  T(��  �&4  b) ^) (T �(1  �) �)  G�2 ��  �E     1       �P) ?I_ �$[x  U?��  �$�  TC�+ �E      �E     .       ��+ �) �) �+ * * &�E     .       �+ +* '* �+ d* b*    G�: {�  ��E     1       ��) ?I_ {&[x  U?��  |&�  TC�+ ��E      ��E     .       ��+ �* �* �+ �* �* &��E     .       �+ �* �* �+ + +    G�k cU   9F     U       ��* -I_ c'[x  8+ 2+ -��  d'e#  �+ �+ (�Y  f�  , , (��  gU  �, �, p�  tY9F     C�* K9F      K9F     
       l+ =- ;- + b- `- &K9F     
       + �- �- U9F     l� Uv Ts     0�7 ?�  Y+ I_ ?'[x  ��  @'U  �Y  B�  2�* G�  8n G�  { H�  2��  R�     Y�a 5��E             ��+ ?I_ 5![x  U 4�3 #�+ I_ #![x  ZJ $!�  ��  &&4  Q  '�0   '*�  
U  �+ )r 
U   ,կ  
@�E     P       ��, 9_| 
3  U��  
		  �- �- ��  
�  . �- UhS @�E      0x 
�S <. :. �S f. d. �S �. �. �S �. �. zS $/ "/ 0x �S N/ L/ �S w/ q/ �S �/ �/ F�S `x �S 0 0 �S D0 B0     ,��  �	�F     �      ��- ��  �	!�  m0 g0 ��  �	!�&  �0 �0 ��  �	!�T  �0 �0 
��  �	oW  81 41 n �	�  �1 w1 
/� �	�  3 3 #2F     1       �- !��  �	U  �t @�+ F      F            �	3�+ �3 �3   ,��  w	pF     �      ��. �[ w	!�i  �3 �3 9LM x	!a   T�  y	!?  x4 t4 #�F     �       {. 
IM 	Vg  �4 �4 �F     �0 Us Tt Qq   &pF     �       
1 �	ao  �4 �4 zF     �0 Us Tt Qq    /Y %	 / �I %	*�`  Mj  '	-+  ��  (	�  2p1 =	  p2 >	  ��  ?	3    'h 	�  c/ �I 	(�`  )x 	(�  )y 	(�  �U 	�   '>9 ��  �/ �I �(�`  Mj  �-+  �U ��   'Q ��  �/ �I �'�`  )x �'�  )y �'�  �U ��   /�H �H0 �I �&�`  )x �&�  )y �&�  ~� �&h  Mj  �-+  2c �  ��  �3    '�E ��  u0 �I �)�`  /� �)�   ,�0 ���E     D       ��0 9�I �!�`  U
ȩ  ��X  �4 �4  ,|@ Gp F     �       �R1 i G!�`  $5  5 9�I H!a   T9�  I!?  Q$� *1 
�I Od  \5 Z5  &0F     .       
�e hnk  �5 5   ,ME ��E     �       ��1 �I �,nk  �5 �5 
Mj  �-+  )6 #6 
��  ��  |6 v6 �w p1 	  �6 �6 p2 
  )7 #7 
��  3  ~7 z7   '�. ��  72 �I �*nk  )x �*�  )y �*�  �U ��   .�O ��  �F     x       ��2 �I �*nk  �7 �7 
Mj  �-+  8 8 
�U ��  h8 f8 	F     �� T0Q1  'iZ ��  �2 �I �)nk  )x �)�  )y �)�  �U ��   /_8 �]3 �I �(nk  )x �(�  )y �(�  ~� �(h  Mj  �-+  2c �  ��  �3    'RY �  �3 �I #nk  /� �#�   ,OB sp�E     D       ��3 9�I s#nk  U
ȩ  u�X  �8 �8  ,al 1p
F     8      ��4 �I 1$nk  �8 �8 ��  2$�D  9 9 ֳ  3$dX  E9 ?9 ȩ  4$�X  �9 �9 n�  5$?  �9 �9 &�
F     u       
��  @  ":  : #�
F     )       �4 
�  M�  G: E: 
�L  NY  n: j:  �
F     ��   ,�g ���E     �       �m5 �I �)d  �: �: 
Mj  �-+  ,; &; 
��  ��  ; y; �w p1 �  �; �; p2 �  ,< &< 
��  �3  �< }<   '�J ��  �5 �I �'d  )x �'�  )y �'�  �U ��   .2 ��  @F            �+6 �I �'d  �< �< 
Mj  �-+  R= F= 
�U ��  �= �= �F     �� T0Q1  . f ��  `1F     T       �7 �I �&d  > �= 7x �&�  �> z> 7y �&�  ? �> 
�U ��  |? x? 8 r1F       �� ��6  8 �? �? 8 �? �? {1F     u Us T1  �1F     7 Us Tv Q| R1  ,�b u �E     �       �8 �I u%d  @ @ 7x v%�  T@ P@ 7y w%�  �@ �@ ~� x%h  �@ �@ 
Mj  z-+  "A A &3�E     D       
c   nA lA 
��  �3  �A �A P�E     � �7 U�T `�E     � U|    '�h l�  .8 �I l(d  /� m(�   /�@ `W8 �I ` d  ȩ  b�   ,�O '@	F     $      �9 �I '"d  �A �A ��  ("�  !B B ֳ  )"�  `B ZB ȩ  *"�  �B �B n�  +"?  C �B &u	F     \       
��  6  =C ;C �	F     ��   ,W �0�E            �C9 9��  ��Z  U ,^ ���E     �       ��9 9��  ��Z  U9Ǟ  �3  T9��  �3  Q9ڰ  �|  R .�: ��   �E     )       �}: ��  �(�Z  dC `C cY �(�  �C �C 
Q �(   �C �C n�  �(�  GD AD |K  �E      �| �Y: �K �D �D �E     �N Uu Tt   H)�E     xF U�UQ�TR�Q  .{M ��   �E     E      �< ��  �(�Z  �D �D /f �(�  wE sE Ԛ  �(�^  �E �E |K  �E      �~ �"; �K F F $�E     �N Uu Tt   U�G +�E       �~ �H ?F ;F H yF uF �G �F �F �G OG AG �~ "H �G �G /H H 	H <H �H �H GH /I +I _TH ��E     F]H 0 6^H ��kH mI gI ��E     uT �; U��T} Q0 ��E     �N Uu Tt      .{> ��  P F             ��< ��  �"�Z  �I �I n�  �"�  �I �I |K P F      � ��< �K GJ EJ ` F     �N Uu Tt   Hp F     uT U�UQ	�T $ &  .dD ��   �E     s      �b> ��  �"�Z  vJ jJ Vu  �"3  �J �J vT �"		  AK 5K �X �"�?  �K �K 9>W �"?  Xi�U ��   cur �3  gL ]L ;�  �s�E     |K  �E      �v ��= �K �L �L :�E     �N Uu Tt   U�S \�E      w �.T M �L !T �M �M T N N T �N �N w 9T 3O +O DT �O �O OT UP KP ZT �P �P FgT pw hT �Q �Q     .; �   �E            �? ��   �Z  �Q �Q |K  �E       �E     	       ��> �K :R 8R 	�E     �N Uu Tt   H�E     :V U�UTt   .�9 2�  ��E     _      ��@ ��  2/�Z  iR ]R #` 3/�[  �R �R �  4/�  �S �S �  5/�  T T X8 6/�?  �T �T !�K 8�@ ��y
�L 9V[  ,U &U !�K :�  ��y
�U ;�  �U xU 
K�  <3  V V 
��  =3  `V ZV !0X >y]  ��y;�  y��E     &�E     zH U@ U T��yQ R��y ��E     �@ U T��yQv R| X0  �\  �@  L    .` 	�  0�E     e      �!F ��  	)�Z  �V �V #` 
)�[  �V �V �  )�  �W �W �  )�  �W �W X8 )�?  5X 1X !�L �\  ��Xcur 3  ��
��  3  vX nX 
/� �  �X �X idx �  |Z dZ 
�U �  y[ w[ 
b �\  �[ �[ ;WD  (�E     ;5- >`�E     ;�Y i��E     ;�  %	�E     $p~ MB !ӱ  '�\  ��
�N (3  �\ �\ 
��  )3  �\ �\ �E     �I U T��  $} F q L3  �\ �\ val M�  m] e] 
�: N  �] �] $@~ C 
ڰ  �|  �^ �^ len ��  �^ �^ ��E     g� �B U��~ ��E     O� C T ����Q��~ �E     9� Qv   #X�E     f       �C !�S  �!F ��
�;  ��  _ _ 
�Y  ��  >_ <_ r�E     xF �C U��Q4R��X0 ��E     � ��E     � ��E     � ��E     �  $p} EE 
ڰ  �|  g_ a_ 
�S  �   �_ �_ 
�Y  ��  I` E` i ��  �` ` $�} wD 
�;  �  �` �` ��E     � �E     � �E     � *�E     �  Z�E     [� �D U��~T8Q0R��~X0Y��~ ��E     xF �D U��T~ Q} Rs ����3$v "X0 ��E     �N E Uu T~  Q�E     g� (E U��~Tv  e�E     g� U��~Tv   1F �E      �} V�E PF CF (a "a �} ]F wa qa jF �a �a   ��E     �N �E Uu Tt  ��E     :V �E U�� w�E     uT �E U��Q3 4�E     uT U��Q0  `�E     �I U��~T��  �  1F  L    '/1 �S   xF �O ��2  ��  �3  cur �3  �Y  �?   .xe ]�  ��E     ]      ��G �O ]�2  6b (b ��  ^3  �b �b cY _�  Fc 8c 
Q `   �c �c n�  a�  �d �d cur c3  �d �d 
/� d�  e �d c eh  f f 
Ku  eh  wf sf ;�  ���E     �| !��  {�  ��
�N |3  �f �f K�E     uT �G U��Ts Q��� $ & ��E     �N Uu Tt    '�Y �  zH �O �2  ��  3  /f �  Ԛ  �^  cur 3  /� �  c h  Ku  h  T�  P2��  +�  �N ,3    ,�l � �E     �       ��I ��  �(�Z  
g �f �X �(V[  �g �g 0c �(�  ,h &h �X �(M_  �h xh !�  ��\  ��$pv �I 
K�  �3  i i 
��  �3  ei ]i cur �V[  �i �i 
��  �V[  j j �v !�L ��\  ����E     �I U| T��   )�E     �I U| T��  ,�[ r0�E     �      �|K ��  r"�Z  |j tj �L s"V[  �j �j cur u3  Dk Bk 
��  v3  ok gk 
-G w�  �k �k |K V�E      V�E     	       �J �K 4l 2l _�E     �N Uu Tt   |K e�E      0v ��J �K Yl Wl o�E     �N Us Tt   |K ��E      ��E            �	K �K ~l |l ��E     �N Us Tt   ��E     �K +K Us  ��E     ;N IK Uu Tt  8�E     �L gK U�PT|  ��E     �K Us   /�6 h�K ��  h%�Z   ,�L ��E     /      ��L ��  '�Z  �l �l Xcur 3  �`
��  3  ?m 5m 
�U �  �m �m ;�  S��E     �E     �N 5L Uu Ts  ��E     �M SL U�`Ts  ��E     �L qL U�`Ts  ��E     ;N Uu Tt   .: ��  ��E     $      ��M �O ��2  �n �n ��  �3  Mo Co cur �3  �o �o 
-G ��  �o �o 
�U ��  �p �p ~end �Z�E     O ��E     '       �	pM �O �O &��E     '       �O vq tq   �E     ;N �M Uu Tt  }�E     �M U�hTz   .�b ��  P�E     c       �;N �O ��2  �q �q ��  �3  �q �q cur �3  $r "r err ��  Kr Gr {�E     �N Uu Tt   .a: W�  `�E     �       ��N 9�O W#�2  U9��  X#3  Tcur Z3  �r �r 
-G [�  s �r 
�U \�  �s �s i ]Z   �s �s �u c bh  Ot Et   ,�Y 9��E     c       �O 9�O 9�2  U9��  :3  Tcur <3  �t �t �O $�E     "       E�O �O &$�E     "       �O u �t    /�b '�O �O '�2  ��  (3  cur *3   ,L1 ��E     f       �CP �B �Y  ?u 9u 
ڰ  |  �u �u ��E     g� P Uv  ��E     g� .P Uv  ��E     g� Uv   Y�; ���E     �       �xQ -�B ��Y  �u �u (ڰ  �|  2v 0v b�U ��  �\(�O �3  \v Vv .R �E      �E     8       'Q GR �v �v ;R �v �v &�E     8       SR �v �v _R w w kR <w :w   ��E     O� EQ Uv Q�\ �E     9� ]Q T|  j�E     g� Uv T|   0�7 ��  �Q �B ��Y  :idx ��  ��  ��  ��  ��  2�U ��  v  �		  / �	    0�B y�  .R �B y#�Y  v  z#		  ڰ  ||  �O }3  �U ~�   4#j hxR �B h�Y  �O i3  �� k	  �  l�2  ��  m�2   G�- J�  ��E     �       �hS -�B J�Y  kw _w -/� K�  �w �w -ڰ  L|  Qx Ex b�U N�  �Le�  _!�E     [�  S Uv T8Q0R| X0Y�L 8�E     g� 8S Uv  j�E     [� Uv T4Q0R| X0Y�L  ' ? .�  �S O�  .$�2  ��  /$3  _| 0$3  )n 1$		  ��  2$1  p 43  r 5�  s 6�  2val E�  b F�    'D ��  uT O�  �&�2  ��  �&3  _| �&3  )n �&		  p �3  r ��  w ��  pad ��  2c ��    G�L ��  ��E           �:V -O�  ��2  �x �x -��  �3  ,z z -n�  ��  �{ o{ qp �3  ��( 1 �3  �| �| (][ ��  } �| (,B ��  �~ �~ (d ��  � � (�} �?  G� 9� (��  �?  � � (�7 �?  �  � �Bad a;��  e��E     ;��  js�E     ;�  [��E     $0| �U Rc �P  ă ��  $ |  V 
o�  �  � � ��E     :V U��Tt   ��E     :V V U��Tt  T�E     ,� Uv T|   GXR ��  ��E     p       ��V -O�  ��2  Q� G� ?��  �3  Tqp �3  �X( 1 �3  ̄ Ƅ Rnum ��  � � ��E     �V �V Uu Tt Q: ��E     �V Uu   G�C T�  �E     f      ��W ?O�  T�2  U?��  U3  T-Ǟ  V�  [� O� Rp X3  � ݅ Rnum Z�  w� k� (�} [?  
� �� (��  \?  �� �� (.i ^�  3� -� (��  _P  �� |� �Bad �B�E     �u Rc }P  �� ��   .�i ^�  �9F     h      ��_ ��  ^!�o  � � 
ڰ  `|  �� �� fi a4  �� �� 
�U b�  � �� key c�   �� �� Xlen d		  ��~
�J e�  5� /� ;WD  ��:F     $@� )_ !> r�_ ��~$�� Z n ��  �� �� ^b �;F      �;F     (       �RY }b �� �� pb ԋ ҋ &�;F     (       6�b ��~�;F     �d Us T��~Q1   U�_ �;F      � ��_ �� �� �_ #� � �_ r� p� 0� �_ �� �� 6�_ ��~E�_ [�_  <F            �Y �_ � � -<F     �c  
<F     ]� Z Us T0 L<F     ]� Us T��~    �` �� �^  ` �� -` � 	� :` ^� \� 6G` ��~ET` �a �:F       � "�[ �a �� ��  � �a ؍ Ѝ �a >� :� �a x� v� 6�a ��~�a �� �� b 5� 1� Eb ^b �:F      P� V
D[ }b o� k� pb �� �� P� 6�b ��~�:F     �d Us T��~Q1   K>b �� �[ 6?b ��~+>F     �c �>F     �d Us T��~Q5  [b ?F     5       �[ #b � � 60b ��~-?F     [� T(Q0X0Y��~  >F     ]� Us T��~   ^` 8=F      �� )�] p` � � �� }` f� ^� �` ΐ Ȑ �` � � 6�` ��~�` ]� U� �` �� �� E�` ^b V=F      � �
�\ }b �� �� pb #� !� � 6�b ��~[=F     �d Us T��~Q1   K�` @� s] �` R� F� K�` �� 9] �` ޒ ؒ 6
a ��~�?F     �d Us T��~Q4  �=F     �c C@F     �� T|  $ &Q@R	��E       [�` I?F     5       �] �` )� '� 6�` ��~b?F     [� T@Q0X0Y��~  �=F     ]� Us T��~   �;F     ]� ^ Us T��~ �;F     �c   ^b �<F      �<F     #       x�^ }b O� M� pb y� w� &�<F     #       6�b ��~=F     �d Us T��~Q1   z:F     �c :;F     �d �^ Us T��~Q1 j;F     �d �^ Us T��~Q1 z<F     �d _ Us T��~Q1 �<F     �d Us T��~Q4  $:F     ]� H_ Us T��~ h:F     ]� g_ Us T��~ �:F     g� _ U}  �:F     g� U}   ks  �_  L    '�U @�  ` ��  @(�o  )n A(�  �9 B(�w  key D�   len E		  TWD  X2�L Q�w    '�; �  ^` ��  $�o  �U �  key �   len 		  TWD  : 'U9 ��  a ��  �%�o  fi �4  kp ��3  key ��   len �		  n �S   tmp ��  TWD  ^�` ڰ  �|  �U ��   2�L ��w  2r ��  > ��_    .k? �S   ��E     )       ��a ca �(�  Ucb �(�  Tkp1 ��3  �� �� kp2 ��3  Ó �� 
v�  ��  � � 
}�  ��  � �  '%L L�  Nb ��  L%�o  fi N4  tk O<3  key P�   len Q		  n RS   tmp S�  TWD  �^>b ڰ  `|  �U a�   2> jNb   ks  ^b  L    '�> 8�  �b ��  8$�o  �- 9$M_  val ;ks   ,UW .��E            ��b ��  . �o  b� \� 
ڰ  0|  �� �� ��E     g�  .�T �  ��E     g       ��c ��   �o  ڔ Ԕ ڰ   |  ,� &� Ǟ   3  ~� x� ��   3  Е ʕ 
^�  �p  "� � !�U �  �L��E     O� Uv T Q�L  .�\ ��w  �F     �       �'d 7key ��  r� l� 7len �		  Ė �� n �
S   � � �F     Ʉ T| Q}   '�b ��   {d ��  �$�o  � �$?  )len �${d ^�  ��p  key ��    		  .g t�  pF     {      �#f ��  t%�o  �� �� $g u%ws  �� � 7n v%�  8� 0� 
^�  x�p  �� �� Xstr y�   ��i z�  +� %� p� len �		  �� t� val �ws  �� �� #xF     B       �e 
ڰ  �|  � ߚ !�U ��  ���F     Մ �e T Q�� �F     9� Q��  �F     #f F     :V �e U��Tt  /F     �f ]ZF     f T pF     uT U��Q0   G�: ��    F     h       ��f -^�  �'�p  � � Rstr ��   B� >� $0� �f Rch �S   |� x�  L�g  F       � ��g �� ��  � `�g  F     i Uu     G�3 z�   �F     x       ��g -^�  z$�p  ߛ כ Rstr |�   ?� ;� $�� 6g Rch �S   {� u�  C�g �F      �F            �g ͜ ˜ &�F            `�g  �F     i Uu     0�Y ^S   �g ^�  ^'�p  8ch `
S    0VJ  �H  �g :a �H  :b �H  8ret �.  8tmp �.   *|K  �E     	       �7h >�K UH)�E     �N Uu Tt   *.8 @�E     D       �gh ><8 UI8 � �  *�2 ��E     H       ��h 3 � � 3 V� R� 3 �� �� >&3 R33 Ν ̝ &��E     -       A3 � � N3 � �   *�+ ��E            �i �+ E� ;�  *�g F     c       �Ci >�g U�g �� ��  *�. �F     �       ��i �. �. �� ޞ �. 	� � F�. �� �. Y� S� / �� �� / � �   *,�   F     �       �l :�  U� Q� G�  �� �� a�  � ݠ >l�  YT�  T�  w�   � � �g F       � �ej �g z� v� �g �� �� � �g ߡ ۡ �g "� �   �g 7F      �� ��j �g _� ]� �g �� �� �� �g �� �� �g � �   �g eF      @� �	k �g �g .� ,� @� �g W� S� �g �� ��   �g |F      �� �_k �g ף գ �g �� �� �� �g %� !� �g h� d�   �g �F      � ��k �g �g � �g �� �� �g � �   �g �F      p� ��k �g '� %� �g p� �g N� J� �g �� ��   ]F     C�  Uu Ty   *(�  �F            �nl >9�  UC� �F       �F            b Υ ̥  �� �   *R�  �F            ��l >_�  Uk�  � � C� �F       �F            p D� B�  k� i�   *R�  �F     2       �m >_�  U>k�  THF     nl 5k�  t   *,�  F     5       �Wm >9�  U>E�  TfEF     5E�  t   *��  PF     `       ��m >�  U=�  �F            �  �� �� C� �F       �F            �\ � �� ��    *Ə  �F     `       ��n >׏  U�  ަ ئ <x�  �F       �F            �Cn ��  ,� *� ��  ,� *�  =Ə  �F            �  Q� O� ׏  v� t� C� �F       �F            �\ � �� ��    *n�   F     >       ��o >{�  U��  ħ �� <x�   F        F            �o ��  � � ��  � �  =n�  8 F            ��  7� 5� {�  \� Z� C� < F       < F            �\ � �� �    *� P F     Q       �p � �� �� � � � F� �� � x� r� �� 1� F� �� � Ʃ ĩ m F     g� p Uv  � F     g� Uv      *xQ � F     �      � r �Q �� � �Q �� �� �Q 4� &� �Q ݫ ϫ FxQ  � �Q �� {� �Q � � �Q �� �� �Q K�Q `� r �Q �� � �Q 7� -� �Q �� �� L�Q H!F      �� ��Q N� H� �Q �� �� �� 	R � � R X� P� 6!R ��<.R �!F      �!F     8       ��q GR �� �� ;R ܰ ڰ &�!F     8       SR � �� _R &� $� kR M� I�   U!F     O� �q U��Ts Q�� �!F     9� �q T~  �!F     g� U��T~      "F     9� T Q}    *��  �"F     �       ��s ��  �� �� ��  � � �  �� �� �  � ݲ >"�  � ��  ��  /�  J� D� :�  �� �� G�  �� �� T�  P� L� _a�  #F     x�  �"F       � !�r ��  �� �� ��  � �  Kj�  @� `s 6k�  ���"F     Ə  ,s Uu Ts  �"F     Ə  Ds Ts #F     � U~ T��  �  #F      #F     
       F�s �  �� ~� �  �� ~�  ��  C#F       C#F            ,�s ��  �� ��  @#F     Ə  Uu T0  *\�  �(F     j       ��t {�  ε ȵ ��  $� � n�  6��  �`��  �� �� ��  � � ��  %� !� ��  g� a� [��  !)F            �t ��  �� �� ��  ݷ ۷  B)F     T�TQw   *��  `)F     i       �u ��  � � |)F     �  �t Us  �)F     $�  Us TsQs��Y1  *8 1F     '       �du 8 s� o�  8 �� �� H71F     �� Q0  *8 @1F            ��u 8 � �  8 A� ;� HF1F     u U�UT�T  *m5 �1F     J       �~v 5 �� �� �5 -� !� �5 �� �� `�5 Fm5 �� �5 S� I� �5 һ Ȼ 5 Q� G� �� �5 ȼ Ƽ �1F     �5 Xv Us  H
2F     +6 U�UT�TQ�Q    *H0 2F     '       ��v g0 � � Z0 H72F     �� Q0  *�/ @2F     <       ��w �/ ,� (� �/ i� e� �/ �� �� 1�/ @�/ @2F      @2F     ;       �\0 0 � ߽ �/  � � �/ ]� Y� &@2F     ;       0 �� �� =+0 O2F     %       ,0 �� �� 90 � �     * / �2F     �       �Ey 2/ � � ?/ �� �� J/ � � U/ �� �� c/ �2F       � 	Wx u/ �� ��  � �/ v� n� �/ �� �� <3F     �� T0Q1   @�/ �2F      �2F     (       	�/ �� �� �/ � � �/ D� B� &�2F     (       �/ k� g� H0 �2F      �2F            �"y Z0 �� �� g0 �� �� �2F     ~v UsT15Z0 s   3F     �v Us T| Q}     *]3 �4F     '       ��y o3 �� �� |3 .� *� H�4F     �� Q0  *]3 �4F            ��y o3 m� g� |3 �� �� H�4F     Ey U�UT�T  *�2  5F     d       �z{ �2 � � �2 c� ]� �2 �� �� �2 � � ]3 5F       �� �~z |3 (� &� o3 P� L� 5F     Ey U| T1  =�2 5F     D       �2 �� �� �2 �� �� �2 �  � &5F     D       1�2 @�2 5F      5F     D       �&3 '� %� 3 O� K� 3 �� �� 3 �� �� &5F     D       33 �� �� =�h 05F     (       A3 � � N3 6� 4�       *�1 p5F     J       �B| 2 e� Y� 2 �� �� 2 �� �� `)2  F�1 �� 2 � � 2 �� �� 2 � � �� )2 �� �� �5F     72 | Us  H�5F     �2 U�UT�TQ�Q    *� �5F     �      �l� � �� �� � &� � � �� �� � �� �� � u� k� � �� �� >� � � ]� Q� � �� {�  �� �� _ �6F     _ z7F     _' �7F     =/ 6F     u      0 �� �� ;  � � F �� �� Q 6� ,� \ �� �� g D� :� r �� �� } F� <� N�g *6F       � ��} �g �g  � �g �� �� �g � �   [� �6F     p       q~ � ^� Z� 1� � �� �� �6F     ,� ~ Tv  �6F     s� L~ U}  $ &T~  $ &Q��� $ & 	7F     ,� Uw �@$ $ &Tv   N�g 07F      �� ��~ �g � � �g 3� 1� �� �g \� V� �g �� ��   [� z7F     V       c � � � 1� � F� B� �7F     ,�  Tv  �7F     s� B U}  $ &Q
w � $ & �7F     ,� U~  $ &Tv   [� �7F     �       � � �� �� � �� �� � *� &� 8F     ,� � Tv  Z8F     s� � U}  $ &Q��� $ & p8F     ,� Uw �@$ $ &Tv   &7F     ,� -� T
s 1$ $ & f7F     ,� E� Tv  �7F     ,� U���@$ $ &Tv    ��* �8F     }       �� + �� �� + �� �� `+  F&+ �� '+ -� +� 3+ l� d� =+ �� �� FI+ � J+ � � �8F     �� T~     *�*  9F            �]� + G� A� + �� �� `+  H9F     l� U�UT�T  *'d �9F     b       �߁ 9d �� �� Sd &� "� `d ^� \� md �� �� \Fd �9F     #f ʁ Ux  �9F     �f Ux   *��  0AF     �       �>� ��  � �� ��  l� d� ��  �� �� 1��  N��  0AF      �� �
�� �  $�  � 	�  ^� Z� =��  �AF            �  �� �� 	�  �� �� C� �AF       �AF            r\  �� ��    =��  TAF     G       ��  ��  ��  &TAF     G       ��  � � L(�  zAF      Ж �$9�  B� >� �AF     l Ut      *�  @BF     X       ��� >�  U<� TBF       TBF            ���  z� x�  �� ��  =�  �BF            �  �� �� C� �BF       �BF            �\ � �� ��    I�o  �o  "~IO\  O\  �g�s  �s  7I:V  :V  �g\P  \P  rBY  8Y  ? rD  D  ? I�`  �`  @vI�I  �I  @�I�s  �s  @�ge  e  �I�W  �W  `I�>  �>  �g�b  �b  8I�  �  AI�?  �?  eI�  �  BXI��  ��  AI�U  �U  @{ �5   2�  &  �n �:  p�F     H      � ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  	)  �  	5  s&  G   �  N   	N  )  A"l  r  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  `  -    �   m�  �  �  `  U    f  �    U   ,  `  -   -   U    J   �"8  >  �  PH�  Ǟ  J;   ֳ  K@   pos L@     N�  /[  O�   �K P  (�R QM  0ڰ  S`  8O�  T;  @��  U;  H �  ��  <v �-   ��  �U    �  ��  ""  �    @   ;  ,  @   ;  @    A  �  	A  �   Z  `  k  ,   v  :-   �  L�  x Nk   y Ok   �  Qw  	�  ~   w�  
  yk   �!  yk  �   zk  H  zk   "  |�  �  (y  M} N    5�  N   `�  	G   _| 
;  
!  5  ?   A  2   A  B  U     �  �  	y  �  (Q�     S)   0�  T)  N5  V�  �   W�   H� X�  �1  ZG     �  )  �  \�  �  �  N   �K  �!   �   pmoc�  stibu!  ltuo�  tolp :  �  �8  5"e  k  �$  �4  S�  x U)   len V5  e� WA   �#  Yp  	�  �%  {�  �  �  G   G   �  U    �  �#  ��  �  G     G   G   U    �.  �%  +  @  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(  �  (�/    0�  U   8*  �  @ �  �  u(  
@  	�  �2  (�  �  G     U      X  �3  ;&  ,  7  X   v)  ]D  J  _  X  ;  @    �3  yl  r  G   �  X  @   U    H7  ��  �  G   �  X  �   �  51  0�  y2  �K   � ��   �7  *
 �_  / ��   $ �  ( 2$  ��  -4  lA  +  �@  �  $8  �A  	G  S    ��   	^  {"  �)  !  �5  \   �G   	�  �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U    :   �&	  xx ��   xy ��  yx ��  yy ��   5  ��  	&	  8  �c	  ��  �X   ��  ��   $  �8	  c   �}	  �	  �	  U    �  ��	  Kl  �U    �  �p	   s  ��	  �"  $�	  �	  �   +
  �� -�	   �W .�	  Kl  /U    %  D=
  uR F�	   �
 G�	   }  I
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @	<  5�  	>k   ��  	?k  �"  	Ak  �"  	Bk  i!  	Ck   %!  	Ek  (2!  	Fk  0�  	Gk  8   	I�  �"   	sn  ��  	uo   5�  	vo  ֳ  	xk  !  	zk  m  	{k   v  	}  J  	�#�  �  �!  �
}L  ڰ  
`   {3  
��  S0  
��  �/  
��  �1  
��  �1  
��#  Y/  
�=
  �*  
��  (�)  
�L  0+:  
�$  8<8  
�$  X�*  
��  � �3  	�"Y  _  �(  
��  Oe 
��#   �-  
�{  ڰ  
�`   U  	�"�  �  �  8
�  ah 
!�#   Oe 
"r  U1  
#=
   ;+  
$�  0 i(  	�$�    l;  �
�v  ah 
��#   Oe 
��#  y2  
�K   {:  
��  (�� 
�X  h/ 
��  p�� 
��  x T   	� �  �  _  �	J  �!  	�   �  	�  �  	�    	�  �  	�   �U 	�  (�  	�  03"  	�  8�  	�  @`  	!�  Hd  	"�  P�@  	$�	  X�;  	)�  h�   	+{  ��  	,o  �
  	-o  ���  	.o  �?!  	0o  ��  	1o  ��  	3o  ��  	4o  �ȩ  	6�  �ֳ  	7J  ��� 	8  �K 	<�  �ڰ  	=`  �^�  	>,  �U  	@=
  �t  	B�	  �k  	CU   ��L  	E:  � "  	 W  ]  1  X	m�  ��  	ov   �@  	p�	  �e 	q�  �L  	r�  P @  	$%�  �    0	\  �-  	^{   ��  	_v  �W 	`�  x 	a�  �@  	b�	   �e 	d  0�"  	e�  pi"  	f�  x� 	g�  ���  	iK  �.a 	ky  ��  	l�  �J  	m�  �Mj  	o�  ��  	q�  ��  	r�  �M  	tU    Z  	u-   _"  	wk  (   	xk  Ud 	zU    �L  	|  ( �!  	F#    Z!  	A[  ��  	Cv   T 	D   �!  	E{  "  	F{   S  N   	�   Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  	[  �C  	H  0  	`)G  M  �"  �
e�  �1  
g&	   H+  
h�   x+  
i�  0��  
k    8�)  
n#�!  h�'  
q4  p��  
rA  t�*  
y�  x ^  n    �  	�)�  �  �!  H
�*  $  
�U    7:  
��  s4  
��   b  8	H�  !  	J{   m  	K{  A� 	M�  �� 	N�  �  	Pk  
  	Qk   ��  	Rk  (�  	Sk  0 �  	U*  x   	�$�  �  �!  0'  ad  )�   �1  *{  &D  +�  2B  ,�  x� -&	     	�)%  +  �"  P
��  ��  
��   �1  
��  �&  
�(  �3  
�&	  ]7  
��  0�7  
�U   @�1  
�A  H P6  	�  tag 	�   Kl  	�   �6  		�  �  �5  N   	
  i7   �&  9  F9  8%  �*   �,  	
�  ./   	6
t  b 	8
   5�  	9
�  ��  	:
�  5  	;
�  Q(  	<
�    -  	I
(�    �8  N   	��  �:   4,  �6  $  �/  l9   �2  	��  �#  ��  �'  ��  �  �  �  L   �2  �      L   l/  �"  (  �  <  L  <   �   ;)  H��  �#  ��   :  ��  �5  ��  F1  ��  ,8  ��   2*  ��  (�*  ��  0`1  ��  8��  �  @ j  �-  �B  	�  d)  s�  �  �  �  U    9  F#  	�  �$  @J�  �#  L�   y2  MK  W� O�  �� P  �,  Qw   M4  R"  (�;  SO  0�*  T�  8 c/  X!�  �  �-  (q�  �-  s{   Oe t�  ��  uK  � v�   
  �/  )�  �  �    �  �   g%  .    "  �   �.  1.  4  I  �  I     3	  73  6[  a  q  �  q   �  �8  :�  �  �  �  �  �   "3  >�  $)  Y�  �  �  �  �  �  �     �6  _�  �  �  	  �  �  I     �3  f    0  �  �  q   ;0  l<  B  �  [  �  �  �   �&  x��  ah � �   y2  � K  H�8  � �  P�8  � �  X�'  � 	  `� � 0  h�9  � �  p   �.  �[  "9  H2%  Mj  4�   H5  5�  (�)  6�  0�  7�  8�  8�  @ �0  :�  T%  �=�  ڰ  ?`   �0  @�  q5  A�  L)  B�  )  C(  Ǟ  E%  �  F%  `Ud HU   � X+  J�  1  1  �  �  �  �  ,  v  �  �  �   �&  &�       v   �1  *    �  ,  J   �6  -8  >  I  J   w-  1U  [  �  j  �   �;  4v  |  �  �   =;  8�  �  �  �  J  t   B$  <�  �  �  �  J  �   2  @�  �  �    �  J  �  A   7  G    �  3  v  �  �  �   q8  N?  E  �  Y  v  ,   )2  Se  k  �  �  v  �  �  A  �   �  k.  ��r  ah ��   #,  ��  H�4  ��  P,;  ��  XEY ��  `/q ��  hZ)  �  p�#  �,  x'0  �I  �.  �j  ���  ��  �� �  �`9  �3  ���  �Y  �5  ��  �U#  ��  � �2  �~  �  8S  ��  �d  �<   �W  ��   C  ��  	�  �&  0�    y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��  *  V'9   ?   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |D   �'  ��   �   �  �   -   �  �    c	  �9  ��   �   �   -   �    A2  ��   �   �  !  -   �  (  !   �   8(  T!  ��  )�    $�  )�   �-  )�    )  !  	T!  3  <�!  �� >%�!   ��  ?%-    a!  #  Af!  �!  �U  
�,�!  �!  �B  
��!  �� 
�-   Oe 
��!   fP  
�,�!  �"  4I  P
��"  ֳ  
��   �� 
��"  �q 
��"  R` 
��"  �W 
� #   P 
�#,#  (�U  
�#\#  0�v  
�#�#  8�v  
�#�#  @�J  
�#�#  H 	�!  ��  
��!  wq  
��"  �"  �  �"  �!  �   �J  
��"  �"  �"  �!   �\  
��"  �"  �   #  �!  N   \  
�#  #  �  &#  �!  &#   N  U  
�8#  >#  �  \#  �!  �!  N  N   �O  
�h#  n#  �  �#  �!  N  N   �n  
��#  �#  &#  �#  �!  `   ;O  
��#  �#  &#  �#  �!  `  N   -k  
��#  �  �(  
�_  �  L  $  @    �  $  @    �  -$  @    H'  
�%  N�  #F$  L$  N  [$  <   :�  )g$  m$  <  |$  �   8�  /g$  �  5�$  V 7N   x 8�   ��  :�$  ��  =$�$  �$  ��  (?%  I_ A�"   J�  B�  �m C%    �$  f�  M%  %  <  /%  �  �   �  U;%  A%  Q%  �  <   ��  Y]%  c%  �  �%  `  �$  �  	%  /%  �   r�  a�%  �%  �  �%  �$  N   ��  e�%  �%  N  �%  �$  &#   �t i�%  	�%  ��  @i^&  4v k :$   �y m Q%  v n �%  Ty o �%  hn q [$   S�  r |$  (��  s ^&  0��  t ^&  8 <  
�/  �  �   �&   @   o 	p&  
�o �&  0  �&   @    	�&  �r ��&  0  �&   @   � 	�&  �o ��&  <  �&  @   � 	�&  �n )�&  Ez J�&  H  '   @   �� 	'  n u'  !�&  	�yH     !�&  	�wH     !�&  	�tH     !�&  	�rH     !�&  	�pH     !'  	��G     N   ��)  6s  �p wm �s Jq �u fq �m qu �r 	Bv 
q �x Qu �v ^v z tz �o �p `t �s  t !�z "�w #�t $0o %�u &$z '/y (�v 0�m 1r @�s A1w QTr R;x S�x T�s Uw V@t W�q X�z `�t apy btr cXz p�t ��y �Es �[p �is �v ��q ��y ��z �o �?m �wx �wn �.r �Pw �x �y ��n ��s ��x ��r ��v �jw ��m ��q �v �up �Bn �0u �t �)n �[x �jo �p �Po �s �u ��x ��w ��o ��r ��q ��p ��p �9p �}o ��r � [  �)  @   	 	�)  "2q ��)  	��G     �   *  @   T 	�)  "�o �*  	 �G     �  -*  @   	 	*  "�u �-*  	��G     #�m �%  	��G     �  o*  @    	_*  #]m Bo*  	��G     $d&  Z	 �G     %�u I�  @�F     
       �+  &ϖ I%L  � � &�E  J%<  O� K� 'J�F     e5  (U	��G     (T�T  %�y <  �F     #       �@+  )sid %�  U %an 
<  ��F            �y+  &�  
#�  �� ��  %Qy �N  @�F     �       �k,  &�B �'�$  �� �� *V �'&#  T+�Y  ��  � �� +��  �N  q� e� ,�   �F     - � .min ��  � �� .max ��  Y� O� .mid ��  �� �� .map �%  4� ,� +Oq �N  �� ��   %�u ��  ��F     �       �"-  &�B �(�$  �� �� *V �(N  T.min �%  � � .max �%  G� A� .mid �%  �� �� +�Y  �#%  �� �� -� +Oq �N  N� J�   %�y ;�   �F     �      � 0  &ڰ  ;+`  �� �� &�B <+�$  �� �� &�  =+�  G� =� &Y�  >+	%  �� �� &r ?+/%  �� �� &)�  @+�  <� 4� #�U B�  ��~#�y D 0  ��~#.x E 0  ��/� �/  .n N�  �� �� +/� O�  � � .map P%  K� ;� +gy QN  �� �� / � V/  +��  X<  9� 3� 0J0  P� ]�.  10  1r0  1e0  1X0  -P� 2�0  �� �� 3�F     r5  (T    00  �� c�.  1+0  10  -�� 280  �� ��   4��F     ��~
/  (U} (Ts  5�F     )1  "/  (U  4�F     ��~A/  (U} (T  3�F     )1  (U   5��F     ~5  �/  (Ts (Q8(R	p�F      5]�F     �5  �/  (U��~ 3��F     �5  (U��~(T8(Q��~(Rs (Y��~  3��F     �5  (U��~(T8(Q0(R��~(X0(Y��~  �  0  @   	 6�w &D0  7gy &,N  7�y ',D0  8n )�   �  6�z �0  7��  +<  7ȩ  +�  7.x +D0  7�y +D0  8n �   9�m �G   p�F     7       �)1  :a �"�  V� R� ;b �"�  T<(q �%  �� �� <-q �%  �� �� <�t �N  �� �� <�v �N   � �  91v >N  ��F           ��3  ={ >"<  �� �� >��F     V       �1  </� L�  ,� (� <<v MN  p� j� ?p N<  �� �� -�� ?c S�   � � ?d TN   b� \�   /@� G2  </� x�  �� �� <<v yN  2� *� ?p z<  �� �� -�� ?c �   �� �� ?d �N   O� G�   -д ?p �<  �� �� ?dot �<  �� �� @�3  �F     � �3  A�3  %� #� A�3  L� H� -� 2�3  �� �� B�3  B�3  B�3  24  �� �� C4  ��F     D4  D$4  3 �F     x4  (U�U(Tt    E�3  (�F            �A�3  �� �� A�3  � �� F(�F            2�3  =� ;� B�3  B�3  B�3  24  c� a� C4  -�F     D4  D$4  3-�F     x4  (U�U(Tt      G�w /@   r4  7}W /*<  7��  0*<  8c 2G   H/� 3G   8min 3"G   8max 3'G   8p 4r4  I`s �Ics WInm �JW4  8mid CG   8q Dr4  8c2 EG    KH�  wG   8q xr4    H  L�3  P�F     �      �e5  A�3  �� �� M�3  T2�3  F� :� 2�3  �� �� 2�3  �� �� 2�3  @� 4� 24  �� �� C4  ނF     D4  D$4  N-4  �� 45  224  � � 2?4  �� �� 2J4  �� ��  OW4  h�F     _       2X4  �  � 2e4  b� \�   PF>  F>  kQ�  �  Q�  �  XQ�s  �s  �Q�I  �I  � �   ��  &  /{ �:  ��F     �      �� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  )  A"C  I  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  7  -    �   m�  �  �  7  U    f  ��  �  U     7  -   -   U    J   �"    �  PH�  Ǟ  J   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q  0ڰ  S7  8O�  T  @��  U  H �  ��  <v �-   ��  �U    �  ��  ""  ��  �  @       @     @      �  �   ,  2  =     v  :-   ~   w�  
  y=   �!  y=  �   z=  H  z=   "  |I  �  (  M} N    5�  N   `�  	G   _| 
  
!  0  ?     2     B  U     �  �  	  �  N   �f  �!   �   pmoc�  stibu!  ltuo�  tolp :  �(  �8  5"�  �  �$  �4  S�  x U)   len V0  e� W   �#  Y�  	�  �%  {�  �    G   G     U    �  �#  �    G   3  G   G   U    �.  �@  F  [  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(    (�/  3  0�  U   8*  �  @ #  �  u(  
[  	�  �2  (    G   .  U   .   s  �3  ;A  G  R  s   v)  ]_  e  z  s    @    �3  y�  �  G   �  s  @   U    H7  ��  �  G   �  s  �     51  0�6  y2  �f   � �   �R  *
 �z  / ��   $ �4  ( 2$  ��  �  c,  +G   N   	��	  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �   H'  �%6  b8  D��F            ��	  ڰ  D7  �� �� ��F     �  U�U  �:  ,7  @�F     7       �D
   ڰ  .7  �� �� !N�F     �  U   "5Q  �J  ��F     �       �9  #^�  �   %� � #+[  � �	  �� �� $g9  �  � � %ʈF     �  �
  U�TT	0�H      %�F     �  �
  Uv T0Q2 %�F     �    Uv  %�F     �  $  Uv T0Q0 !(�F     �  Uv   &�{ �@   ��F     V       ��  #^�  �&  m� c� #�  �&@   �� �� #_| �&  o� a� #/� �&@   � � $g9  �  �� �� '&�F     �  �  U�QT1Q�R !:�F     �  U| Q0  ({ ���F     &       �>  #^�  �$  � �� )͇F     �   (�{ �`�F            ��  #ڰ  �7  R� N� #*�  �U   �� �� h�F     �  U�T  &w{ iU   p�F            �)  #ڰ  i7  �� �� #wO  j-   	    #v  k-   F  B  #*�  lU   �    {�F     �  U�RT�Q  &�{ GU   P�F            ��  #ڰ  G7  �  �  #ֳ  H-   �  �  X�F     �  U�T  *<h <h @*{ { A*�{ �{ [*){ ){ �*�{ �{ �*�{ �{ Y*�{ �{ �*�I  �I  B �   M�  &  �{ �:  ��F     A       �� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  �   �  8"U   	+  K  �   	%  L  	�  M  '  ;  �  �  �  \   �G   
o 6
 -&| $�  ��F            ��  idx $C  U �   | C  ��F            �
�{ X  ��F            � �6   J�  &  �| �:  ��F     �      3� ,  i   �@   �  int �  �   @�   �  �    p   	4   �  #	4   X  &	4   �  )	4    �  ,	4   (�  -	4   0/  2G   8�  5G   < �   �  	�   �  8"W   
+  K  �   
%  L  
�  M  '  ;  �  s&  G   )  A"P  V  �   ��  �  �U    ��  ��  <h ��  �I  ��   �  X�  �  U   �  D  -    �   m�  �  �  D  U    f  ��  �  U     D  -   -   U    J   �"  "  �  PH�  Ǟ  J   ֳ  K@   pos L@     N�  /[  O�   �K P�  (�R Q,  0ڰ  SD  8O�  T  @��  U  H �  ��  <v �-   ��  �U    �  ��  ""  ��    @       @     @    %  �  �   9  ?  J     v  :-   �  Lz  x NJ   y OJ   �  QV  	z  ~   w�  
  yJ   �!  yJ  �   zJ  H  zJ   "  |�  N`  N   �"  �T   jt  �C  �H  �H  �K  RR  Zs  WO   �  (�  M} N    5�  N   `�  	G   _| 
  
!  0  ?   %  2   %  B  U     �  "  	�  �  (Q     S)   0�  T)  N5  V  �   W�   H� X  �1  ZG     z  )  �  \�  �  �  N   �s  �!   �   pmoc�  stibu!  ltuo�  tolp :  �5  �8  5"�  �  �$  �4  S�  x U)   len V0  e� W%   �#  Y�  	�  �%  {�  �    G   G     U    �  �#  �!  '  G   @  G   G   U    �.  �M  S  h  G   G   U    �8  `��  .   �   �; �  �1  G   �5  �  �+  �   `(    (�/  @  0�  U   8*  �  @ �    u(  
h  	  �2  (!  '  G   ;  U   ;   �  �3  ;N  T  _  �   v)  ]l  r  �  �    @    �3  y�  �  G   �  �  @   U    H7  ��  �  G   �  �  �     51  0�C  y2  �s   � �   �_  *
 ��  / ��   $ �A  ( 2$  ��  -4  l%  +  �h  �  $8  �%  	o  {    ��   	�  {"  �)  !  �0  \   �G   �  �N   }  �-   )$  �@   �   -   c,  +G   C*  6U   +D  C4    :   �V	  xx ��   xy ��  yx ��  yy ��   5  �	  	V	  8  ��	  ��  ��   ��  ��   $  �h	  c   ��	  �	  �	  U    �  ��	  Kl  �U    �  ��	   s  ��	  �"  $
  	
  �   +B
  �� -�	   �W .�	  Kl  /U    %  Dm
  uR F�	   �
 G�	   }  IB
  N   ��  10   �(  Q;  �4  �(  �0  *  /  d2  �+  	a0  
~5  �0  k*  �,  U5  l1  �.  �)  �/  l,  a-   .  !�5  "-5  #�%  $�*  %�-  &_:  'N*  (�8  0a#  1(  @�$  AI,  Q.  R6  S^6  T�9  UL3  V�(  W�:  X�7  `Z'  a�,  b�7  c�%  pU.  �I8  ��,  ��5  �+  �r'  ��9  �U$  �-  ��4  ��4  ��1  �i$  �@-  �#(  ��0  �/7  ��+  ��+  �E:  �x0  �+'  �'  ��'  ��)  ��%  �,  �
8  �9.  �0  �|;  ��:  �54  ��5  �+-  ��2  ��-  ��2  �+6  ��3  ��9  ��6  ��%  �39  ��$  �8#  ��:  � �  @<<  5�  >J   ��  ?J  �"  AJ  �"  BJ  i!  CJ   %!  EJ  (2!  FJ  0�  GJ  8   I�  �"   s�  ��  u�   5�  v�  ֳ  xJ  !  zJ  m  {J   v  }I  J  �#�  �  �!  �	}|  ڰ  	D   {3  	��  S0  	��  �/  	��  �1  	��  �1  	��!  Y/  	�m
  �*  	�"  (�)  	�|  0+:  	�"  8<8  	�"  X�*  	��  � �3  �"�  �  �(  	��  Oe 	��!   �-  	��  ڰ  	�D   U  �"�  �  �  8	"  ah 	!�!   Oe 	"�  U1  	#m
   ;+  	$  0 i(  �$/  5  l;  �	��  ah 	��!   Oe 	��!  y2  	�s   {:  	�p  (�� 	��  h/ 	��  p�� 	�  x T   � �  �  _  �z  �!  �   �  �  �  �    �  �  �   �U �  (�  �  03"  �  8�  �  @`  !�  Hd  "�  P�@  $�	  X�;  )�  h�   +�  ��  ,�  �
  -�  ���  .�  �?!  0�  ��  1�  ��  3�  ��  4�  �ȩ  6�  �ֳ  7z  ��� 81  �K <�  �ڰ  =D  �^�  >  �U  @m
  �t  B�	  �k  CU   ��L  E]  � "   �  �  1  Xm�  ��  o�   �@  p�	  �e q�  �L  r  P @  $%�  �    0\1  �-  ^�   ��  _�  �W `�  x a�  �@  b�	   �e d<  0�"  e�  pi"  f�  x� gz  ���  is  �.a k�  ��  l�  �J  m�  �Mj  o"  ��  q�  ��  r�  �M  tU    Z  u-   _"  wJ  (   xJ  Ud zU    �L  |;  ( �!  F#>  D  Z!  A�  ��  C�   T DP  �!  E�  "  F�   S  N   �P  Y   �  bmys�  cinu�
  sijs    bg�  5gibF  snaw  ahoj�    bg�  sijs=    bg�  5gib�
  snawk  ahoj�  BODAt  EBDA�  CBDA  1tal�  2tal�   nmra �  �  0  `)j  p  �"  �	e�  �1  	gV	   H+  	hz   x+  	i�  0��  	kY   8�)  	n#�!  h�'  	q\  p��  	r7  t�*  	y�  x �  �  1  �  �)    �!  H	�M  $  	�U    7:  	��  s4  	��   b  8H�  !  J�   m  K�  A� M�  �� N�  �  PJ  
  QJ   ��  RJ  (�  SJ  0 �  UM  x   �$�  �  �!  0
';  ad  
)�   �1  
*�  &D  
+�  2B  
,�  x� 
-V	     �)H  N  �"  P	��  ��  	�   �1  	��  �&  	�P  �3  	�V	  ]7  	�z  0�7  	�U   @�1  	�7  H P6  �  tag �   Kl  �   �6  	�  �  �5  N   
5  i7   �&  9  F9  8%  �*   �,  
�  ./   6
�  b 8
5   5�  9
�  ��  :
�  5  ;
�  Q(  <
�    -  I
(�  B  �8  N   ��  �:   4,  �6  $  �/  l9   �2  ��  o  |[  O7  �� Qo   �\  Ro  red So  q  To   �[  V�  �#  ��  �'  �[  a  �  p  |   �2  �|  �  �  |   l/  ��  �  C  �  |  �   �   ;)  H�<  �#  ��   :  ��  �5  �<  F1  ��  ,8  ��   2*  ��  (�*  �O  0`1  �p  8��  ��  @ �  �-  ��  d)  s[  a  �  p  U    9  F#�  	p  �$  @J�  �#  L�   y2  Ms  W� OQ  �� Pw  �,  Q�   M4  R�  (�;  S�  0�*  T  8 c/  X!  	  �-  (qK  �-  s�   Oe tK  ��  us  � vz   |  �/  )]  c  �  w  �  �   g%  .�  �  �  �   �.  1�  �  �  �  �  /   c	  73  6�  �  �  �  �   �  �8  :�  �  �    �  �   "3  >]  $)  Y'  -  �  K  "  �  �  /   �6  _W  ]  �  {  "  �  �  /   �3  f�  �  �  "  �  �   ;0  l�  �  �  �  "  �  �   �&  x�6  ah � B   y2  � s  H�8  �   P�8  � K  X�'  � {  `� � �  h�9  � 6  p C  �.  ��  "9  H
2�  Mj  
4"   H5  
5  (�)  
6  0�  
7�  8�  
8�  @ �0  
:H  T%  �
=  ڰ  
?D   �0  
@�  q5  
A�  L)  
B�  )  
CP  Ǟ  
E�  �  
F�  `Ud 
HU   � X+  
J%  �  1  7  =  �  `    �  �  �  �   �&  &l  r  }  �   �1  *�  �  �  �  z   �6  -�  �  �  z   w-  1�  �  �  �  �   �;  4�  �  �  �   =;  8    �    z  �   B$  <+  1  �  E  z  �   2  @Q  W  �  u  �  z  �  7   7  G�  �  �  �  �  �  �     q8  N�  �  �  �  �     )2  S�  �  �     �  �  �  7      �  k.  ���  ah �B   #,  ��  H�4  ��  P,;  ��  XEY �+  `/q �`  hZ)  �}  p�#  ��  x'0  ��  �.  ��  ���  �E  �� �u  �`9  ��  ���  ��  �5  ��  �U#  �  � �2  ��    �&  0�Y   y%  ��   �/  ��  �'  ��  �6  ��  �+  ��   �6  ��  ( �7  ��  *  V'r   x   �0  �*   u�   |#  w�   �#  x�  � y�  C4  z�   �&  |}   �'  ��   �   �  �   f   �  �    �	  �9  �!  !  !  f   �    A2  �*!  0!  �  N!  f   �  P  N!   �   8(  �!  ��  )�    $�  )�   �-  )!   )  T!  	�!  3  <�!  �� >%�!   ��  ?%f    �!  #  A�!  �!  B  �(  	��  <  |  "  @    N  "  @    z  ,"  @     H'  	�%C  !�} &�  (                                        "�O ��  �"  #�-  ��  #.a ��"  $ڰ  �D   �  %,~ k�  @�F     �       �V#  &�  k*�  < 6 '� (.a p�  �H)�U q�  � � *&6  t�F       � t9#  +36  � �  ,��F     =4  -Ts�-Q�H   %~ �  ИF     �      �E)  &�-  &�  � � &�|  &�  � � &f| !&�  � � &.  "&�"   � &�| #&  � � .�u  $&7  � (�U &�  ��)ڰ  'D  � � (~ )�  ��)�; *�  V R )�k  ,z  � � )�| -z  [ Q )�} /P     )�~ 0P  � � )�| 2J  %	 	 )8| 2J  �	 �	 )�| 2%J  m
 _
 )C| 21J  L H )
} 3J  � � )} 3J  � � )!~ 3%J  V P ) } 31J  � � )=} 4J  � � )�} 4J  4 0 $�} 4#J  $�} 4.J  )G} 6N   � � )w} 6N   � � /x 7-   l h /y 7-   � � 0f,  ]��F     1� �&  )`�  �G     )R~ �G   a ] )_| �  � � 1� �&  /p �  � � /q �  > : )�} �  v t ,�F     �6  -Q|   2E�F     �6  �&  -Uw -T��~���~� $ &-Q�� ,4�F     �6  -Uw   1@� $(  /p -  � � /q /  � � )�} 3  ) % 3J�F     C      /r 9  e a /s :  � � )5} ;    '�� /aa @G   / ) /fa AG   � � /fb CG   � � /fg DG   � � /fr EG   $ " /ba2 GG   S O 4bb IG   /bg JG   � � /br KG   � � /ba LG        5&6  ��F      ��F     8       Y(  +36  7 5  5n"  �F      �F            b�(  +�"  \ Z +�"  � � 3�F            6�"  � � 7��F     �6    2̜F     E)  �(  -Uv -Ts -Q��-R1 2ٞF     n"  	)  -Uv  2w�F     �6  ))  -Uw -Q�� ,��F     n"  -Uv -Tw   %�i �  @�F     �      ��-  &�-  (�  � � &�; (�  p d &.  (�"   � &J� (�  � � (�U 	�  �L)ڰ  
D  P J /s �  � � /t �  $  10� v*  /pad "�  � � )l~ "�  E 9 $p~ "*�  )^% #�  � � ,/�F     �6  -T1-Y�L  1`� &+  /i W�  L B '�� /ss ^�  � � /tt _�  H 8 /j `�   � 8��F     `       �*  /val f�  � �  3��F     (       /val z�  � �    8`�F     P       ~+  )5�  ��    /i ��  B < ,��F     �6  -T| -Q~   1� .,  /i ��  � � ' � /ss ��    /tt ��  � � /j ��  M ? 8 �F     1       ,  /val ��  � �  3��F     (       /val ��  ,  (     1�� �,  /i ��  j  b  '�� /ss ��  �  �  /tt ��  z! n! /j ��  &" " 3��F            /val ��  �" �"    3�F     �       /i ��  �" �" 3(�F     �       /ss �  F# ># /tt �  �# �# /j �  4$ 2$ 9�-  C�F      C�F     U       +�-  Y$ W$ 3C�F     U       6�-  �$ �$ 6�-  �$ �$      :�} �o  �-  #�} �8�  4a ��  4l ��   %�} 4�  `�F     f      ��2  &�-  4#�  C' %' &.a 5#�"  �( y( &+} 6#J  �) �) &R} 7#J  J* >* )�U 9�  �* �* /p :  n+ h+ /i ;�  �+ �+ /x ;�  c, Y, )`�  ;�  �, �, /y <�  {- s- )�| =�  �- �- )}~ =�  �. �. 8œF     |       X/  ;tmp W�  ��*&6  œF      �� [	/  +36  �/ �/  2�F     E)  =/  -Q��-R1 ,�F     n"  -Uv -Ts   1P� w/  /tmp �%  0 0  8P�F     3       �/  /q �  X0 V0  <�2  ^�F       �� w+�2  �0 �0 +�2  X1 H1 +�2  *2 2 +�2  Q3 ;3 '�� =�2  ��63  ^4 B4 63  �5 |5 63  ?6 76 6+3  �6 �6 673  97 -7 6C3  �7 �7 >O3  ��F     �       1  6T3  �8 �8 6`3  9 �8 ?l3  ޔF     c       6m3  @9 89 6y3  �9 �9 6�3  �9 �9 6�3  ): %: 6�3  g: _: ?�3  �F     #       6�3  �: �: ,?�F     �6  -T0    @�3  �� �1  A�3  64  ; �: 64  E; 9; 6!4  �; �; A.4  2��F     �6  j1  -U -T} -Q|  2ȖF     �6  �1  -U | "-T0-Q�� ,�F     �6  -U -T0-Q��~  >�3  G�F     w       j2  A�3  6�3  w< s< 6�3  �< �< 6�3  `= ^= A�3  2X�F     �6  #2  -Uv -T0-Q��~ 2��F     �6  G2  -Us -T} -Q|  ,��F     �6  -Us | "-T0-Q   27�F     �6  �2  -U��~-T~ ����-Q0-X0-Y�� ,�F     �6  -U��~    BN| ��  =4  Cڰ  �(D  C.a �(�"  Cd~ �(�  C\~ �(�  D�U ��  D`�  �N   DR~ �N   Ebpp ��  D5�  ��  D��  ��  D_| �  F�3  D�h ��  D�| ��  GD� ��  Eend ��  Dm�  ��  D�� ��  D/� ��  GD�  ��     F�3  Elen ��  Ein �  Eout �  D��  �  D�� �N    G4len �  4in   4out   $��    $�� N     Hh} @�   �F           �6  I�-  @%�  �= �= I�; A%�  => +> I.  B%�"  ? �> Jڰ  DD  �? �? K�U E�  ��J`�  G�  @ @ Jֳ  H�  �@ �@ J�} J�  !A A Ju| J �  �A }A 1ж a5  Jp~ k�  �A �A J\} l�  VB RB ,��F     �6  -T1-R} -Y��  1 � �5  Lp {  �B �B 8�F     I       �5  Li ��  �B �B Ls ��  C C Lt ��  TC PC ,<�F     �6  -Qs   ,(�F     �6  -Q}   ,�F     �6  -T} -Q��  MD~ 6&6  CUe  6�"   N�X ,@6  CUe  ,�"   O&6  ��F     -       �c6  P36  U On"   �F     V       ��6  +�"  �C �C +�"  �C �C 6�"  GD CD 7�F     �6   QBY  8Y   R�`  �`  vR�s  �s  �RCs  Cs  �QD  D   R�U  �U  { %U   :;9I  $ >  $ >  & I  :;9   :;9I8   :;9I8  	9:;  
9 :;9�  : :;9   :;9  .?:;9nI<   I   :;9  .?:;9nI<  .?:;9nI<  .?:;9nI<  .?:;9nI<  9:;9  .?:;9nI<     :;9n  .?:;9I<   I     &   I  .?:;9I<  .?:;9<  .?:;9�<   . ?:;9I<  !.?:;9I<  ".?:;9I<  #;   $.?n4<d  % I4  &I  '! I/  (4 :;9I?<  ) :;9I  *>I:;9  +(   ,(   -! I/  .4 :;9I?  /4 :;9I?  0:;9  1.?:;9n2<d  2.?:;9nI2<d  3 :;9I82  4 :;9I82  5/ I  6.?n42<d  74 I?4<  8. 4@�B  9.Gd   : I4  ;.1nd@�B  < 1  =.4@�B  > :;9I  ?.Gd@�B  @ I4  A :;9I  B4 :;9I  C  D4 :;9I  E.Gd@�B  F.G:;9d   G.1nd@�B  H  I.?:;9I@�B  J4 :;9I  K4 :;9I  L.?:;9n@�B  M.?:;9nI@�B  N :;9I  O.?:;9nI@�B  P I   %   :;9I  $ >  $ >  .?:;9nI@�B   :;9I  4 :;9I   I  	 <   %  $ >   :;9I  $ >  ;      :;9   :;9I8  	I  
! I/  & I  .?:;9nI@�B   :;9I   :;9I  4 :;9I   I  &   .?:;9n@�B   %  $ >   :;9I  $ >  :;9n   :;9I8   :;9I8  .?:;9n@�B  	 :;9I  
4 :;9I  4 :;9I  .?:;9nI@�B   I   %  $ >   :;9I  ;   9:;  9 :;9�  : :;9   :;9  	.?:;9nI<  
 I  .?:;9nI<  9:;9     :;9n   :;9I8   :;9I8  $ >  .?:;9I<   I     & I  &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  .?:;9n@�B   :;9I   I  .?:;9nI@�B    :;9I  !.?:;9nI@�B   %   :;9I  $ >  $ >  :;9   :;9I8   :;9I8   I  	:;9n  
I  ! I/  & I  9:;  9 :;9�  : :;9   :;9  .?:;9nI<   I  .?:;9nI<  9:;9     .?:;9I<     &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<  .?:;9n@�B   :;9I    :;9I  !4 :;9I  "  #4 :;9I  $.?:;9n@�B  %.?:;9nI@�B  &.?:;9nI@�B  '.?:;9n@�B   %   :;9I  $ >  $ >  :;9   :;9I8   :;9I8   I  	& I  
;      4 :;9I?<  9:;  9 :;9�  : :;9   :;9  .?:;9nI<   I  .?:;9nI<  9:;9  :;9n  .?:;9I<     &   I  .?:;9I<  .?:;9<  .?:;9�<  . ?:;9I<   :;9I     :;9  ! :;9I8  " :;9I8  #:;9  $ :;9I  %>I:;9  &(   '(   ( <  ):;9  * :;9I8  +I  ,!   -! I/  .4 :;9I?  /4 :;9I  0.?:;9n@�B  1 :;9I  2 :;9I  34 :;9I  4U  5  64 :;9I  7  8.?:;9nI@�B  9 :;9I  : :;9I  ;4 :;9I  <.?:;9n@�B  =. ?:;9n@�B   %  . @   %   :;9I  $ >  $ >  I  ! I/  4 :;9I?   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   4 :;9I  !.?:;9'I@�B  " :;9I�B  #4 :;9I�B  $��1  %�� �B  &��1  '1R�BXYW  ( 1�B  )  *4 1  +4 1�B  ,�� 1  -.?:;9'@�B  .4 :;9I�B  /.?:;9'   0 :;9I  14 :;9I  24 :;9I  3.1@�B  4. ?<n:;9  5. ?<n:;9   �� �B   1�B  4 1�B   :;9I8   :;9I�B  4 :;9I�B   I   I  	 :;9I8  
(   U  ��   :;9I  ��1   :;9I  4 :;9I   :;9I  1R�BUXYW  ��1   :;9I8  4 1  .?:;9'I@�B   :;9I�B  4 :;9I�B  'I  4 :;9I�B  .1@�B  1R�BXYW  :;9  4 :;9I   :;9I    1  !:;9  " :;9I  #4 :;9I�B  $1R�BUXYW  %  &U  '4 :;9I  (4 :;9I  ).?:;9'I@�B  *4 :;9I  +& I  ,
 :;9  - 1  .���B1  /I  0! I/  1�� 1�B  2'  3(   41R�BUXYW  54 1  6.?:;9'@�B  71R�BUXYW  8��  91  :���B  ; :;9I�B  <1R�BXYW  =.:;9'I   >  ?  @
 :;9  A :;9I  B :;9I�B  C :;9I  D.:;9'I@�B  E :;9I8  F4 :;9I  G�� 1  H1U  I.?:;9'   J.?:;9'I   K4 1  L4 :;9I  M
 1  N1R�BXYW  O :;9I  P4 :;9I  Q. ?<n:;9  R$ >  S>I:;9  T.:;9'   U :;9I8  V.:;9'I@�B  W.?:;9'I   X :;9I8  Y <  Z.:;9'I   [4 :;9I  \
 1  ]>I:;9  ^:;9  _.?:;9'   ` :;9I  a.:;9'   b.?:;9'@�B  c4 :;9I?<  d.?:;9'I@�B  e
 :;9  f�� �B1  g���B1  h.:;9'@�B  i:;9  j :;9I  k :;9I  l4 :;9I
  m :;9I  n(   o4 :;9I  p1U  q.?:;9'I@  r.:;9'@�B  s :;9I  t1R�BXYW  u���B  v1  w.1@�B  x. ?<n:;  y%  z$ >  {   |&   }>I:;9  ~4 :;9I?<  :;9  �5 I  �.?:;9'@�B  �4 :;9I  �
 :;9  �1UXYW  �4 :;9I  �.:;9'I@�B  �
 :;9  �.?:;9'I  ����B  �4 1  �. ?<n:;9   %   :;9I  $ >  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I  # :;9I8  $:;9  % :;9I8  & :;9I8  '(   (4 :;9I  )4 :;9I  *4 G:;  +4 G:;9  ,.:;9'I   - :;9I  .4 :;9I  /4 :;9I  0.:;9'   1
 :;9  2.:;9'I@�B  3 :;9I�B  44 :;9I�B  5
 :;9  6  74 :;9I�B  8��1  9�� �B  :��  ;��1  <.:;9'I@�B  = :;9I  > :;9I�B  ?4 :;9I�B  @4 :;9I�B  A.:;9'I   B :;9I  C4 :;9I  D
 :;9  E  F4 :;9I  G�� �B1  H.:;9'@�B  I :;9I  J1R�BXYW  K 1�B  L  M4 1�B  N1R�BUXYW  OU  P�� 1  Q4 :;9I  R  S 1  T��  U.:;9'@�B  VU  W1XYW  X4 1  Y1R�BUXYW  Z4 1  [
 1  \1UXYW  ]1  ^1U  _ :;9I  `.:;9'@�B  a.?:;9'I@�B  b :;9I�B  c1R�BXYW  d�� 1�B  e
 1  f :;9I  g :;9I  h4 :;9I  i. :;9'   j���B1  k.:;9'   l>I:;9  m1U  n1  o1R�BUXYW  p.:;9'I@�B  q4 :;9I  r���B1  s.1@�B  t 1  u���B  v4 1  w. ?<n:;9  x. ?<n:;9  y. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  #:;9  $ :;9I  % :;9I8  &>I:;9  '4 :;9I  (4 :;9I  )4 G:;9  *.:;9'I   + :;9I  ,4 :;9I  -
 :;9  .  /4 :;9I  0  1.:;9'   2 :;9I  34 :;9I  4.:;9'I   54 :;9I  6
 :;9  7
 :;9  8.:;9'I@�B  9 :;9I�B  :4 :;9I�B  ;4 :;9I�B  <��1  =�� �B  >��1  ?.:;9'@�B  @ :;9I  A.:;9'I@�B  B4 :;9I�B  C :;9I�B  D
 :;9  EU  FU  G�� 1  H.:;9'@�B  I.:;9'I@�B  J  K  L :;9I  M :;9I�B  N�� 1�B  O��  P4 :;9I�B  Q1R�BUXYW  R 1�B  S4 1  T
 1  U��  V4 1�B  W
 1  X1U  Y1  Z.:;9'   [.:;9'I@�B  \4 :;9I  ]1R�BUXYW  ^.:;9'@�B  _���B1  ` :;9I  a :;9I�B  b4 :;9I  c1R�BXYW  d 1  e1R�BXYW  f1U  g :;9I  h :;9I  i :;9I  j.1@�B  k 1  l4 1  m.1@  n.1@�B  o1  p. ?<n:;9  q. ?<n:;9  r. ?<n:;   %   :;9I  $ >  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  # :;9I8  $:;9  % :;9I  &4 G:;  '>I:;9  (4 :;9I  )4 G:;  *4 :;9I  +.:;9'@�B  , :;9I  -.:;9'I@�B  .4 :;9I�B  /.:;9'@�B  0 :;9I�B  1  24 :;9I�B  31R�BUXYW  4 1�B  5U  64 1�B  71R�BXYW  8��1  9�� �B  :��1  ;  <��  =
 :;9  >U  ?��  @4 1  A1U  B
 1  C1  D�� 1  E1R�BUXYW  F 1  G1R�BXYW  H.:;9'   I :;9I  J4 :;9I  K  L4 :;9I  M.:;9'I   N.:;9'I@�B  O :;9I�B  P�� 1�B  Q.:;9'I@�B  R :;9I�B  S4 :;9I�B  T4 :;9I�B  U
 :;9  V.:;9'@�B  W :;9I  X.:;9'@�B  Y�� �B1  Z.:;9'I   [ :;9I  \4 :;9I  ]
 :;9  ^  _1  `���B  a :;9I  b :;9I�B  c :;9I  d4 :;9I  e4 :;9I  f
 :;9  g
 :;9  h1R�BUXYW  i1R�BXYW  j1R�BXYW  k.:;9'   l
 :;9  m1R�BUXYW  n :;9I  o4 :;9I  p4 :;9I  q���B1  r���B1  s.1@�B  t.1@  u
 1  v4 1  w1U  x. ?<n:;9  y. ?<n:;9  z. ?<n:;   %   :;9I   I  :;9   :;9I8  'I   I     	$ >  
'  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I  $ >  & I  4 :;9I?<   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !:;9  " :;9I8  # :;9I8  $:;9  % :;9I  & :;9I8  '>I:;9  (4 :;9I  )4 :;9I  *4 G:;  +.:;9'I@�B  , :;9I�B  -���B1  .�� �B  / :;9I  0 :;9I  14 :;9I  24 :;9I�B  34 :;9I�B  4.:;9'   5 :;9I  6  74 :;9I  8.:;9'I   9 :;9I  :4 :;9I  ;4 :;9I  <
 :;9  =  >! I/  ?.:;9'@�B  @ :;9I  A.:;9'I@�B  B4 :;9I�B  C.:;9'I   D
 :;9  E4 :;9I  F.:;9'@�B  G  H��1  I��1  J :;9I�B  K�� 1�B  L��  M.:;9'   N.:;9'I@�B  O  P
 :;9  Q :;9I�B  R4 :;9I�B  S
 :;9  TU  U��  VU  W�� 1  X1R�BUXYW  Y 1  Z 1�B  [4 1�B  \1R�BXYW  ]1R�BXYW  ^1R�BUXYW  _1R�BXYW  ` :;9I  a.1@  b.1@�B  c1  d4 1  e1U  f
 1  g4 1  h
 1  i1  j1U  k1R�BUXYW  l. ?<n:;9  m. ?<n:;9  n. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I8  #4 G:;9  $4 :;9I  %4 :;9I  &.:;9'I   ' :;9I  (4 :;9I  )
 :;9  *  +4 :;9I  ,  - :;9I  ..:;9'   /.:;9'   0 :;9I  1 :;9I  24 :;9I  34 :;9I  4.:;9'I@�B  5 :;9I�B  64 :;9I�B  7
 :;9  8U  9U  :4 :;9I�B  ;  <��1  =�� �B  >��1  ?  @1R�BUXYW  A 1  B 1�B  C4 1�B  D1R�BXYW  E1R�BUXYW  F�� 1  G
 1  H
 1  I1  J1U  K1U  L4 1  M1UXYW  N1UXYW  O1  P.:;9'@�B  Q.:;9'I@�B  R :;9I�B  S4 :;9I�B  T1R�BUXYW  U4 1  V4 :;9I�B  W1R�BUXYW  X1R�BXYW  Y1R�BXYW  Z��  [ :;9I�B  \.:;9'I   ]
 :;9  ^�� 1�B  _���B1  ` :;9I  a
 :;9  b.:;9'@�B  c.1@�B  d. ?<n:;9  e. ?<n:;9  f. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/   :;9I   4 :;9I?<  !:;9  " :;9I8  #4 :;9I  $4 G:;9  %:;9  & :;9I  ' :;9I8  (>I:;9  ).:;9'   * :;9I  +4 :;9I  ,.:;9'I   -
 :;9  .  /4 :;9I  0  1.:;9'@�B  2 :;9I�B  34 :;9I�B  44 :;9I�B  5
 :;9  6  7��  8�� �B  9��  :��1  ;4 :;9I  <U  =��1  >.:;9'@�B  ? :;9I�B  @4 :;9I�B  A.:;9'I   B :;9I  C.:;9'   D :;9I  E4 :;9I  F
 :;9  G�� �B1  H.:;9'I@�B  I�� 1  J :;9I�B  K :;9I  L.:;9'I@�B  M1R�BUXYW  N 1�B  OU  P4 1  Q4 1�B  R
 1  S1R�BUXYW  T1U  U1U  V1  W1  X4 :;9I  Y.:;9'I@�B  Z���B1  [ :;9I  \4 :;9I�B  ].1@�B  ^ 1  _ 1  `  a4 1  b. ?<n:;9  c. ?<n:;9  d. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  "4 :;9I  #4 :;9I  $4 :;9I  %4 G:;9  &.:;9'I@�B  ' :;9I�B  (���B1  )�� �B  *4 :;9I�B  +4 :;9I�B  ,
 :;9  -U  .  /��1  0.:;9'I   1 :;9I  2 :;9I  3��1  41R�BUXYW  5 1�B  6 1  7U  84 1  94 1�B  :
 1  ;1U  <�� 1  =1R�BUXYW  >4 1  ?1U  @.:;9'   A :;9I  B
 :;9  C  D  E4 :;9I  F.:;9'I   G :;9I  H4 :;9I  I.:;9'@�B  J :;9I�B  K4 :;9I�B  L.1@�B  M4 1  N1  O  P
 1  Q. ?<n:;9  R. ?<n:;9  S. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !:;9  " :;9I  #:;9  $ :;9I8  % :;9I8  &4 :;9I  '4 :;9I  (4 G:;9  ).:;9'   * :;9I  + :;9I  ,  -4 :;9I  ..:;9'I@�B  / :;9I�B  04 :;9I�B  1
 :;9  2U  3��1  4�� �B  5�� 1�B  6��1  71R�BUXYW  8 1�B  9U  :4 1  ;4 1�B  <1U  =1  >�� 1  ?
 1  @1U  A4 1  B
 1  C.:;9'I   D :;9I  E4 :;9I  F4 :;9I  G :;9I  H
 :;9  I4 :;9I�B  J  K.:;9'I   L4 :;9I  M.:;9'@�B  N :;9I  O���B1  P1R�BXYW  Q :;9I�B  R4 :;9I  S1R�BXYW  T  U.:;9'I@�B  V :;9I�B  W4 :;9I�B  X  Y :;9I  Z4 :;9I�B  [.:;9'@�B  \.1@�B  ] 1  ^. ?<n:;9  _. ?<n:;  `. ?<n:;9   %   :;9I  $ >  & I  $ >     :;9   :;9I8  	 I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  ! :;9I  ":;9  #4 :;9I  $4 :;9I  %4 :;9I  &4 :;9I  '4 :;9I  (:;9  ) :;9I8  *4 G:;9  +.:;9'I@�B  , :;9I�B  -���B1  .�� �B  / :;9I  04 :;9I�B  1
 :;9  21R�BUXYW  3 1�B  4U  54 1  6��1  74 :;9I�B  84 :;9I  9��1  :.:;9'I   ; :;9I  < :;9I  =4 :;9I  >U  ?1R�BUXYW  @1R�BXYW  A  B  C4 1  D4 1�B  E1R�BXYW  F 1  G1R�BUXYW  H1U  I1  J�� 1  K
 1  L��  M.:;9'@�B  N.:;9'I   O :;9I  P4 :;9I  Q  R4 :;9I  S.:;9'I@�B  T :;9I�B  U :;9I  V4 :;9I�B  W4 :;9I�B  X
 :;9  Y.:;9'@�B  Z.:;9'   [
 :;9  \�� 1�B  ]
 1  ^ :;9I�B  _ :;9I  `.1@�B  a4 1  b1  c1U  d 1  e 1  f. ?<n:;9  g. ?<n:;9  h. ?<n:;   %  $ >   :;9I  $ >  & I     :;9   :;9I8  	 I  
4 :;9I?<  I  ! I/   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   5 I  >I:;9  :;9    :;9I8  !4 :;9I?<  ":;9  # :;9I  $ :;9I8  %:;9  &4 :;9I  '4 :;9I  (4 G:;  )4 :;9I?  *4 :;9I?  +4 G:;9  ,.:;9'I@�B  - :;9I�B  . :;9I�B  / :;9I  04 :;9I�B  1  21R�BXYW  3 1�B  4  54 1�B  6
 1  71  8��1  9�� �B  :U  ;��1  <�� 1  =1R�BUXYW  >U  ?4 1  @.:;9'I   A :;9I  B :;9I  C4 :;9I  D4 :;9I  E
 :;9  F  G4 :;9I  H4 :;9I�B  I
 :;9  J 1  K4 1  L1U  M1R�BUXYW  N��  O4 :;9I  P :;9I  Q.:;9'   R���B1  S.:;9'@�B  T.:;9'I@�B  U :;9I�B  V4 :;9I�B  W
 :;9  X4 :;9I�B  Y��  Z
 :;9  [  \
 1  ]1  ^1U  _.:;9'I   ` :;9I  a4 :;9I  b4 :;9I  c.:;9'@�B  d4 :;9I  e
 :;9  f�� �B1  g :;9I�B  h1R�BUXYW  i :;9I  j :;9I  k.:;9'   l1R�BUXYW  m���B  n���B1  o���B  p :;9I  q1XYW  r1R�BXYW  s.1@�B  t 1  u.1@�B  v1XYW  w4 1  x�� 1�B  y1R�BXYW  z. ?<n:;9  {. ?<n:;9  |. ?<n:;   4 1�B  (   �� �B   1�B  4 :;9I�B  4 :;9I   :;9I8  (   	4 :;9I?<  
 :;9I8   I  4 G   I  4 :;9I?<   :;9I  U  4 G:;9  ��1   :;9I   :;9I  ��1  4 :;9I  4 :;9I   :;9I�B  4 :;9I�B    4 1   1  1R�BUXYW  4 :;9I�B  :;9    :;9I  !U  "  #& I  $'I  %I  &  '4 1  (1U  )4 :;9I  *1U  +! I/  ,4 G:;9  - :;9I�B  .:;9  /(   0'  1 :;9I8  2 :;9I8  3  4 :;9I  51  6 :;9I8  74 :;9I  8.:;9'   9�� 1�B  :4 :;9I�B  ;1R�BUXYW  <.:;9'I@�B  =.1@�B  >. ?<n:;9  ? :;9I8  @4 :;9I  A.:;9'@�B  B :;9I  C
 1  D
 :;9  E.:;9'I   F
 :;9  G1R�BXYW  H :;9I�B  I1  J>I:;9  K$ >  L :;9I  M1R�BUXYW  N.:;9'I   O���B1  P!   Q4 G:;  R.:;9'I@�B  S 1  T. ?<n:;9  U:;9  V.:;9'@�B  W�� 1  X��  Y1R�BXYW  Z:;9  [.:;9'   \
 1  ]
 :;9  ^ <  _>I:;9  `4 G:;  a :;9I  b :;9I�B  c :;9I  d>I:;9  e(   f:;9  g.?:;9'I   h.?:;9'I@�B  i4 1  j1XYW  k1XYW  l1R�BXYW  m%  n$ >  o   p:;9  q&   r4 :;9I?  s1R�BUXYW  t.?:;9'   u��  v.:;9'I  w4 :;9I  x1UXYW  y.:;9'  z
 :;9  {.:;9'@�B  |4 :;9I  }1R�BXYW  ~ 1  . ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   :;9  ! :;9I8  ">I:;9  #(   $4 :;9I  %4 :;9I?  &.:;9'   ' :;9I  (.:;9'@�B  ) :;9I�B  *4 :;9I  +4 :;9I�B  ,4 :;9I�B  -1R�BXYW  . 1�B  /  04 1  1��1  2�� �B  3 :;9I  41R�BXYW  5�� 1  6.:;9'I   74 :;9I  8  94 :;9I  :
 :;9  ; :;9I  <.:;9'I@�B  = :;9I�B  >
 :;9  ?U  @1R�BUXYW  A4 1�B  B4 1  C
 1  D
 1  E1R�BXYW  F1  G1R�BUXYW  H1U  I�� 1�B  J4 :;9I  K1U  L 1  M  N.:;9'I@�B  O :;9I�B  P4 :;9I�B  Q.:;9'I   R :;9I  S4 :;9I  T.:;9'@�B  U1R�BUXYW  V :;9I�B  W4 :;9I�B  X
 :;9  Y.:;9'   Z :;9I  [4 :;9I  \
 :;9  ] :;9I  ^1R�BXYW  _1R�BUXYW  `��1  a1  b  cU  d.?:;9'I   e.1@�B  f 1  g4 1  h���B1  i1UXYW  j�� �B1  k. ?<n:;9  l. ?<n:;9   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I   :;9I8  :;9   :;9I8  >I:;9  (   (    <   :;9I8  '   I  'I  &   :;9   :;9I  >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<    :;9I  !4 G:;9  "4 G:;  #.:;9'I@�B  $ :;9I�B  %4 :;9I  &4 :;9I�B  '
 :;9  (��1  )�� �B  *��  +��1  ,.:;9'@�B  -���B1  ..:;9'I   / :;9I  04 :;9I  1���B  2��  3.:;9'I@�B  4 :;9I�B  54 :;9I�B  64 :;9I  71R�BUXYW  8 1�B  9U  :4 1�B  ;1R�BUXYW  <! I/  = :;9I  >.:;9'@�B  ?.:;9'   @ :;9I  A.:;9'I   B4 :;9I  C4 :;9I�B  D4 :;9I  E1U  F 1  G
 1  H
 1  I1  J4 1  K1U  L4 1  M1R�BXYW  N4 :;9I  O
 :;9  P  Q :;9I�B  R
 :;9  S  T :;9I  U :;9I  V  WU  X�� 1  Y.:;9'I@�B  Z
 :;9  [.1@�B  \4 1  ]. ?<n:;9  ^. ?<n:;9   %  $ >   :;9I  :;9   :;9I8  & I   :;9I8  >I:;9  	(   
:;9   :;9I8  $ >   I      :;9I  'I   I  >I:;9  (    <   :;9I8  '  &   4 :;9I?<  I  ! I/  :;9   :;9I  >I:;9  :;9   :;9I8   4 :;9I?<  !4 :;9I  "4 G:;9  #4 G:;  $.:;9'I@�B  % :;9I�B  &���B1  '�� �B  (.:;9'I@�B  ) :;9I�B  *4 :;9I  +4 :;9I�B  ,
 :;9  -U  .4 :;9I�B  /4 :;9I�B  04 :;9I�B  1��1  2��  3��1  4  5��  6�� 1  7.:;9'@�B  8.:;9'I   9 :;9I  :4 :;9I  ;
 :;9  <���B  = :;9I  >.:;9'@�B  ?U  @1R�BUXYW  A 1�B  B4 1�B  C1U  D! I/  E.:;9'   F :;9I  G4 :;9I  H  I4 :;9I  J :;9I�B  K  L�� 1�B  M :;9I  N
 :;9  O
 :;9  P.1@�B  Q 1  R4 1  S
 1  T4 1  U4 1  V1  W. ?<n:;9  X. ?<n:;9  Y. ?<n:;   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<   :;9I8  :;9  :;9   :;9I  (    I  !! I/  "4 :;9I  #4 :;9I  $! I/  %:;9  & :;9I8  ' :;9I8  (.?:;9'I@�B  ) :;9I�B  *4 :;9I  +4 :;9I�B  ,��1  -�� �B  .��1  /4 :;9I�B  0
 :;9  1U  21R�BUXYW  3 1�B  4U  54 1�B  61R�BUXYW  74 1  8�� 1  9
 1  :.:;9'I   ; :;9I  <4 :;9I  =.:;9'I@�B  >���B1  ?.:;9'@�B  @ :;9I  A  B :;9I�B  C��  D.:;9'   E
 :;9  F.:;9'I@�B  G :;9I�B  H4 :;9I�B  I  J4 :;9I�B  K.:;9'@�B  L :;9I�B  M1R�BXYW  N1R�BUXYW  O.:;9'   P :;9I  Q.:;9'I   R4 :;9I  S4 :;9I  T.:;9'I@�B  U1R�BUXYW  V1R�BXYW  W1U  X��  Y1R�BXYW  Z :;9I  [  \4 :;9I  ].:;9'@�B  ^ :;9I  _4 :;9I  `.1@�B  a.1@�B  b 1  c 1  d4 1  e 1  f
 1  g1U  h1  i1R�BXYW  j  k. ?<n:;9  l. ?<n:;9  m. ?<n:;  n6    %  $ >   :;9I  $ >     :;9   :;9I8   I  	4 :;9I?<  
 :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I  & I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<  >I:;9  I  ! I/  :;9   :;9I8    :;9I8  ! :;9I8  "! I/  #.?:;9'I@�B  $ :;9I�B  %4 :;9I�B  &
 :;9  '
 :;9  (U  )4 :;9I  *4 :;9I  +��1  ,�� �B  -��1  .4 :;9I�B  /1R�BUXYW  0 1�B  1U  24 1�B  34 1  4.?:;9'@�B  5 :;9I�B  64 :;9I�B  71R�BUXYW  8 :;9I  91R�BXYW  :.?:;9'   ; :;9I  <.:;9'I   =4 :;9I  >.:;9'I@�B  ?4 :;9I  @4 :;9I�B  A1R�BUXYW  B4 :;9I  C1R�BUXYW  D
 1  E.:;9'I@�B  F
 1  G1U  H1U  I.:;9'@�B  J :;9I  K
 :;9  L  M4 :;9I  N  O4 :;9I  P.:;9'   Q
 :;9  R
 :;9  S.1@�B  T 1  U. ?<n:;9  V. ?<n:;9  W. ?<n:;   �� �B   1�B  (    :;9I8   :;9I8   I   I  4 1�B  	 :;9I8  
4 :;9I�B   :;9I  ��1  ��1   :;9I   :;9I�B   :;9I  4 :;9I�B  1R�BUXYW   :;9I8  4 :;9I  'I  �� 1  U   :;9I  :;9  :;9   1  4 :;9I  4 :;9I  1R�BXYW  I   ! I/  !4 :;9I  "& I  #  $U  %'  &  '.:;9'I   (4 :;9I�B  ) :;9I  *.1@�B  + :;9I8  ,.:;9'@�B  - :;9I�B  ..:;9'I@�B  /.:;9'   0.:;9'I   14 1  2  3(   4.:;9'   5�� 1�B  64 1  7 :;9I�B  84 :;9I  9 :;9I  : :;9I  ;
 :;9  <1R�BXYW  =1  > 1  ? :;9I  @1R�BXYW  A4 :;9I?<  B��  C1R�BXYW  D :;9I8  E
 1  F1U  G.:;9'I@�B  H���B1  I. ?<n:;9  J :;9I8  K1U  L1R�BUXYW  M:;9  N1R�BUXYW  O>I:;9  P:;9  Q :;9I  R4 :;9I�B  S$ >  T
 :;9  U1R�BUXYW  V <  W>I:;9  X4 :;9I  Y.:;9'@�B  Z>I:;9  [1  \ 1  ]��  ^  _
 1  `4 1  a4 G:;  b4 :;9I  c :;9I  d4 :;9I?  e
 :;9  f���B  g. ?<n:;9  h4 G:;9  i4 :;9I  j:;9  k :;9I  l :;9I  m:;9  n4 G:;  o.:;9'@�B  p
 :;9  q4 :;9I  r. ?<n:;  s%  t$ >  u   v&   w4 :;9I?<  x:;9  y(   z 1  {�� �B1  | :;9I�B  }.:;9'I@�B  ~
 :;9  1XYW  �1XYW  �
 :;9  �
 :;9  �1UXYW  �.1@�B   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   (    <  &   >I:;9  :;9   :;9I8  I  ! I/  4 :;9I?<   ! I/  !4 G  "4 :;9I  #4 :;9I  $4 G:;  %.:;9'I@�B  & :;9I�B  '���B1  (�� �B  ) :;9I  * :;9I  +4 :;9I�B  ,
 :;9  -U  .4 :;9I�B  /U  01UXYW  1 1  24 1�B  3��1  4���B  5��1  6.:;9'   7 :;9I  84 :;9I  9.:;9'I@�B  : :;9I�B  ; :;9I  <4 :;9I�B  = :;9I�B  >  ?4 :;9I�B  @1R�BUXYW  A 1�B  B4 1  C
 1  D
 1  E1XYW  F  G.:;9'I   H4 :;9I  I
 :;9  J  K  L.1@�B  M 1  N1U  O1  P. ?<n:;9  Q. ?<n:;9   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I  >I:;9  (   (    <  &   >I:;9  4 :;9I?<  .?:;9'@�B   :;9I�B  ���B1  �� �B  .?:;9'I@�B   4 :;9I�B  !��1  ".?:;9'I@�B  # :;9I�B  $4 :;9I�B  %��1  &.:;9'I@�B  '���B1  (.:;9'@�B  )�� 1  *. ?<n:;9   %  $ >   :;9I  $ >  :;9   :;9I8   I  & I  	4 :;9I?<  
. ?:;9'  . ?:;9'   .?:;9'I@�B   :;9I  . ?:;9'I@�B  . 1@�B   %  $ >   :;9I  $ >     :;9   :;9I8   I  	& I  
4 :;9I?<   :;9I  'I   I  '  :;9   :;9I8   :;9I8  :;9   :;9I   :;9I8  >I:;9  (   >I:;9  (    <  &   >I:;9  :;9   :;9I8  I  ! I/   4 :;9I?<  !4 :;9I
  ".?:;9'I   # :;9I  $4 :;9I  %.?:;9'I@�B  & :;9I�B  'U  (4 :;9I  )4 :;9I�B  *1R�BUXYW  + 1�B  ,��1  -�� �B  . :;9I  /4 :;9I�B  0
 :;9  1U  2��1  3  44 :;9I  51R�BXYW  64 1�B  7�� 1  8  91R�BXYW  :.:;9'I   ;4 :;9I  <1R�BUXYW  =4 1  >1  ?1  @1U  A4 1  B.:;9'I   C :;9I  D4 :;9I  E4 :;9I  F  G  H.?:;9'I@�B  I :;9I�B  J4 :;9I�B  K4 :;9I  L4 :;9I�B  M.?:;9'  N.?:;9'   O.1@�B  P 1  Q. ?<n:;  R. ?<n:;9      �  �      /home/user/.local/share/lemon/sysroot/usr/include/gfx /home/user/.local/share/lemon/sysroot/usr/include/gfx/window ../Init /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include/lemon /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits /home/user/.local/share/lemon/sysroot/usr/include/freetype/config /home/user/.local/share/lemon/sysroot/usr/include/freetype  graphics.h   window.h   main.cpp   list.h   types.h   stdint.h   fb.h   stddef.h   cstdlib   std_abs.h 	  cmath   c++config.h 
  stdlib.h   stdlib.h   math.h   math.h   surface.h   types.h   stdio.h   ipc.h   unistd.h   ftconfig.h   <built-in>    freetype.h    G 	�"@     
�ff!.  tt!.�  	#@     �*  	�@     �K�"
�' t �	�K t�C�#��<tKxfftK� ot��K�"
� t�KA�#�( t ���<t���K *�t%����'��= k�u4� �&tC<O JC �c XC � < =, � � E:0!='tD< J t X. = �? �M   �^ t �m / !�ut<�t<hKfht<h�g\$��(�6X�f$��(�X9�@�<B$�2tR�$<<U�cXi�<f/�5�$<�;�XK�k�<B0B�4�B �<RJ�>�P.<_Ja�<8�:�<(.*�<.�0&�N�h0fhti� ���1u<6:Kf<f(<�
v'9$0
u�$Y4�K/Z/�.�t/gt.g�u?,$!
>,�, t � / �kv>f�.�f�.�f! J�f! J�!ffB J3 fg!ffC J4 fh�u,fftJg,fftJg�& J( t��& J( t�tf � ��"u%�* f�/.���u�<f5 �; t& < �.�"�.<fE JR fT �9 <d Jq f �s �� .X <L�13$V,f!�8.Ef:�J�u[�t<K'f�J='f�JZ'f�)J<='f�)J<" >4 <; t f6 u � K 3 . a.$�� J	�w  �" t f�	u5ut$ X X J t X�ut���<K)f�J=)f�JZ)f�+J<=)f�+J<!>3<:tf8u�K46t# X X J t X���<K'f�J='f�JZ'f�)J<='f�)J<>1<8tf6u�K6��'�t�$t<�t' X �; J�tJ" X' t <Y���.��K60tg\+tgZy.mf A'XfMJfC�RfIfY<<4.t��, [�� f�}���<J  	8#@     ����  	f#@     � 
�u  	x#@     � �  	�#@     � �t J tZ��/ t+ �$ t; X/ tF X �h�t! X �0 XF t' �K�! X t0 XF �' t=" f tut�tf% J ��
�K  	�$@     �  	�$@     )�#���tY��Y����  	�%@     � �t J t! X t7 X> th�/ t+ �$ t; X/ tF X �h�  	@&@     	 � t J / �    �   �      ../src /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include  fb.cpp   types.h   stdint.h    - 	m&@     �B��K �   b  �      ../src /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include/bits/posix ../include/lemon  filesystem.cpp   types.h   stdint.h   stddef.h   off_t.h   filesystem.h    0 	�&@     D��=>'�"3LH��=:>I��=3>?��KB>K��K �    �   �      ../src /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/lemon  ipc.cpp   types.h   stdint.h   ipc.h    , 	�'@     ��	�K2>������    �  �      ../src /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/sysroot/usr/include  runtime.cpp   cstdlib   std_abs.h   c++config.h   stddef.h   stdlib.h   stdlib.h   <built-in>      	P(@     �u��2�u��2��@��@��@�� �   Y  �      ../src/gfx /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/gfx ../include/lemon /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits  graphics.cpp   types.h   stdint.h   surface.h   fb.h   graphics.h   stddef.h   cstdlib   std_abs.h   c++config.h 	  stdlib.h   stdlib.h   <built-in>     ? 	)@     4� Y�	V2 ?0=tY Y�	V5��� Y�V	x. <0=t+ X tY	g[��t. X tY��#u	��E1,���tgXuXuJ�Xv�K01�!<b<, J9 <G <; <# .R J` <I <k Jx <� <z <b . J t 
Y>��X t f . =E0&�h>(ggwgg)w5�0t;.f�� t% �5 � tK0�$t<A.�5tI J5 t X <	 >g:f/�� w��]>8�J/<J&JJ�U>��
XL%K(�.<�4�6<%=��vu t �, � t� t �- � t.�$� f2t�Z JP �L f_ Xb X9 �� J� �| f� X� Xi ��(�-tJ><C�J<Y2�.f@t��@f<@/6�2fEXHX���H< <@/6�2fEXHX���H< <�F  � g t w<�o>�ggwggw t$ �4 � t� �� X� J� t� J� t� J� �� J� t� � Jn <| Xq J� t� J~ t� Jn �� J� tc � J6 JD X9 JS tH JF tU J6 �` J\ t+ � J .�_>)+w>�ggwggw#�*t6 J* t X < > t% �5 � t� �� X� J� t� J� t� J� �� J� t� � Jn <| Xq J� t� J~ t� Jn �� J� tc � J5 JC X8 JR tG JE tT J5 �` J\ t* � J ,�D>
= t! t. �> t5 <! J �)<"t8.?tG JV t? < f t{ = f[ .k �e tp Jb f  J> �4 t, J6 fP <G <' � < ��V>#%6<%<@.FtN Jd tF < f	 <$ =7 <& <A .H tP Jg tH < f	 < = <2 X9 tA JP t9 < f	 <
 = t, �< t3 < J� Y f[ .w �g < Xy t� <� f� <� f  t> �4 t, J6 fP <G <' � < ��O>�
� t! t. �> t5 <! J� t! t. �= t4 <! J�tf"t$<KuEtQfTt�<"Xt(<5X,<6JT�8.2I  �� �   �  �      ../src/gfx /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../include/gfx /home/user/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0 /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/bits /home/user/.local/share/lemon/x86_64-lemon/include/c++/8.2.0/x86_64-lemon/bits /home/user/.local/share/lemon/sysroot/usr/include/freetype/config /home/user/.local/share/lemon/sysroot/usr/include/freetype  text.cpp   types.h   stdint.h   surface.h   stddef.h   stdio.h   cstdlib   std_abs.h   c++config.h   stdlib.h   stdlib.h   ftconfig.h 	  ftsystem.h 
  ftimage.h 
  fttypes.h 
  freetype.h 
  <built-in>      	[6@     �K��>���X>K	%[hLu	%[Y"�K(Y��!�&Zg	#!1�@g	#1�v���X>K	%[h<u	%[Y"�K(Y��!�&Jg	#!1�@g	#1�`v+�K�f' JYf�L t+�1�f� tgJK ; 9	 c	�)�5�0t;.f���?g#��" t0 � f�	��U�\�If#�u.it<=& t4 � f���(�=tK�1fQfTtf%K �)t+� �.�CtQ�7fWfZtf(�6�KtY�?f_fbtj�J:5�>t�&Y<'�f'�f.�;@X;�4J&JTJafXa�ZJLJnJH<�.��X���JyJ�Ju<.%= �)t+�vt	 � �%�'tKqh(f J t' X$ t@ XYfYut���<t�K	U)65�0t;.f�	�ut�	t�t� K Y-["t	�Cg#�[& t4 � f9 <? �T �[ �H fr t9 t#�Y�`�'fytth* t8 � f�,�AtO�5fUfXtf)K-�$X7t9�$�2�GtU�;f[f^tf,�:�Ot]�Cfcfftn�J>B�9XLt�*Y<+�f+�f2�?DX?�8J*JXJejXe�^JPJrJL<�.��X���J}J�Jy<.)=-�$X7t9� uX	 ��-�/tJ�_X	yX	<!  �    *   �       ../src/gfx/sse2.asm      	�B@     !>==ALLKK0=!#!>==?LLKK0=!#!>>K0YLKYKYKYMKL1="#!>==>K0YLKYMKL1=" �    �   �      /home/user/.local/share/lemon/sysroot/usr/include/bits /home/user/.local/share/lemon/sysroot/usr/include ../src/gfx  types.h   stdint.h   font.cpp       �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftinit.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftmodule.h   stdlib.h   fterrors.h     	�C@     � u uX	RxX�
BzJZ	x<
XX �tXtXtY�<�
�m	 Z  � F�	fNZ��	K	�	 Z  � F�	fN���	K	�	 Z  � F�	t\�JJ7 J\�O
 Mf J J6�������v
�Y	X�X=M�~J	[�
BzJZ	x<X���.yf��qJfJ<�[y'?[�/ utX c�   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  fthash.c   ftobjs.c   ftutil.c   ftcalc.c   ftcalc.h   ftrfork.c   fttrigon.c   ftadvanc.c   ftoutln.c   ftcolor.c   fterrors.c   ftfntfmt.c   ftgloadr.c   ftlcdfil.c   ftstream.c   ftpsprop.c   ftsnames.c   stddef.h   stdio.h   setjmp.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftlcdfil.h   ftdrv.h   autohint.h   ftserv.h   ftincrem.h   fttrigon.h   tttables.h   ftcolor.h   tttypes.h   sfnt.h   fthash.h   ftstream.h   ftlist.h   ftoutln.h   ftvalid.h   ftrfork.h   psaux.h   svprop.h   svsfnt.h   svpostnm.h   svgldict.h   svttcmap.h   svkern.h   svtteng.h   ftsnames.h   <built-in>    string.h   stdlib.h   fterrors.h     	pF@     3=2Ju/<JJ<IJ��"=	=t0<	<=t(f=I0J	<=th0	<?�x��Kz^�<	XK�<Z
�M
K
	Y!fyJ<X� .�f�H>Y<1�YZ�xJJYXJ���x�f  �x.. 	�G@     �LX	JL	vJZ
<	�=J%u.J
<�JKX?X	zf	u��$�u<�
�u<�
X�uJ<<�
v�� �.�jL��j�
JK
w	���j�
F�J��jL
w	��J��jL�
�j�K
1	�N�J��jL�
�i�K
1	��J��i�W
�j��<<� z 
 L+ W ]�  =?t.w;>r=7�Dt	�J	=	=2r<<f�>
�	ZJ	=	=2y<<f==a.�<?q=7�t�=.�=?t��
�>
V<	JJ	=	=2y<<f�>
�		XJ	=	=2r<<fYN8N= U.	
w.	Z;u<	=	t�&�&:	K<,tZ:fJ>= �~t=>X�ZZ&Y;=&�u=;==�&X�)tmttjJ�J�M�JY<%<<
�M�<t`v_Y<X�yJCy C ...y.JO8Xp�J	X?Gi  ...+a�"XX ....EX��X�<�L<]�t�pJXJJN�~IY� <XJY�<�~JI[�J�<�~X��pX	<<�	J�>
Z	v	IKLJw<$�.�>
�[/���xVX	`Xt�+Y	<	�l�
X		f	K!M=F	?	L;	@�=uvKut!u	JX=KKLaX;;-.=KKL� tmXt�~�<X�LV)�"X�=W)�"X�3z<�"�M3<[)+LK)H2KK)GK)K2K2NZ�
J	J�	�
	YNXJJsZM
�	�b*<�
Jf.o X2�	�|L	�t�| 
�K
�J
wL
K	=
�M	��|L
	�<�| 
GML"	^<
�<
GM	��|	�.m	�|�J 	^<�J 	�.y^
vJWKJ>�[X�JZ  �}Xz DHu�Y!tu!���X	<t�M����YZ�e�J��lX�y
t�xYt����J�y<	L�>YNKG>K �	=LYNY�>[K� Ju	=>K
	Y��}�<�vXu�X��}J3 =�'t=mg� �=>w	X X < Y X < . < X < . < � J = - < =>�	X=>w	X X < Y X < . < X < . < � = - K>��L<
<K
w	� J
.(>xn X < g X f <% � < K% - < =>�� #�|L�t.�|f�J�| �J�| 
�!
K;J�	L
��L
?
GM��|LL��|LL
	=�
��|<	K�J
�F
�J�|fIK
�	�|<
��J	�|<Z
�J�|<<	
�M��|LL
?
GM�	�|���	�| �J
�J�|<
�Jd@,	<
u 	J
C
wJR
yJQ����|tL��|�<
<K<
<K�L
M	��J�|X Jf�<i�|>�J�%iK.�<u�|�JL�v�|�J��=�|�J��Lu�|�<K�%fKZ�K�|�J<����|XJ�J��L�|�J'�f�|�J�<�L�|<<%iK.�<u�|�J�J<J<J<�L�|Jf%fKZ�xJ<�=�|�Jt��z [G1Bw
	Ȑ<��
�Z�
�Z�0
�Z[
yVNT^8LT
<
yR
zQJ����u <t.KH?Jr��sY�g
�
<Z
X F X>
X<t H	X��<=ItKI =I.=Iu;'=;=L Y WjYJ�6.jf�{Ju���{�K-K>
�[�{�K-K><��{�K-K><��{YK-K><��{YM+?f>�xJ=-=@�6.�{fJ=-=@xJ=-=@�xJ=-=@xJ=-=@�z�[G1Bw
	J�<XZ�>
>i
B
<O  .��=Kf=0 J < gym J �
��`!f � . />)=X<-=).)<<�>�	g	1 � < .
.v � "  = - K& ; K ; =  3  " < <" J J	 < �! t	 I Y L	   >�%<<�=%..�6J7O2<<ttY� X])	.A.)	.3�X	K;gx<
	KJ� � H� < . � . /�	J=	/	.#�M	+1.1fN*J@$fJ..
tg<KLt<�< � J u  � < � < X J u  X < � < < X �  <3 <' J � yX � J t Y J t
�wXZ�g6d�,y��`	�[fktXk<�gM�YtM  m�
	YvJp . i��.�[-i#g#vvfX��o�Yt � �4�uHvS��G?<Y<<@I�;YfAI�:YfBI�9YfCI�8YfDmwHv��n ��j�l��v^,tX ��?Y"\t$J\< $ . 	 c@     S���.�~(X!�Ju!��~(=IK(KHAEK.(XJM0ABw%Gw%t��~0*<�t��['JFK)'H-L�� K/  < :]��~�W[�=Kt	 �  K<  Yf	 1# s J�IY�3�fJf� �luJ[=t�Bzef[=t�( >
�_ottt=�sK�K�Lt ttt=�sK�K����[W[>V>y�`�}�S��<*tJ<	Z�LKX foJ..o�.nKK=u��yQ@XX 	0g@     � W�~f�tM�~Y.�
	K�� �  �.��   .J8�t, X <W&��~�X�~�<<���n r�tKI=uGMtY1�t[
t^�|���  .	z �|<�t	� �~��p��=J�<JJfA	� �<tXXYZU=A=y<K$O=y<KA$zXK]SBz<$Pz<=B;S$Pz<MZ�:�� KGJ'LKHKK9=x<K;=>��Jn	px<ztukxJ�t4� .wtu47��� .puvD�~X�.t�a�KeJK]�!��S� I'K;=IJKA
X K's=eKI=>
#XhK eJ=g�!��	^�#=/;XhJ	�#=/IXhJt�J�Jh,��ZvX �.�"iK{ytK	ZJ	�J�	<nXfofMtY0��|�J�|J�f �| f ��f�o=NYt.kWt\�z�Xt��JY[J�3XY[�xt�~X�X�xJ[�~YX�
����Z�xX���w�f  �xff	� ��	� �f[vv
X"��!v`!<J��!Kc�%u%8�%�%�& �P#�#���[	tL~]C x� R tZt�
-J	m��l	K�EZ
f�	N�l�fJX�k���z 4 �e Xe�X� ��u
�=�u��k	u�EZ
f�\�k�ftX�jt�
�r�.f�`J X..	u�s	�Yi Xd<�"�j���&X�NPzfZtCY���vJ3JLJH'�J;'=3;2=sK2fK( %JIu+K4I;JJY4;JJZ��jvY�%<%J<=X�L�j�%<M%+<?>�
JM�jt�%<%J<=��L�jYV�#8��,:K,-�,KL�jJ�<��j֐�MsJ�jf�%<K%-<=�<J
<MX 	0r@     jvHL]ct�� Jf��� 	��"�s	�<	=��? � &  �   ?
 	��i��%<%�<f<�	L��i���L�
X	K�	K	K�	4��itL<
<K
KfM
	K��J	��iLJ�1KL8cKIYZ..x.	��&t t.	=	=�	ua	�Ks	K	K7��iY�%<%t<�-�J	K�<yfK�<�i��%<<%J<=<�%<<%J<=��%<<%J<=����i�%<%�<f��Y 0 D�.�   Xi J[��Zt�z%XX��jJkX-.`[ X! t u /4 VwXJq	J4t�v�Z0,XD<<XH�
�'�	f�}NW���
M�`f$�V�� �zP
ZwJ
Lt]z<uYKZYq�)Yf�<..zP
L]�H�^]z<uY�YX���vu�Jtp�.<n<�.2
	��5�gtLJ
JK
1	�JJJ
$J<�K�gL
1	�J f�L�%Xg�fJ��K<<�N�L%Xg�fJ��K<<�N�KIKIKJ <.�J� .  J��� .Bf>XE�X�f�X��w�f���[[t u� X X u � < u J .   [BzJ�  .z.zxJ`  ..q ��`�\Q�	K[JLZ
<�
<VJqXX' f. =' W	�	u.ht��X6< X <#[<K
Jt
J4 s .�5w �J X tT wt	<=
qX. l�."�� X �  XvK i	   J �Z$ f fq-.YLtJN��� � t  XvY	J.=
	Y�	�mtK
xJ.Yvf*��'$tm<�	��Z)/'�IJZ
<	��Z/-tIJwX4X'c�-n�?�a X��% Y�� uf � u J X  J	YFj � w�  t  <��t  wX X .  X��t���>
.ii� lf t l J X  <YE] ��G[  nXXt<w� �  t  < � X J .  ��et�[� tf J X  <	YA S  t  <��< v. t  X��v�t�� Xht y� C X y Q < y Q .  
 	YNF\ �f  �� Xit y� 5 X y Q < .   [!  ..-z.�[ ...9[
�W Xit v� 
� X v 
J < v 
J .   [/X ..JG[  ..�[C X <[t< v� 
  � < v 
J .   Z
�MKXJvJ
. v�
.� zX � <[t< � t   Z
�MYXvf�
J�z<�x	�K��LJZ
 Y1 �	i<	u�YX .. qJX mfX�n�tX q<	 toJ&�JZ
<�@W	h@X tsJ.  s .�X Y9 sY�[f�J<Y
	Z		J�y m y.t . .	�T�zPJ<[
	Z		J�yJ5 y .�  �TPt[
	ZJ�t. W�T�zPJ<[
	Z	J�E3 Jf  ��T�zPJ<[
	Z	J�zJ4 z Jf  ���[
= X�v.z�_u<�[	vZ
<	YKwZM
�M
`JsqX	fY�
� ��~[	vZM
�M
`JsqX .�  ��z��;tL�JY<$<J
�Q�<.<sJ.�zPZ5 X < K5�/���w	t
t	Y.h
	�	K	K,<	M�<ZtZY!wX	JXm%.f.t[X�%.n�Z(;K(<M	Z	�VJXYoXo.o<�=K�KIK�~X=�t��}K<X�NNJY[�[��$�E3 <..�~��c�yJ�XJ�f��_	��EZ
f� wJM
��_� ��^t�!�B	�JsZM
�<f�t��{fCI	�$	J<�~X��� 	P�@     � 	`�@      	��@     [vF]/�ZKK?Y>Y>Y/n�-;��� ��.gx��uftl�X	@�!J	<ZY,= Y> �N
fJZ�J�J!o	<X�$�g�XJ�V��)I/. B��c� � f��(.�mZzP�
	Z	�Y.i�.if.� Y p5 [Y�5pf�,.�?./J/>V=<=�L�o �2��\i�Yf	�U���d F=Kh�
v�

��X"hrXt>"<�WY;=;YzXZTJK�X=w
�
���
M	hX	K<f�kS�NT�uJ���~�.=<oX=	<�#=0;=;KI=;=;Y	\	KJtJm:��<J�O�J@ ��cK������RxX�QyXCyX�uj�J��Ig;=;=;Y[�FKIqK;=;t;YZ�XX�X�KUKZ�Y�Z��[(=B2yXC2yXus=;Y2zX<Zu��<=8
 � �~ �X �~f < �J J �~ <����
��9�~�YIY� �Y� �X� �~��X <XX_<</� �Z#K#K
i.�
�J+	�	M	 �  J x.X<��Y��VjuX�rJX^J\9?9@ZI/  ff��v�o��f��v
f>�h�}JY<<	�I��}Yf	�I��}Yf	�h,�fm��Xu��&�	�[	VLX Z*  > =  ? K
  F^5�v�60v<f )�< \)Ju; 8	@)J	=Z<KIH��zX	J	K	?�=>KGK=wX,XJ(<XJJ+�Kf
.[[�(XR<�4�]wJGK5:�5���[[�� JsXX�<�� �������# ��{X�JX( �5 X! X�.myJZ:�,h<L^zJ=<Le<fJ�'!M'9?!t=I=!h	 '  g �	 =  h :	 >  x 8	 @  w< X  < l<�W
ZPf4.-Y�~X�=v<	.wJ
.vJ	.=v<	.=v<	 w<X:YY/� ..�XXK�[GL�<kfX[@xt�$Q)~��[x.�Cz'<>�'Jt<=I=IYYZV>X		�X	:.u"�< � �	���W�	Z��MU_�zL<
<�
JKL
�
<�
w	�	H"�`< J	�<?�N�K�w<"!y<A�zY Y	�L�y<JX	�<M�yL
XK
<KwL
	=
�M	H�J	�� ��yL
�u
Iw Y	�	�J� X��&G�H. � � � <  J �X < � � �9f�zY Y	�9[K�X�z��X�X�
Y
Wv�� X�~.� 	��@     �y	twX	�wX	f.��

� =X # J	 zJ	X .	K-X	#X.P
=
K
 � L- M�
 v�9 
J
z�H'	J�-�� Y Y Y Y Y Y Y Zu�X� �
��t	J
	��oX.XK"� �Y�J
J�t
JtL
		�>�Z�S
	J%#J�	Vf ;C�"�		�%	!�A�A.�
Jf
JfLY0XoK0�hJ/uuuuuuv�Y���	�|JZ
�X���,<,�J�JuJh�
	[��}���JxJf�...�|JH tH fu�=K����� X JY/��JZ
fXMG1  
sJfoJX  �WN\]J#JW<Zt
.XJrJ.  
h�fG[  q[AK��J	X�Y<
<hJ.L
XX ..x�F\mt=ft�`XfJX 	��@     5�JJ[�Y<<<
<Nu=w<f<<X#� = XvH</XRJ<<8u l��
zXo�.#��~��~J�X�~J<Y
	��F@	�x<>
	Z�Y�	� 4E['K	7u'KX 
�~���~tU4�J�
'K�~<.�'KJX Jmf]J
#X Y/ ;X%fK'=';K�� .�	�~���~t� ��YL!JM��X � �
r rX<0�~<�X�~J<<�t�� �I/g(�?�K0Jgt�L�K0Jg��L�K0Jg��KAK0Jg.J./K3K0Jg.KKl�Ha[JZ
�fuI/  �u��	X p�
	gt<x�hJJht
	Z��	^��	X z�uI/.	m�m
.f�|�wy{J�..<<
.�LP��(X.TK� � W�W�e�W@{cyJ%U>1yXN%.X%<1S@%;1%W.X%<1S2%;?%I<f%J:B��!
f
�%�JMd"�JM;#�F<0JM:#�-<M;�B>JK���
f�L-nJ�T�hX.K�W]�YYtEm.lCW�J�..
��f
� ~N
XJ
JL[9�<J�
�XL� =tX.
�X�� �J� X t.F<!
f:��J� X t.
�f�
��
�tx�hJJht
	Z��	^��	X z�uI/.	m�m
.f�x�hJJht
	Z��	^���	X z�uI/.	m m
.f�x�hJJht
	Z��	^J3�	X z�uI/.	m m
.f� �j
<XXJLK%Xt<]t
�JN�zW�J�
��J
�~�
XJL[J�zt
�XJ�	�%pJ��
J�
	X�zJWJJ
Xf��yJ�X X
�z��	��<�+�	�<	L�}�yCu[<X�]�yCu[<X���x�hJJht
	Z��	^3�	X zJuI/.	m�m
.f��w�0:�t�JvL�<��X� Y�{v�~J�X�~J�J�����f..	R��	�
�
	Y/?<.2'K	I=�	<@J�J	� �	Ks�	�	Yx.	/-	Lx�/-J.	/x���W	=x�t�W	=xf	=W	L]�	�	�	K	i� �	/�	/�	=��k�R��X� -J=.��f��fJ�|�J><<XEJ0<<XSJ@Z��X>X<YX<.<X%W<%J<=Z�>|	�zfy	J	VK	;Y<Y�Yn��#xn�:Zi�<<Ye/Y�}J�.��t?�}XL��}�.�?tL��0<w%fK%<I=;-<Y;=-J�}�.��t?�}XL<��}�.�?tL<�
�K(=;=(LX���x`1
\�.sJ<s <wX��;/Z�}J`.�?tL�M*./*I//o�<oJJo ��}�.�?tL<�K&<[G0<10<ihX.�}�	NK	:ZY��fix�tv:Z1�<<Y;=Z�|J`.�?tL� XgV>K��|�.�?tL<�: X X [=:���i�e�e��|.k�Z<=
mX�Z=� 
fwu�=��Xz�OS�
�JL=Lf  ��
v<O�/X</<Y
 ��X=Z!:!h>1HH[)g��� ..x��kJ.<...�~�w 	<wX	�<Y[K,vX JzJ^  T�w 	<wX	�<Z[K,vX JzJ^  ��y)_y<�qX)_Z
��
XJ
J�...yX�;=�=�
.y)_y<�qX)_Z
��
XJ
J�...yX�;=$=��$��
JrXJr
J�<JM�>Lv�LX iJX�X�z�v���
XX<�[L.M�~JL�KK���LM� .J
b.
PJ0 ����>
xJRK�6 �IK JJ�J� f�..�� OJ1fL 4fuX���y�YXV�X/M�}X[���}X.��{Z�~J�M�~YX�	��	� �t��}JX�..�<x
XvX6><Z[�Z��{��Mf...oOX ...�vJ
X....J�x
XvX6><Y[�Z��{��Mf...oOX ...�vJ
X....�~�x	XwX6=<Y[�Z��|��Mf...oOX ...�vJ
X....���s�u�X�P�rZY�[. t�ltZ�~�X[�~�XJ�
	���	� J��kJXJg�XF�[wJZ8�uYy�_�n��Npu<K�}tY<<��g� .�� ��tu��pJLJ�<X
<J
JY�X Jh�Z�}
	w�u�KIK
L:L
���
<<[��[�K
Q�v
	�
JX .._�!X\��{�� �~
XJJ��K	��|�	��{�W=>���J���z.�f�tf
	� f��}[	vZM
f�M
�JsX���<�~ 	J	L�	��	]���tX.X�M1�c�
tvtAi>YJ�	�u(z��=9 �
��}f�	v
	YNX�Js�M
f�X	� f�l����@ X J[vJX�X�`� v� 
' � t�}�<�.�}�['+�t�}����}J���y�}.���}����}<���������h<?�;Y�� <Jx
�
����6 ��(�!J�yJ�J���M!J�yJ�J<���J��
X	M�!�eJ�ftKwXYN	v�Js�M
X	�e"&MU�	.�	�}X<� sK ?4 Jh4f�[
< 0 .�
<	/iJ< ti.	v�X<�}t���;�J�9�7��
 �4 ;	� �y. �J	��y����y��EX �	
f�AW?�����	:�	/	���~����L]xJKZ\zJOK<LxXR<J���X �~<5 f � X
�4 JiJ	��	2 . tXu�	�vf#O	[#}D>J#@�	2#<�z�J��<�wJ<��<�� 	�e���	�|�t	�{�	v��*>=?K
F�9��tO\FFIK
X7Kx
XvJR<LX��	�}X��z� tw��tX	��.�&Xf��
t�X�<�</
�
�W�u/��<	f�:JyJZ�
N��`$X	f.�f�_J!.JJbJ�r,XW�)�֐....X 	��@     ���v�sJ
t� XZX�</
M
OX .. r� <�I�  .-p�X	y<�� ff..�i���T{xRtY�	J>:/X<�kIY Y��w	fKM
sX
JJ<s<
�X
J<�uTuJw/�
JJ�x-��# J	v�01IGX!H��OoOK��
J	YY�vY��	�vY��	�X ..ut�}X�f<X� 
Ji�tK� JLK�X?
JJfX
J
J	�K�v�t��tn��kJGvw
�<X
J<J�jY��JX ...7 cf4  7 J4 <J�jY��L
 �LJYXMLK�K�kX�
J�aX&XT<������Wof�X�8�< GZ=<<
�	MKW	ۭxUKX�5
tJN
z<K;K@	JKwLJ��XK
�*<.fXJ. ���.f�{K
JJ�?#u;K?
u;�	[�	K	�4�	��K�_� t�RB	vX�Js�M
�
,TJ,t�^��!�<K
f�|�^X�!�K<Z
JE X�EI	Z&	J<�Z��%���=��{Xt�_�� AZ=�/ 
xfw�/ u%<)Jx�)R�!X=�
_J
�&Z&VX
\J<�<>,JL:=s�#L4.�<<JJZ<:=J s JWf�
D)xU�X>
J J�K�..a<�>t A�Of
<JL.g(X"JK*(e<=I>JgJ(KH><Am<y<.L"XM]B(x<AOoMBtX <)JLtJ=�'.0X+JI=).>�X<.Lt<>
�
'J
J �= � K= I�
�+XE@=).<>�JL
��
�MMY�.(XuIK(KHA(GHK0ABw%Gw%t� ��XX�OJ1X X�	W��JJ	N�@$J+�#	fg#;x<=�/u.Ju�=sW=�t
�M0�� <>�*�  X �.oJ<X<r��aJ=v	wX��XL�����=X	LX	�J- r . X �`<�@G[XJXP$X<J�5E<%O7JZXY5%?qRZ�M��YZ�e��/X ...x�t��(   <���<X<X
<JL�I?GK
	Z�	KO
+O(J,tNYLf....�\J$X����YZ�e
�f�d<<�� xJ	�e��x�>#%�W?
.�X<X
JJ
 K; ��	K�K��eJXf
r�;��YKLgX X���:�Y�==Xjt<Jkt 
JL>=L
<Q	��O
Zu�K�K-=h
t�Mr�<�
J	Z	�J+7J	XY�sJ	� �	� �t� �X 	��@     	0X 	��@     �j8\Y�~J��~X�..<<
.�L
� ~�
XJ
J"J�. �) � K) WL)��
 qX <Z
<� Jt
�~����� �	��rXsXJ;	�J	��~J�
�X��~XL�8	���X	<�<�~�
��J���XJ<��~JWJJ�
�XJ�	� � i  X t J �  g	 <Z�JJL�~W�J
���	8��~Y�	�
�~��
�	�	t�	� �3 + <3 X+ J	 W Y J	 I[Y�	=ZX�X&���;`XyXKX>&Jt^J.�J�.�@  �1<[U[�<uu�JrJX�pJ�..<
X�
�J�p���
�
X<���.]o<Oj�p�J�pJ�
��
�J�p ��
�
X<�p�� �pX��pt<�Kkeg39�pXu���
	��h�}J��}���o�Jf�rJ
�XL��X
X�
!�2X!X6;�XfJ�>�r�J�rJ
Xf��rXf��pY���
	�
�o���9�p���	�~
�rX���X
�
��8j0VZ
Z.����q�
�L��
X�

�J
<�
7�
	f\
	�XJ	�3$;	K3$J	Y3$t	Y3$t	Z	�J	�	ZH>	Y	g	g	g�
)�J��q�J�q<��K
J�X�>�q�J
�����q��X[�� �p��sf �f� �pX
���
�pX��X�
�q�	�<�� X�NJ� 9�pX��<�<���GYhZ/ ;K/~N bY/ tY/>/, JL�X�� �q��t�<X��J�Yh�t!.a<!.a<�e<�!JfJ�(M �  X J  X K ��<2 �+ J�
<	��K	M$,	L<�<� 
<��nX�tM�n�X���K
	� 	K	�X�
JL
�	Y�
	K"��J  "5 t t < s	�<Y	YJY	uJY	wZ//�K=���~��<
X:�X�nZ�~�JM�~���
	���	� �
ZXY��~�
�
]��U�K<L��� �KM�L�<! Y <( � <I �K<�RJ	�fZ�;�I�X�~��mXJZ
������XP�l.X��^F	<<�~�~��oJ�
��1c����o����'�>'����Jt��
t
<%JJLXX� 
<����	KX��n��~�JM�~YX�
	���	� ��	����nX��;j�	�X�X;���~X� ��~
s�=tf	f�[z.!5.<fX`X
�"��6���Y
J�
P��pXZ�~�JM�~��t�J�	�fJ	� �
�!�TJh�rpCy.��
�rX���X��b�w%nfu%�%�%�#�#�v#RgX�6�|f�;� ��E�X�
J	Y�ot	��G�X�5�	��~�XX���~X�~X� ��nX��~�JM�~YX�
	���	� J��w [xJc[8u�Yy�_� <O�.
i.X\c<
X��<J��t��sX=K������YZe�XXhKJ�J  ...zt�sJ�X<<��t��X ...�Y<�t��J....Y��t�
� X� �xn<
�<<.`Y<L�s
�JX�sJ��
XJL�� �&	�rJ�
���	�J<�If	Kt:&
��
�tL�sJWJJ�
����sJJ
��J�e<thX.f<X<w�	�
t"h�<�
<�s�JWJJ�
��J�(��AWKA;(�%��
	�	K	K	K��
�st
��
��	�	K	K	K�.*&��X<%xJ�
�%<%X<��r�J�rJ�
��L
���
<��s� �st.�K43J.
�r�t��sY����	��~fS�b\9[7u�Yxf`��� 	P�@     �m/� �h
t3L.	�.3J	@�& X	�	u	�	�KK:	K.gtuw�XJJ zJ Q sJ   Z
��Lp+JT�(�XUEI
fo�� Y��!-�!�fo�/� �h
�
W1
X �D e�	�9J	O.�& X	�	=	Zk�uw�XJJ BJ ?J �J   Z
�XL(sJ�p�XEI�)Y�S!-�!�
I�f'Y�'� �wJ	<`<r��iJ=vT��XL	�d�Y���� ���<<=
 � t[K�.F�
��w{� �tX>% W < YM�  -X 	��@     f<� f <LJJ=^
>�wfB
,>g.[	=Z
�
iEc. `���>sK[>=S����=UPLY@;uK=<z�� �y��sX&F\^	�^t�!�^t�EZ
f�!Z��X]EZ�
QX �XJ(.  JI^J"X.r�HvLXb�(X�_���x	(>��MY
Q  .ti . .o�X
�� ��   ,  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/truetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  ttdriver.c   ttgload.c   ttgxvar.c   ttinterp.c   ttobjs.c   ttpload.c   ftcalc.h   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   tttables.h   ftcolor.h   ftmm.h   tttypes.h   ttgxvar.h   ttinterp.h   ttobjs.h   sfnt.h   svmm.h   svmetric.h   svtteng.h   svttglyf.h   svprop.h   ttdriver.h   fterrors.h   ftmemory.h   string.h   <built-in>    ftlist.h   ftoutln.h   stdlib.h     	P�@     �wu�xX	JfZ<;.w�<�; YO swX <p&JK�&7K&K�&GY[
M
OG�=�
	0	K<X�0�uWJ�"ggg�/�	�r���	fK4*�u�  u/  u+ u' r J u #  �nt t Z   " H >   �  u  �4 0 X .4 t�.�|�5�	<tXb9	<t<tp�	<t�u.�	
<tft�	�tf\> � �Xt�	*tXtX<tX<tXz<Y	AtftX�X�0 � �^x6 � �Yw	. � �zX � �u � �u � �o � t ty�y5 � �Xt�tv�tn�/ � ��X��r #<<Oy	�K�<u��X�X��X
f�][J=# wt�>H�=�ftj�J=2 yt�
��<Ju6<J� <Z��<Xx��-/	&J	u� $Jt�<i6<fJJ�LIsuud�.�<�	\J"<"o.Jo<	u� t�<g$w� <�<�	d�"�	u=��w&��=<IKKw��J1��w&��=<IKKw��J1�A�A��
�!��)J=K)J@IB=�
���
���q���!f���Stz�z��g<
�	�	�]f(ty�	�	�����rt�ZtJh"tg
Q<
<]u	u�J	Z2'X<ti<
<Y4�Xk.*�=t' t�
 J st
 J3 I�q�suX�f�u�L�<����;-iv;9?;qM?Y�=t�p@0<�J�
	��	L�[��Z
	�t9w:s$�v���Xt�~�
	��tv�~.� ��]<Z<J	�"��]f<�(�p�<g
M�H.fX	iXL$rt	>
�	�t<> WX J
Z�H� Y
	� f��~�J�~t�XK X�t=JJ=-K� �<� f�t<� <
f$J<���K	d��	u-	�� K X.. k.�K �*�% �I � I  �PXWuwx.���!	t��v�t<�
	2=I	=1c	/>�tZg.	i�2.	=?G�L	=>Y��	Lzt	=AX[*
J XMJ
�.� .1z.B�<.<��
k?�}v9W2 �# J���w�
<K
w	� �J��w
�K
w	�!�J��v��
�wtK
<M	��J�-�/fPXvXf
XK!u:u!Z�v��� �k�K!ve�u!Xp�?<?tJ6�JrL?<�v��	�M�v
�K
1	�#�	J�w� ==v	fqMi
	K� n�Zv�. ��zPJXZ���
$.X^<V
$�\.%)	(�+�+ �H s&�( �� <Z
f^#
�_
`
	X;J9 Y? W	XY(��� <�X� XX<...wX	tAJ<. <...� � X� .��^�]X ..t��<�]}yY�<X�f..��j�X
�
���[
�+ f	��X�X>f.% ^�		��< X+ ��.z
	yxt�
�XX�JJ���<-�L	J<�
�	>
X
Y;=
<LI/  Jkt
X�<t.�;��
	�u.KtJX.f.�	�yt�$�� J
Jut@P3�	��6U�
� �KX$ �. ��_!J
	Jwt>P3�$g�<� J�'/JJ.JK
t	Z�u?X .f	�J�3�i,
f	���Z
	Z�9Ks�+� t5�	\�L�31�L<<<
fK
K<w	�3�L
M	�3�L���3J�L<�3J?@<��	s� XA5t)	\�L�3?�L<<<<$�3<
�L<K
K<w	�3�L
M	�3�L��3	�L<��3�?@.X�	s$`� <t�LX�NF�<X���X���X�zf��vXX 	@A     �~g?Zt<X���������r�f�f �>rvZY�����X1p�wZ���X � ����X �t A[u ���FuZf	 � / d	 L   K ; �  �  �^��JZt	 u 1 e	 = �  �[��XX<.hw�zvr0X������H�
	Z� �  � �	 IZ��
J	Z��K;��K;�X�
J	Z��K;��K;�X�
J	Z+	I��K;�X����e� r� �a�
Cy.`sf_y<'yt'J<yXQJ�
�L@X . �y�=L��������!�ytuP��	!t	J!	�!Mtt������i~x�#1su1	K �G	WY0p���X l�g �q�Y]�M��b8#vX ���=tO��.0 � �z   
 J K 
  w	  � �J g '  f�
v���$�wt�wt��y*�*���y*�*���
6nXkz���t�������| � � z�h��<h��f..W��y���y<����t�~�.$�w�Y��Jt�	�3<JK%Iu%y�/KN��#ttJ!u�W��p.tX .Mp�"u%q�zt*"�t*�z�u�"�zT"�tv�}�|u����uv�j<Kus**��������f�
t J�&f;�
 � t
 i.�X .��%��%��{�
6x<�L
<XQ  .& yt# �M�Mv .�JX 	00A     �~zlKa�	Y��Nm<	�
�J�>//��.<
J	�nJn<JX<	/	Z� JZ=;�/K_�Q�d�)��	yJ;�X	/	[� JZ=;X/K]�
>
�K	;K
?<� �
.v.�K�Y�
�X<X<J�/��v
�		J� � 2 ; K X <	 ��1
h�!J	m�J � 2 ; K X <	 �z J �  �2 ; J	 .�	��	;X]��	�tZ
t	Y0ttp�#�	Ytjf	JfZV	>	Z:!@Xw �  /��tvX Jk��=XtfJX=..l ��uX�
�ut.�
JX
�u K
1	��
J/g� =�uX�
t�u 
.K
1	��
J�v�&UuuK&= ���YJ8M#t<��0YL�xJRZ��Y
�J�=
� 3* x JX�Y
Jf C�	MG����zJ�
f
�u"jqIY�t�
�!J
M-:
v!Uu!v
	/��S><L�
J�JJ=
�T
J�JJ=
z�XYJ=�z��;	�J	[;	=�<<!h)JJ�?
	f<	0J	[JJJ<t��~#FY�XZf...�~�z<B�0 r� � �  � <. � � Y 
� �	�J	�	g<	� �  J	 ; X�;<X	��� .	
�J	�	=K;<M<!e)JJJeZM
	J	LJ	�JJJ<J<X
g,h��	�����zfy�
�vJouuwYt0Y��|/�t�}���~��X�����Y�8��Y�X JX�|�.oX�uv�qXK;gfK� JX<.C�
M�;=X�6��X<.OX,X._
J�
J�NjrY;K)
� �H ��	 �  �. W � :	 � , W K	 �  y JJ-aXJJ	�<	X�JJf �  � �	 I[����<otL�`�f�fKq����}�r<>��������t�K��}�
�
K;=
YX���~<���~�
�
X<�X�}<�<[�}y��
 =.; �
 Y; W�X�}<�<[�}y�
= ;��X
�~<;W�Y;gE�U?&�A�<<
�b�<Z
�ta
�J���� ����;YX0
�.X	
�X		��
��X
��vV�J�
		�� J � �
 K!J	3<�f.<	�X�>J��f
XK
w	�0�J.<X	 uJ"X����<@ �~X X J X�<tYs. /  �' ; f\��n�
	��X�~��<[�}7	���� �   �, -  = �	 J�� �  �, - =	 � �X	�X	�	F�J	. �  �, - =	 �(� �X	���. v   �g   
 X K 
  w	  �+ �J) < X+ z	 f � X�H�Ld>h:��

<s�[L
RxtVZ
�xX
RxXM
X
�<v�X�*��X���}�iJ
.v<�KX�KL�+�'X \� 
Z <v
�M
fNut[	 Y  ; K f s X��6.=u
zr<L
XJ	Jt�<�� ..
 �~�# ��h�
�XJ
 K1 �
 Y1 s�	J
�
X<��L�
JX
<- � tm
<�
�
XX
 �3 �
 K3 s�7JX� J��X
�
XJi ��
1X
<jLdLf	v�JX �% � K% W�%�	 �$  h J/ t J$ J J/ t$ 
< L! tJ$ 
X	 K$ 	 �  t �/uXX
�
XJi t�$>$rJL
��
�X
f g6 � Y6 sh6�Y6sk
	�

�
�X
JjL	�X�X<	i2 � < JJ�
 X
Jl+ . �L^GX �   J, wJ  	� J, w J	 J- A� J� X�X� Jf4w 	JJ4w<	 < �g�
fv<�9uuKOK	"�B
<�
X	���Igf
	�
p@�2J	K<y<K�� <KKL�f!
�
J�-tJv��K@82
\
0e�
�	�@
<��hJX..��	�=
vJ	<��K;	Kv.
.JJ	h�<�$�Ig$g���=��	�?G�IK;	K�WK�	Ku�KI	KtJh�=$XJ�B-
Y;�$%:tJFX2%JX5z�'=��{�@�.�JYp�O0r.�#	t.X
��2�=�<.�Ny�4�=�� f�y�<2
 �L V �	 Z   �  � xX/�o�
XnLX�	��~!���	��y�- gt��tZ
	Y(./
	Y(J=
	Y(J=
	Y(J<wt
	Yg
	Yu
	Yw�l��t
Xt^x)uuhv uu�u�/�%eu JM$�JZ
- X	ht-�&?q	t-hd	v	/&	N*	K	�	L�P<X�	�/	��um u�P u��JZ<XJJz<Xtt�ZMULJJj<tXZ�JJ��<tttJZ<XJJz<Xtt�JZ<XJJz<Xtt��Z<@fJ\<?L:=t �ZF=.;N<JN<.w>:=t�	�< Xz� /B s6L:�@ImvklJu�
�	�v���
�	i!
	Y��
�	k!"
	Y<t< jX+����
m.�3�tt���uM8=t�<tY0t2I0[2e\%J	���
	��.,<,t<tfwu���X�<
	�� ��^<�f��!	�t��uM0tp=�
J	��Q�.>�Q<<<<
<K
K<w	�.�Q
M	�.�Q���.J�Q<�.J>?.<��_<��!	E�	��Qt
.K
1	��.J<�ktȬ.�ft.)<9=>)JJ/�
�(�t�	x(F�<�	\(<<	jf�eX��BJ<	uJZ>ZY@�	uJ�dJ+�X<Jbf
	v&	w	��e��e.
.Y
w	��J.<&tXx<=&Cv<=&	<f<f<�fu"qtwj�L�� .  � K  � X G^z. � t, /1 : J
	��<tX
<X
�XPX������u�}t
 �/ � Pt
 1�/ W
�/�
u/I�
w%:#IM
� 
 @= �
Np�
X
tX
 �; �
 u; W
�R�
.�;Wt��;gX? �2 �A ;
�iX��
�
�X
g3�
�3W�f� ��X �  � K  � X G^'� .�~�'���.� f'�����;KX0
�.X		��
��B
���V�J � f L
  <		f17�N7r�Xj]!fa�!< ��	� �. 0  =  � �	 G�	.�b�<	�0".w�JL�b�XJ�b<
JK
w	� �J<=�b
�K
<M	� �J<( uJ	 <��|�u�&�Y"X/J"<J�	�;Y6<�X�	�(3=;K3J% t <	 J�YTKLK[
�k��6 ��5<JX�}y���������}�y�?����}��.
	��� � � f J@ �}� � t X �	�� .  M G � K  � V J Z  J . =  f zJ
X��	�~� =   �, ;  K �	 <Z� =  �, ; K	 � �AH�d> X < < L  i G [   J Z � J M  
  � ��
 � � Xvf
Xut
�3W
�3W �	�wX	< �  �, ; K	 � �����}��X���}�"�X?		LX��.�<qJ���tt.� f�~,<X,J<!Xg!���YJXG|Y"U<J��f.<X��3=;K3JJ	 t<��b�XKL�b�
K
w	�N
F�J=�b
<M	��J?
����6 ��5<JX4 �  . �6 ��5<!J/ xX �6 � �5<!J/ xX �	�~	���	�~f
X�~<t�Y�~J� J<XX��of�I9�Z
+tL-tLm�K�stKJZ@J<�Xw
���{<nt�o�JX0I��<� X[�������szJA/";#=;�~"��#�FX!�:t[���v=�
J���mJ=�g�=f0K<���@8  J�[�
4 �	�Xh�$�l�?Jg�	�	�
Jv�	�	�	�	�	�	�	�	�	�	�X	y	�	�	�	�	�	�	�	�	��Y;=I	>Y==If
	��sJJ
XK
w	��J	g�s
tK
w	��J	��s
tK
w	�x
F�J	��s
w	�x
F�J	��s
w	��J	��s
tK
1	��J���yut�J8J<��{X%��=�:>�	w<wJY��
tXw
��:vh
A  � f 8 s	z	���yX.;
=	�OS	�u�g$Mp	�!�#tz�	z#	g�
��1,zzJ;�{J#�X2�{t#�f,�{t#�Ju�{;fv2tv,6i,Gtu.-uK<u�w*uut�/�";�M>�v��w
�}�[	�#w���u
���xK7�#
~jvXu<#J�#u#u#0#!Z�!�!�!�8N
�i�5<
�<�+L	3!�FJ:<!JKL	���<>�x#�<
�yJK
w	��Ju�x
JK
w	��Jq
X
fM�
�
��.r�y�t�u
���
�}X0�}�tv�v#
vt
J�}Z
.
�&
O7X��
X	�	��=�v�
�t
<�gfX�X
<uJt
f	YD�I>
	YF�Ii
	� �
�z<	�y
	j	uxZ����x#�<(J
�yJK
w	�3�J:<��x
JK
w	�3�J:<��
��<	 � ( I J\�
X	
�
J5\58KIY5[fu
�w9[g
4 �	�(X(uJm�(x�	NFCyJ	�	�	�X �: ( �: ;h:#�:Wh:#�:;sfX	�	� O! . }! O K!  �  Y  X J f	 xt t J"XX	i�"XJ	="J	K[F	K	>"<tt	="t	K
9	Y	Z"Jt�	="t	K
<u<F	Y	Z"<tt	="t	K	w�	Y	Zz���	�XXtt	n	Zr	v0htYe=. 7 J	 J	tf&�=JKV	K&=I	u	vZ&V=I	uzf	u&=I	u	xY?�H	?Y?�H	k�X��X��X����
J	��qJ
JK
w	��J	g�q
tK
w	��J	��q
tK
w	�\�J	��q
tK
w	��J	��q
tK
w	��J	��q
tK
w	��J�
	�[G	uz<	L	Y<	M[�~��<��z�u	J;K
��!)J=;K
I=
>	=I=	J� ���	 AJ�vwp�F9
XxX�F\Hzf`v.JK`w<uZ[ZXx�[U?JZYVM�Ku[TuxFu�Kw���xK5<��7t�$JJ�
�
�4�
J	�)	��w
JK
w	�N
FJ�	=�w
w	��J	>��p<tgJLJJ�M�~	�	ux�}Xd���~~v~vuVuuVuu����'�J�'XX.���{���X�X	�w	uxX�	JX	�W	K��X�	�� ]X�X	�	K	�	�.�j�yM��f,X�,t�,u,u,*0,VZ*K*f�*f�*f�K
X	�tXX	� "V	> �w�
<J �	\�w��wX
.Jw	
�?
G�J	=�w	��J<X� �w�	�	�	w	��zX�+�o./n<.oJ<nJ�JKL<<H?IHKK=:K=>��@�<<z	<h<hJX	>%f	M[Y	<h<hJXJ <..Mt	Z%f	M�	Dr<rJ	Z%f	M[�J_�J�5�J<�5<�J<
.K
w	�5��Jf�5JX&�W�&;=WXX��n
����	�sgJY�Y�Z�=9L�&:�0�/'�/X4t"<4 �" .	�;K*<K�& ���
 ��
t	�{� X��sgY�#X	>:	>J�~�
-JXX���.�tJXv<h�~�-M<�tJ	X\$I�~<M
-J����K�~<[
-J�X���~X
�Jf��~��	�<I[	K"-=��J	��y�K�y
�<ht�0
	�X��
<ft<M<��
	LL	$7�	\.|t .	^f�"^J." X�
�sLqX<�JX	j�(dJJX>F[
��<
J	Y%I<(j%J;XtjJX<!XJ%tI[
X:	Xh"X:2h.5t2�J�25tJ3�	J*V0JJfff	[�$;<XȞ58*wJ0J	J(�BWSCqz�^��>� t�tYuY�0��� X�<� <p<XXpJJZJ�.�.t�����
t�	mZwX>	^	zJZ9LM>%�	 �& 	 =% J 9^1�>�_���	 � 	 K
  qJ	ZG	?�xJ	|
qJXX<t�|t�f
t	N�	J
����@X
t�	w 
X�t��st���1�}xXJ\1�1x[yXQ�
t�	U	OlXt	_>lJOm�>xNLMXL.%M	 �& 	 =% J 9^1��>	 � 	 =  J G`�
X�
ti	�K	hf	��	K,�E	K�	K�	K	�
<	/,
J,<J	=,
J,<J	=
<	u
<	L�	ZJ" fiK	J
I	KI�:�
.�
!�� .
	�	vJ	��K	i�L.�$XJLGKv= � 3 I. J K I X�vutp�L�u�
��[
X.
tJ
��
Gw&
J
�Jj
<
�<:�
�:;
h:�
�:Wj�G�]GXx�
"�
�Jj
<
�J��*�;K<J�0�;=Y;YZVZ
.�9<3=G�!z�JtXt, �$ t�YIu=U�9�G[� �� 	i<	��;	u	Z	= ! * ; K X	 I\w	 0�2 ��	 � J8 �J	 � J �  :	 Z! �X � � X��
Xt
t	� �	�9	?Z ���tu� ��X�w	���&K;KJ?0�
	Y<J!zJX�	�trnt�Z	�L�L%
��%
� �X ��JX6X	fJ�	�	"�% � . <Vz�<
X	�O6JJ;	��	���	HX
		�	�J�JK�� � J �z<         �.<=JJIwtJ�tI[��J	JhJH.Z1<.�J .1tJ3�	<#VJJX�JLl..	g�r��rX<
<K
w	��J<t zJJL
�	Y�r�X��X���z�5F(@IERX�����Z	%�	��X	K �	�z��	��	��1�	J����t
J� Je 	� �	K�X
#��
&�o��w�
c�
Jc�
X�J	��
�
Y��C8JX	�Y/WJ=e
�*W*g)J�#0L
_vfu
x�K
0y<
_Jy�
����
J��..<	�1 �/tX .	Lt3�X�
	�	���z.X�<.vV3e�.J�x�
J�JJ��x��
J��..<	h1 �tA./� X	L�
)�
t�K���<J.i	.�+�Y I/ I6<;<9H?K	Q,v<X�<X\J�
J���Xwtp��LxJ��dֺ<
J	h	KX E�	.
t�?	��	�JhKXEX"�
�JMt���KMK3�KX<.W�	�K	�JZ=/S*JJ��tt
JJ
fJ
Jh<Xd.� t�fx`t�MMxJ
J'y.u':JJZt�
N�[�M[
	M�X x�.�6/I>C�vXI�.
X��z&t����K�	 <"  J J I 	X t J   t I[/�.xJ	 �  t Ib�
t��
�~fz&t����K�	 <,  J J I 	X t J   t I[/�.xJ	 �  t Ib�
t��
�qfo#.o.#.oJ�JKIY*<;X�t���5XB5zfZ5L<JNy�_�!at/X7JJJ	\%<J$Y1I\(<(<J(K�[0J�\H(�<�4�z�?M�3J�z�
JK
1�	�z��J1XI<<X��Hbt.k.t3DJ;. ��x�.�
t&KIKJ>w�-�0WW)���X!_JXL��=&I]
	Z,t	[<�!cJXcXf'�(��7q�F	�)�3]��(!C*�F>)�F*HF>*,D*x.�F!X��b�MX��a��z�u.	�vuXJJY
��
X.�<1P+v���iu�tFm�XN /� J���~J��}JY
������~��z�vfdWW\�ft"J)+fX#'��
X	gY
X	uY
X	uY
c�"rXXnJiX���	�Xh�<�h����~`x�KfKJX��
J�
t��
 J��}u�����~u��-��
t�~�J�w.� � � � � ��}�~�
 �.UX
#f
]XXMy�| ;KX-��.Y,�)s=,<.-t[��"�[=X"�`gX�� 
X�uu�n�J)<%�'Ig�
!X_f!X
�
�t_�&XZX&<
.<
J�&#fKz<	XWgsuJ� ��� �� X�~�����	� �{�
��
t	��uV��h
�ytX!AJL
-�

�X
�|�1	� .	��|..X	��	/	��X�}Y�uX1�
 ���
�t�t�Y�uX1�
 ��{����,WW��}
�yt�	�/ ��~��=?��
	��+zfJ�Jh
��	�{	
.	.'�q#BzX	?!J	>#	YT-
X�w!X<J<%	JX	^ZAKAWJuX	��� �<.'Hu.!��	�	K@� ���t$T/�YMK.X �p�=u�LZL�.<J� X�f��L�.<M^
�M
X�
 Y �) sNf�
J
 �+ �
 Y+ ;��ZX�
J�XN�X
t	Z!z<	P!	�!z<	P!xMXX�
J�~�t���~�J
�~<u<Z
Xf� J� 
�~�*�
K*;
L*�
K*sN�
|�
�M
%z�/,V<Y3;
<*w<=-.n�7
.	�XJ	�$xJ`<x�$x<J`.xX.0
	�J>:>8J
J	�&VJ*J<�J� 
���y5 x�! � t�L
�
�XJXM
UF.f\
	�#.!X�
�^JZ"=[GM=<��J� .X�	H�	Yo<	Yz�#X!X� X� 	�A     vt 	 �A     �|y_yX_X=XJ .pXZY\�Z<K
	YjJ*. 	��A     �{gwX	 wX	J.�'JY�tZ<
	
J.

�`f.	v�%
<f.	`X(Xt�Jr	�K	:ZZKW�;K�>�J- ��<JuJv	=I=	JC	y<C^�i�r<�Xaf
	��cXtJX*/Xi ;<�r.���"[#*.V.
% ��zt4z��Z�<f�Z
�����#�V�D�!I	t�Z!�u���������T���X�!�+�|<f�t)Ji<.t)�
t�.
<�<�<Jf<N
f
J	�4<BJ"�<O
�%[J�	$�	K�J�ZL��
6���<;�L
�
J�t
t
��	�z�J	�2'fJ����dJ!��;L	t	�zJ��6$.J	J
�}��X��J	�zJ	�K f , �( �, < .	 �Z�J'!�# ����� �f, s#�,*�%#��U��s��[�wX�S�wX�X�X�-���
	��-su(JM%�J�  f�t�'1u*qJv'/1N'*K'�'L�I<Ȃ�6�.�~��~��l�
����	3tr.��I����4�Z����y���)�t
LUK-*
Py�-Qw -
J
�tJXJMc[G�L�L�zwX?q[g�BS�z<=z^�]X Z�>vX
Xv�
f
X�
XuJ<
�<ut3�X<�	�	uH�J�?	H��OJ�
�c�����d�!�IK��d�!�IK��d�]J
tK
w	�"�"J���dJ ���VJJ�)�VKKIKJ��)�V��)�U��)�c%</-KZZ�������X��dHK�q� pLJXX��dHK�q��pLJX�X��c
f���c
f�u;u���WM
�	��J�(�WM
����'�z��nJ�k.Z �t�	<�	f<J��J���^t��<
Jv���Iu��$;L�~X�W;9�u��<X��
J�'�W;9t��(�VX�*�WKGKKf�'�V��*�c����c����fKJ�J<v
S
A�.u��
�	�'%J.��c����Y��&�cJ����[J�2��%�d����rt3�.mt	��j ��$L
	
�	60�<	<t���mL
�3�
����G�9?9y��������l,t�
=�=
X>	(� �� ��$L
� �
�(�	�IX�G�&�!�E��X���k���kJ��
%�-[-�$���	��G�
#���k
%�	{�j �$I�L
	��f��`!
vr��R�u�I[����n*J.t�1Js�)tW<)Xt�.h<�<<r�L	��<<<J�����`!
vr��xJRv���k�#K1W8<�.��;��� �cJ����w?U
uNE=	�oJ
��H�	Y
	
�L$�<J	>
�	��>�=;JJ?9Kt>t���iJ[��~K8���V ��(�_
sK
f�!su�.JL	�I!�<X�t��#rCy<Jv/%�KKIK,v�l<Ȃ��!
	�J��uJ���>���
�eL�	#(Jf(t<x�)��eL
��
J	�t<J����XM����'�XM�֐�)�]t�su<JLY&J
J�
JWJ\[
��N�sK!ZpK;KJY���t	�}	��� '%J[J�	$�	K���y=
t�J�	=�JI���w$?
��X�	CX�	
<X�		< X�	C#�	��
#X	�	<

$�	�� f���dL�*M	�%<%u;KI=%=%t?9?�=
Cy<C
��?�m��uw��
>:>
�<h?�m����dJ���e����T
��tJ�+�eL�)M	�<t
J	�&<JX��\� t	�suI<JKZ
Jt
JVJ^[
���#uU=#WIKKr�Yt�� ���!�^
sK
f�!su�.JL!X<!t<	YI[
��t�!rCy<Jv/#u#�LHK,v�m<JJ��X�!�U�sX�+�<��y���Y
��
��	���%�U�J�*�U�J�*�U�J�*�U�J�*�X�)��V��'�c���VJ�)�VJ�t�)�U��*�U�� fJ�(�d��d��d
�w�<qf
��	�	K.�#�hJp���hJ[���iJpX��e����c���g
��t�	�	�o ��$L
		�<t<f��WJ�J�&�tK�*L��t:�H>)=;u)<fJ���WM��ht
JK�
�htw	��Jf�)�gJ>
��5X#�K�#X��#X��5X#�K�$X��$�����gJ�+ ��h
��K
L/0)D�;=����h
��K
L/0)D�;=����cJ����U>����*�U6�><���)�ZJ �
�����~�UJ��*�U��*�U��*�UJ��+��T��+�WJ��'�c��U��+�����^
>rZ
<�.I�	�f��KX�		�W�J	w�	KX�
	��W��J�hXKI�X	�z5���&�gX��!���J�VX
	���)�l�
� �����{X��Q�<XxXJ�*��f��	�	"	�J�s
%�����	��G�
#����e�[X&�����m���[XapX�
	��W��J	�eXpX&���t�u
�X�~�n.<Ȃ��&<JJ	�	��	�|	��	�t<MX	�	� ���� ���[X��=	J2K,<�X���JY�t��<t	�!�L!�.!<>ZHh.�p	J2K,J�X	�~	���	�X�"��dXX.Xi-X.X�r > �<�	V>\!J!J��	�2NX	�1�	��fX�X��^
h���L���j�#K1W8<�.�[�	KtI��p-�.X	�z X
�4tpKw���Z�%/�Z.<�%<=�Z..�%
�Z<K
�%J
�Z<<w�%�Z
M�%	�Z���%�=><<JX
�,�!��-t�X�t�!t;L�IX��X��#�cXsKc?�<JX
�X�X
n<
o�<
oXX�?��Y[X�t=I=X��X�X���Zt
.K
1	��%J<X	� �;<�mX	��;<�m�o�ym�M
�X
J<��}K
d�
X
JtO���}<����u��X �}J���/��z	XoX$	tJ�z�O.A" f�XLx.=KKL��X .J.lXZ�?���}�
f, �% f�L.Nu
�
<	<!� t	�.�
	$��	fh��	J	Yu�
	�
��sut	�~f�u��Dt	�X�u�XYv���X��XW��Xr��XY���XZU�&�X
.\<v
"&^��& v&�h o�u
toX
td.�x	$�$�$�$�
X
�t
�M�
�Ms
�M�
�Ms
�M�
�Ms��xX
�9��
�x�Xw
�xU����x<�JZ�x�
X��
X
�t
�6(
�6s��`J��Ki	X�}X��T�v
�}�t�}��<%�1D�}J�X1�u�}�X_y<��}J�<+t�}<Y�
X$X^bXtef$fsbt�$\<������������z*u*t��z*�*���z*�*��f��| m ytg ��������z��f��
t�uXvv	V!	�!	�!	�!�E	Xt�	Kt;[�%:iXtV�ZJ�	�
	Zzz<^� �!� � X1.t�)uh'�	!�~�� t���	���rX�zuu���X
t�h�X
�y6�
�6s
�6�
�6s
�6%
�6s��X�x��u���v
.vX
fvt
J2 �
�2I
���|J�J�|J��Y�|t�JmyJC�!�X;u��;X�9G��9G��%G��9G��9G��%G��
	�*	g*	f�	?J�Y/�~��,�T$�K$N,u�j
XK
w	�*�Jv,��j
<K
1	�*�Jf� �J�{���
<	:���d^�M����X=�
 	mQy�	3	��
<	0��##"u��y[��z�w��t�X�&'�Y&UL#�!xJK!K!PIl[9�s�fK
t#
W����KP
2�	��	Mg(u7s.	Bf�		�!XtZ"HZX"T�"GY2�YX M
	��nX<<
K
Kw	
�w	H��	=�n�JB%#LK%G#<L��~�� �- I�- � �- d�z @� �{�<��
��f	�=I	g�{./u9s.<X��"u	�z�M�*	M*� �� X���!<t	���/0/6t�YZY`j�j!tJ�XX����kX!�f��kf!���k
K'�
�k�J<f'�$�
�k�;$�Jv
�k�M	%���k����k
w	���k<���k
fK
w	����k
w	���X#�n[xJ	{<� J\	�tg(0<�	�*	g* �"v�l�?K�� Y3 s�]K
�\ZfJ{ X H O  fr� � H O  f	o�?�Jg�X�X�"X �K   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/type1 /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  t1afm.c   t1driver.c   t1load.c   t1objs.c   t1gload.c   ftcalc.h   t1parse.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   t1objs.h   tttables.h   ftcolor.h   ftmm.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   fterrors.h   t1driver.h   t1parse.h   t1load.h   svmm.h   svgldict.h   svpostnm.h   svpsinfo.h   svprop.h   svkern.h   ftstream.h   ftmemory.h   string.h   <built-in>    ftoutln.h   stdlib.h     	��A     � Y-J=t?>�@�u*�LP�k�=�?+>�uZ"K0,>+=	 �  *  �	 Y + � <	 Y/ + � X X J xXnfX�<u��<(uttt	 <? ! J J IXoJ
�n 	<�KX	 </ ! J J I[�t	 <!  t I[
J	Ky/ 	bw/ efX�u�
.<^.Y�. <-  J J I� �  t I[
>u�=X}X��$K-$=J<<f �f"v
��	J>	> X < <Zi9?@#t>
  X <	Z:	u-	KXXX.yXz.ZxXX.�vf!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��|�kKv]t9�Z
	Z	g%���~J�K]urt�"t	J8�zz�JXX�
	�>!Y	s�#Z#r	�	�O8N8~v�f�% � Jv�I��YI�Z�LVZJ?)'�K)'�K)'�Jt  ....	@tp�0�=<tw
�  ��Y_LJ
�	Y:J	t�QX�.sJ3ww<$�J�	.wJ	<�"c�"p.�u����h�v��
X J	gH E <
�J��...	�u.<ft��$JJt�	.�"q�"�u������	z<vxJZ�
	K�xfX).OJ	 � 	 v   F`�~�lpu���
.J �IY <.J	Et( �D ��D��D%	�=	� 	� us	u 	v �=  �! s ==  u! s u= ! J	 p_f�Z!��=" ��X<f��XX<�
JM(�3�
�M�	 K@ 5 � �\�t.tX�yu<X�LVO	t X <
QuX!�=��SJ��
LsJt=ZJJNX 4.  ) N � =  � ) �' ; u I M   wJfW=l�I=Z�}�^uX X��LLV�
�
<~�oYJY�	�	Z�	g	KW	KL��	��t	
J�	yJ �  ( L � =  � ( �& J K  	 x
t&M�f6�"X="�Kb<�Q�  XuX(w<vX�U[L���?UYJZX.K�Ev���ZgK;KM
t�
�
&�.�>t	 L  2  K! L t2 � M G	 =2  J	 L!  K W	 = ! J J <	 >   rt!HX�f;���Kf�x��JX�rvX�dvXX 	0B     �.�w�z=AE=<X�	 �  t I\���X��X�	  	 � 	 �  � F`�$��	 Y  � �	 z   � X �  J z	X��a.���X��X�	�	�	����ArL<=	=	�
J<��
J � �H W	�#	���~f�
	�u��LQu
\ct
�	Z���Xs� X�-u�u
J	�	K�J  ....l�J YK ;	M#	�#�~X��X J..s�J �N ;	�#	�# �~�? '�?s	�<�<	 � % - = ;�v<	�f	t�t	�	�<Z� u ;=M%<�J�	0�t<	�J! J JZ! �� Xu�	/	�X JJ	�~�IWhAx� �H>/ Xy�"��DL!;=K<��2�$@2�@$"�L�#-�3.�Jh�& X�&� �!�!���Ku./%��v"�KY� Y8 s
�<?���
<Fj!v<�2�."�s<B"{s<Z"�y<	�wJ	<�"d<"u�fwXu"qJxf� p��������yU��Y��W!�
kE=�
	�ʀ	��G	K.v.V	Li?A� IL&	
J	� X�"	�)  ���}J
XK
1	�N"�Jh�}
XK
1	�"�J	jX�� K 	N5 tw ���}
JK
w	�"�Jg�}
JK
w	�"�Jf	�+%X�G	K%X?L%EX	L��J� J��~J.0��	� <~	wZ�	�%[U	�%YI�I	K%X� �)�2�Z8J<���� o�X�~��fB��Jy� 	t �}   5 �<
 �}J K 
  w	  � �J u �}   
 J K 
  w	  � �J q Qʀ�) ��}�z�	XwJytuZ<X���x��X��X��X��X��X��X��X��X��X��X��Y���X��X��X��X��X��Xp�Y
���X ��~�!fF&�z.&P. H X>
�	KF2  �I/  W/� z �yJP=yX7Kv><�d�;� � � . � ��'	� JYJE<
t�~<Z
J J � . � � � X�JX��~f J � f � �	�tK(	�J�f	ZuJ�f�$ J JE � �	�1W	=1�t���w$ J JE ��J$ � J	�	L;	=/J	�&.<	h"< Y)xffW?�J�=� g9 ��9��v��Z�<G-��v�t�JXX�xy�wt�K� $�M��(�<�vXY-Xh7>
d>
:	3t	+tu.X�-XA.
	Z	u.3Z-W�!.Z-WYwXY-XsX
	Z	u.mX
	�	u.�v�z4z.=vXX
<JL
tlMX ..	x �JK��	.wX	�w<M��L��	��K�FuwXY
	Z�
� M  . � t Y  J ^h
<	Yv%u
fc3XK����AO=zJY	tw<Z=�X.'<Ok �_�+tUtYtYt)XS�� fv=
�
J X �	�J	� J�u
<�
�
k	�	�7���	�.x�WJ.u�	<�t	K	� �&X J&<	[ uG e �G �  	`&� �2 ;��JJ�!KY��=;Yv�LX	nJtI�� �wUw<
>f�[+��M
�"M
��K
�XXL
��M
�"
 �  �f.J�~�<	K	M
J��	�J ��	�X�K�J�}�$XJ$�<.L
M$<L
P$<.K
 ��G ;
���M
�"M
�X$M
�$M
�$M
�&M
��M
��
�|XDoK9[??93 f�JK�,J<+ Y <C .H IX
�L
fu��� t�<� XN�$X$�<.K

� <
J	.�	��J	�!KYst=;	Y	vd	LXJ
	_�[w<L 
J �C ��vv�>5t
��u
�v <
J gD �	Muy
t	Z�	;Y
�$
�	�J���ff.�~JKu
<6 f	Z��ff. XKff.	� ���	M�	K�t�&�<[Jh(
Jt�(J
X �
X�s ��	
Jt< tf
J,=K^,yJ;NK>ID
w<(<��.uXL	uXMu<Jh�Z�
��'�rvY�KY�YY�YY�YXY)JZMNt/tu��XR�u�uX O�u0X �z<XX 	�3B     �}�u��.		�J<) w <v*f�
i
JZ�	Y)u<<tI/J...	xtA"H�hJXJ�~�.hV.Lvt���u�E�
	/2tx�
	/1tx�
	/0txX
	!/t;��
	�<	Y�!r��
Xw��
Xw��
�w��
�b�
	/2txX
	/2tnX
	�/A .AX �o�
	!2t�
	/1fn�
	!2t��
	/DtxX
	/Ct	[Xt�.X\�/		 X ��$*�<=�J�,X��� .�}�
	/#fp�
;  	�6t.t	YW<K���*r
	/,%fq�
	�(.�<	=".oX
	�/t.x�
	/#fx�
	/1fu��
�z�
	!$t`�
	���u.�<�~�
	!$t��
	�/t�|X
	���u��
	!2to�
	!2tu�%
t	�/A .AX �#�
	!2tK�
	/1fr�
	/34�%
t	�/H .HX ��
	!2tu�%
t	�/A .AX ��%
t	�/B .BX ���
	!2tr�
	/1fo�%
t	�/A .AX �v�
	�2t4�%
t	��B .BX ������|�uTuTuXu]uTu�~�J=.t.<JZ� qu�Y�|J7..OE@!:L<	XJoZ<<"t�J=�>
`
	[JmX�	�|�KI	=	L��|J
�J
��	�#1�?JLJ$=1<><g#1�?JMJ$K1J>JIL#1�?JMJ$K1J>JIL#1�?JMJ%K3J@JIMj�"u"��
�"/J<<g"/�<JJK"/�<JJ��gv�t<<<\� �  � IL�X !  t I\I/  �lJX.�X�v�t<<<��� K  � X IZ�f /  t I\I/f..kJX.�|J!uwXXK0J� R�
�<JO%IL�~,LG=L� /I KI=K N p9K;K=U?FM
[
J	�� q�X�\ �  X J t � X Ix��fntJ	K�J	�.�s.oX�N�<v�
��Y�t<*\	
�	K=;=	�]	��~
.K
<M	�J�JX	?Z=zJ�
	h!	K!XJ^�X..�R�.X��u�J�y�KK
X	�\J	�	�t�	�	N	^J	 � 3 n JX	 `  X J J N5JYMJ�y�<Y<	<	g�1J��t	8HJ�X�t<Y�P��t� �� Y   IM�fJ�~�= @tYMK.  ��J. 	GB     �{'�uJZ,�!<Y>Z. 2Xt ><[ c?ZY6J3 <.Y� �<�2Z?Ys�
	K'�XY�JbP<Y
	Y6	Jh%� ta�z�y<l�f"��HX>�
X�0�v0�Jr���>Ko�Z<Z�
 
J<� J�KX<f
 �� �) INxp%��J�.O
JL
J b: N �	Q�b"tT	Ya("XG	�	=W	K 	J@
JJL,;�K;�L0;��0;��8C�Ju8C�Jv
	�	Y7	u[c�:;	��~JsJ�YJ�J<�<YJ���<>�J�J�=<<��
�<
X�j	<w<�ztBYLJ>
r>
J�XZ�LXY;/��	[G�s.KxX��K�$�� ��~X�� JȻ� t��	�Ys	Kf��z
^z.
�XJX .jJ!P � �M�L�Z:�XNX .��yc.�nt�.�mX�.�wT5utV�X5wt�P�<<*�m�<�m��<w��m�J�m�0Av��������XK�
� ��Gf�N��~~�X�ȑȑȑȓ���n�����n��i��K��l� K
�
��JK��
��X�3�to�H��N�n���
�X
��6;��!��/�n�HYY/[��L��nz����� f��=J	�	Kn�	uW\����!#H<ZZ	�	�pX	�YI[fggh.��:ZuWY7X<7<<�#�,:�,X.;#�9�
��Z
		f	�	�	�	�
�
J�;�Y%�"�%X�;�Y%�"�%X	�%J;	Y	�#[	�#<�	��=�K�K�L!/��Y/IY��K��L�zt�+ �F �M�t �J eK\.�B&Ku�t#�<	K	$J � X

t���v0{y�u�����wt��s��u��!��uB!�B�!<u7f����n�L
V����mgX�	
�Z:	��u�	�	K	�X
	�����n�2]27K���
����t/7�t6��6�[w�	�Y��yX	�.\*	N.	�.	��Y.� X X>M�6v�6�Y4�2F��ȺX�X"�"�"��
	�	[�Jt��t�n
�B��\	�<	�s�	�	KL�X��	�nJvXX	� XW*�	��~<s�Xq�vtXXVs<t�v�t�z<w���ffu�K
�oO
	/�
	�
�u�K
	�	u�L<���tJJ�


��
t	/�
	ZJ �2 ;�<upu�<KIK1rL1u<s1KwpK<Jw
#0<Fu*/9v
u<	4yu<�		[� �!�
	�	Kr�	M	Z	� K9 <	�c	�	�W�WY	Y�.<�t	�~ttYM	��Q�
PP�JKJ�JJ���~J�f < .	�t�� �W�WY��~J�f fJ�</�%J.��$P�zX�.� W�WYk�-�IY �Z   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/cff /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  cffcmap.c   cffdrivr.c   cffparse.c   cffload.c   cffobjs.c   ftcalc.h   cffgload.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   svpscmap.h   pshints.h   fthash.h   t1types.h   cfftypes.h   tttables.h   ftcolor.h   ftmm.h   tttypes.h   cffotypes.h   cffcmap.h   cffparse.h   fterrors.h   ftstream.h   sfnt.h   psaux.h   svcid.h   svpsinfo.h   svpostnm.h   svttcmap.h   svcfftl.h   cffdrivr.h   svmm.h   svmetric.h   svgldict.h   svprop.h   ftmemory.h   string.h   <built-in>    ftoutln.h     	``B     %zB���1�fM�12h�		�	K	Pt	J�xJ/4f=?uy�v1J[<t�X�`�=wt< 	paB     =wt< 	�aB     �wu�xX	JfZ<;.��<��tw>Z
	�<.�	vz4Z
�
V4
^f
.	Yt	.J�&�t< 	pbB     t< 	�bB     t< 	�bB     t< 	�bB     t< 	�bB     t< 	�bB     t< 	�bB     t< 	�bB      t. 	�bB     t< 	 cB     �y=
_

X�f.v<C	2	J-�.f5X.pX
J	Jm.	��	-X� #tJ <'.<
.WJJ	+	&J-�.f.+J5XJ.J��	-X� "fJ&<J.� � .���J[1�C>.Rf#
X		�)EO}	=f	K[WKJ�L�=J>
J	>X�W
.K	�	K h+#;K+=#=��t< 	�dB     
wYK�v�!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��w�":A�X�u ���JZt	 � . e	 = �  �[�G�Zf	 g , e	 K �  �[��XX�z�gK�]t9�Z
	Z	g%���}�>�>*#tK Y  � IM*#tK �  � IM+$tK �  � IM1*tK �%  � IM��� � �*#tu �  � IM+$tu �  � IM�!����<W[
QUM
	/tZ���f ��6Jx� %<XuJuO<%zJY�
 X <	YzJl z �iJ.  [�<gu(�ufrf�,�Y �
 X <	YF@ . 	�iB     �}v
YXqf
	L
	M�~	-f�Ke=;K
h	��gJ
	L
	M�~	-f�p<�X <�~�X	��� J;KJ�W)< �� ��� <�<LJ�=
	��ifZ!�!<>Z�g�<YI.g	2K�~�� �zfqf	LM�~	-�	�Ke=;	K	��$J<iJ	�fS.qf	LM�~	-�	�Ke=;	K	��kJ	�� J;KJ5 �
J	K�zB	9�#<�.<��IYI=AX�� �fPX
h
�
x�<
m
		X<	�.<T�=IYI=TX<XX=<1<	� ��e	=	#<�X	�<X<	oX'<=;.	���w	�ut��X<�J�	�/�f�J�~
[
�(tJJht<L
	w<<`�+J��
 X J�<�X	`� `J f  `J. 	�nB     ��z<�z�fXD�H^
�X�P=I u" ' J1 I Ji=jr�
�X<
.X�� 	<wX9 .X9t X9v.GO.J<J7W
X�~�����X�~<JJo<X��
j<8Jw
�
u�W	X<=
JX��+M�.t1J<=

�
J	>	g 3   �J �>
	Z	��% V �/�tXii	�	�%<J$ Y1 I \(  <( < J( K�X\-J	    �uJ   �
 < K 
  w	  � J . �
tZ�2X<LHLJKWKJ[X�
6��wXh	<uX�I�vmX� JJ t A� � M
 X J
 X8 -KU8���JX<..hXl<NA�WX�1�	��*�LZ���L=IY	   f& < J J	Z-J	�	��*&qJJ*J�		f<X�
	Y=
	��t�X���	J�X�w<K
X�
t�$�X
JdX�
-K
A<9�u9I0d\~N9�u9I2�KL	�Y-(JJ/	e\�X��� <J^N\X)<f���J��<X>X	��;(JKf	����	I
��s(JK�	�����t\fyfmfv.t
.�{fu).tM. 	@wB     ��wZ
f
	Zt	[M
	Zt	[R
	Z	�V0.X�\$Xc<.����}��u� X �X7�a<t�<
JM ��L Z�L Z�L Z�L XL&�&�(�(�Jf�u� X �>Xx���t�X<
JM0�>[
	Z�>[IC�`!Xv�<{#�#t�H\�X!\#.= /ut�|�$xTu�Z,�!<Y>h. ��L<Z��Qy�uvuxt	 /�K�	 | J n	h7�	K_J.	��~t.�w%yX<wz�
	Zv	ft �	 � XHh..,�f��y
C<ht
�	�����Qy�uvuxtt	�/�K�	 | J n	h7�	K_J.	I/.J	Q�/�X �~J ?;� [�K	wuX
�X�gt��L
Mt�� J	h!t	LH�X	�z�&�w	�<�1O<	�'XJJ;J=t.��/� � < <�o=
	�.	K�.J Q S    >^ �
J	�j
X	Z<<	>J�'�tX<K3J7I	X	uJ|X<J.�J	�&9M9?�J	MJ	/J	� C � �   =  Z f*J � �3 iX7 e=�w	�J[��KM�JL
XZZW*t� jt.�Xf�X$� 	y �|�^Jz.LKCyXX�=�bLZ
X�>	tX9JX J.	T�	�'��X JB�
X�LwZ
��
<^=/J*>:%LFK5:>5:LX
J��
�
�JL
	[�J�X J.	v<�O�}���ZDJ<<3u�X z.(ttXX {xR�Z?HL8<9K<�w��tX�|� ��KzPv �: s\
	L���z�f�
�|��dֻJc�J�ZXXou	�
 � K4 x��� ���~t�X)�t[.;$kf�.nJ<tJ��-K<p<�pJZr�g<�
	��	1	�[	9"I��
�JK
	��	��"
�
t	�"	�!�	�O�;ZOs[ď���\&�&�&��
	�*	w*U	K*	�*�	K*	K*�~�.Jt\t
<	K<>'�u�~�XKFM�W!IYZ
	�ȟ�	u�V	v��t��	D �(*��?u��(?��=K��=K��.K��=K��=K��.K�NK8Lh.g.
f-t�)� ��/t�+t�J�	�z�<HvG[8�	� �'p/?FY�i�)YeK)K)		J1	� �	��7�F�$.".	Q'	LX	�#	� X	#�	it) .���|J
XK
1	�\"�Jh�|
JK
1	�"�J	jXX�� K 	M5� ���|
JK
w	�"�Jg�|
JK
w	�"�Jf	�+%X�G	K%X?L%EX	L�:9�k ty� 	J �|   5 �<
 �|J K 
  w	  � �J u �|   
 J K 
  w	  � �J q �2)�K)� �<g�J� JX	��'p/1TY�[�!rf!�K!) J t	�~t�6DJ$�v$��� >�H�$.".��}�6�+�/-c..g. �#?�-�/-j�~�[\[
�v�
.r�?�
Xf�#�
4Gw�J
�	�- ZJ V		�	�� � )  � �    �	 q �� 2�r�<
fv<>RxJJ^t�zJhK
	J�.J	RJ- `XJ  X	�	�� � )  � �    �	 q!X��Oo�Y���X��X��X�X �w�z�	�w
 suY?w
	��
pKYtYJYt\	M�}��J�����x��xJ���z�t���sJq�r���X��s�����Z�|�t��q�����q�u��X��X��X��X��Xr�Z����	�t���	�tX��wYf�|�  fX�{�T|X?
X'y
_�'�	f��f	��Xr
�'��.wK'J�~f�X
J�~<X��~�����~X��~�����~X��~�����~X���
.�}�
<
PJxXK/I=7;07I9/C<9	Je�zP�4eJJ�<�	u�tJJLHKLD	w	��	?�������}"^�tt	�X	�	=		�NVZtfX= :	 J��J�}�fw.Jf�~f+;JJ	J0 ��.�y��� X	� J���y���!K� fg��+	J0���`Y�f<<X�~J��,7|>�tJ"MJ=h�J�=!�J%K7%Y�$K.�}JmXE]�gWYZ<bK;Y�<J�t�Xw.�� =_!=X� vJ
Xf�}X<��-Xw�Kuv .� �t.�<t�<�yt��t���gw�
Jd
Zf �q<   X � = 
  7 yX A
  y. Y
  � z� Y    \
  X
 J X�K[�
X
 K �D - �+X�z�����q�f �
 v J d v�q����qJ��^�/�#91Z�~�
Z/!���hmf#�x�"K X t^wU5�h2 ktX <�"K^�v.� TsX �~..vK'J%hwJ	J%<Ys�%[q�	X�		.�tG'[JfVX �m<J[G?
T	n8�	u8)J<	v	K	LX�X4zX0K'Jf.fttt	JY
^��
^�.  .Jj X � �K w� 	� t
	��v
��O�
�/��xq?�EK3IK3M7Uw�
sY.t< �:vv��57yoKXZ�JtJ	<;JA�J;K;.;�(t��=t.�X=t.�X=t�/t�.iJ�'J��}��JZ�&X�.uySOX
�O=u=�4<�4<	#,F	gZ&<�4c	J�}&X�}<� .�X�M'Jy�	J<D�w�`K������	M��%�X,	KZ�t yJ	h�J��
	�	�,Jtt�YX�;.
Jh.ff� �������/�~��� +y�%�$f�!2<.<J jJ	h	K	[/�	�	hZ+J�!2<.<JqJ�#Q<�� JK������
Xk.%<.<Jy�%<.<J��tF��F��F��Jz^zX^X=XJ .vXZY\�HX=g -f 	p�B     �yKuf�	wO)ZY܂..P<+uXJY�
X'dJXJ..Yf<	Y&ZJ&�  .Z.. 	0�B     ��p�X�
Xv�t7x�J<sf�pXX�y�pt<��
�p<�<Z}��p<*=
]tXA
y<Y
tz<Y
X
JX�Y[�<:�h<>��LL:{0::kX�:l<������v���<��t��\� \�o��xX�����o���<J.�<
� K <5 ;�J[N<�Jg�J�
�	�	u� �  . W ��
�t�
���~�.�~t�.�~<�<�=
�.<�s���	�	b.	�,<	u �  ! e ? ��s�u�wrXJMrX<Z�<X"�X"["[Z�vX
SX
X���u�

�<u
	��	u�J� Xfu
	��ydfT��f��{�
<�JW;� Xy�YX
�[��stu�ytQ<yf_�/��Z
]w�Z=
z<KKKM
X
tti�
%���
��
f
ttft< &+)�\/9)Iu/w
tt
tj
$t
t4�vVvi�
X	�J�ft/x.|�
 
tt�rf�Jt�rX�tYsuj([�utK��Y� ���X1�	�
�t
ti
�su
k
t�u
�$2	��Je.	��JX		ts.�XX	�
�rX�<�r.
X
tt&f#�1u���
X�?
�(,<�	't�z�Z
.4�Z��q�
�	E�	v}X���
�t�
�%X

X�
�
tt&f
Jt
tf
J@X
�
�t
thNeuNsiN�uNs1N�uNs6
		��t�Zt�q{
�
J&Y*Xp�uWuv(��*	?�' zt w1 N'z�	t�<u�� 
	�. � �	tzt	u �	�	<I	�wt����xb. f( Xg���#;X	Y �	�	    �	 g  X �	�.	K�us)�"Zt ����ZY�YY�YY�YY�YY�Y��~
	�fv
]�KX<	�X	�J	�X��u
	"	��A!t	y@Ft@vXsJ	K5@r;JuJ	L5@f	�5!�w@}L0�?<y<	v?9	�F'K;.2vtF;	=;04zt0BJ1�xt	�1J	�	
<		�>O"M<�'&��{� �{Z�	�	��		<.	Pp28�T@\��f K0 ; J	6,JYJ K? ;L	>zt<P
	�,Jo	��J?�v�.�?�J> v�	 < J �	y�y�	�	"	Z �9 <��	�	�  .g/�	��rW���!���X�
�Zt
�qyt{
f�
�|�<��
	�,	J� �}�<Z:v�Y;u�Y;u�Y;u�Y;u�Y;uX	�~	�	�X�� ��!��X�~!���|��J�|�"��%IKwXJKKXf"" <Mg�|+�.K
�	�@	�XMf	+?/	\	[XhY�;Zs<
Xt	�5�A��{�"�X	"��!��X�~K�{X����{X��{J>��|$�;=$Z�>k	L+-;+u;�4<f<	t�r	
X"	\"2</+<h�\7+K	� X	��+�|J��
�	Q��	v�X	�~�	��Z�
�qy��
������vX�	X�vtZt
�	px
�v�Xy�
�t
tg�3Wu3sk?[c[
X0
J	h	�X�
vrL[qwj�J�!w�s��JM�stY�� �v	#	�t	�XX�t	j(/� X�	��
�
�	s�y���y��	f��G���	��.�
�	Z�Zr	vf
t�x�tL�Z � tJ	t�(�
J � �	�y�"�	�� t�	zX�z�t�	z	�z�t��~"&[9[&<w
Xt
tg/��/��?' �y��X<���tj��<2?�t�X�;1-�w;,X*w�8<<J%nJ$X�����
�	�X�ti	����<j��&<�0�ƞ�#>#dZ#vXttiL0vJ[9M+�w9*J%ut<<J�X	� �-u"lXX	�z	�t	�XX�t	j'��%[9[%Jw
Xt
tg.��
��
tjZ�����<2vd5X�<3&t&J<Z<\s/ <>I9J =In�X�<.XX<� �Y��XY�zt����
v
	�t� �sX�	X	ft	�XX�t	j�X���	�tttX2 < �XJI�[ 	� ��f�XX� �
X�
Xg�0��
��
X�X�<	0X�<,d<��X
��
tg�:��:�h:��
��
ti��X<	8M�w�	Mt�J�7O7LX��g)��)�h�)W��JHLHK r	��.xXXI��XX�|j�uX֞�<)XX
X�
ti�	"%.�	M%�[J	�<�.rfJ	X�	���J1	 Zf1�<.�f��<,jX<�  !   [  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/cid /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  cidload.c   cidobjs.c   cidriver.c   cidgload.c   ftcalc.h   cidparse.c   ftsystem.h   stddef.h   stdio.h   ftconfig.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   tttables.h   ftcolor.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   cidparse.h   cidload.h   cidobjs.h   fterrors.h   cidriver.h   svpostnm.h   svpsinfo.h   svcid.h   svprop.h   ftmemory.h   ftoutln.h   ftstream.h   string.h   stdlib.h   <built-in>      	p�B     �t  J#�zJP-#,�v-<+<u+v t
��}�!�� :
�gXXL�:�tq<w1q<L+y.�+"<1
L�}\��|�w Y��LO�fYt>Yt>Yf0^Y>�Y0��kKv]t9�Z
	Z	g%��ZJ=KRqu�KtZ#tO�<J�L
�3's�W�"JIK9^`t>
�	�<�
�0-tu/K��.yz�g.Jvus1�0;AzokA=
<�
	�X�
 	��~t�<(.�<J-%  <��I��YI�Z�L��<<M)'�K)'�K)'��	�	���<�5�Kt..J�~�<	�X�0��#ZX#V	�(JX	Q�9N�9dv*�<��~�	&6/I=�	YYI	=�:Xt5<�X�6Fx<6Tut
 t
Jh�D��#3Y#sK��."JIK9^>'�t�"JIK9^?=�JIK9� X��� �
t2 �
	�<W
X0�� <
�J�
(��� �
t	\	��7	� <�X?.�X.pf�Kz�fXJ�7"w�u h 4 F j � � .    $  X$ <, Q y., _ yf � 	< wJ 	< �"0"� ����{XU~KtL�,�J>���	ʀ�	�-�@#�B�
O#zfL#L
	/!�
�' .	���}J
XK
1	�N �J	h�}
XK
1	� �JjX	��	KM3	#y��Jy� 	. �}   3 �<
 �}J K 
  w	  � �J u �}   
 J K 
  w	  � �J q	_�}
JK
w	� �J	g�}
JK
w	� �Jf�)#X�GK#X
�:GL
f�~�r>"0)v"�6�	~w	Z��	�#YI�HK� #�._� XXJ `� t	�J	� JX' B��}�y�
�tJqw]	h	�JZ�K;uX�J x������X��X��X��X��X���X��X��X����X��X�XXf��y�t  �"u�<>
�Z
�	�
	�)�r	�Y�	KY�	YY�	YY�	YX	Y+J%XX+�%UJJ+<uUX-tru�
X��u�x	tJ	u��u7u�=-Xnt-zw�f..gt
�J
�M�	 & - 	 u- t	 �- 	 �- 	 �-  � wX��XX 	 �B     �'�uJZ,�!<Y>Z. 3X @<Z�Y4J3<W� �<�2Z=1N1p�xX=
	K(�XX�JbP<Y
	Y7	Jh&� t��ufvrJf�
�� J�����{X.0�X�zt�<t�~t�{�=�fY�~��z.J.0:�
[[
X�
�
y<<.�Y�����}�|�<��X�{���u�K
�~N
	/�"v�L
	�	u�L<���tJt
��
	/�
t	ZJ�2;=u p� �=KIK2rL2=f�2�=�Jv
�%9<F�0/9�$2p$@p�X�}YX7h�T�A	>%J	�c>	u�	�	Z~	Z	<X'w�	J�g�FeN%��!J
Y;g
X
�9�$��s<�2:YY2��u�
;Yu�YZXX�
J�JJ���XX�
��B
DfZ�DWM	 .X&����|� � �<oJY�w		Y�X�	y$�	JZu�GeO�$w	J	w���<
�J�zXM
<
Xt�f�&
s	[�
�X
��
�~t���~�
��=�d#�\J$<<	w�<.
	�<<C�
�JD<�
�
�Z<�<	�<��{CI�%��	�J	�0XJ	(t]Y���� ��~A;����M��|JKJ�JJ����
�~w�$M�.���\��Mt	�}	f�t� �'�f� Y�	M��X:�+J	�!�J�0Kh:L�-ttn]�&JbK�Y:�zu��eX�\�|J
���7>S�>�kw&�M<X��
t�~��	X�	=
J	P��F	=<	l��X	��&�;=<t�� Nyt"�t	�
<wq���f.�
	�
t�
L�L0.IfJW�tN�
	�'i
	�&w
t��|�'����l�fJ�X�{XX�	�
	KX J=z����{���#����zX	"��#�	� t	uX�Wt�{tX�t�/�<3� J.�<3� <?:
��|

tf+
wv�K[
X
���-�	</g
z�

<vJ
J
t	L<	?	�#�<�
��J��.�K	��{f�JvJIK9^1�=eM�	J	�t�`.f
�	�>�Z
<�<
�g6��6;j
��<�!�	b3�JXJz
t
�t/�ffX�|�KXuSuXJ�X�z<t� &���}���5���t	� <tXY�	0�X���s��t��|�
� JJ�WYWK�<	z��X����� f �0   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pfr /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  pfrcmap.c   pfrdrivr.c   pfrobjs.c   pfrload.c   pfrgload.c   ftcalc.h   pfrsbit.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   pfrtypes.h   pfrcmap.h   pfrobjs.h   fterrors.h   ftstream.h   svpfr.h   pfrdrivr.h   pfrload.h   ftoutln.h   ftmemory.h   <built-in>      	�B     >%gs=O	Z<	� f H Xq�y`��u&?@Z/I#<.u
Ji
v�#X.u
Ji
z..zX/t 	2F
4	KJ�4zJO;4	L=I'<<	uJ	f	pt'X.	gJ	fp.:X
>	ZL2=Jt=X yPKs.<=<�/=` =Htv]M>Z
	�)J	�.��y�u�K>f�?'qX� .��ff6up<J<2	�" XV<�fo;/'Jf.q.��zJ<
X �A �	�	K"TW	K'G	K	g.0J><X�JNM0.��.J2MsJZ/.>�[t<		.tY.J	2LJY�@'J�tXJ�t.<%Xt.
��T�.fJ�>=<JL>X<�
�tXX<JM-#IK-�J =  f I�~ RxJ�=���Kc? �J��vKv=v=vJ�*�. JJX  � � : @  v  � � � < @  � � � . @  �( kJ J J � : l<�>J W � =:2 � J H @  v  � � � < @  � t � < @  �( jJ J H l<�
�.JpY�.M�9M�
�O�~#�~��~�wq?<X	w����Xq����Xn.Lr�~<t�?�~&u:vX���
zzX�
?T�
<�J��JK'�9KJ= 'K)sB)z<N��Y�]�
.	�I<=>:�>	Z<<�JL:<.>X"su"="u(!Jff..zt�IY...��6t�J	f�<	h=L<.<�~��S�.�
wfX*z<B
<<X�N��X<��
P7�Y<X� � <�
t��
< W	J�<
JM�=�KX ..�`J.Kf..hJ�{tXX 	� C     A�@wY#f0Y"f0Z)J1f<)�Jc?1<�YLYL . ...n�WZ.�ZsX -<KY (JJjL(J=sJ=?
�	,J2�L=tt	�KI	Y�M=����O[*ffL
J]
JXt 	zXOt 	u<\FN
� .VwX�pJM��tXrt�����z
�zJ
4z<�
^X<� J .
 �� �0 ;NKJLt X� ��{��M���K=<IKJ��)��SJ
*./	X�<f<XD>,LkJ�>
	Z�<?
	m�JfX��~J��M�~
#�� f)���|
�
n�	<JYtt��?M\<FN0�|�LLJ�J<�<<�f<��#JJ<.�JX�
�X
���J�VLh�	��	=	@ <�	��	=	@=?
	�J�<�
	�� ��*�� JX���?q1
	hJ�1<��
	Z�1��@�j�	�}�[
�r<���	� �J��J)�
���X	�	=,	L	[	�K�I	K<	1f, �� w�{J �� � �{   0 �<
 �{J K 
  w	  �= �J � �{   
 J K 
  w	  �= �J � X Je�	��� t��|XJ�)<LJh�~�>��J<��<<�f<.���~�����~X�X	�	=0<:	LXf� XY�XN")f�XN<��X�y�Yz<l��� ���<K")f��<��	��� JM�	�� ��<efoX�(Y;Y(�Y=o.�(�Ytef� X K�}J���}���X
X�}U[0�[�K���<�t����&J&<JK����&J&<JK	���<K�	���<<	=���<<	=��}M�?[�X
t��)����Kt �  = 0 G J �J6<XXX��|� ��}��1=MU?1TJKK=!�WK>L�9�}�f��}X!�
�<X�|=�X��X�|�2�MX�W�)Z��|.�Kh �_��0Ju��w���|tG[��Z���|J�tX<�|�tJ7=
Zdh
	/�uo��K
	K�
	��"K"M��
	�!p	x � �~   5 �<
 �~J K 
  w	  � �J u �~   
 J K 
  w	  � �J	 q_�}<
<K
K<M	� �J	g�}
w	� �Jf��t�/)X/Y)W>HK)Z)H<K��� f� �su�J	2zJ	�gBWvZX.twX1X.%J?9?g=]<#t?q]J&X
X�D��}��X�}.%�<VJJ*X�}X�<%<VJ*X�}Ky.PK;K=-K=v!
�,J%��}J!H�L
	Xr<$t	<��$o<	<�9Y�@���X	+{�h=;/<>?
G	YJ�@
Z	/<f	�	�+.f�� ��X�	�|
fX�t����X��
�
Y,tsK
	u��%TN�p\t
��K;��2�}J
�L<��K=&<;KIKYt<�^�-� �t<�<K��	.;X.;XJAJ,<t�	'9h1C:U?F:3*;,O:8'F?s:A1KH?19'yJ2f1w<K
<1v<'yJ1m,KqX	�,HK,I*L,�	�*#M*q	M2	h�?��Y�=��~f$�f��|$*ug$>�>%<=%-<=�J�~J��.<�{<;nVX<	)	=	Y@cfJ.Zt<�
�
	K>
J
.<	0	=gHX	� .(�.JJ�~��K;/;<=	X��WY�=X=wX�KYX��YXY	X��I�;=�tYwX���KX�4X�J$<<�`���<.uyX�JX<X�X�<�SJXX�~JY	>x�X#X�	�<���|	�X�|@wfk=<mXy-DZ	.	/	K,dqf<L
X	KJL
	g>=
J
.<	0	/hIO�t��z<<��z.x<;
f*XR<	*�	=	Y:VfJ.Lt<L
J
[
<
.<	0	=hI	nX<j�[JJ=K=;K	jXX<f!.��~��xR{�t�ztM���<X��X��X��Xz��'�)�)�X���X����Xyt��	�	=�8^!��zJ!�<���zX�XXt	�0�.�~�JXJ�~X�t>�N3f�~3��!;j�~�,����~�
 J
�+�
�	<!�J(J9e�<9;��~�<���
��~��t
XJ
�+��X�
�J
�$�
�$��
KfX
qlX
J�%��KL����\*hv
	�Y	�g>
	�If�<�
	Z(L&J(eJ&�$:	jg#�?
	Z$>&��$/":k
J	0�}�><2�<�%f<J�	���g�
	Z� >J<�9�X�~X&�JX�x�J�}P���zJ
�f!:�z��t
z7hv�K
�J
�#��MLEv�$g$u$u$�$�$�$�$�"9ihJ�$J���h<d@*���Jm	Zt<<	hJ	��	K#�J	�I	K	��XtXL�� �t���uJ�xM�.eK.V:<�	Kt��J3 s	 <P�!�

f	gZO
iyf2
	K^&tK
�D
tS qw rL9zzJu�r2KeKu.=<:v=D<%K;D.=0<I�
�
	�&�:#rIvXo#vXvIfIsX&Xu&f&t.	�	�\
	�	^�	g	w�.�*�	J^&�	Zw��	�<	u �*  = +4 J L K2  ; K2  ; K  K 	 zJ`"�	X��J�f/�KrX��{XZX.X���+L+�>!�v�
��
t	�$�I���%��%�(8�'t\'F&sO)u>
	u>��=�>=t>J�
�X
t�
�t�DvX		<	L�J�:	@���. g<<J	�ZXW�/@zX	2�s��z�Z otX<>Z�ZX	�Vv>H'J	JX%fJ'.\<Y��MX�zXt�<�z���Xt��J	 j   G  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/type42 /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  t42drivr.c   t42objs.c   t42parse.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftdrv.h   t42drivr.h   t1tables.h   pshints.h   ftserv.h   fthash.h   ftglyph.h   ftrender.h   ftincrem.h   svpscmap.h   t1types.h   t42types.h   t42objs.h   fterrors.h   svgldict.h   svpostnm.h   svpsinfo.h   tttables.h   ftcolor.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   t42parse.h   ftmemory.h   ftcalc.h   ftsizes.h   ftstream.h   string.h   stdlib.h   ftlist.h   <built-in>      	�*C     � u�LP�k�=�?+>��,�t>=JZ�K(t?  ._�t>=JZ�K(t?  .� �tc�KxJq<J��XwXtzt.��x ��YW/LZt ��y�
XtJwtY[���X��X��X��X��X��X��X��X��X��X��X��X��X	w�	�X� ��X �� AJ�^<L/ zt^ �|.!f~	�w.&Pw� EZM
* X& �	Kk�.tI/f.;/�X�b<��J�><> �' t�g<�
JW�Xb<< <�]f%�f!�<	Z	�	��	:	>K	" >�	L��
	�
�

� Z :>	& � J� X��~��
J�J	<	=X�k�wf�b�&�Xt�&/X&�J#� JJ�<� ��/#Xt&�J#� JJ�<X61!X&xJ%RK!x<�tm1EX!X<&0,K&!<fv��XJXt��1!X&_JJ%!fK!_<!!�:t ��X/ 
'2 ! J < � p�f./5 Y= e X��?��fJ  �X- f  Jg<	��	��K	9CX9<CfI<	�<l�	X�X<	MY�	=	KXS� .�f	�XJ	=�X<X�~<����{f	.w.LwXMw<	Jh�Z�
����KY�YY�YY�Y�Y)J[Wu\&tru�XR�u�uX YXu&X �<XX 	`6C     �~J=.t.<JZ�  �  �fqKz<K><�
��
uIu
�
�7)<<).A<
J	Z(t
�"��<� t�"��<� t�"��<� t��� X/�����X
Mu
<�
�
J�\�
v=
\
J K# IYuv#�� �LVvn
�	��
��?
�Xt�
�t�
��
�t�
Mt�
Mt�
�~�$X�XK��~fu
�u>w�t	Pu	�st<	Z<K<Mu=	� X!	�J	�	K!u.X<	K?	�	�� X&J	� uG e KG � �	�vu	v>:	Z	K<	�.Z.r	>�	u	�&t �&� J&<	Z�LfJ	�.;	K!u.X<	/<J�z�ArL<=	=	�
J<��
J � �H W	�#���~��
	�utX@
�u
\bt
�	Z���Xs� X�-u�u
J �: '�:s	�<�<	 �   - = ;�v<	�f��	�<Z� u ;=M%<�J�	-�t<	�J! J JZ! �>�ufJ YK ;	L#	�~�	��X J..y�J YN ;	L#	��X J.	�~�	K�J  J..	�~fIWfr<CK
� �H>/ Xy�"��DL!;=K<��2">2�>" �L�!+�01H�k�' X�'��� �!�!���K/.�*=.t.� 8OJ�1;.�X\p@T�'fY<%&Z<&XZ<�7"]J�!_t��������y�t@1 JK1 JL'fgFF+fg+fh-fg-tv-usuwf....��y"'y<CJttYZ�� �|�w
<vt�XoJXoJXXUXvt�v���w��~�	.
�v�v�u�	=�v
�
Xt� ��ȑȑȑȓ�w��YX�X/���xGu�K�pN/�yt	<w�QL�u
��<Q��tJ�<LJKJ�T�f�}�� ����� �0
mX����
�.��Gf�~N��J.3
t	YN	wtuxX������
	�uV	����t�tq�&(tv%tu%tu%tv.tu.zz�v�/�gZg[
	�	Kr�	�	�	� K9 <	�c	�	�YH��t[YH��		Y�<��~JJ��
e���
h�����zXPf
�X
��6��!�~����/?�~��7��v�2�$�J	�	L;	�/t	�&.�	h"J'����
��JY?;	� �YtJ�f�y<�~��H��~N��YH��kX/H��f	�Y�	��t��v�Z#XJY�;e	JZ����	�=t�vL����"�	f`
.<.X)v<�[�9�Z9��~J<�X�~
���� 5�J>X� �J� <�t>Vkx"� w��v��h0��st�u��!��uB!�B�!<u/ft6��6�[w�	�Y�yJ	�.\8	N.	�.	��YJ�>[�6v�6�Y4�.X� ��
(X�� �"��"�"�" '2O27A7���
��X���X�x��tbX�uX� �   0  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/winfonts /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  winfnt.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftwinfnt.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   winfnt.h   fterrors.h   svwinfnt.h   ftmemory.h   string.h   <built-in>      	�PC     ��J=,EJ�B=2[>B19?UQK
	Z<2/kt-./�.@t�+J>�~X'y.�=%vZ'0J*u0IK!5/�'3Jvt .X�=��
vXB ���@�g)vzBB/ f J <��Xw��L&�:nx�)w
frJ=973nw<�w = K K �3L[fjF�u+�Ku
# / f fC ; �J� X����hXj/8Bl)dv�J� �mt 
�k�	�%f	? � + ; K> ;5 t	 < X)J	X��xt.1w[x�|/t��d�X���XX 	`TC     �~y<=J J %  , J L�q�
XXxX�.�o(J/�
JvX�z�x
�<<X0JX  Jt
 Q@ �O#JX|J i nh��n
�
KO
E� 
�e �YJ'X  ��.t.Xt<�tf�|t�t�|J��Mu
�|.�?�|
<X����u��t
�
MEL�
�
	gZ
	�[
't
t�%MvJ	�xX\wX	K?9L?:O9G:	L�yJ	L	M	�,
vJ:
Jv<:
Jv<	
J	�	�	�	�	�h�	�X	xP1J
JR1916H�
t�����~v����t�~��t�
�{.C�s��fM�u	6��P
&�Fvu�Xv
	�	����|
�E�W�
� ���
<�
�
J���� �K�3SAoA<
Xt
t��&�
:�KH�
f	��	�{+w-Y`3w<.	<XJ�>�	�		��Z�'<<�X	m	�o</X	Zb����X	��	�|�K�	�
N"	%�	vfX4;uX	<�Xf�t\���X�}�"KXt�.tIZ	6y	�x<�	Z		�t	�	>	�	��	�J�H�	�*=�X*u ;=<	�*=XJ	x 8=<	�	hZ�JX� v�	��HW	���	Z"�$��;X	.���DW�X��7��9[XJ�J��$<&��=J.���FW�X��7����L��1J@,&;(��?<.���HWO��XKL�OX%�>��J<hXfXJ�� �����~X"M(K�K7F�(�?(vXK�JJ��S`xRvZ��uX X 6   o  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pcf /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  pcfdrivr.c   pcfutil.c   pcfread.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   ftbdf.h   pcf.h   pcfdrivr.h   fterrors.h   svbdf.h   svprop.h   ftmemory.h   string.h   ftgzip.h   ftlzw.h   <built-in>      	�aC     � �LA��K%,;J0J6<.% K; X0 J6 fH ;NL&�)y2D/;B=/;A<H= --LVwt.�K=(1=J2X=<8<<w�	�Z'=JHL28��+=+;J=
hJ	h	K@6+96?+93>F/$;+HEL1:>L1=VM
x+>9>��t=t>�)�%���|�)�?<Z4�K5�K2Bt�t Bmz<=J J %  , J L�/q�
XXX<xJ` f;N.<Z4�K5�K2Bt�'I/  m�(J/�
JXcJX �=�V�t,�JL0TYZI[vc9pCCS:v7h�07<><�s�.4<�2H\9=wt"zD,PwJCh;>";>9>?9>Pttu>"xtK"zJK"L\tj-th:L��
�
 �2 �
��2t.[	
��|t�J�=+zJP=G>K=<u��� ..�I 7X ...A<07<><��07<><�� �� � X j��{t?&O/..6.f<//.<6<f<//.<6<>0<w�	��|t�<�=+zJP=<y�X.���PI)
P�
t  e JTXu	k�%JJ^	�X~	
�KW	=J	>Jd.Xu��XX 	�hC     �{	w	�v�X��Xq�]<tJ	�	�Z�e�/�����s�X��������Xq��XX�Y�XXP<+���xJD�
�JH
X/<.	y�<M [..;/� � @p@f<X=dXZ
	�	gJ2 	l�	 ?*	g �}���<�X XdXXX
XM3EXg3EXu3EXu3EXu3EXu qfX�tz4z<�tt�P� JX �J
�M	�d<tyX0
	J
��;�u
��=�uZrJM�Zr�M�
��**kXr�M
�Zr�� ��
�ut.�
K�u
XJJ�Qf3t�s�

t7�N�+s\Jk&-J��w
'���#tN#F<�
<� J�I��	K�u���x�uXP�
�
JX��e�XY�X
�
XJ�4<�
X<JM.��JJ�A
yX	vC�#X�\y<�<��J�K��w�Y
�K
t �JX��K
�w�.��yz uXP�
�
JX���M�	�
	���Z!
<	��	
Z�
�VJv
X
Jt�Lf
&�XXA-	M#+===Y*	Y#	K#	Y#	Z'j2JJ��L�
J�G��K��z%P��K��:Y�X@�X�%
��%J�	��f	�\
�	vJ"mJ�
=
e	1Xt�|�� XXf�
	�X<�	�%<��zHv!��A>	>*�'<<*J<'J.tJZ;<K�>dt�	M8�K;�r�
'cXXJ6�L
J$�<5;�M
J$�5e�'w	<'wJ<XJ�<gJ�	��vt�X�!
<	q�X<	yXX<X�A
e	�[
�uJ.=X���{�w��|uXP�
f��b<tyX0X�
J	�tt'��t's�� K
>*c=
0:qK
>:-<M
.��K�xb�)fU)Ng[(<E(A/<�)J$;=)e4K$;6<:="/,	WOt�#\
f >&
<�XJt[q<J1		]�4tJJ.tX	�;wX5���K��
�qM
	/��~��tX�v�zX�YXg'J<=��13>1V3>�]�Xg'JGeMY��Xg
JH;
LH;L��tg
JH;
�H;�H�^�
	ZX	Y&zXJh�
�<Z�X�
�J
J�	>	[	Z	\�<	L�@	
X<dJf
?J� 
J�g
 X	� ��w�u�L
XJ
t	�t	qft ��ti	�	g�J���		�_ ��			��J���	m	��� .^J�V�JM	�	Y�J�	
�� JvX
fK	��J			/ V= ���X�}.�Y<H�	�|X�XX<X]��
�yX�
��
�e�[�X� <�+���
`J
�X
X<��K�
��cvh?
o�<�	�	C�XJ�		XJ�M
�C
�X
<�(JL
J	�f��K
2�}�JXXH�t�y
 	�	���!�}��JJJ��xXX�(� �f	?�[X?�t�0�	u�Z JK.�w	Y	;=
X�Ȑ��֐	�t	�X��X� JKxX��$.֐� .Xth��{#XXX� �<�	�|	�X�X�#��|L,f
�v<�v
JYL�&� ��		�	�
"�u�vY
�.
� .	�uu
	"f �- s�-s�K�f K> IL�*eN< KA ; f	x�	YQ�~��~XJ�X J	d�	Y	�.X	��	�
� ��~X��HZ 	�~ &�f	Y��
 O1   V  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/bdf /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  bdflib.c   bdfdrivr.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fthash.h   bdf.h   fterrors.h   ftbdf.h   svbdf.h   bdfdrivr.h   ftmemory.h   string.h   ftstream.h   stdlib.h   <built-in>      	�C     � � = -�	=�
�X.Xv
	YJ+qMG�X�kJ.zf��q�JeJ/  � = -N	=�X.XZ
	g"+qM<9�X�kt.zf]�q�JeJ�W�j���v�=(usKM*K%���	zJK	h	p�M<<hZ
X[�>
`
/A<<hX.	j<J<	�J	gf-%	2yJK-M	h	�.�M<<hZ
X[�>
`
/A<<hXZJXr <=J�f	ZtJ<	�kJIcfv.Dx
.I�tt=t>�~�,�<wZ6�K8�K-4Jvt 0�/=�9l�!t'fJ�!J�XJJLOag<gZ�tWuuw";9M
JtJ=j":v)?j"=:K"d7�:"9K"9K"cK9"<P6>�;��� .�t_�uj�t�u�u�{� f.\G�Z4fY
X�?J��
tMJ�vXX_� =MZ�� ��
^zX
&pu
��
��Ov�LMxX ..�XX 	��C     �}

��.�
	Y+9MJq[G.�z &��.�
	g+9M+<q[9.l^ g�y<=J J %  , J Lx�t-q�
XXx �.�n(J/�
JvX��u�vfXqwZ������)�J��
J	g)q	MX��?9XXG��#r-JLX��X�m<XJ?rJLX��X�m&{y<X���t��t#�+JI��
e�
	/��w��X �oX�`xRv�t��p���X��Xs�X�������X J� �vfI�Z<u����q. � J �  > V��	AvX�	�J,.)<L
XgcJ	.0<;.pf��X<���	Y/J<N
�;tJ!�L
�
XA�L�
���!����	k�<LX��_X�J�I%<s	<�<��0IJ	JRX�	j�	��
;��MxF2Jnt_! _XY$��[�<���	w 	ftZ/#X</Ju/K/W/ �t��t-�:f�t��<Z"�XY 	`tI	g	K3 Y 	o�L		g!	=3 	e�L		g 	=3 �Y��yfytuz<�X]<
J���J�.��(t�=	�t�
�qg�tJL<=<K>:L�
�-
Qy�{
/	�.����	
t�|-X��"�
	�.���
�Kt�t<�
�	�t
��|-X��KnJN
of�K
�0
u
�<
J�%
�	�	���	K� JX ..���}
yfu�
X XJ�K
��	�� t��|t
2�	w9JK�	
\�K
<���Odq�:LXK����� X	Y�	��
p�yfi
tr.��L
XJ�Jt
���q����q��#�
X<J��j
�sJ�<K
�sJ��YK
�s�~�
���~<���JL�q�J�qX��r
s.Y�
�
�<�]:@yX�y�=u�	�	�	=
�		���YY��<��4�t�JL���
	g�	
J'g	�XX<.1<XZ 	ih!	M&Xh	M'Xh#!-K#	iJ<1<XZ!j�
t	��Jt	�
2J �r��/��	�I!�/�])MFK4��JkT=
���
��pK�����X�:<X	�:<��	wtY�<	 �
"X�^�.�Jo�pt�.X�o���J�pK
��xJ| J�u�[����p
 X	����p
 � J	�����~�u0�����nX��t�oX��t�oX��t�oXy���o��o.f�
	ZX	�&zXJf
<Z�X�
t�<	�	M	�	\�<	L�@	
fdJf
?J� 
J�: Lu:qJL
�	�#)J��	*Jt�	7�.�p�	Z�.	�p�6Jt��	��	�q�*Jt��	�tX	�q^'Jt��	�tX	�q�J	w�� <^vd�t	i�X	�q�	MX	�Z XYX	b	K.	�	�	J'�z�6 � . u J	 ��+%>#H=�#��}<KY<H<t	��=&�>r>d>Z��}HI�<
�H;���?�A�� SI I)�g	��~GI'�g�Y1>1V>�<HI�<
�H;�u<GI'�Ge�Yt��	�r�"	�r��	�r�;�����[9M�1ztz�~�)M�Tt	
�� XvX
fY�<	�!���~���J�ktJZXJ�#eX$.����p+;J?X*.�	?�B�&f n���� �X�X5 -�'�5I���J<s� t  �1 s �1s�K� KB �L.�N� KE �P%#x��%�Xf�xX
� XY� #�#�.�}J.�vJ[=.;=XZwJJ	�JIX�
J	Y�JwX�L=n .G�J[m�Z�yt���tt
pX
�pX
Jp<
�.  t��J�t
�{		��J�t
�{		��v*�JZf
�
 �"
Y	KfY�/
 t� (	oJ-	Y-W	K-	=�	2�.f	�J,	Y,W	K,	=�	>�
jf�y�X�yJ��f�	I<M��~�/t�
���~f
t-Mqg��g?Xf��
�L:>Y��/��y<M	�Y;I�J:Y;I����y�?�~�1/t���?M@=
IKJ�	H<+��	�
�JTX�lX[�~�zfX�~<���~f�x�fxJ�Yx
XX<. ��(J	�L	Q�	/���~�J�f tr
J����
J�HL#txfu	�X.	K�f)�1J	I�M�L�
 ��
���.K
�&J&J�uJ���
$HvHL
	�	��
 ��
���.K
�0J�vJ�	.�vJX��	IY�v;X�<�	Z�Y�Z;?;+[ZZ�
 ��J��.K
���
�J�Ldv
��x�wJ�J'����wJv�z��z<���z<X�>	XL�������Z�~�KJ��
 ��
���.K
�2J�uJ�
.�uJX��
IK�u-X��
IK�u-X�
�
UM
	f�Z�
  ��

�*Y*�K�JL
� K+���L
���	�$����	
"	L	��Y�Q�
��1JK
�&JJ=�=�xX��		�g��K�.�wX	L	u_	uS	u	X���y�t
�hX
�Xh<J
Nt.�w
 � � <J� ��<K
�$�z����"�tM
�	�$J	K
�
	�J	��
 ��
	�	� �f��|�L	K
��K�<��.�}�
 ��W�L��x�	�<	��<��	�|�
	KJ� �( ��
 ��
	�	�#�
� ������J
X	���~.�		�X
fJ
JJ � ��
	�	���|�Z'�(Ii<k�v �vHX���K
���
�X
�J
J�>
��}XZ��}J<K
�(J�N
�
i
J	��	J��
�-�-I<K=1�M		�0h���~�
 "�
=sK
i'�x�X�<�Y��X�� X
 ��
=s<K
i'�x�X�<�HZ
�u� �~XK(:JL<	h=-	/� � J/	}u-	/	� ,<= I<f	/XB Y
 �3 eZ3I	w�Y�*�
 ��<K
�0J�xJ��<�IY�x��<�Y�IY=X[7=2SYb\�YL/LHLYWK��KZ
	�]
J��	�~�� �
	��	
�;(��	KKI	=	��J	���J3	w� Y
0�'�<	>.�
�� X
 ��
	�0 �'X,>6V<<fLK!	{Z
fX
Ji��X�~XJt�� �	�}X�	��	�X�~XXtk"��	� X7)�4z^�	� X	�X�x���t	� t<.�	��Z�	 ��   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/sfnt /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  sfdriver.c   sfwoff.c   ttcmap.c   ttcolr.c   ttcpal.c   ttkern.c   ttsbit.c   ttload.c   ttbdf.c   ttmtx.c   sfobjs.c   ttpost.c   stdio.h   stddef.h   setjmp.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftstream.h   tttables.h   ftcolor.h   ftmm.h   tttypes.h   wofftypes.h   sfnt.h   sfdriver.h   fterrors.h   ftbdf.h   svbdf.h   ftvalid.h   svttcmap.h   ttcmap.h   svgldict.h   svpostnm.h   svsfnt.h   svmm.h   svpscmap.h   svmetric.h   ftbitmap.h   ftmemory.h   <built-in>    string.h   ftgzip.h   stdlib.h     	��C     � ��u'5p0. �h�u uw�7 �x�u#5 ��.�f-[/.'.X/<<'t!./� � <��Xgh�.( f < JZ
 f	v	i X: tY(u.<J�.� W u w� t< �Y�{�;=W
�2j�K� �3# �& J3 <K�=�0K
Jq<�<=�M�%�h��1�
)Ku
<	3.	=tp<	�.	>^�"Xt	?[.t&zJBX=3Z	wJK�?>f<.A=Jf<.
A�zJ	�	Y<	�</vt+
..<Jf.�*=KK0�
	Z@F�	K�	='JJ�qffY
<f
	�JI<�	<Z�dX� >	y�<�t�<	!f�.	A	Ya��f!XJ�<0-.=-yJ	JXJi�<	Xm�*�M�%�h� �L.����HK�rXfr<$.o<.. 
�<V�0<Y�:��:��:��
.Y	i T# @  ��u	0.�. 
 v.	 K  6 wJ	 = tY	vf0' X0 < < .	Y	�y.�<z�	<<<��.t|� <�
XM��K
EL	OZ1$f.@dJ�<qJJ�<02.=L$K6$J K5��Z,LW�=Jz�N=��<4<b�;<?JL"K"m K�1 ^J�'.
.��r.�KqfqXX�hJuf.hh�fKtsYX..X�Z�gW��KX>
	L�
�ZV�HL%_y<%QV%>V	u.�� ���0JL X	<��=�
� r� � �� .w�X� � .�	DJ	iZ$1$919J?��KJh0<K��\;��X.l�.	p���\�� .�/ f��%..#�t.�K0tiut.��J�aX	Xt	�u<ZX/&<Y�;hHK�L
zX:X�.�
	Z	=�
�	�	�K	D��~>i�
.	2���~�<-�t
X.
X	Q	�X�	?��~�.�~X�sY+tUf	+�<YKIWh:LV	K�<	NJ�K�% � �Z	z�Yy	�.�	�~�t^�"XZJ>$< \�4�Y�:L�xJ4XYL�BYJ�;h:K�;>H=�XLJh��X4��,JY�=Hh�9Kh:K�uK;Y�t		�$X<[�~��.�t=<h0X<=���X<��0L0V<> f0�;�L;VL��~X[�>�	o�J��X)X�v��H\X �0tYu=Z:v�<>��<fx�H�HZ:>,/u:=J8<C=/pJ�;>H0:=ZHLJltt��~�t� �<Xc�<X/ � �%..�~Xz<�)�XJ���XvJt�����L,K�sg[�Y'�M�%�h� �KJ<�I>1f<+1@L	.Y�@�Y-u�PX�KtQ	gJZZJJ�
J4
y�J�
<4
�t<Xm."./hf.qf</] ..�M�%�h��Kft/	�
wJZ�Y/
tJ.4x .	.&1&+1XK
/��>vn�.�&<u��gY<>
	[4&.<4<&J<	[X0�=q
	[4&.f	[M.0<[X9.,/	s�b��p.9.,/�E 9./�M�<.Z� �KoM	0XL.Y�@�K
btO.)=[>[	gJ>ZJJ�
J1
�J�
<1
[w<X.=i�.ay<
<=s Z�M�<.Z� �L>dh� �J�u.HLs(JJt&<t��=./X>N
	[&t	[1�0�=q
	[	�Zf�=q
7 u� J J+�-K�	t�	i
w.	J.v.	K	L�
.v.!LKu�	<�nd	<�	�uJZJ/"fZ�>
zX:XU+.L
	Z	=\;KKh	�flJ�
iJ	f4<<&J	J�Lq<KKKh
	��<JK-KXY!�M�<.Z� �L>dh?�J�(JHLt�7  J JZ�.0hM	v
.X XhKKLPK�
.v.!LKu�	<�nd	<�	�uJZJ/"fZ�>
zX:XZ&.L
	Z	=\;KKh	�flJ�
iJ	fZLq<KKKh
	��<�K-KXY!�M�<.Z��L=�0�K� �g�V�>�	@<foZ J=#�YKMz
Bz� J/#tYgI=
zJ<X/s.B#<	YJZ
�	@cZJ=!JY#.1
�J/!<Y#f?
E<X/r 
Ah	KJ	�JX
f	@cZ!J=%�Y��
A�!J/%fY<<?
E<X/ttJA	KJ�u-/�JJY[�>R]�. pt
 2 .I �OX|�x.2qJ<j..*�Y-/!JJYW[�>Nw	X^J tJ
 CD � 4D z. 4D z. ^ sX
 2 . �I V J��=DztuJ[4�?t< 	��C     ?t< 	��C     ��Y?�c�Yu%�J���t0<F J/hDsNY +Z	�<%XX	Z$
<%Y.,(X%X<X	(,@ %S<< -%S<,fJY
<�V *. Z���G?T	�JwZ#+f�=.�>1
JZ	g<�4"J�v6 � u W�+.K*�?U*h:<2Vf\'u's.KL�yE=J=J=J>y
X.ifX�<1uxp
 zf?�J"�Xqct,<
[J%f�axX�<DJ>w
�KLc�<
t	Y-�Jk<���L[1���M1 � J v �"�:</	� J�<� � JJ��@Z%J=%f=J0]t�%J/%<.=J0]t.<X��!)<h�J�!.a<�J��� <  ��=J�zJPK����L
J[XY� JZ
,K	=tt,�[,K	=��KEKY j� .( �@ J	J(TJ �JJ"<)<t<�g&J<JJfK<��A<� 	yJ �0  J g 	 G(�	4<KA2<AJ5...* s < JU.� .�� � X] 7�tf	1� �, * J6 K ; /6  06 : . =  K 	 )(X	RJJK7(.7J&<7J3@>+z<<	@3f	hZ6=XJ* f < J f	Q9	1�`J	]3X3<.	Z�G� X	Q<� �t�Ks<EKnXK( �@ J	J(TJ �XJ<%J+<f<�	 _&!J<qX&;J.<q;!$JX3Wx<�efK	tf/!<l.!J3.J3-23TNtJn�
	����	`�:23FJ	>@�	 �  J K I	 /  > : .	 L  t	�
<	Z�Z<uJJ/w93<</W=<>( J X JJf� .`�.Xg;3./;Y�	� � XT�KXtt=;Jl<J.X� XX 	p�C     �vv
.v<
�vX
��=�\b�
�<�r"G>J���
J�KIKI=W/L
t�Zf<"./'.]� � � & � <�?G?
��WY�L
�hw
J2
 �( I\X�!f<<
�	Y/<tZB
	�J	L!f	<Lu<�g<� ? K 	 v J.<��<".� �ggx�� J$p@tY�� �~.�� ��tJ>!�J\
	ZJX:
	Y>J<�X	t�huh.��#}k=�u�XIsXXJ;Ke�"1T=?
�t�?
^<.<twX� f�..JXJ<��
	�2	�./ YA �*[s*gWXA;�*	JOe�w.�{�� �t0:� t�XY�1W
�1��!t�w =�gI== :L/
> JJ.I�.Ix�J"&;"KxsEuEu�	�zRxJ<�BX	>vX
X�f��+zh�� �Yl�t* � X* � X, W�W�Y��Y�.	uXuX�XYJX .qJ�
	L6 tfE\  .w.�
�wfy�LurX�<f/MY;KXMt ..r urX��x.fqt#RyztutstXu;@LZ_<tB
	��	=J!�/-Y\Z��
		X<Y	�JY �  �  �X<...	o�JY	�J�	Y�I<	=J�	��tJ g*  �* W	�<YI/WJ	=J�o�	t�fJ g*  �* W�*�*Wf�JX�Ji��~�
	JwX
	 wX	QFK
<��LJL
�SJL
JM
<�v<X>X<nJ.  
t�M�
	XwX
	 wX(_FK
<(V	<L
�����>
��J��>
[
fwv<XL��nJ...
tf��g=�
J/�w<>dLtX<��M��udn�*�=IK^
dL
XMX�#��1 �	  	 /  I	 =  X tX
h�<mJ.JZ<
XXMX<Zy	�
<XM	YztJ �  � Y �hJ.u . .x���-2�JJZ�f=V0�J;
�w<	<�
=�J�� �~�~�=IK^� 
�
�t<
X�YHKz<[YKai9uW/-g/>	<X�K<J[K�<KI�/f	<X� ?  . �[���JW�=�~�� 
	K� �Jf� <��f� �J� .�	��f� �J<� ��-��� 4  .	 s � <M��W/f =  . e�y�Jv�\t
	]J	=X�!�K<<�~�
�y<�KK
JX�Xy�Q<J	<J wZtY1
 F 3 �H �	�t
�sJ�	fqX
��Jo�5Hǂ�t�<[� �KK
<XMYwtJ    �   tOhJ�u . .x��p�	.wX�LXfK+JXX�
M�;uZ:v[��eJX  .hX�
%
 �= ;�v v   � ; K   X L  X�u�l�u�	uv�		t=x.9;; �   / G< J�
" f	v&  X��K;��� X XX(K<�DL
��JMX$J=5��~.�.Kf.M�F�=�u!<(f
X
�h(K<����'X	'�G	w�<XJJ K? ���-�-K�?;�X�� \wS{t�Hh �X� � \wS{t�Hh �X��z.��yt{
�	�uX	i��	0�	v� � - s = � 	 ���	-�	��	-��<�xpKZ%tJ?	 � # s	 K X �����Z(!�JM	 u # s	 K X �������f.���	J�u[
�	Y1
�	Y[
�	ZY�	�u<�
�v��	�v�����	X���X-�ytw�yt���n�-�wY�������� v��X��X��X��X��X��X��  .	�uf
	��v��J�
���Xs�X�u� @J�v�� ��Mu X JSP<X� .��":A�X�u �c��t�v�i�X�KMXrf8����KX .R�
<oJ��
�Z
�J��K�[U�Yf0�= ;= ;X��/�Z�5J<5f<�[G==HKKv
�IJ7XJ�..s<�sX�v��KMXvf�����E�X f�~X
<sJ��
�Z
X
J<�J�Y�./�.yX,Xu.,�v\F/[U/?9.Yf0"5.i2qXJK<v�1
I�,	fL�
�	BX	�s	�XJ	�'�\8NV<:	=YJXJ�	[*�?
h�	<J	� u.;�	��	�'r\r:	=	>YJXJ	[-�?
�
Oz�K
�w
��
���X	.<	� u5;�	��	�'r\::	=	>YJXJ�	[3��ym[�|t��|tJ>X�X	�{fJ!zXJ\
X��� X <
X
t<v�>o�K
Xt:
<X 	�D     �/�w�.�J�mJJg�K<.t
>MxJJhJ�IKf<.
>	�-�~1�=J����YWYL�w<	t=
J[Ju�/.0
���f...frJX X.rtX� J	�	[L�	JZ�	M1�7�9	1	��w�s�.U<.M+.?��J<�?�* 	 J .KJ	�G	[3 � <9 f b@ 2F I	���JJ<.?}��? �* t	 J �f<	<=
J��gWY�=X>
� ��}�����}	<���~<8;y�J
J�
�>�����~��X�~J<WY#.�J	�	�v�Z<��2M12U?	�	K<�XX�X	W��	�\f
�
�fW.p�$Jvf;K3(;9=<?1<@0K<Y�e��<3>=�H=�=	 J	%<X�}X5K�XyX� t_�t	'�zlvJ
J;K.>=tvJ%�+;K+=g
JM�[��M	��{�K=gw.-;K3/3e=w.-;K3=3e=w.-;K3=3e=XX��t.0JDX��tXtK�<-t�J6f������ �ZK�z�zz�^z<=_
JJ$euKVY$K$�$�$�6&JK;K&D\��z�u<u�f��X2*gsYXeKcM�,�J\
H,L
J>:h	�+I
X+v�	=+.=�+x.	KKX�J	�Z["9(g"e,	u�(K�;=:-;	@ �1 � L � >  u ; =	 �"Qph�	g	�	�"	K#"!��KYY\	&[J	9w	+Y9J!.M!Qf	;@���<	 L   X 	< : Z z< _ L tJ K 
X I ; Z = : K = uJ	 �    	 0     t. J = s<. J K sJ. J : M G. = I	 K t. J K rJ. < K rJ �	 g t t � / .0 l J J	 /  l< -gXXtY�-f<J�/��
		� t5 � �H xf�;;	t�	�	�	���X"[?wA"7#wxJ"zyXu"u"*�"8�XK
�$� 2--tJ�XJJ�� e--��@t�K
e\D�	� �w�	-<s�	t�X< K �: ; �,� 	�~�6t�	Z,J	K,=J	L,V2>t	K2Jf		J	Z��	"��	J1"IQ_"t<6H/48p	�[�	MX	N�?�~�yf
m'<t�J�21=2I1=";K"�02�;K2V�"Ȭ	� �;	=	ZD	xJZ	�	YE	Z0�	LZtc	L+%t=.7t.��	M\�	O[�	MX	N��4"=4�"�K"��XX 	�#D     �~w.u<�uX���U�g�
���X
	����X �~��f	4��	��;	=Y;	=	Z:	>Z		�,J		t		X�Y+1J	L<	�#��	uX	� vf�~�Y
	M�	r<Y
NY
	��	Xf	�r	�.</	�C � Zw	�	
�h.�JY1+�1J	� f� f��\Wut	�W���
LY
	KY
	KZ
��	�	r��	u��X���	�b b.<b< bXtgRX �sJ
|� 
X 	�'D     �{1.O<"KvX�K� JX<J��y�
	t�>
XJ
J/(tfY�X	X(�
"
 �> ��su�	�XfJ	2X	\1*t<	�" YH ;		t	
�b�J.�<t"<Mwz<w[��<
� �7 � K7 ��
" �F �	�tw		<*#tJ	��?3,t<�+ Y$ JJ ;x!%vf	Jf�) "�! X�"X= �K �j�.��i i.<i< iXtgJX u�\J
t� 
u X 	�+D     �{]#.]X#X]X#�f/2Jt<��%t
�.M't�0'v���v0
�	J
	�%�
	�'lX'.N.
�z�a$ \.��<0Uw/
J
�M��fm�u
Mt��uusY>
^xXK � ��
#�*LJ ��� �7��J  � ��ZV'%Y�u6.v
.0 f t0 . �	�7(X	Y1(�	K(	�	X .�	Xh�YXJZ'�M Z VtvXP"t	J./t�t� XZ�X���O*�g.sfvs�;%<X�=(�E	Z<%�cX
 �<yk � t���7�m=�K�],��
��eJ@bJ=eJDxXJJi�J
	� .�
� 
	�J���
	M�tY �      tZ�eJ �          � e J          = � J          
< � t� J    .  	�. w� R   ' f�
	�<�
�
�=ytQ=
<=Y	�>
DxX�x
7 X	��
	�M
	�M
	�O
	��x���xtJ>!.J�
	���!zJ�
	�t�	u�x����
���|.��<K$J�
�tK#J#J�
	�< �x �� �zt        J > �!�J\
	�!z�JX<t!J\
	�X�	�z�!z�J�
��	�	#o�#�A �D ;�1=��	�y�!ztJ\
��� �xQ
	��	��J	�%�zflM�yX�X�y��J�0
	L.<�<�A�fJ	 tf�	 	v�u�� � � f�, �= � J5�tX5<X�<�w<*M�K<F#	X;X<wJtC8�Y+t,L;:;[,g$,XfMM �(,X(X,J� kJ� @�#v"#K"I�#��yX 
�} 
 
 
X 
X 
< 
t 
k 
X�J
	��	*+�*U�	K*	�*	�*	�	'�+ f	�-���>��>���	�7�!�-�3!-3/!��	"�"	� f5�"x�	�H#�H�#�	�X�{;  ��	��	�<Jt5X��z<Y[Z K; <�� 
	�}<�
�XgXX� -���>��>�X	�}<�<��#o�#�	� �J ��n�,�!��D!��D�	�}�<���{v
.vJ
 J� J(��
M<t
tXtwZJ�F@
1 X	K�r�.)�J�Jl�Xf�H=
<a=RyJ�x
�vX	� tt4 <  tK X�r
f	h<	Y2 t% J <u	�JJ" _ J5�fJ...m ,X=aXX��ZJ�<0,.=gX�Xy�XJX�X<!����w	.wJ	 J� \F�8@<Z
J� J?�H>f[
���J[!ZW���=!?
�K
 YC ;	��)t�=IY�JZ#	�Y�
f ��6'tY.6'�	hJ<XZ<�#	j>9<?�* u6 .* � t? ;Z�.<	 �   �X = b �	>ZYJ�YY9M+=�;�	KuW	K��f�� $�<8 X��X]��* �5 .* J t= ;�<�C�fJ���<<t =�ZJ�<0..>YxȺtWXy�J�n�� ��= T� < J	��K��H>f[
	K�atX<8��<J�QBCW!s�/�Cs	w�XX�K
��	W� J<���JJ�i hE��dL7 X S( AN<O�J	Z	KJ<�=Y�XJo�w�X<�ty5yt#'J�%-tX71)7�SK1�7t � �e,� �t	J��=	���	�J�@F2: K> �Z�XL>�n4..4<<f,XX.xJ<v+19?4X,<XKJL�	� �%BJf�� �Je�tbX'  �.�<�04..4<<f,XXKy<�X��X.����JJ�$N,�8/<>6�J6;Z�XOXJ..��J	0	KJ<�=t�kX<��z�zJ�J�$k}0,0:L6��J<6IZ ς		�XY	�JL2F2: K> eLX��	 % i M 9	h��	=	=�XXJJ�Q�X<��z�zJ�J�$k}0,0:L6��J<6IZ ς		�XY	�JLX	 j% n M 9	h��	/	/Y�X�%q�J	[q9fJ�VfX<�tz4zJ#�zJ^�$[,�cY;Y6�J�6�Z 
Ȃ	"	�	"��M	��S	!�	X	[	#u	�	��Y JJ�-5�c>?GM � �^�t+t [  J( t Jh�iJ��Y�J(t
JZtf	JX�]EYJ�1C�9�UC19MCJ � ��� ��:L uJ J7 t �* r J��׹./u�XZ��<��� �*p�JXp�X��� tgX�z�te�Xz�tR��it�t\K
W[!.J&t<=&J=&J�uX�
�
.wj
	`�q�.ef	�Y	=K<<  ��3 f .fn Rx(Y
z.	hI	=<	.�.3 f .fn Rx(Y
z.	hI	=<	.�r.$8@p$TxgRX S
XK�X �zXw.tX	�w�=JlX
�"}X>w
X<N
�c�#ww��~

v�K
XXX	X� f��
�X
X��7s�-	��I� ]�	\	Y�Ih�vJX� 
XJ
X����~J�X�~<��w+�1e�	f�JJ�<7	��X_�	cX��	�J�4C4y<[<�X��
	w�K
X��3/J,J3T�
&J
K5�
u5s	.	�1	Mt	�1X<MZ����~�����X	���t��
�X
Xjft� ����X� �wX�fXX�%J<M! N	8XXX���tl�u�<.XLv
�
��I/  ..W<
�
t	Z5t<	Mw3t.i
	��-JI/  ..nt
�
t	�XQI/  ..	\ 	��#FJ:XJ	s�	��t[t�?X�<�}�z�J
Z���t���}
M
�	H y<yX.mf>��K��g[t�X�X�g��.�df��}��[uetX.X<�}J��� ��J�}f�X�h<�K
Z�Z
��JXX
 �~t> WJX���
�v
�M
J
 �2 I	�X�/	���+ n J��;=Y;KY;=\!
JZ-<(X	�	�J V`	'+<'J<J+<���~
Xp<
Jp<L
XJ�,l�<�k.=� ��.,�<�
X�!X
J]-X�	_	
 L
	Z		���2�	�	�e��	��<	]� n��� �� ��:<>�3��J�~X/� �fK_.<! _<!tgJX vJvJ
v� 
x X 	@^D     t 	P^D     ut 	`^D     �5	�� .�X� X�X� �f//Jt<T�	v
�.M"Z"v�����v1
�M
	��	M�rJ� <r.�m.�yf'h

tttLK��wf��~JxXp�Y�?
��>
X<J���
J��}
,T�K�
��XxX�C��JC��-J�CI��?gC�!��
�JB��z<�<���Q�Nu�[���t
M
t�� �X�C�{�!�
	f8IJ����	-19O%V<0NFJ�����
	JvXK
	wXK
x<J
y<
Qx.=
��
� �<J
�3$
�3I�
��
tJi�X��tb<�XJJb��;KY;YY;YY;YXZ

J	Z��Z	������JQK
 � X�=
�u<���"0�T��&� U� �
.�#?� ���M�?U
ltt
�J��K�Mk�vM
�C J�)X
K�;X� ��
< K; ;L;;�
	�f�pNK��~�>.�d���q��<<J��|��
�J � J� 6� �@ � K@ ;��;!�	�!6X	
X6v�	
<6v.	Y	KfrJJ� �   1 I : L 	  <�3�Z3:<	Z	t	w�� 	� * wX	 J��NXJ�X��~<
��
$�
��.	�!'t!<'�%XI��J� K<�..��|.��CIYC;�C�YC;��CWuCIh�CW�C;�C�C;hCe�C-�Ce�CW��f�
7v"�J"X7�"L;7�xue,e>,;7:	z!e<!ftW�f� ���~X���~��\��U(<J(YJLG�Zhw
J�$JAW(�Ae�$JA���`*KFM0=;=<kZ?
gAI(ZAeZA�-ZAff� ������X�<X��}�Z
Y<�t�[#J>
	X<w��,.
	��f�
�
�<k�N����z<����������������
��0��X&X
�	��	[X	M	���	�	YGJ+HX�+JJ�  .Y!MH�qK�vX	I�����X�XJ�~�3E�J� hH�(f�<L	Yt�	Z	KKY�XJn��z.X<���&�~)t>���t<@��D;@
� 
��.-��;=Z:>Z�g6e�6s/6;�
��
��K-����w
X	h	�;	KYV�tY@<D��>��7�X� ���X�X	�wz�^0)q)�
@t)8
NX.MsxX_Yu�YwoZqYvVZ2,t�/�
J�	Z%J#.Y%X#.Y#J\
&�F<JH�	��8�tg�wU?[��/
	KX�t�XUXX�	w�	\T	K	Mq	K	�Y+֐�~X�x�z�o<
�pJ
XXpJP�
X
��
XJ
K0�NHLq<	�J7GMGZ
fJ�zz<�/r�KX�JJ `��
Z���z�o<�
XJpX
Jv<�
�
��
XJ
K0�N%HL%<<h
�<	zX<GMGZ
ftJ�zz<�0rK�X�JJ `��
Z���t$X`X�6 .4�
� YNJ^JY9:90�XBvr�7:70�]�n�}q�vv� fl
�2��EHvEX-K.>�
e	J	��	��J<	��f	=>V	L<�fX�.KF<	P<	L��HL
���e=	>�}."[�	�	�	=��}<���}J0K	-K?8Me�"	."J�=-=Q�.K	JJ;�\
?GMML	.Jf<>
XixX\<KJ	�X	uXfX�t	K<	KXfX�t	K<	KXfX�t	K	/Jf�<�/i%J7</JX�<<��z�CAC)OC)<> t<�W��
g
Jot=
f
=of0
p=
q<.s<9v
s<g0
st=

<�t<v
g>=
/�V.�X�.J�~�<<f	Q�</�=	JIqJ
#t�)�	Z�	�<�
X	�	>:X	ZX�{	.X	/	g	=g	@#X	[#X<	1"X<	1X	/	g	=g	@"X	["X<	1"X<	1X	/	g	=g	2"X	["X<	1"X<	1J	/	g	=g.//=>==0/=�~�.0�~�/.gg�//gic=wv��~<>0��~J=gX0��~\.��~</��~.g<J=gt>�
��{X02H0-P�
k�{JP	��{<J�JMv	L�.K;<�	XJ!�J.�z.K�		.#X<.uXu	Q#X<��	c<<<#�(	�	�E.��  \
�
X	Y9H9�r9v:�
X�4
	Ze	['u'��?X� X	�;H;�r;v:�
�	ytX�	;l
	�l
��{eeW� x�   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/autofit /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  afangles.c   afcjk.c   ftcalc.h   afhints.c   afdummy.c   afindic.c   aflatin.c   afmodule.c   afwarp.c   afglobal.c   afloader.c   afshaper.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftoutln.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   autohint.h   ftserv.h   ftincrem.h   afblue.h   aftypes.h   afhints.h   afglobal.h   afblue.c   afmodule.h   afscript.h   afstyles.h   aflatin.h   afcjk.h   fterrors.h   afwarp.h   afdummy.h   afindic.h   afloader.h   ftdriver.h   svprop.h   afranges.c   ftmemory.h   ftadvanc.h   stdlib.h   <built-in>      	@�D     �x
�x.`�&�	@	 [  ;	 �  J	 �  J J yt XHXByJ5/ � � :ZfJ
t	
X�y� 	X  =  t	 G�	�Z;gj���
	g.<<� G^u 	 `�    </ x<	 
< ��X��Y0t>Y0t=�.,0rOo0H+1LGK�w%�JJQ�wX�XQyXY�w��w<
.K
1	��J0
��h�V.��=[	�f	��.CLuI=;=;=;KI��ZJj��v
<g
w	��	J=�<J X0�
	YJ$HJ:���z�*�zJ;u
�z<K&J�ztf�K���JgAi� (JuWb<6i*gnXg<#���h	=�K
[
9< vJXJL_
Jyr Jv
J�t�*;uf�z����&�X 	P�D     �Y0t>Y0t=�.,0r�:0K2,J�=K&<���MtO�r=<E�6�J�
Xm�8  J	ZG	[)�(X<>\&N.bXi�9Y&J..�?hKM�K�
L
	Zh�J6 wJ JX...� 	wJM�qu*
�<z<K&J�qtf�K���JgAg>
XE f�@ (Jtg?g+he<g>Y	<Etv�Y	<�n��s�M�w����	�|�z �  f I[	EL;E	JK�tJ@LK�/>#-t�nftb<J<���?	!�X,`
� XK
w	�	� 	:��� J	�J,;>g,	 �,  t � I � X w X�<1 y� . J z	Z	KM\ = JH= K JsX/v t<�BHQztF�YK@oY!z<u!u!�!��
�!,X=!1�
�="
	J.9"ztB.�
XZ0u0�VKKKZ�LG��O&,J&uJ	JKvJ5M,	ttJM:,	JG,[wJ	t"x<1<	y�..	[9X�<W=���#J#KI.?�J."> �<YLKK<�9 Z@ JG J	 J�KL$=IK�z
<�JK�z
<Kw	�"�J?< <JK�z
w	�"�J?< <JL.�=IKL��X�

<�J
t�>�:<ZX
��!xXR,=!1�

<�J
t�>.�>:>X
�M	� �	K3JJI=	=X�J�~�"XJ"<<�!+W=!�Y�	X�	K3JI=	= z� . | 1 H8 J L J �( 	 XJ� X��	Z4fX=L��
uKWJ.Xv<f$
<�"<<u�
%uX%/W<.Xv<f$
<�"<<X<<?oJX
�i+��K�Z�LJf=J>:>H>$<<$<J$<"�J^&f�Kv�|f�
d�f�X�t�KJ�}<� �  K 9 G J]L(?(9<�Kv.�J �	 J� �q�-<J9 b	 J�<[�&IN&GIKIN+IK&zX? X? S& J X [  X( >],>9b<JL,<�K	at� ��i,XXJ9 W�	 J�JMN�|�
	`	=f
x�<>fX�`(9Q(yXKIKIK9(S-PWS�:2Z-,2g:-X2<.�	�.f�Kv��~<<.X	�~us	K!,X=!1	n�	�	y�us	K��.<uX��J<�5J�t�U<1�[.=!+�! i����	 � # V L	 K  � X��t�!���rX�X"��IYJ
��	S&<gX-1s�xDq�84
fq�;X��x�fpXXrX	��	
t K8 s6�	7�J�}	�v�	^	8JJ�}	KtL<NK[<>[f@hvx.Xt�A X  J�6IKB <Y6Bf <].�# gE ev L!
7xf$:Y� 7�.$;Y7Z!h� <!�<�i���q�X��
J'�2<2J<J?�	�z<KF�!JIt�L�!K�!s�;CgtX
�q�)J�
�XY
�X	��
J	��XX��M2[<GM2JJM��)�<@!sf;n<	�q�Ys	K$J2<J2J<M��~�.5 geY��'XK'Z'XX&X!�!+j;�qJsfZ ,Y!h<!fX <Y!e<lf%�Z)u<�~�X�A�XB0X%zXK�z��0t% �G e�'jC+�YC+�Y�2"TK"Y2":Z' KI ev$L;(,Y%;zX(-Y;[!��%�!zf��%�!U$%��L�'
�r�X�� 
�q�YfX-�����1+JJJ?
�Y7@<;;M�Y4?<;;J@ l J	Z	K	K	K	MJJXY4@<;;MJJY6?<;;@]JJX\�qȂXXX�	�.	%�2<GM2JJM�� �~2 X	x�K�L�XH	 � # V L	 K  ��t��7��J
<'�<�L "
 f�
��IHu�ZJ �
 f �X�=X ..." t�
T�&J�<�
�X<Y
X<�X
�		XX�ZX&.���	^us	KXwX.XXf\.X	�Xa.�	��	N*2px8\K-'J�yfY�/t�I(K�<� ��	AX	�	��IY		Y	�Y����uJ' � J �\�#Y	���v�	�v<.
<K
w	��	J<	Y	NJ7 �~ J ��fJo��JQj�IYt JQ
�;.ZJ=�YL�J=JJYLT:XZ@�YJ/�6�-��(hQ`XX�z y
�
.z.KE���tQytuvKM��, � J J��{<��|J
<K
w	���|JF�<y.
�|<J;�.
�|<�JKK�{
w	��J=<<KK�{
1�	�{��J
f	�M9J	MAX	Kf	1�{
<K
1	��J	>-mJ	K)
J)vJ<	Ld�	�{��{<
<K
<M	��J	0��# M� ȞJmX	KJ<�%)�/YI� X 	 �D     �z. 	�D     �/-=4�qA�Jz<
XvtY2�wJ<,ttw�Y=* � Q  "  < X ^X" "XD�p���X�p��p�X
�K�
�p<1	��J0�X?�� dXxJ��J3 T J�
� Y3 WZ3Wl
 u; I ] �	�<J	=	�- X � J vX�y		\	$X%X	K	KJ	=X	=�o
g
w	�J�	K	KJ3DJ�3 � � JZ
���J z	Z<X	=	�X	' J	Y 	� 3`JJ�:�#N#8JK2J	Z	K �   K  L2wXJ	�yJ-D	�rJJJ � @  ��K<�Z. J'<<=*�HL$X<=�XL�KJJ	�X�tJ<J�XvKs	5��	J tu2 �� J � .� ��~�	' J	K 	� ���1 W�J.%� �}    
J v< Q* q < X ��x�yfl<
�2KE����<�{f	L�	�$f. � < J� �L�$K$ R t . � �& - ,& > J w �w   
 < K 
  w	  � �J . K  L   xX�v��w�
tK
1	��J;
�����}t�	�w�L�wJ��
�w<K
1	.���wJ=�Js	=	K4ffZ4VE		X<	L
��5KL$K$# ���tf9 ��;h�O7O7K+x �J	��v<�	�vJ�	<
�v<K
<Kw	�
=;KM	H�	��v.=�	J
�v<�	<x<	K
�v�	JyJ	K�v	��	J?<<	K	K	��v	�	��tJ� � J	�	>t	 MZ<Z[. ��g.R��~�$d> �   J < < � G^�w��w.<��w<
<K
<M	�J���<<uv��%).�&<=.&<K.&<>YI� X 	�D     �yk
<�Jo�
	Y<X�Jr�
	Y�u�tr�
	Y��tr�
	Y��   J tY��Jq�Y���u
�}JWi#�	�XZ2"s$@�YXZ�� sJ�h ,XJXX 	��D     �p�	 
X�X+�%ft<.Z	�X?�X��*X%X<<Xr<>	kWfJJ�f=i�y
	Z.t3�J
�
h	�	g�N�J�<<	�X� X� <<� <�YJJJ�i�JJ���� �J<U�KJ� tx3SRf.�
- �	�X$JK�-<=X@/J'�/s'=;'=<=Kz<g<���h
j  <$<��;?;;=>=>�<v
t
<<
Jf�y�
�X�ZK	JX ..J	�Xtx
6	Z[*VX*f\�<O_KMX ..J�<.�x
��<J�{�&<�=	�!z<(J/JJZJ=JL
<L����2��n
 v. �=[�Y
�J	h�
	�'w'9	Z�	L		��#6EJtM��"JJ� ?[M<t��'XfZ	�W'fJJ��~l
+�
�<� �'ft<.Z	sX�JJ��J�� �i�M9Kf<L�XjJ<��?9=�y�Jp��8(�#6EJtMZ�'�X%.J<>g<U'X%.J�<�<X^� J|xX&-IKqMf�?<<X&%<L.�i�y�<y<QYNX q��LX �	f�|J��|�<��|X�u2=Y2z�,<�<hz<KK8=0	Z	K<>,	L		K	h<,	AYX3mJX��|3u��tX2uKP,ytQN,uJ[rC<�6�J�
X	�.�J�*XM<j%#vkJ<+��-YF;1YhKKM#+J�-YF;1YhKKt8[J6�J�8>�J	�	KX4fAX,X	iJ:Xt.	JZ&J�KX.fw'�J+X]'�<�;vJZMZ��	���	Ptu�2�J�.� �3�|t� �L
	ZhH�JX-JgJ6uJJX��}2�q]7Y2F<,ytFYK,J�*��yfX
<K
1�	�y��J�.
�<V�S�J<�<l�	L	i<J.	=�:	L�OZK-=
�gXJtXMZXXtJ<X1 
	�' J	K 	� J3�XJX� �#��YKA2�J	Z	KXgKL2wXJ	�	K�;�zJPXhJrfZ. J'<<=�HL�hXLZKJJ	E�[FNZJZK!�r��		L��~	�	�t#X	K	KJ	=X	=�x
g
w	�J�	K	K.�~��*4�!XX<�\J�&����t<JJ<CKK=;=>��	BuJuJ	Z	LZ�	NuJuJ!XX<J.of<<X��uX.��
	BuJJ	Z	LZY<v�u�
�u.
<K
w	��
J<<f.�IKG'L/L'HJ=K�	 � 7 H L	 K  _�=K	:�-�J� X�	 � 7 I K I[�� 	 � 7 H L	 K  X�=K		�J�	�<	[xJ	XX� 	 � 7 I K I�~<<� J Y6 I � <J	\�J�[J�	xJY
	��~'<	���~J&��-�J*�	��~���	��
	��~MJ�IK<I"[J�"IK<I�X-�J��<X� <�x<.n<�vTLX>.�=KK��|��|J�
<K
w	�J�<c�< �h-?�lT.,.<b�K==J`<N
<J
�X
�<<	�	=	�	�x.=C$=I�e=WXtP"J<�<<������	*�1c	�	[J	#x.YCx<$	<I�e=WX�^�|
<K
w	��J<<�"<�L�?<U��[
�x,Y;`x<D"�X;"=J�X
�}Xv.

 v�

JX��J JuJ.�c�.�~J(�t)=@(uqL(K(�(�(�(�(�(��~YJf��[��#fuX�J��
_
m	;\�rL/1�JKwXhKI���>JoJI	;X�	;��ZrL/1�JEwXh"tE�Z��ZV>JoJI	;�JM�� ��
"J.	gfJzf�!�J	0<�KXEX1�)"� �HY���z��&<��~�Jt=�z���|X>���}J����~�|��}rurKY<ZX>*ftLX_'�='((�5�~��tG�q��~����
� Jc�X�0�\t�UJ���	J GKL
	��	v�$JYZ�t�6XXZ^t�bJ�1M�w�
t�<�P�|��|�����Z J�
HXX�~<,;?�J��JZ�.>
�Lr�X=��(�u�� �f]�}.�J��}J.�.K�}
K
=w	��Ju�}
JK
w	��Jw
�
������KLII�I.�:H��.K."=$M.T">$MWK
O.v�K$K$O
/MI�
F��	� JY5��|J#�JM#�
�}JK#�
�}Jw�	�}�#�J2��X�
��~X�4P8s6g4g��}ttX�z�Y1&z1zXM1�Z)[&�Z�;Y^~�Z$f;;?��	�E �	�*	�%	HX8<J.K
5XK
1	�GJ�(�*Y(Vu*(;*K(��	*	%�X^	U%f	[X?
KX7.
|1	�ZJ�*,�	X*iXu,*;,g	J,k<*W�	,k<	t"W�'Y;����K�����u�u
�N� �f�|�X�=
	�"��	v�� f
	K�	t^�~J���
�~��J���~
�<
�~�M	��J3/
@}�
k 
J	Z�	y�
	��"���"�IE["xJLgP�L�KIKI��)��,��+;��u�
JK5I�	�}J�J�
�}�K
1	��J	3`fyt/JP���u;KI�)L:	�);	u)t�	��� 	�I�	�J�}GW�� S�x-RtYXiX r.XY
	L"�X	vo�X��Mv�
�.X
�f
�f
	�<
�f

�f
�f�Y0��M�Z� X��f�
	KX�� X��J08X�X3X0�nf�
	KXh�J/uuuuuuv��}t	�wX	JwX	X.�L
+J%}� J �	�? Ji"=t
	tL
J� *X�
�~�J
JtM
	�XfP J>��.�~�
W�t�/
	�$��
!t�

 KX#J	zJ	X .	K-X	#X
K
Y
�Z-[�
v�9
X
xJZ_'�-�M = K = K = K = >�
tM
	J%#X�	�t	�Z��� ����	� t	�%	�~td"�^XJKMNKYJ XKxJKKIY=?�K�I1M.>.<yJX�I<<
�K
J
Yw	�
<J
	-&J	[J�<	&J @y<=H	-$> NFK#NFGLM xz<KM#z<PLx<L=LLL�K�NKO
&
f�&
J�$(J�Yv$(J�Yt^�..�	�F@Z fu#�
	�$<O�Y9O9K�~	��~f
<g
w	�	�~�	��~<	�J>X�R.f�
�	�sJ<�<=�KM�~	�W�~X
<XK
1	
�\
F	�J��~
1	�	�J���JJ	fXJt	M	��o"KIK
>���6x<�x�XK�
t	��j"�
XLX��
'X	OHYH;	��{	�X�{�K,&<J&jX�K�	��|JKe	KX	
�t2OJ	�J	M	K	L\!XJ	_Ks	K�~��J]�%�~f��f��
	JJ)UX�
M �w�w��|X;�<�XqX�<���~��	b��}���}JH�]%J��}JL	�X0RJ�
XjK
�
Y0I.�

��
f
�
� f.XKY0�~��JY�~�<X��0�@�#�0�Z��/
J[
J	Z�|,�J,�|<�J�|J�J�|<	�J0wJX0�J�
�J	geJY	�eJ\
	Z�|,�J�	�X�	���|,JJJ�'�	��{	�X�{�K,&<J&jX�K����M
J	 �	�Jw�;KD[pJ<_;K?^J	f0�JX	��e���$J	f�Jw�;KD[JpJ<_;K�� �,�{��J�zJ%�=	��t8�X
�tJK
w	�2�JsX�<�	��~�,&<�K�<	�~t���}��
J�}XH�]%J�%�}J<L	�
�� � �	��~X�~0@�#���~X��
�	R	�twKsu�L
�_�	Q�;	u�Jt� 	��~�^%<<YJ�}<<��(;8M:0L/,.%��!�%I�!J%J	0"J/<tKI	=Y	MZXu	w	Y	x�Z�	w	Y�p X 	��D     �y��y<t�XK�
t�&�x�<�
XLl��M
XFuYFW�'	M,�{I
JzX	�<�{�&J;Y&�=&l� X���� �
X�K
	�
�
>	� X�"t� J		�	LGt�JX<.0�~J����.��	��m!2,J�=	�	K	[	K	KKIK�	xJKLX5oJX	��f���JEX�wX�X�w<Y��
V*JQ��wX���wfYL3��wX3���wtZ��
N$2J
J	��w+su%V�r�
�<�nX<��nX
.K	/��J<&r��m��VZ J	�<	Q3E	L	u��(J=�L�m
<K
<M	��J="�8<,�%i�.K�L�m
<K
<M	��J/�K&@�'�	��{t	�<�{�<,Y&XJ;Y&d<�=qAu<<��'�v$M�;�<			KX	J;K;	K@�	{t2�J	�J	MuJ	J	��	_JKI	K�X�{3��wX3�t�wJZ��
�	�| !	O*� �1:J*L<<�
Jv�L�,g,>ffL,=<fL+>:L+t!<+=;!=;u!L�	�~X	�	�	�	�	Rx�	LX�~�	Ke	K�G�\�+K>A+y<;KK<<L�g=<<L7�K��}� <#��.��V��	,�	�J�+JK�	M��|Jt�			vXG�4JX<
f	��	� �m!2,J�=�	�	K	[	K	KKIK�	xJKLX5oJ.����J<J��J�#�"'J��J			vF�!lJ�t�GZ�U�tY<;eJ\Y<<�JXJ(J7J>J%IJ��}WX/f=JL,g,>ffL,=<fLv+!�"=;K"�F���	� �m2IK,�=��
	�X	K	uwKsu�L
	�"J"J/<�	=	Kt�	M�Xu	w	KJ�
����};�<	 �J�'-(	�	�t��y
	Z	KYJ$�J�	�h,�q	�J�q�%X�=	��t8�X
�tJK
w	�2�Js�	���	w	KX��m!2,J�=X�W�k����.zz&<�I<M<J f  �   t � f�JJs<M��	wJ	� . r�  � � f  J f 
< 
f 
J 
� 
J 
t �   t J J t �  � .  < f < 
� 
� 
J 
f 
XjJ<�gF� . rJ  J �   <�{�u�.�{t.�t2�{u��X<=C�{�<X�{o	<��<	�YI		X�	�	��Z	�{X��|�
 � ��><u��v��{�������{Y
�	>c	�	Z		��I	K�	>.X	q�.<�sM X* �!�	J�:	W�:u.�	;Z�N�	 8�  * ,�*�	M.'=.s'�.r*�.i	uv*,J*�	M.'=t.g<'�.r	Y�*c��t.e#JJ.=��.&f.J8 p.�=oX<�tLzXuti�JgfJj.X<J�I<		J		���W	=	2�Z	�}	^	!	u�tn.
t-X�^A<M��<t�<' J t1 ; < J J8 o < < X�<' J t1 ; < J J8f<<9X	�.<�~X<��
>�1�~J<���~�K?� ���' J t < I
 �' J t < I ��}&xtDzf	><	[	KJy<XJ�X�J0xtDzf	><	[	KJy<XJ�X��M�	��t
�	Z�Z!<)X�)�<�w
�WB��tX
ZHv
	�'.tW	$�	f�'JKs	��X��p�2819�\Tt���tZ�
�W=
1!KZX�M
[
X	ZXk�i.9X`!*=X J.r .`!*=X ...n!xp=w!V><XQ� <.y<���{�!yo>w
!V>
<XK�� <.u��Ru�.�{t.�t2�{u��X<=C�{�<X�{n	<��<	�YI		X�	�	��Z	�{X��|�
 � ��><u��v��{�������{Y
�	>c	�	Z		��I	K�	>.X	q�.<�sM X* �!�	J�:	W�:u.�	;Z�N�	 8�  * ,�*�	M.'=.s'�.r*�.i	uv*,J*�	M.'=t.g<'�.r	Y�*c��t.e#JJ.=��.&f.J�  7t<XXV>)�,q�Y,Z<{t�<D�u7-:AJ�KI	ntZr	>	PX�~����~t�<X$ �	 J����~^!v,t�.m<8m�t-h�s B[<' O_twJJh�L �zJJXJ<J: S J < X' "�_t wJ Jh�L ȺX�� .����J$�|�JX	�|�J	���"�t�|J 
�<�<
� �1�{fX.���}��>��LJ2Z	��K� G`X�~t$�}�#<��� t
�vX
Jv<Y#Cm.<�Xi.�<�g><JJf���.X@XXJXXX�ȐXtXk<�<�g>�J><J���<J2XtZt1@X1X@J[@�<?q[J.i& Y( /& s? .B ; ��"I�z � ^ z� <�t)"tX�XX�XX.JXXXX�|!.t�}��xtDzf	><	[	KJy<XJ�XDxtDzf	><	[	KJy<XJ�X��JM+	��t
�	Z.cw[!<)X<t)J<�w+[+M9M+uvi
	K�
	K
	�DX
ZHv
	�)f�	
�)KI	u).���t�~.v�t@$<���[/~B]X'JY<'<Y�'Xd��* f�Xg��5wf/�J<M<�����2<��.=J�<�J	 
�  < ��zXJJf��z<v<8	@Z	@	[	KJ<j	�<j	L\	LXmf� X�J�X�J	RJh	NZ<J c	Z<	f<	>Jj<.tX#�~JXX��v��8@J��g.
X��@JJC.��J,XY!<SX�J��;��!v!V><XJ�JJ .s��
���s�<�Tt��vtX�h�
�W=
1�|KZX��
[
X	Ztk�i.9X�{�*s�J$�|� �>YyQX.<_Yv�  �;     �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pshinter /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype  pshalgo.c   pshglob.c   ftcalc.h   pshmod.c   pshrec.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   pshglob.h   pshrec.h   pshalgo.h   fterrors.h   ftmemory.h   string.h     	�E     � <#U.�
J
<[zJr<  EA�\�<=�C<<	� 	>�.HYH;� XKY*.tL�)p�J�<.tu}_�t
<K
w	��~J=IK�K�.	L� �~<
�<K
w	��~J	/�	L	�(rJ	KJ�qX��Y�A& ��u<,v[& ��u�vY�|t!���w�~J<
<K
w	��J�~ 
;=
;M	��J	Y<1wXz$-K�	h�}'�J
�~JK
w	��JA<	u�}
JK
w	�N�J
�~<A�J	u�}
K;KM	��}
w	��J	w�}��J@xȐ i<Z�t��}�-� .�}.�<owt	�p?u�f	�Z"<f/�}���}<
.K
w	���}<�Jy�"f/�}���}<
.K
w	��JX,w	J*yXJ�jT�.<	�	wt	=u�X&*nJJK&JK&JK&JKj�|<u�u�u���}uv�}#u#u#t��}#u#u#t�)��}uv�}#u#u#t��}#u#u#t��w�K��y�>M��YJ�z�����z��������wv��������wv�J<X�qu�X��r��X �J�=Mt!�%� t�JX�uut� ����fJX�~t�K%MqX�s�#Bw.�vf.
�^
	Z	wJh�Y $f�SJZ
	L	KXK*�AX	v	K>&.dZJMY	xXX���.e y��v֐�m<�'�X[
-�	[�	��&�JZ
<[zXP
	`t��=*<M?#X <Zg&`JJ=_�XL��=*<M?#X <�zJ	!X��L�?(fYCe[Kfe�=$*<$J:<Mi#X <�zJ	Xf���=$*<$J:<Mi#X <ZgI=�"eK=��v�eK=�u.q
Xq.
Xq<
.q<
Xq<
<qX
Jq<
J 6JX
K�6$
�6�
K6Ij&�/{&x<LrKF��	>(,0JL	=<	=<8
X�9ML�<	/�ty5y<5X
ZP
M$uJZ
	L	YWJ\
	K$wfJ		<X>uX'� J�`J
�J	� &e	KWXKX.e��9ML�.! z�/<
H>Q%fY,gu1KX J[ft]�E��q.t
J	KL�f��w
	JfX=X �}��<	A�}eL�t!J�X	�	M�}e<L�t!J�	�JX ��y�*37%7*\0*�O)K_�g<;<ft�J
J	K"<?$Jt3	J ./%. W.=
;K%.
.1  t��JY
M�JzZ:l�YxK!M?$ �, < J	L Jf�|KQ#JJ[��
M
	Y<f...Jf.	�{
HL_ A EJY	�	/	KN�|KL#��|J!Y�
�f...Kt
Wl�{�]�1=�=<W�t
J	��	�;i���	k	.kX	X��A
J'uJXX<.	yX	YX<.� <YI���}��X .%����� 	 > 	 Y   U �	 |%  t I\�}<��k<�t�{�=Z=(u(�*�*�*�*���~�fz�(�f� X&�} �X�HJ�~<�L�	��~z�K�
J�
J[	AK	zJ	XM(� f� .5 H < J X :	M�.� �tn<@�
J�\&tK=
&yXJL	C	�H	KJ<>u	FX
u�.f�
	M)�	Ix	8GX	[\	�@�Jf<t<��~��� ������}[/&< -/= ;=&J�0�J		�� .��=Jp�y�}J<�=�}�~L�tX�%J<X�
	L�}�~<L�t�%J�<  �}.��  .�x�y�/x(=�Xo�
<	�0Jj.@	>	'aJ<	0X�	J.�2;[=L
	YAJ�.� �/=  	K�>H	0vfA	mXKL	?<dXOQKz�f=>��EA�u
t�<<+wZ�K?X�X	M	=J	uJ�h<g	  	 =,  X s XJv
�gY	w,;	K,<	uJ�	 m,  ;	 K,  < s Xcf		 X   � � < a< �	h[@>���:54yJ<Cr<ZKh�N(=?(F=(Mr<X>:	L�9<�# X.��=t� f<���S�XX
<J�*xt	N*�	�s	u "  > I I = 	 _+	t1w
<X1v	�+	Ys	u 0  > I I = 	 _2F AI2F\ Ht �zJ �E$	&�~Xf.�80.�)<J	X	��~X�h80.�)<J	X	��~XXJh80.�)<J	X	��~XXJh80.�)<J	X	�J	�'#��!�!)>���!��J=X .�}�<z�.xR�}.�<t�~X
t<��~<
tK
w	��J<�J�}J
K
w	��J>
 � �& MCw�� ��MZ��}B�.fB,.fNB+�}J
<KB�<J
�}<w�	�}��J(=<<<<��<��~0�08[�L
	hX�
	�	gdy����~�X�~JKWKI2=;=?
<
<J
J<<���;K
	�I	K�J	v�K<<�JL!<KmJ <8 �~��&MCw	
�� J��� J������
��&�
<��Jg
[&
f%z�J
���JJ�Z�K;=
f[)
tȺ�J=
[)
t%z�J
[.��	�)W	K)	uXd�Mz	s<	[:	L9	K�X .	]����JJ�~�Mz+<�	e�)X	u�	K� �_-Y-Iuw�XK	ct(���K&J�	g�)��tX^f�=W��&I&gX�k�X)P)zfPz<K<K<�utXXX	�~XJJwXJ���x.�.
�x<�<%�x��<#X�x
��X�xJX>
�X
�xXX.%9X�
JJ��v������X�
�xt?�
K?��YN}�wa	"f	K<b.X	L<	=	L!JK;	=0#/#I*J��Z#JKK<E_	M	K<b.X#KA.�<	
�J<<KI<=s	g�~;=IK;=;=;=��,|�,	LJ<=I	=	>�~=;KI����,��G	M�h,t5<J	�0�0)�I=;KI	K0	KJ��~��U	M[�9W0
�~�JJ[)��U	M[
�~�JfJ�)�W��~����~�J>-z<&JLu�		KJyJX�~�� �,�XJ�
�j>�		K	[	�L:LȂtt<	K[�	L:	ZZ0t<X�	v�f	<K�JgL:hZ	0Lt<<	<.	fgX8A\J�X�"V"�H�O�"V"�H���$��qX��q��t�q��<
�qX�JY�p
1	��J=L
J	"m�<	>	��y�X
�!G�!<�!9w!<v�|��X�|��	��w���K�	
�-zP	K&yQyJZtu�
	_-uJ	K&tJtJX�X�<
8�,BJJ� X<ZtK
<�*XJX	��u�J<!%�K�W�	�
�{&
X&vXJK=4Z4VKx� \XJ��JiYX�	</pL:	�	�Z@b=,.JM�%�<�}�z�		=3J>		�K�(J	JZh	X	=r��KLSKL����!Uw
�y��)J	Jz�=��f	�t<Y(dJX	��pf �(J	Jf&`J�M
	Zt[]&<v�"���s�*-�s<
<K
<M	��J:;��<J�<	#f�|#�y�/(tJKx�
Jg4cJ^n��W�u
<<4uJZ
i<X	Z(JJ	�J	iE7J_=4pJJp>X� 	^J.X	\4t�J�
J�
<	JK.t+�	<X�!<J�f!XJ�-H.XJ�!������	��~���wJ�rJ �"zJ=JKX9/	whw/z<JX
��w<	Y� X6�JX	��w�o�XKM.	�@
	K�J*gJ<�
X	[L
	K.�	�Kl$X�	�=;=?��$�q�.�[�q(��q<
<K
w	�(�J<DLLgXv[�q
<K
w	��J<?LLX	>�sf�q
<J��
f<��	F/�rJ�
�rJK
<M	�"�J.	>�Y�r
JK
w	��J=.1r	J.��gf.<��wYLZ ��s
<K
<M	�,�J*<�� �r��r.<
<K
w	��J'-J	+J�D����{X�0�*W�	�}<`zfK�
)X	���~��.f	���.�
JJ
<�� Z�r��r<<
<K
1	��J*-J�$J���<2�{�J�
tKCsO
i	pMv	�!t?q	i��	G!J<	?	[!�Y6�%tZ LHK1sJXt=!JJZ	�qM9	?f�	�J	?	�$�Y5�%tZ LHK1sJ��|W���~Xr�U	M��~��U	M��$� KfW ,��� <<8.! t� f� 	PNE     �u��i
Jp�<`4�=;Y:4gKH4=;\�	zJ4X	JXX�~�&KI=]+�{�4X.4f+<f+<4<f4J<+�4<<4f<+t���{.M
���{�[/���{�[/��(�	X$X$�XY
O��
N_��X<X.�~�Q_Z�	���~X�
�z��XJ�|K���zJ���}�J��|���t�|<���}YJ��|����u��zX�itqJe<LJJ�!J�<X	JX<J.o�}[=�#JJ[!M6+=<S@+6;>I-=\	�	>Vf<.	y+	00K	[.0KlX<.�X ....�}t�Y��X ....��vx.nKN!
JJJ.�a�<fnXJf�
Mv
J=  ..��vx.n=N!
JXJ�a�<�n<J.<fZ
Mh
J=  .. �%   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/raster /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftraster.c   ftrend1.c   stdio.h   stddef.h   ftconfig.h   ftimage.h   ftraster.h   ftsystem.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fterrors.h   ftrend1.h   ftoutln.h   ftmemory.h   ftcalc.h     	�SE     �'�t��K��vXsJ�WgM/eX
	K<o�t/^�ux�uu 0�Jvt50oJK
	ZKkHvL�LK<XmL/xtuZ�u>KI=<M9?<".J<<" J XY-J�
kK#<<;=#+m�j.��<?< 	   q	 1   	x�	u� IK;K;==;=K:KFKHLIK;==;=K:KKN�HKJ;K:==g;K�=>9>@GIHKFLGKIK:==g;K�===9>KGKKK� v�u<.uJ	
�K	IW	JK
#<<
<.X>w�h.t<KM�X<"��f	�J	K<<J��= X_XL
L
	X0K<JLJ	>>X�i;K-KX��t=;
X=
@	�	j�<	P>H	>".$<h$:<$J"�vJ<f�KWu,X f.��KJ� ��KKKKYL<:Z<fZ Xg!tLK  .�fyo�IKruLru;u�
&	�#�@t
	_
	t Z  : h @ J K+ ��ւ	���N�K,LX<	N�Y	./f	g Z  /��IY <+�o�IKz`ruLruuuu�
�f
�
&	�4f	i �  J � � J K+ ��ւ	���NX�.
	�Y'�ZK,LX 	U��	� �  : h < ���IY  �.=�"J<=�W�E	X
L�	�	K	LXlJZ
	
�	=J	K9	L?lJXJ��v�<JJu	�
O
S�
7J=@ g( < J <: ;Z�
/> � G < ?��
	Y<<0?#X:>#/+M#X
9;K=+0
r1+-
=;
H0
<	L<	A��YJ;�	[	�<X	�_!f	�;=	=� tX> X JZ6?<U&M6�&.2��
<!S	�(���<iX<	
<.Z.&�J�	 B 	 Z   ! � J �6 @ F N J6 t <6 <> s!��<	� X!�<3 `X��!<J; 4 I�<h!<J;9f�u 	�J<<<Zt
.=
>X	m�.	>/ X fZ<$t&/$;0J$J&K+-=WK0.	 iJJi<.it i.	 ;=	=� tX>+ X fZ9!t#/!;-J!J#K(-<uv2�.
<!S	����<wX<	
<.Z.8�f�	 B 	 Z   $ �* e:�"t3F"e.J"J$KX);*@!B <	6�!�<3 `X��!<J;4 �Jh!<J;: ����f�ufJ .J>`>J'JJ< 	@dE     �fX 	PdE     �nw	.w<	.>u�t� l
�
.=;g<
<1��-=
�
	�*X�*I.��	=
..h��i
fKt�����=X
JY
	X	=W=��JL
=
<	0	=>uXYI/���
Wg
;=
?�
�	h	��\X<<f
�Y
�K=0��#]J#X  .J.hJ/
YVgX
JY
	���1�
JX�}�ZX Ztg!tL
�PK,LX .	]�$J$.X�#�EJ;X  .A<
J	�/&f$ 
f ID W Jf�
�df
J	Z$<$.��$ �	n $t;<.�t$ t ���f��@.!�wJH|�<;�JK!�w�F;���wJXv��J~LJL�wuKZ�NB\�~t<����~H��muHt><uKHKKKU===>�<<?<<t?<Y�>?�M
X	�!=.;=;KI=;	=.@KMKL��JKL<��W==�<<��p9�� fJ>��KKKG�KKG===>���Xz<<<y<<=y<<>�Xk�J��� �
�	���I�I	=	>�<<	�<�&L,:&�,X?,9�XJ	c��>K9KZtW=>t=<<��fX	�	�xt	�J=su>+	/ .	v 	(0	u%9?0:	�9	vXt4�I/��wf��W=h��	�(X�	�vtI<<ւ	� X<�� +t[M/�?
<#Xg	ht0Y2�[�
J,�	�wJ
��
t	YJf!Z�)��vYv�f�0W	.��0�	�JXd.	M+u+	�Jm4=4;/�ut	�	�t
�	#�t��|�{�u�{f���{���{�<<Y�{J��<<Z�"K	GL"..>
fh
�u�{�
�
hKE`K<�qX��q��	
�	&����}���<xZ���	G`J�.&JJ/Ih
�{t���	Zf�	�I	K0�zZZ
�
�BwJX�<��zY�
�
ZKEXK<�<���*J3J&<3J%JK$��f	NW	Y�3&�<�Jf�NKTJ�Z=LXfCMc=U/W<=;@���=8M sJuKT	2�	�fv		Y�	�W	K/�zZZ
�BwJZ
^	F	=<�`	Y�	�W	K/�zZZ
�BwJZ
^	F	=���zY�
 
�KE`K���Y�u�/YZ�
	v	x�KpJ�X�z�	F	=�ZX���fu�y.XKs�XK�X�X�X�X�~X����zJ^ <..t�<�wXw<:?:<�.<�f�<�X��V��l���K��J+ �! J�J ��ew<7
X;�Wb�!<�< ���S-t/;K��$����~-�l.�u
�KKJ���<2/ytz�<�u�y��8�yt�$Yy���ZK4<J�����1w��;�z���;8��;�X�t_J!.[f��!.t�~t��lt;u�J�uX
�JL=N4?f  �g���et<X 	PzE     
Lr�Ru<���3�
� �t�[K�t.DJU_��
�L�)�[�
&�	&w�L";gJ";XuZKW<YX�I8t\D�8X�<M�i�s�T��Xs����4zf2Yt<Zt<Y�t[ �   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/smooth /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftgrays.c   ftsmooth.c   ftimage.h   stddef.h   stdio.h   ftgrays.h   setjmp.h   ftconfig.h   ftsystem.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   fterrors.h   ftsmooth.h   ftoutln.h   ftmemory.h   <built-in>    ftdebug.h   string.h     	�|E     ���q�#NNx<sf������J .J>�>J'JJ< 	�}E     �fX 	�}E     �zw�?UZ���1J"t1JtM
>p=Y
.<b<	!<t<X.g*� B�� <�@Dt@<D<<��	�.	M<	M<	M<	M<	M<	Mct<X<	"XfX 	�~E     �z < J9? .K<Z
[
1xJJZ
	Jtj,J,Jt�/<=>H>>	oJ<=ptn.� 	�E     �X
�XmXL
	�Y
KI/
M
JtJ	l�Z
	��J<�;K&9L&<=i�J<uW=.j%�8�Jh�FL�4�	ֺ/�|J
�t/�}<�<�NW��v��	�.	l;	KUL<�h��r	b	gZMa	�	�	L	YL�|J"$<$JXKX*		�%f	=f.	�"uJu<	Z.XK.�
	YL
t	M=�,cJt.��K P��	�X��=Wt�J�J+ �! J�J ��ew<7
XIf�td<<8�
J[�K�E�LHg�/"�# JG�=.C�=.�f �
\
<- J .M
J[
<	M$*JJ>&|x������K@�� �����v�t� tw:�;�=9& � X > X9 � � > X �w�X��zBuy<_I@	+IKX �5 s��W{zf;B	9:IK	7Z	L

���*<<(JJ= f = � <. J pJ � T. <fX	�����[2FGvVK.&.>V/-K	�t.<�u	[F=	L9	KW=� 	YL<K( .<MYsu���
��	 �    ? K T < K & 9, < . K   V	 ? �? t[^zJKWKM&,;g/WK�? �[ZjF?)�@8HK.&.J/-K? ��.ZiJ7�i&,Iu/-K��Y<;�JXY�	 �    K  ? K& + M, c < K   V	 i��J=t<j�y=L9�L)<<)JJZ�,�  .���uX
�JL=?f  �r���et<X 	�E     Lr��G�<��u.;
�<P[K�.��~<Z�n.;
�<L�XtW�M���~<
��
����].;�<
�~�$
X
��M�rLYW;A8;O9r=/,@Z=N�C>tBX>X� �
� �-��<���~<<X��t..�� tjBr�K	fw�KnxfL[
��K
z.
�v�	Jw�	J�Y[�
��Ku
iK��.�1�
�,K
(%yX	<u��q�9g��
��K
�su�Y[�
��K
=-u
iY��1�
��K
i�uvu�Yeg��z�uyX
��
<�J..�gf�Ȃ�	�	� �!  J /!  X J Y!  X � J	 T^!w�		JXwXX��XX� ��� 	��E     � 	��E     � 	��E     �
.KuJ.KsJ6x��uzt�KW$	�y<_w<YzJYYY[Y,s$�.eZ,sZ,sZ,s�
"�M��M%�M%��
�� 	y�=K
Jz<=8=>;<q<?L=AzJGzJK� �JOLz<Q?8t<K9@9;MqJKtJ>KKKKKJ:_�,s�,s�uu.�K;=�J<<Y�~�
.I�u� o< oJy$x9qYKYYY[Y,sL,s$�.;Z,IL,s�
<	J
wf=I
�t�hK9f^<+�f=<�	;�=QwJKzJ===<ME=IK>z<K;>;IK8I<:JEJK	:4�Jg�..ptYJ]�uu"t� �J=�f<Y�w.4zf2Yt<Zt<Y�t[ `(     �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/gzip /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  inftrees.c   infblock.c   infcodes.c   inflate.c   adler32.c   ftgzip.c   infutil.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   fterrors.h   ftzconf.h   unistd.h   zlib.h   errno.h   zutil.h   inftrees.h   infblock.h   infutil.h   infcodes.h   inffixed.h   ftmemory.h   ftstream.h   <built-in>      	�E     � e .`<�a�G`�� !� 	  J �YX	�.K�f� Iw0
Xgt I <1y.j<�Np	<:�n��qKfI?j�.J#.J" � .[.f�N	:�	<�=JJ	IX�<K
J<JJKY_=�y<x��7<
��� �� tmfDJ<.J�3�� J���#J =X8Y=;=I==I:>YNJ\�	�<
z.	K..e�i	`JJ	��IJ	�
�Xf�<Z � .<� J<.L@*X
X	cJA � XZ.h
WW=
�f	�
.J=s</�	 �
 ! ;
 / J �NJ	 � ' - .L	1g;J=.�	�=
:	=J.8.��XB�Xu-g	� �X�	��CXXJf� �)��X
.f�N�	<���YJ=.<YJJYY�2��~GguJKH�Y�J0KX c  X JW.Or.�,�.
-�.I</'u
/yX_� X J- X) JW[MJY��Y��0���}g%�
I/ yX_J</KH0:hY��	uX�-	=	g�tg�I���<��<ft�< �ffffff��	t	��W�	�s&�YIKI=s�X � 3   J J = 	 = ��n X���uKM[�~M[���~f����uv�u��X"�v..��� .�|�X 	@�E     kX 	P�E     q%.-KOXY�c%..hJOXY4�
%)
�XJ� JX
 A<$ WP' �uu|XJ�	�J	M�!	�J	��[�.
J � �% I  #��~tzCMFK( X K2 ; = Y   J <[/s=JYJX.JM�;Y?fK8MX J.Pt�
IK<\=Y�"J�=
GM���JM�;Yn�Mw<	<Xu��s 
s����WJ���|<�%btJ[%b��[�%f�GJ��J�=MTK:4uY	+_�
/ g�/u�$��vg��i���z��g�*X` .t � J �- �) <�#� f#�XL#:Y fX'X � )  u2 e � A � *  u3 e  J K A J *  u3 e  J K A J *   t �  K  W g� X�<� f � *   t �
 	�	g	�	u�� yJ_�� � $ " t
 <	�	g	�	uw.;X �  " g ;" � ;- g( X - =-  .
 <	�	g	�	udX<�gV�u=X�<� X � *  u3 e  J K A � *  u3 e  J K ��<�=��� X � )  u2 e � 3��4��
J	h	g^<,<�JJ�J����<� <X��<XX
� ��2�� �JXX�6M
	�	��~	��~<���JJ��,#MJ:g<=q2ff�J�f<�f#J
<�JYI&	�vuBX<�JJ��<JJ�~
�
��$X,Y:.@<,<@<4.s	�	YXX�J�f<�(X�	K;	Y�0XI<0=W<4�;XX;�%<<	����J�<5<"X	u5;DX	=DI	g;X;X%<<�	><�5<5X"X:tsX[2�X>XA.�2�X2X�<�X���0h����/�

X8��<� JJ��<JXX�~��JR.�R<.<JfY<�X�/	�6
	�}X���}��X�}<��}X;"UK�J�}X�J��}XgK3	�Z=#�~�X�~<�XXXtJ<Y�}� ?�t,� �JKX'*<f�J�f<�>:Z:Z
"�(<<	�)u�)
<�
XkJJ):��X��B	;<A
�X�X�X�J��	Yu=	JYV=	<=	<=
Xy��f�JJ�
��~�='	���<Y
	�@�@[	_� J�Jt�f<���;=.�gY�YY�֐J�Jf�/XX��J�Jf�'	���;<
	�<	Y=�	Y�� 	YX�J�Jf�1/Z#�#;.�L.[	=	I=Y	�;Z�	��Jt�f<��t=	I.	�	bd	h�X�<<X��<XXX�r<
	i	K
	K
L.XX
���
	�<	Y=�	YX;	YX �J�Jf�'/YdwZV?V;Y@�X��
3�Je1JJY
J	v	g�	� �
J	g	u��!'<
<	Z	g	�	up� �	yf 4�.	�J��<J�gqf0�JX<��J�<JXX�~� X�~ ��	�~��<�<f�� �eXXeJX\�	�	�	�
iJ�<�Xj��Y&�	Z��=�	Y��u<	$J��<J�<�~<<X�<XXXY	3�J�� ��K����J�f<�hX:<�&<tj<<�	�3.t3J<.�!%JKK�	(<f	�~��J��<X"��sJ<JXXZ.�J���B	;� ����~X,� .�4�}�Y;1� XJK�<gWL�3�!� Y�^X*<JNp9u�NNJJ<Xqf�X�&<�� X��/��	�u	M��X��<XXX�+�
	�vX!<	��X�	��<�� �zֺJ=�	S�<<�<J<XAX
	L	Y!<	���<	��X��~<
=�		gL� XX�� <3�}��JJ�<�~J�Xt	9	u	�X� XJJJ=[�u�JJJJ<X����fXJ�	ft	u	�X�t�zY
��t
Z`�	JtQ�/ p�	
q�tt���~g�9XXtf<�<JXXN<<3�J� !8�JJJJ�	� tX<�<<g��.3pKs.t�uKvVt�
�.LK>	�
�Jk<�
	vF=�Xu
�
zJ��	-	�XX<.L�t1	&J	u�zJ4 <.
C�YXX0XMXf� �y'ytC��k��+&t�
	Y:�us<v
 <Jo<g=:Yu8:vY
P < .JUt�~t���3< f.]�>M<Y+t&tg
	Y=;uv�;uv
<i�
�<�MZsuK!�tuu)u��� JX 	��E     z �n<JPXK�?�=L�J<��}Ku<=N�LtuuY
�l�
JyX~xI�Ls�L
X6����"J�sK�	J:!MfM�u��X<�Y�<
�Mb=
M[:
J	�.J	J��}��K	�S�[:!c./X��	��}t��".�}M[���}f����������X(���=��X	
J�f�!tytXtJ;_VZv<KZL��YM�/Z�

J[[�G?  V�*XXfzJ^  qXZ:>tcf*Xw� 0   [  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/lzw /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftlzw.c   ftzopen.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   fterrors.h   ftzopen.h   ftstream.h   ftmemory.h   string.h   <built-in>      	��E     � 
%)
yXJX
 v�$ OzF\  � � XY��zJ=f }. A�
	h<	=	�/ � �dA
�C�%�I\;Ks�=u���,>XH=/>NZJJ/s0:/KtJ/JJ1XVt
	�	u%Y	u.n�X  ^�<,�#t<c.Z((x<((<Zvt
JyJu
`
<	��XA�X
J�v/�	m��	�zJ.
�5X�K�uuuzs=J#uL�vrvK�c�K�uut� tz �	k<J	JXKM?�=L
�JJ��u��X .�Yn<�}H	Js<KKLtuu�YQ	�cK	X�~��[�"�~�&zt�\JJwY��uut Y<X����f� �KKUP�~<JZ���~<u��~<��X"����-�:KK?[.f�X:KK>J<  J.	�t  ��u;9M	k	�J� gUthY*�LJy�<	J<Z(J�*,JY*,JL	M	g	M�~��X �D �	�&u�=;	=.f	�	[=,	u=y<A=�;	>�	@	Y	wY	>	�n��� _ �.  g��	.�	< . s	 = h i�l<��  �  J zJ�� � � ��~u�f
�
�
JJ�/L/VLrL\�X�f�<i � �  �	 � � � ��~Y�� r� tUpf�5t�gM�t�1t:<t:<<
<	Z=s	�bf�<t� &=
X	�=;Yuv2�X	�t���(!W�+tK��u�Q�uu	� ��� �5�0t=� t�<0?w=;uv<	��
��nth
[�
X+�=@7Yv�y<Ov�tJv/u -�   A  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/psaux /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  afmparse.c   psconv.c   psobjs.c   t1cmap.c   t1decode.c   pshints.c   ftcalc.h   psarrst.c   pserror.c   psft.c   cffdecode.c   psintrp.c   psblues.c   psread.c   psstack.c   psfont.c   stddef.h   stdio.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   t1tables.h   pshints.h   fthash.h   svpscmap.h   t1types.h   tttables.h   ftcolor.h   ftmm.h   tttypes.h   cfftypes.h   cffotypes.h   psaux.h   afmparse.h   fterrors.h   psauxmod.h   psobjs.h   t1decode.h   t1cmap.h   pstypes.h   psfixed.h   psarrst.h   psread.h   psglue.h   psfont.h   psblues.h   psft.h   psauxmod.c   svcfftl.h   pshints.h   svmm.h   psstack.h   <built-in>    ftmemory.h   string.h   stdlib.h     	��E     �Y-J=t?>�@�{�>;E<[tll
fJ<LK
\X
<wJ<sX<.=�>Xp�~>K�Z�Ybf..=
���	�frJZJ< ��	v
 � J�
 X	iJ<ut�>J�  6xX�CyXYZX[XLX< r<ZMZZ
X_pJ. <�  ?Z �n
vJZ<	ZjX�
<XZ
FX
vJX=�=�2���QX<>
L
		J	\	J�K`�>X>g�Z<V A/  A E�<J	DJ	�JhJL8� �K=�J�<�
X[
�J
< N  U^
lJ.= x�<Xz��	�	�> m� � XL	QJ	�>z�� X�>X	p<	��~.�
<JL
F�	��J_Kl.>XU 8��IAX7YYT2�
<<������ 1%
y�� �A�� .D�
�; `�[I=X JV=KfUf
�
 ���PX�
J Xf
�	p���
�Wf�3�.<X��;t �
�z�uu�iJX=IY[<�K:�=Y
;=
	��^=X .��u�L
X	
J3�Z�F.u�L
XJ	<JHJ6<u=B8HXX=<ZXx<n�	
X	=���	� <lX X	x<YJMJ0JK (��iXZ tX .JbJWKK"JN%�WK%JZ		��	�Jt	���<�	>IKZJ.....l ���y��� 	 �E     �y��y�J��y<X�>J�Z
�
M�x��yJ@U +.k��x\<x��.�x�<ffZ�i
[!	<u
[</
	ZJ	Km<Xm<<<�<Y<��A>�
  ��d X�x�	X<x��y>�x.�y>�  uKK=Kn�� �MY:� �K[�$ f, J$ J X @1  J��]�2`v6$I-J=;KI=Y
�\'t
<	P4J q� J	gJ� 		=I	=efg�.MY:�M�-oJ<qJ-IJK	,Lc	=t�� �K[�$ f, J$ J X @1  J��]�2`v6$I-J=;KI=Y
�\'t
<	P4J q� J	gJ� 		=I	=efg�.MY:���p��pJ[.wsX<<>"=;="J?.g<y&zX=yX�%X/X/Z1�l�u����  �=wgs=K���  �=wgs=K���   =2gg2s-=Py.=����91& K8 ;LfMl0H<'yJZJ.K
t�K
JA._1/vXD/y.,�#�KB=DztuJ[4�?t< 	��E     ?t< 	��E     �
,y.uw,�y<uuuuw� ��f<J�� <	<� �X<	� �%�K�K��&�	���J� <��f� <<X	��J	_\	f�0	?%X	*<f	
�J	gt�~�	/�	�� �	<� �X<� f�JJ�JK%-f<J�%-f5<<t�	5  �%�%����s�J ��?J* /. f7 Ih,]2Jֺ�t2 J J	�-M0X:vJJ	.�~��~J
XK
w	��J4Wt�~J
<K
w	�J�	.�~J�.�><<�JY�|��l
X�|���7" . t�&?J
J.&J
<6�<+X
�}J��|f9�2�C
���<
�	�mK
����h9X��
�~�N
N
J J]�| �.J
J�
�}J� �|f 9 ��
	�r	��|��|<�J�|.
<K
w	��|�#��|.#�J-.	K#f�C�K4<J < L 
 ΐ./	��6N"+!�
	�('u(I	''
J	O�tJ�	[J" Xj�
�}J��|f9�X���y<";K3y_���tv�1�t<<��tJ1<;=9;�.NL
	�J�.t	��u
u
1	�J�
<�t
tu
1	�J<���;.� �
.	\ J�.t	X�t
u
1	�J�<�t
tu
1	�J�<��u� t	j. <JP%.t[Yf<	��<JP%.t	X�t
��u�+<yf�t
� �� �OfXu�����X���}f�J?�}Y:�t�t/��f�t� @tX� �~t":A�X�u ��.i@zX	J
�X
J<	J�yX��~(KH>H=�
<	Y#cJX�KeKXX�
�S
O7
OXX<JM#J=Mv=K��X ..�|�
37
]S
O7�K
.<�
JJJ��X .
 oJ1 ��WKKuu��(�X ��&
v�&
.v.Y/QG�&
<	Y	�J� 	�.Xgf� Xa�	JwtC
XJ
J	L	K
vX	Li	�JXgf� KtJ. <� ��Jf2K8KMYXX n�J
���M
�u.�w<-=-�JKY;��;Kfhu  ..�t��<Y
�tf<�j<��WZV>
�
g
e� XY�e� .J' X f��� X>����
О	V	�t<�qJh
��
	�X<���
\J
<��
.�~Xf�\�70e	$�4`<$<' 9Z
X�
<�>;�vX��X\�7+.�	�J�P&e?�Jm�	�< �	+	�	�"XL�J<X80�	�J@
<iuJ0�
	�ftXJW	�<�����<X��~<X,XP<e� .�t��.�;Z:�Y��
�W�
�u��
�
�"�	Y�-UM
	��
X]J_�Y
X� �N�
+�<XR	�	K�f.c���y�J�y<J��yfX��HX 	0�E     �|ufXuX�Yt�
[:�Y
M
�d����2$�\X2#X�.�~:X-XA:S<K�f�Y���^z<Pz<YX<Jfk0-v  k� fJ#� >  U M  X =.  X � K.  t � K.  J � L   vX�	�t���=�K�K�L	.�~$JJ	t	�� 	]f�YJX
	�JtY
� �XY	� �=	n�	��0[�	Xwt0KfD��KsY<ZȻ.J��	J	>��	��/�/�J
�
�Y8�  I=�~���J<3$]KLx�=N$=$:LY
=Lj�
�	h	
�
go�	��X��}���J��y�M�<$XXX<ZJ�'<�E=N4 ., < R X�"X4sJ+J�L?�=�]
P=N�.fSJ.�A	Km���P0X� <�y��z.�< �yJJX��z�<�zJY�=
��[
��u<�
�
�X"�7Y"I	u>
X	^L
t]JZ�
XX =��J�zf
+�<XR	�	K�f�c���y�J�y<JX�uIX 	p F     �s=J%�g����LHLL K LnJLY�� �K�f ��� 
�t�v
��)Jt
t�NK�KKLX k��}t���LXL�
h�
J(d<J
�	�~�
�
J�{��  �<O�� i	�~J�	�~.X��,XL��>
�
�$�
	�m6C�iKHJ<KZ,!U� <�f� A? .A�X
	y�� �J� f6MKKM
l<<
K
<M	�J=� 
	L� f6�� X=IKMZ,!W<	�~��	� f6��	T.7f6�XX
	Lf6�X	�f6�X��]J�]�g1*$Ju �  � IM*K$-u �  � IM+K%-u �   � IM1K+-u �&  � IM�����*u$-u �   IM+u%-u u    IMySg��vrv�<\g
	 �  &   X /  X /  Z 	 V��6�wX-.=$�h�~�!- =J)�f\"� ���������!�!�� f�X\0#tu%�#� � � � � � �#�!��'�'� �y�!K^�J
J	Y&4I&K4;�� q<K.  u� � 
J ltX �.%pK4J
J	Y&4I&K4;��  u� � L
Jy�K. �|��xo�KK>Z�?IKK�Z.J=�u
	Y/t�������XX� /W�wrKK>Z�f?IKK�Z��
	�	�Z"<u8"t�������XX�r�xy�/.u<
tv/JIJ<?f-LȂ H X>[
/ X�/�	LF2 X�oJXfo X��/-gJ;J�Xy���X
�wlKvqgN�gZ�v,ZX ...XkJX  ...�t�%4V*%�� : < X�
f��X$E	.Z �Y	ft.�|�
�
�wst�
��
�Y
�\�_�w@J	L	X	u i< �
 ��]�Xk	�	u$	u��
� <�<�� -[A	E�	
X	u uJ �
 ��	u�	u��	�w.�K
=
;	�X\
[vHL	X. �	 0 R<J:X�...	m��	0 W < JZ
=
;	�X	(J��	pf�	>uX�X�<��	� f � �	 0���[�$f,J$JX@1J��]�2`v6$I-J=;KI=Y
�\'t
<	P4qJ	gJ� 		=I	=efg
�n.u MJYK ��v�y�#tu2rg�pt-�tg�p
0W
� �j�vrvU/.  "Y��3.t@?
U�!>��!	�<\ <X�v.w�x<��x <��x<�t�x<�<�x �t<
�x<K
K�l	
�M	:���0V>:0�x
�K
K<Ml
	=��
�xtM�J	�x.��
FJ�
�x.�Jy�x
wl
	=��
�xtM��x �J	�x.��Jy�}���9�Y X �{J ���z�J�8�D�z��z��  	�qX	�X�Cy<
<	i	K2 Xf J�
	[J�"�zX�J g3 I / �zJ 3 ��".�y	�<X.Kf��z
�	�Xig�Jt ���!ffr�,�t	Cy<<iK4 cf J	�ZJ�"<�<O
: J-v:s>��z��z�~��t	��z�	?��z<� �zJ	�	��z$	�-��z��z�~��� �X��{�N��~J��L�~
�	�%D�uf�s	K%_y�	M%	�	v"Xf<.	1"�="�5I�$YKf$;K9:�<�~J:��	<"$<"<$J	L�$�
	�:<J>JJ><<><XK,�&�X�~����J�|�6�}� �6J ��}J<[	�~J�����	?sK IK ;=
�	k"	M�}�h(IJXi<X��z��M�xX��
X	L>JJ><J><JK,t&�Q
�J<$YK$e=$;K9:	3t"$<"<$J	Z�$�EtX�5
��otw)�]X�~X<yX_���}Xf��~X�0�	Mf[B�%z<J�
$f�}'�	Z�[Br^ Jg.�K�}
�		�	K�}��f��z��zt��0LcK6LVL9X�u<I]o.2X-<t��z��X�<�z��z�~�����N< p t	��yf�j�yJi	�~J�	�~.X���,XL��y�����~�z��X�z<$�\rXI�z<�f�z�v���z<$�X9�}�<�~.:��%0�Z%LXf��|. J/.�
5KX�~.!�JPJ/(�}	��}�X�}
��<��f��.J�X.J��.J�X	X�}!�J	L�}X��}�~�	J<Xgf3�	�JXgf� v�-&<J&JJ^/IuK��-&<J&JJ^/IuK��Jl��0�[�	�Jtg�t�J#� �P. J���s�	�~Jtg�t�~J#��O.Ju~	�~JXg
<�T^zP?tX���X �=� � U�J(<tJJ�
fg	 u�o�X
P�� ��
z<Y
X
�����XY\(KHOUME=Z
<	Y#cJXX<�X�� ��L?KJ)J>)dKKIKZK.f.
��<X� t�ZJ&X��K� X .f:f�~�#�~�J��	J�~<<�?����1v<C-M_~Z�-NXoX�Kf....%`<g�
�<�{��s.pt�qt�|p.�t<JJJ! X\�~"KYYU/==9=;>KH=KG/===�w
K
K<wl
M	��.f� <'.v�<� �	
T	��
�	j"=	s�
	$�	�G	[9	[hx�X ..�f(��9�]##J���+��XX�~��w�/	Cx<=;=;=
�w<K
J�l
M	���	.�<�wJ.�V�wX
<K
w	���wJJ�,L:>�w
<K
<M	�J�J<
YH��
YH��J
uH��J
uH��
&s
�L�� 	xv��Jf� �	
UF�	�
U	f|
�	��	2$
3  "��	s.
) �dX�Xf
�{Xv#
��YJ<<
.�ZuIL$t1Xm..:u.s.KM�	�	w uf 	<v�
� -u v v 	t<%�	I�~���~���~t�<.�~1=AG1q�u1tv�u�
 �s.6 � �0Jt�! < X�~��E���v�		.�I�J����X .pJ��
�s�.t�<t �� f�	�KIgh-;-3q:=>9YYt��u���`uu�. �t <& �8<tJn%#Is�Z u v+�zBz.Pz<�ff�_	��r.=;<�<�rJ�1�rX=;=�<>�r<<�>1�r<<�<9�rf�.a@IK0?zJ0H=>?0vxt:Y>y.Y���u
or��u���q���uuXt�Y�Z[ ztu vwk#=Iq%�J��s�y
fU=0vtQYM:-K. J XX>
WY
	/<J��`��%9�[	KI	K  J � X � �   � �  �  K X   .W�[	I<	K�

	x
LVL
	2J_X	��
�SA
O	/��	&J�t 	@1F      � ��\J!�NX .� XLX .+��oX
��Y
J  .	F�  *X 	2F     �=�t 	@2F     8	EM�-cJ<cJ-IJK		=Ltt(X
v_�+JKR��4JJ�
X	Y&4I&K4;�t	���� XJ=X<.[�Yd�.�< VJX).
�oXYuXLj�t<`
�o
	���
�p��M$�t
�p�$<X
�p�$X
�p..w��J-cJuIK	KI	=LtJX
�p�6�
�pX�J-cJ<cJ-IJcJK		=L<JJX
�p�6�
�pX�J-cJ<cJ-IJcJK		=L<�
�p
X	�...� �} J�t 	�4F      �.�NX/� �KQ�[X0J-pJ<-oJJK	<	=LttJ$�	�rX�uY
J  .	p�  *X 	�5F     �p� �<� X� t#�g�f�t=<<�<� .T<`</K
� TJf<K-
w	�Q1XJO=-w<
?	�Bz.B
<Y�I?H*JW<M&<ZJ&J�f�?��[Xw-y;R(�<;(=<:�X�3<	�J^<
".K\
#<<M	�JZ
	�$J<�#�fN?cK[�x-KCxf(	<I�e=:WX�	$J$<<�L�11<	�	�	[	$x+=Cx<Rx<D&�J;&=J8�X��r%..s%fsJ<K?<!L�JHX>	fX�2�J
cJ. �bJ��v[Bz<�S�
RK  .o.1K <��K	s<u<	Z	�	�(Yt]�-?�Y#�?��.�K�u�<cY �
 � �9 Wv�f�Z�	�X�~
rJ��Yb
X��f	���rvX�vL�o�	b��	�X	[	�s��	�X	�	���~����J��}
��
X�Z��
��
JU	��
 �X� �	Q�	�X	�	�[�	�	�	�	�X	�	�	�	�	�a��}
��
X�	��f	���
�J�� �Y�~
X�L� ��,4f�X�i�f����}�L��f��~f���	")�	K�f�<�	�}
V	L	�Cy�JL�QU~	Z	�	�X	�	�	�	�	�	�X[�
��� �
��z��Bz���Z���Y��V/uJm=,�	@JX�	Y�	K�$,PX.y.u��]1xJ!xJAJ�<˯4seu�pt-�tg�p
0W
� �j"Vv"u"�  .�n�Zm0LUK6LHL`�CJ�<?Y,Jh�J�� Y,JfIX	�<X.Kf
� �u�Lj�t<`
�o
	J����X� M
�o
X	g1X<J� ..X 	@BF     LJkh	�Jtg�� L:LtX	�Jtg���Jy<yv>v<4X��
�~���|4XcXs�
�J�}tL��X�{�_Y
��}�|��g$�|������z���.�x���|���������|���������|<��Z�yXF�#o����y�tiJ��w��&�tTu�yJ�t&w�y<&�t�yJ�~t������yu���yu���yu��v&�{�t��&u���%vyt�%�y.�%�z<�%u%ud%vC%y�)�%�
�}.%�X
�}X#��%�{.#�Xy�{
��}t�
��~�
�~�,�X � �{   � �   X t <M=XN
�
tJ�K� J��K�
�|m���|�
J
���~.�
���}<
���~Jz<^<�J� ���� X��W� �K�	�{�	��
	Z u+ WN);	 ) �+ :	
." t/ f f .
t
�
Xl	�.<���jJ�	�{�	��{�<	� � 	�t�	�x�J��q�w����X���h���X���h���X���h���X���hZ?������lf7 ��}���f�j���<��i��<�#A7.AX	�~�%�kJ#��.=0�� �k	�J��<><<A�;=Y;KYCx<=[�KZ��h�5�yJX��B%�kJ#��.=0�.f'X>;=Y;=ZBx<KZ�LL��h���><<�A�k#�<���lzJZHL[Gw.wYJx<X��;uY;�Y;KY;KYBy<KZ�L>�upJ	V	�k#��- X	�V	��	Z.	�l#��	�V	�	�	��df	L��	���lJ#�� �lX0 �		�5	M���mU�?��l���v�~����m<u�~J��u������lV�����l�\XJ"�q��3J.tfO&�t@� ��X!�
f�	�hJ	�	�X����	 �   >v�n��X�mJ� ����m���m0���6�nJ �y�����n<[	�~����J�<
�'�f�'X�L�s��yJ#���y<.�AJtJ 2  �* t J < X t��Mtf�Y�zJ#�.�J >  � : L+  @ [ G w  . w yX J �(�{X	�J��	�z#��- X	�V	�	��d�	v��	O���z�		� . X �* `  ;	�|��z�		� . X�2%�jJ#�� C y<Q=;KQfq<Z,K�=XK;KY-K	XwJLy.�XZu<uP�t�eYrfY-�XK;KY-K	�w<>����q	��yJ�	�~��	�~.X���,���y<�Z�Z% � �Z.X@UY�
�~<X�%
�~��!tfL�
t	�4<<�	�����x�Nt�y#���y�<�0fY;uY;�Y;KY;KY;KZ�L><�up.����m	���s(�x���X���k	�J�j �
XX��<���g=�i.�O��	�qu�y.�	�~��	�~.XgX.�,���	�- ����l"��.��iJ��	 �@ 	 � at@ 	 ���
�|��"t'/";JIL"JL�	VX	��
�!�!X.!J=�Z&�E�iX�Jf��k �0X�~��kg<��{fX����g=�i�XJJ<�/]73�
�o&!<J��X���t�h���X�w���[��XTX� ���i��<��iXJJ��<��i��J��i��<�&=<.lX&0.I=.�l]7X��}.X�rt�!��6 � J����m�X�s.�:L[Gw.w[�{X�X���}#�}X�J#�}f�J#�}t�JM�}�=L>LwcM[?.f	u<JJ�~XJ.�
�~<K
1	�J�;�B�~�J#� �^t=t�J�ft�	��<t�
5>�+Y>;<	u&J�������n#���� -M <.0<X.��#�i	��m�.<[	��	�	��{�	� �m� # + ���Zdl�X0XuZ�LX=��
�q���`
�q8Z�8>���!-=�'
�q8Z�8>������1v�x�ւXX��
�u���W=YW=\T>�xX�J#� ���<�x<�t�xf �  � �xX   �J #  � ����x<�t�xt � � f � ' ����uXL) �v< � X X X X����XY�{���X<�sJ�����*X;th�X/D�|�<X/ZO�|.�<f�|�0�|X4���VX�!X=!X=!X/!Zf..NfiZE ��@ts�\�X>E ��1WY1-uJ0�}X���XX�$X=$Z�.<Wt_�#X=#Z�r
.K
1	����&X/&Z...X`�$X/$Z..X\#[#Gw�Z2 �+ <B ;�$7X.$��X�X#�	�2$�Z>f#�r�$���< K @,f$�,b@ /#  � J �rX    . <D �
 �sJ K 
  1	  � J! � < I _ �s   �J #  � ��t=tJ �.�<<�0�~X4��Y���tJX�
�� &8f<g&<���X�|�> � L* / <* K/ ; = - u/  � ��0�P�-�����X�|�2�<XJi��s��� X���s���r<0*�X�r����X�. t X=��tY�0WX2(��X�&7�h�X/@�}�<X/ZK�}.�<f�}X_�X=X/Zf.Xe��.�h�Z�$��z�+)�+X).+JK+)X+JZuZ�>���X�K��~	�&]v�L&�&X0#XK#X=#]#SMmX��9�?-t��'K 'S�= �Y �=l�tX� X[#/-	#w<h-#y<�#K#�-%X�X-� X%J�-,\%T-X,M%U?,I�,u,�5�X�"!��� J �  <3 W5 ; < . < ��z%�Zd0%X<. eXF s�9�?� X�����&X
'�z���
�zJ�'>rv<JY8J<�J�5	X5w<K"I�JY"<6Lu"`"x�ZX?�X$`
'�zX��J
�z��'>rv Jg8J<��&4X[&94J�&4JX0�X����Z�o
.K
1	����Zf��X�� X�m.�7<= �7 . < .=-D�"X=\.X�z�w.tK"�"Z*..X     0 % : X	t"Y;="[*fWtL � Z*.X:�e0�0Z!tD�w<���uX�X>Y<X�w��hX�Z.�fX�Z16X.J��X <X�X0�o�X�~JJ#J��	�;[>��M<4�:	X2)n<)JJ<KulfZ
	Z	K:>J<M/
L	K..N.<.x.	�~JXYfXX�X
���U� X�
t?�)yJuypvY#�l<�X� Jm�Z#��%r� t��
f��� 
�Lu
 J7 X	wL<utg�����=@agj�~� 
	L�}J(�X��)<�"tJ�4�~�zt�<��~t���}xt��x
��~�uii
��~
v-�
���~Z=j
@Ffx
��!
�!w��!y�K!z�P�L
L	-xw
$
��~t�
� ��h
�
t	�#	}�}f:��.�
� �t
� J��
'J<	���!�|�::�<j��tJ
u
WX�}����}e.t
�J�|X��w�|
��
�1qi���|
��|
4�t��|
�4��|
�4��|
�4��|
��|1f	<5.f5rt0/e	�		$.ej'R�J�	irv9.<	�
C	y<g+i
<4|
�	$.c	v.�
7Ct�KCt<�J� 
�L	�~X���	g-.<	K.;	M:g	+;i
.4,
<�"h,9ifaJ(X�<J�
G1
	.flxfhlG�)?>��'/,qt	JX%IJJ� ft'�t���t	$�~%�+JM�Z
�	m�~%�wtJ	JwfX� �wt�
�t#���}t	�
�
\
�
�t��}�<M	�{�
�
��}tgft���~f	ZXi�:>��'/1t�	JX���LX�'%U.JJX�7�t
PD(�XX<
�X>
V�vH>>
	Y9t��3� �Ju� �t��.
�<�f�	�� <	n�}	���}f:�tt
��
	� vL�	�vJ<��v�~<
�%�t� z.���
� t	�~J
��~X	x
�XX<�~	?	�+t.��b�	Ow	M	�	�J
�~��	��}fV��.	D�}:�	��.
TA�~�?Y�=��=��=��=��(&s�&^
"�&]f
#f#iJ
fn<#p
�u
w	�(TJ=��'Bet#b<h
K
1	�%`J:����	�{�
�g�	.X	,t�X
�}
 �
   #  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/psnames /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal/services  psmodule.c   pstables.h   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   svpscmap.h   psmodule.h   fterrors.h   string.h   stdlib.h   ftmemory.h     	p�F     �/-/-g\Jx
`03p�
0.t��	K>!:�<0#JL
.#qJ�
[
	KJjZ<#<JL
.PZ
M
	�JhX+\�L�'72%�/	�%	/.	L<t�.	�/o<	Z<%..=I	=<	^	hY<	LpX
N
>	L	Ky ;	=t=f<`XK=Y..XX��$g3�2.$��11�XX 	P�F     �u K	WA)J/+6\�	�v
g
]
s�)J/+6\�	�v
g
]
s..� X/�.J
`	�=
�	L
W9tJ
	Z)W. Xv(XX (t
HX	/Jp� �g�JvL	�<�	v�t	9<��	vf�%JX�t�_�< � J �V�	 ,  �HJ
J	�XX��`X[ �f I6XMF7<W	4J	KZ K[	M	 [  <- m J J . m <	.	Z���`. e
��	fMF	4J	KZ K�	P	 �  <- j J . jX	J	L�..u<�u.�u�uXXuXXu<Xu<[-�
tJ
��	�	�X���
�Hf� �	�XY�% k < X��	J]hH=u wJf<L
	
�!<.	
�\��	�~���g� �<J� Z��Mt
JHf9=I=	J�4>IK<	�2Xo	,�!�� �   �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftsystem.c   stdio.h   stddef.h   ftsystem.h   ftimage.h   fttypes.h   ftobjs.h   stdlib.h   fterrors.h     	��F     � =JZ � � u "� Xbmy
QLi�Y -�.<Xi�~�<X 	`�F     ;<X 	p�F     c<<X 	��F     � ��y RP yX� u � � �X=S`�#�K_� Ky.��X p �sJX  ZX&X<N�Zu����X  x   I  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype  ftdebug.c   stdio.h   stddef.h   fttypes.h     	��F     ���    �  �      /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base /home/computerfido/.local/share/lemon/sysroot/usr/include /home/computerfido/.local/share/lemon/lib/gcc/x86_64-lemon/8.2.0/include /home/computerfido/Desktop/LemonTest/build-freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype /home/computerfido/Desktop/LemonTest/lemon-freetype/include/freetype/internal  ftbitmap.c   stdio.h   stddef.h   ftconfig.h   ftsystem.h   ftimage.h   fttypes.h   freetype.h   ftobjs.h   ftgloadr.h   ftcolor.h   ftmodapi.h   ftglyph.h   ftrender.h   ftdrv.h   ftserv.h   ftincrem.h   ftmemory.h   <built-in>    fterrors.h     	��F     ,Y'<���#�=0;=;KIK0L�$.a>yJ=.
XL�t4.<XL
���IK
	�(b	Y/<fJ	>� > � : X >  	 7 J
J�J.B�&
	YZ:.	[X�XJ
J ��J� X�.� X^��X	��(���OJ:�</��8KK3X	f=Y3f	t>#WXlf	<#H$?#+.$2!8M=A!wJ	>:LJ/	�.X�	�; � L	��,	�Z<Jf. >  w/  = ; K  Z   wJ ��K1f 0  J =  J <	 h < f;KX �~�J<	�:	��<��>�}lz.=X.Ygf2oKKHuu<r=<>q.J<..�LE�<=J<	pJ��:	��<Xf� �  	< I/ E + 1/  ? 9 K/  / ; = = : = ; K     u�<fJ=J<	[J�h:T	K	L � � >  J =  J	 7 J �A:	��<Xf �  < I/ wJ + 1/  C y< K/  ^ z< u/  X u/  X u/  X u/  / - = ; = ; K     q �J<.J=J<	VJ�; f �8<M �  0 I - g   �� <M Z  0 I ; u   �� �}J�X�}.�X�~�<�� �2<��p. X� pX; se.	 �x�wJ��w<���wX$�Y
M<tNX6[yX
J<JXv,� xJ`u<�y�� ��H(ZJ �( J> I�n<.?j.
.m<
f[k.J
+K
L
h�t<� .Ztu% d J J �0XJ.	�	� u  f	 I �  z < 
X	 % �< J% . <� �uh/	���}�X�}X-	�	Y	M�1�~J:�J�~J�.�~J�<�~X;/;=>.�ci�~�%I%gX=��$I$�JM
	�7*===7cKZ9	=��*.8<	<<hvKLY�.S%I%gXKX�J�~X��J�~�/;=�%I%gXKX���~J:�J�~J�.�~J�<�~X;/;=>IgKX��2y�~'�
<�J�f�+
V�<t	,���	YYyX
f��9M�J� 2�"	�D�� t+rt	�\	F��<,<Xf,<<<�</$J0<<" e�	 <�htMY X�tJJX\	�=<+<	J<�X<.J� �Xw�Y��>X	"��	YYwX�
m<���* J%X:�	w.�=-& �
 <�0QzJ7Py�=7<<�81�:8>:>�J! � <j�1JJg�J
`�`< <2>^t J
<^�k<<t<�
 Dt~�X8�}�x	w. k3 ;8�;C-=IK-X��J� J! � <LY\
�, J�&�Vv��<Lt&<
<	�pX�pJJ�X
J�
X�
J	rJI$Jft$�-<	~-M99H	\;	@�<XX<��:X>7��	XX�
L�K>
	KJ�~JX�J��~J�X1;�xX3�
YeK
jW�J��~<$�Xr.�J�X=E$N?G5<-<FL=:�;��wzXjp��;�V8P:�	t-X-J?	?K	X zJ@[K!v�JuX�0 t,<Ks<,JKsJ,J:MG,=IK!t,<!sJ,JIsJ,JrJJutfs.�g<l	XJK;	KXa�#�2#t� �u"u"�OJ�}t� ��T-M?�Z .7]z�=YKZ*
<�<
�#������}X
     fdim _ZSt4fmodee _ZSt3absd _ZSt3abse _ZSt3absf _ZSt3absg _ZSt3absl _ZSt6scalbnfi _ZSt3absn _ZSt7signbitd size_t _ZSt7signbitf _ZSt3absx _ZSt4fminff _ZSt5log10e _ZSt5log10f FT_ENCODING_APPLE_ROMAN _ZSt4fmodff __mlibc_file_base sqrt lldiv _ZSt9nextafteree fmin _ZSt6lgammae _ZSt6lgammaf strtold _ZSt5atan2ff _Z13PointInWindowP8Window_s8Vector2i strtoll closeButtonBuffer _ZSt10nexttowardfe closeMsg _ZN8ListNodeIP8Window_sEC4Ev at_quick_exit _ZSt3fmaeee _ZSt9nextafterff _ZSt6scalbnei fbInfo _ZSt4tanhe _ZSt4tanhf _ZN4ListIP8Window_sE10get_lengthEv _ZSt5lrinte _ZSt5lrintf windows __mlibc_uintptr ilogb FT_ENCODING_NONE atoll __buffer_size _ZSt11isunordereddd lastKey 10win_info_t _ZSt5log1pe _ZSt5log1pf FT_ENCODING_UNICODE nexttoward atof atoi RemoveDestroyedWindows recieverPID _ZSt11isunorderedee wctomb _ZSt9nearbyinte _ZSt9nearbyintf main fb_info_t signbit _ZSt4fdimee _ZSt11isunorderedff replace_at mouseDown remove_at _ZN4ListIP8Window_sEC4Ev _ZSt4fabse _ZSt4fabsf uint8_t nearbyint operator+ _ZSt4atane _ZSt4atanf _ZSt10fpclassifyd _ZSt10fpclassifye _ZSt10fpclassifyf windowHeight isinf _ZSt4log2e _ZSt4log2f compression mouseX mouseY fpclassify _ZSt4erfce _ZSt4erfcf environ unsigned char __int128 unsigned _ZSt4modfePe ownerPID _ZSt3tane _ZSt3tanf islessequal _ZSt8isnormald _ZSt8isnormale _ZSt8isnormalf fmod linePadding 7lldiv_t add_front renderPos _ZN4ListIP8Window_sE10replace_atEjS1_ closeButtonSurface mouseData windowYOffset _ZN9__gnu_cxx3divExx __dirty_begin __offset _ZSt4sinhe _ZSt4sinhf _ZN4ListIP8Window_sE6get_atEj isgreater windowInfo _ZSt6lrounde _ZSt6lroundf log10 hdrSize 5div_t _ZN4ListIP8Window_sED2Ev vector2i_t decltype(nullptr) _ZSt8copysignee _ZSt5isinfd _ZSt5isinfe _ZSt5isinff islessgreater FT_ENCODING_ADOBE_STANDARD _ZSt4asine _ZSt4asinf _ZSt3fmafff __mlibc_uint16 mblen atan2 FT_ENCODING_PRC stdin log1p windowFound vres _ZSt13islessgreaterdd __io_offset _ZSt8copysignff _ZSt5expm1e _ZSt5expm1f _ZSt3sine _ZSt3sinf atanh FT_ENCODING_MS_SYMBOL _ZSt7scalblnel exp2 strtoul FT_ENCODING_ADOBE_CUSTOM _Z13AddNewWindowsv _ZSt3expe _ZSt3expf keyMsg _ZSt5hypotee _ZSt13islessgreateree ListNode<Window_s*> __mlibc_int8 _ZSt7llrounde _ZSt7llroundf FT_ENCODING_JOHAB AddNewWindows __mlibc_uint32 _ZSt10nexttowardee _ZSt7scalblnfl _ZSt9isgreaterdd floor log2 __dirty_end RGBAColour double_t _ZN10win_info_tC2Ev _ZSt4logbf _ZSt13islessgreaterff _ZSt5frexpePi PointInWindow closeButtonLength fabs _ZplRK8Vector2iS1_ getenv __priority optind _ZSt9isgreateree mouseDevice add_back _ZSt4cbrte _ZSt4cbrtf 6ldiv_t _ZSt5hypotff operator[] _ZSt4modffPf _ZSt5rounde _ZSt5roundf this active char32_t erfc uintptr_t _ZSt9isgreaterff asinh _ZSt6tgammae _ZSt6tgammaf __float128 FT_ENCODING_MS_WANSUNG FT_ENCODING_SJIS colourNum List<Window_s*> _ZSt5isnand _ZSt5isnane _ZSt5isnanf __mlibc_uint64 __initialize_p keymap_us _ZSt5trunce _ZSt5truncf long long int _ZN4ListIP8Window_sEixEj __mlibc_uint8 mbtowc _ZSt4sqrte _ZSt4sqrtf mouseEventMessage senderPID rgba_colour_t renderBuffer FT_ENCODING_MS_BIG5 llround GNU C++14 8.2.0 -mtune=generic -march=x86-64 -g -fno-exceptions isunordered _ZSt14isgreaterequaldd __io_mode importantColours wcstombs ../Init/main.cpp remquo FT_ENCODING_MS_JOHAB _ZSt5atan2ee FT_UInt32 _ZSt6remquoeePi FT_ENCODING_BIG5 __buffer_ptr current _ZSt5frexpfPi redrawWindowDecorations _ZSt5atanhe _ZSt5atanhf _ZSt4acose _ZSt4acosf char16_t _ZN4ListIP8Window_sE9add_frontES1_ fbSurface cbrt _ZSt7signbite __gnu_cxx FT_ENCODING_ADOBE_EXPERT isgreaterequal scalbln __valid_limit _ZSt3cose _ZSt3cosf strtoull qsort long double float_t _ZSt11islessequaldd FILE data2 _ZSt4exp2e _ZSt4exp2f get_front _Z10DrawWindowP8Window_s atan _ZSt4fdimff bsearch optopt _Z22RemoveDestroyedWindowsv _ZSt11islessequalee long long unsigned int surface_t PointInWindowProper _ZSt8isfinited _ZSt8isfinitee _ZSt8isfinitef ldexp uint16_t frexp 20bitmap_info_header_t _ZN4ListIP8Window_sED4Ev DrawWindow acos expm1 nextafter _ZN4ListIP8Window_sE9remove_atEj _ZSt11islessequalff copysign opterr mousePos asin FT_ENCODING_GB2312 __cxx11 _ZSt3divll _Z19PointInWindowProperP8Window_s8Vector2i trunc quot acosh FT_ENCODING_ADOBE_LATIN_1 ~List tgamma __int128 get_back FT_ENCODING_WANSUNG get_at drag _ZSt3loge _ZSt3logf _ZN4ListIP8Window_sE5clearEv _ZSt4logbe fmax _ZN4ListIP8Window_sEC2Ev isnan _ZSt6islessdd _ZN10win_info_tC4Ev _ZSt5asinhe _ZSt5asinhf _ZSt4coshe _ZSt4coshf strtod strtof strtol stderr handle_t short int scalbn uint64_t _ZSt3erfe modf isfinite atexit _ZSt6islessee _ZSt4rinte _ZSt4rintf colourPlanes llrint _ZSt14isgreaterequalee _ZSt5floore _ZSt5floorf backgroundColor get_length _ZN8ListNodeIP8Window_sEC2Ev srand _ZSt6islessff _ZSt4ceile _ZSt4ceilf FT_ENCODING_MS_GB2312 FT_Encoding_ windowHandle _ZSt5ilogbf _ZSt3powee _ZSt5ilogbe _ZSt14isgreaterequalff mbstowcs _ZSt9remainderee /mnt/e/OneDrive/Lemon/Applications/build __dso_handle uint32_t _GLOBAL__sub_I_mouse dragOffset _ZSt3powff lgamma isless optarg _ZSt5ldexpei ceil _ZN4ListIP8Window_sE8get_backEv _windowCount title _ZSt9remainderff short unsigned int stdout closeInfoHeader hres FT_ENCODING_OLD_LATIN_2 _ZSt6llrinte _ZSt6llrintf __static_initialization_and_destruction_0 _ZSt5ldexpfi __in_chrg _ZSt3erff _ZN4ListIP8Window_sE9get_frontEv _ZSt4fmaxee _ZN4ListIP8Window_sE8add_backES1_ __mlibc_int32 FT_ENCODING_MS_SJIS closeButtonFile _ZSt6remquoffPi __status_bits remainder _ZSt4fminee wchar_t mouseSurface _ZSt4fmaxff isnormal _ZSt5acoshe _ZSt5acoshf GNU C++14 8.2.0 -m64 -mtune=generic -march=x86-64 -g -O0 -std=c++14 -fno-exceptions -fPIC /mnt/e/OneDrive/Lemon/LibLemon/build ../src/fb.cpp _Z12lemon_map_fbP6FBInfo lemon_map_fb ../src/filesystem.cpp lemon_readdir _Z10lemon_openPKci _Z13lemon_readdirimP12lemon_dirent filename lemon_close _Z10lemon_readiPvm off_t _Z11lemon_writeiPKvm inode _Z11lemon_closei lemon_open whence _Z10lemon_seekili lemon_dirent_t lemon_write lemon_read lemon_seek _Z11SendMessagem13ipc_message_t ReceiveMessage SendMessage queue_size ../src/ipc.cpp _Z14ReceiveMessageP13ipc_message_t _Znwm operator delete [] _Znam operator delete _ZdlPv _ZdaPv _ZdaPvm _ZdlPvm operator new operator new [] ../src/runtime.cpp surface DrawBitmapImage _Z10surfacecpyP7SurfaceS0_8Vector2i _Z8DrawRectiiii10RGBAColourP7Surface _Z15DrawBitmapImageiiiiPhP7Surface bmp_buffer_offset size_aligned PointInRect rect_t bmpHeader rect _Z10surfacecpyP7SurfaceS0_8Vector2i4Rect colour_i memset64_optimized _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface memset32_optimized _Z11PointInRect4Rect8Vector2i reserved srcBuffer DrawRect 20bitmap_file_header_t surfacecpyTransparent srcRegion _Z12DrawGradientiiii10RGBAColourS_P7Surface _Z18memset32_optimizedPvjm _Z16memcpy_optimizedPvS_m _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i srcHeight dest DrawGradient bmpBpp rowSize _Z8DrawRect4Rect10RGBAColourP7Surface pixelSize magic CreateFramebufferSurface memcpy_optimized surfacecpy _Z24CreateFramebufferSurface6FBInfoPv bmp_offset _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface _Z18memset64_optimizedPvmm _Z5floord _Z8DrawRectiiiihhhP7Surface destBuffer ../src/gfx/graphics.cpp srcWidth colour DrawGradientVertical yOffset available_sizes finalizer FT_Vector vertAdvance FT_GLYPH_FORMAT_PLOTTER oldB FT_Slot_Internal oldG RefreshFonts FT_Glyph_Format FT_Library FT_Driver FT_FaceRec_ extensions FT_Bitmap_Size FT_Bitmap_ underline_thickness style_name face_flags FT_DriverRec_ fontSize FT_Size_Metrics FT_Encoding FT_Outline FT_Glyph_Metrics_ xMin FT_String style_flags FT_ListRec_ FT_SizeRec_ DrawString yMax _Z15InitializeFontsv FT_Size_Metrics_ FT_Generic FT_BBox_ user FT_StreamDesc_ num_glyphs InitializeFonts character FT_Glyph_Format_ FT_Outline_ fontState oldR max_advance_height face_index descender descriptor FT_GlyphSlotRec_ FT_Face_Internal DrawChar bitmap_top sizes_list num_charmaps y_ppem autohint FT_Long FT_Generic_ num_subglyphs ascender FT_StreamDesc FT_StreamRec_ fontBuffer FT_GLYPH_FORMAT_BITMAP underline_position _Z10DrawStringPcjjhhhP7Surface FT_Glyph_Metrics FT_Memory font_default FT_GlyphSlot control_data control_len FT_Realloc_Func FT_Pos FT_ListRec mainFont bitmap_left FT_Vector_ FT_UInt FT_Alloc_Func LoadFont font_old FT_Size_Internal FT_MemoryRec_ max_advance FT_Bitmap newColour _Z8LoadFontPc n_contours rsb_delta palette_mode pixel_mode FT_Stream FT_Face FT_Int FT_Generic_Finalizer FT_SubGlyph FT_Stream_CloseFunc xMax FT_Free_Func FT_ListNodeRec_ tags _Z8DrawCharciihhhP7Surface FT_Fixed units_per_EM FT_GLYPH_FORMAT_COMPOSITE num_grays x_ppem FT_UShort vertBearingX vertBearingY max_advance_width fontFile FT_CharMapRec_ horiAdvance FT_GLYPH_FORMAT_OUTLINE FT_SubGlyphRec_ yMin FT_CharMap oldColour FT_LibraryRec_ num_faces platform_id FT_GLYPH_FORMAT_NONE FT_Size_InternalRec_ encoding_id FT_Size FT_BBox FT_Stream_IoFunc num_fixed_sizes xOffset ../src/gfx/text.cpp lsb_delta linearVertAdvance FT_Short FT_Slot_InternalRec_ _Z12RefreshFontsv FT_Bitmap_Size_ linearHoriAdvance horiBearingX horiBearingY FT_Face_InternalRec_ FT_ListNode ../src/gfx/font.cpp FT_Incremental_InterfaceRec FT_Err_Corrupted_Font_Glyphs select_size FT_Err_Too_Many_Extensions bearing_x bearing_y FT_Raster_BitTest_Func ft_smooth_lcd_renderer_class done_size module_flags FT_Span FT_Module_Interface glyph_size FT_RENDER_MODE_LCD FT_Data module_data FT_ULong FT_Raster_Funcs FT_Size_SelectFunc FT_Err_Debug_OpCode FT_Err_Too_Many_Function_Defs FT_Glyph_Class_ FT_Err_Corrupted_Font_Header FT_Err_Unlisted_Object ft_smooth_renderer_class FT_RasterRec_ /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base/ftinit.c FT_SIZE_REQUEST_TYPE_SCALES FT_GlyphLoaderRec_ FT_Glyph_DoneFunc service_POSTSCRIPT_FONT_NAME FT_Err_Invalid_Size_Handle FT_SpanFunc FT_Err_Missing_Bbx_Field FT_Err_Could_Not_Find_Context FT_Err_Too_Many_Caches GNU C89 8.2.0 -mno-sse -mno-sse2 -mno-mmx -mtune=generic -march=x86-64 -g -O2 -ansi -fvisibility=hidden FT_Int32 FT_New_Library FT_Renderer_Class_ FT_ServiceCacheRec_ FT_Face_DoneFunc FT_Incremental_MetricsRec glyph_transformed FT_SIZE_REQUEST_TYPE_REAL_DIM FT_Err_Invalid_CharMap_Format FT_Err_Invalid_Horiz_Metrics ft_default_raster FT_Err_Raster_Corrupted FT_Err_Divide_By_Zero no_stem_darkening service_METRICS_VARIATIONS get_glyph_cbox FT_Err_Invalid_PPem FT_Module_Constructor FT_Incremental_GetGlyphDataFunc FT_Err_Out_Of_Memory FT_Err_Table_Missing FT_Incremental_FuncsRec_ vertResolution bit_test FT_Renderer FT_Raster_Params FT_Err_Invalid_Version FT_ModuleRec_ FT_Err_Cannot_Open_Resource psaux_module_class FT_ModuleRec FT_Err_Nested_Frame_Access FT_Incremental_FuncsRec use_extra FT_Renderer_RenderFunc FT_Module_Class_ max_subglyphs init_size FT_DebugHook_Func FT_Raster_ResetFunc incremental_interface auto_hinter t1cid_driver_class FT_Err_Invalid_Vert_Metrics FT_Err_Invalid_Composite extra_points2 clip_box FT_Incremental FT_Err_Invalid_Argument module_interface FT_Pointer FT_Err_Invalid_Stream_Handle FT_Err_Invalid_Glyph_Index cur_renderer glyph_prepare FT_Err_Invalid_Slot_Handle refcount module_init FT_Incremental_MetricsRec_ FT_SIZE_REQUEST_TYPE_MAX FT_Err_Bad_Argument FT_Char ft_raster1_renderer_class glyph_loader transform_delta FT_GlyphLoader bdf_driver_class transform_flags FT_Err_CMap_Table_Missing FT_Err_Invalid_Offset FT_Err_Name_Table_Missing FT_Done_Library service_PFR_METRICS black_spans FT_Err_Invalid_Post_Table_Format face_object_size FT_RENDER_MODE_LIGHT FT_Err_Cannot_Open_Stream FT_Error FT_Err_Invalid_Pixel_Size FT_Err_Stack_Overflow FT_Err_Invalid_Character_Code property_value glyph_copy FT_Size_Request_Type FT_Err_Raster_Overflow FT_Size_Request FT_Err_ENDF_In_Exec_Stream FT_Err_Glyph_Too_Big FT_Err_Too_Many_Instruction_Defs FT_Err_Invalid_Handle FT_Slot_InitFunc alibrary FT_Err_Missing_Font_Field FT_Err_Invalid_CharMap_Handle get_glyph_metrics FT_GlyphRec_ FT_Module_Class autofit_module_class done_slot target FT_Err_Invalid_Stream_Seek FT_Err_DEF_In_Glyf_Bytecode FT_Err_Invalid_Opcode FT_Driver_ClassRec_ FT_Err_Invalid_Library_Handle ft_smooth_lcdv_renderer_class FT_Err_Invalid_Outline FT_Raster_BitSet_Func FT_Glyph_TransformFunc FT_Renderer_Class FT_Err_Unimplemented_Feature FT_Size_RequestRec_ ft_property_string_set renderers FT_Glyph FT_Module_Requester FT_RENDER_MODE_LCD_V FT_Err_Too_Many_Hints psnames_module_class bit_set version_patch FT_Glyph_InitFunc FT_Driver_ClassRec service_MULTI_MASTERS FT_Err_Missing_Bitmap init_slot FT_Err_Ok FT_Renderer_SetModeFunc version_minor FT_Err_Array_Too_Large FT_Err_Post_Table_Missing FT_GlyphLoadRec FT_Err_Missing_Property FT_Err_Horiz_Header_Missing max_points FT_IncrementalRec_ FT_Err_Lower_Module_Version FT_Face_InitFunc winfnt_driver_class FT_Raster_Funcs_ module_version faces_list module_done FT_Err_Cannot_Render_Glyph cff_driver_class transform_matrix FT_Size_InitFunc load_flags FT_Err_Execution_Too_Long num_modules property_name FT_Add_Module FT_Slot_LoadFunc pcf_driver_class FT_Face_GetAdvancesFunc FT_Incremental_GetGlyphMetricsFunc FT_Err_Invalid_Table glyph_format FT_Err_Missing_Size_Field FT_Module_Destructor FT_Raster_NewFunc FT_Driver_Class FT_Render_Mode FT_Err_Missing_Startfont_Field FT_Incremental_InterfaceRec_ FT_Glyph_PrepareFunc FT_Glyph_GetBBoxFunc FT_Err_Invalid_Frame_Operation t1_driver_class version_major FT_Raster_SetModeFunc FT_Raster_DoneFunc FT_Renderer_GetCBoxFunc glyph_matrix FT_Module FT_Err_Missing_Chars_Field FT_Add_Default_Modules FT_Set_Default_Properties FT_Bool FT_Err_Ignore advance_v glyph_transform pshinter_module_class autohint_metrics FT_Err_Nested_DEFS FT_Span_ FT_Init_FreeType FT_Err_Invalid_File_Format t42_driver_class size_object_size FT_Err_Invalid_CodeRange FT_Matrix request_size horiResolution FT_Err_Invalid_Face_Handle extra_points FT_Err_Invalid_Glyph_Format max_contours FT_Err_Missing_Module gray_spans FT_Err_Invalid_Driver_Handle FT_Size_Request_Type_ FT_Err_Code_Overflow module_name FT_Err_No_Unicode_Glyph_Name FT_Err_Invalid_Stream_Skip FT_Err_Missing_Fontboundingbox_Field FT_Parameter_ FT_Err_Invalid_Stream_Read ft_default_modules FT_Size_DoneFunc FT_RENDER_MODE_MONO FT_Parameter FT_Renderer_TransformFunc service_GLYPH_DICT service_WINFNT FT_Err_Missing_Encoding_Field FT_Face_GetKerningFunc FT_Err_Locations_Missing FT_Raster_RenderFunc glyph_delta FT_SIZE_REQUEST_TYPE_NOMINAL sfnt_module_class FT_ServiceCacheRec tt_driver_class glyph_hints FT_Err_Raster_Negative_Height FT_Err_Raster_Uninitialized FT_Data_ FT_Err_Invalid_Post_Table FT_Byte module_requires lcd_geometry FT_Err_Too_Few_Arguments FT_Done_Memory FT_Face_AttachFunc pfr_driver_class transform_glyph FT_Raster FT_Render_Mode_ FT_Glyph_CopyFunc render_glyph FT_Err_Too_Many_Drivers FT_Raster_Params_ FT_SIZE_REQUEST_TYPE_BBOX FT_GlyphLoadRec_ FT_Err_Bbx_Too_Big FT_SIZE_REQUEST_TYPE_CELL attach_file FT_RENDER_MODE_MAX FT_Glyph_Class raster_class FT_Incremental_FreeGlyphDataFunc FT_Err_Invalid_Reference FT_Err_Missing_Startchar_Field FT_Err_Invalid_Stream_Operation module_size FT_Matrix_ debug_hooks autohint_mode FT_Err_Hmtx_Table_Missing FT_Err_Invalid_Cache_Handle glyph_class FT_RENDER_MODE_NORMAL FT_Err_Stack_Underflow FT_Err_Max FT_New_Memory FT_Err_Invalid_Frame_Read /home/computerfido/Desktop/LemonTest/build-freetype FT_Done_FreeType slot_object_size FT_Size_RequestFunc FT_Err_Unknown_File_Format FT_RendererRec_ FT_Err_Syntax_Error FT_Slot_DoneFunc glyph_bbox FT_Property_Get version_number CheckSum_Adjust ft_raccess_sort_ref_by_id font_program_size FT_Frame_Op_ vertical vec1 vec2 glyph_locations FT_GlyphLoad FT_Set_Char_Size GX_BlendRec_ num_layers FT_Sfnt_Tag_ rdata_len isFixedPitch instructions maxInstructionDefs TT_SBit_Scale FT_UInt64 ft_glyphslot_alloc_bitmap FT_Properties_SetFunc usWeightClass p_index xMax_Extent xAvgCharWidth hash_str_compare TT_Get_Name_ID_Func SFNT_Interface_ block2 TT_MaxProfile FT_Properties_GetFunc TT_GaspRec result_offset ft_frame_schar FT_Stream_ReadUOffset FT_New_Face panose debug_hook min_origin_SB reset_face TT_SbitTableType_ num_kern_tables FT_Service_TrueTypeEngine glyf_offset ft_service_list_lookup FT_Stream_ExtractFrame FT_AutoHinter_InterfaceRec_ hori errors file_size ft_frame_short_le hash_insert first_point FT_GlyphLoader_Add access_glyph_frame Mac_Read_sfnt_Resource strstr result_file_name short_metrics FT_SFNT_TableGetFunc error_code doblend FT_Get_Sfnt_Table kern_order_bits kern_avail_bits FT_Get_Module_Interface FT_RFork_Rule_linux_cap FT_Palette_Data_ FT_GlyphLoader_CheckPoints ft_frame_end driver_name palette_index max_profile FT_Outline_Get_CBox ft_frame_ushort_le FT_Get_Font_Format ft_hash_str_insert nouse padvance TT_Post_20Rec_ FT_LcdFilter_ test_mac_fonts map_len raccess_guess_apple_generic _ft_face_scale_advances FT_Hash args2 kern_table_size pixel_width ft_hash_num_init face_index_in_resource ft_hash_str_init FT_Outline_Transform var_postscript_prefix FT_SFNT_HEAD yshift FT_Get_Kerning FT_MulFix ulUnicodeRange3 FT_Face_GetVariantSelectors forget_glyph_frame advance_Height_Max FT_GlyphDict_GetNameFunc maxCompositePoints set_palette maxStorage p_arg2 subg xshift langID anoutline FT_RFork_Rule_darwin_ufs_export usWidthClass FT_TrueTypeEngineType maxPPEM FT_CMapRec_ original_name engine_type FT_RFork_Rule_ ft_glyphslot_done Line_Gap FT_New_Size aslot in_y FT_ServiceDescRec astream raccess_guess_linux_double stringOffset structure is_sfnt_cid sbit_num_strikes FT_Get_Postscript_Name FT_Get_Sfnt_Name_Count FT_LcdFilter FT_PIXEL_MODE_GRAY FT_CharMapRec FT_GlyphLoader_Done pfb_len left_bearing FT_Vector_Transform __builtin_memset languageID p_arg1 FT_Offset fsSelection SFNT_Service apalette Fail agindex FT_Vector_Unit min_advance_SB v_prev hash_bucket ySubscriptYSize entry_length maxMemType42 TT_Loader_StartGlyphFunc angle1 angle2 acmap FT_DriverRec FT_Stream_Read FT_Property_Set ft_frame_bytes ft_cmap_done_internal vcmap TT_GaspRangeRec_ FT_SFNT_OS2 pfb_lenpos TT_Postscript_ FT_Matrix_Invert service_id numPoints FT_Stream_New aminor raccess_guess_linux_cap FT_Vector_NormLen FT_Set_Charmap achVendID ulUnicodeRange1 ulUnicodeRange2 ulUnicodeRange4 head2 FT_LCD_FILTER_MAX vert_resolution FT_Get_First_Char last_charmap horz_resolution get_track FT_RFork_Rule_darwin_hfsplus new_count FT_ServiceDesc hash_num_compare maxComponentDepth palette_entry_name_ids minMemType42 TT_TableRec_ FT_Angle_Diff ft_mem_dup Index_To_Loc_Format FT_Stream_EnterFrame FT_Vector_Polarize FT_Hashkey_ FT_Service_GlyphDictRec_ hash_init hdmx_record_count TT_SBIT_TABLE_TYPE_NONE FT_Stream_ReadUShortLE caret_slope_denominator FT_ValidationLevel_ usFirstCharIndex FT_AutoHinter_Interface TT_Load_Any_Func p_error is_cff ft_hash_num_insert load_eblc FT_Set_Transform FT_SFNT_POST size_index buffer_max FT_PIXEL_MODE_GRAY2 FT_PIXEL_MODE_GRAY4 padvances ttface FT_Raccess_Guess is_owner d_hypot sfnt_data get_table TT_Header desc theta FT_Atan2 Modified FT_CMap_ClassRec_ FT_Stream_GetUOffset get_global_hints FT_Face_GetCharVariantIndex linear_def FT_Get_Charmap_Index raccess_guess_apple_single variantSelector char_height rfork_offset ft_mem_realloc TT_Header_ v_start destroy_face TT_Post_NamesRec FT_LCD_FILTER_DEFAULT exec FT_Cos Load_Ok FT_MulFix_x86_64 ySubscriptXOffset FT_Set_Pixel_Sizes end0 FT_Load_Glyph FT_List_Iterate num_locations FT_CMap_DoneFunc right_glyph variantchar_list TT_Blend_Colr_Func FontNumber var_postscript_prefix_len TT_Get_Metrics_Func external_stream TT_Face_GetKerningFunc number_Of_HMetrics stream2 FT_Frame_Field FT_Error_String FT_Hashnode min_Right_Side_Bearing ft_validator_run FT_SFNT_TableInfoFunc maxContours FT_PIXEL_MODE_LCD TT_Face Mac_Read_POST_Resource usWinDescent TT_GlyphZoneRec TT_SBIT_TABLE_TYPE_SBIX glyph_indices ins_pos hook_index swap FT_Vector_Rotate ft_open_face_internal render_mode file_names palette_name_ids FT_Service_Kerning language ft_raccess_rule_by_darwin_vfs FT_Stream_Seek temp2 TT_Name cmap_size memory_stream_close TT_NameTableRec_ allzeros FT_Matrix_Multiply_Scaled usMaxContext ystrength ft_frame_skip jmp_buf FT_Get_CMap_Format FT_List_Finalize FT_Get_Track_Kerning TT_MaxProfile_ usBreakChar FT_ORIENTATION_NONE acbox strncpy degree char_width sTypoLineGap magic_from_stream cvt_program_size FT_Hypot pads TT_Get_PS_Name_Func CharacterComplement FT_Service_TTCMapsRec_ frame_accessed FT_Outline_ConicToFunc FT_GlyphLoader_New FT_Remove_Module new_max FT_Attach_Stream FT_Stream_Free Font_Direction FT_Outline_EmboldenXY FT_CMap_CharVariantListFunc FT_PIXEL_MODE_MAX darken_params cur_size resource_cnt FT_Load_Sfnt_Table is_light_type1 ulCodePageRange1 ulCodePageRange2 FT_CMap_CharVarIsDefaultFunc maxFunctionDefs rpos ft_glyphslot_init error1 error2 FT_Service_PropertiesRec_ numLangTagRecords FT_SfntName_ FT_DivFix FT_CMap_Class FT_Vector_From_Polar maxPoints FT_Palette_Select null_palette_data FT_Outline_MoveToFunc FT_TRUETYPE_ENGINE_TYPE_PATENTED advance_Width_Max free_psnames Table_Version ft_corner_is_flat old_max FT_Stream_Open TT_LangTagRec_ TT_Loader_EndGlyphFunc num_sbit_scales font_program FT_Get_Char_Index FT_Service_SFNT_Table ps_property_get n_base_points caret_slope_numerator TT_Interpreter langTags horizontal x_left set_property FT_Request_Metrics FT_MulDiv_No_Round FT_Select_Charmap FT_PIXEL_MODE_LCD_V TT_Post_25Rec long_metrics missing_func FT_ValidatorRec_ num_tables numRanges v_middle vfs_rfork_has_no_font FT_SFNT_VHEA Destroy_Module FT_KERNING_DEFAULT nameID Calculate_Ppem FT_Get_Name_Index FT_RFork_Rule FT_ServiceDescRec_ FT_Stream_GetUShort sTypoDescender IsMacBinary FT_ORIENTATION_POSTSCRIPT ySuperscriptXSize FT_GlyphLoader_CreateExtra xtemp FT_FaceRec TT_VertHeader_ FT_Outline_Reverse FT_Open_Face FT_Service_GlyphDict cvt_program raccess_guess_apple_double ft_mem_strdup read_composite_glyph FT_Get_CMap_Language_ID d_in FT_RFork_Rule_linux_double numGlyphs platformID ps_property_set FT_PIXEL_MODE_NONE TT_SBit_LineMetricsRec FT_List_Insert d_out hdmx_record_size FT_Set_Renderer FT_CMap_CharVarIndexFunc FT_Select_Size FT_AutoHinter_GlobalDoneFunc longjmp raccess_guess_linux_netatalk FT_TRUETYPE_ENGINE_TYPE_UNPATENTED Magic_Number FT_CMap ft_mem_qalloc FT_SFNT_HHEA FT_Get_Renderer char_var_default TT_SBit_LineMetricsRec_ arctanptr FT_GlyphLoader_Adjust_Points FT_GlyphLoader_Prepare raccess_guess_linux_double_from_file_name TT_CMap_Info_GetFunc FT_GlyphDict_NameIndexFunc FT_Raccess_Get_HeaderInfo FT_AutoHinter_GlobalGetFunc hash_lookup number_Of_VMetrics FT_RFork_Rule_vfat TT_SBit_MetricsRec num_palette_entries sbit_strike_map TT_OS2_ FT_Set_Debug_Hook maxComponentElements x_shift top_bearing yMax_Extent FT_GlyphLoader_Rewind free_eblc ft_recompute_scaled_metrics ft_lookup_PS_in_sfnt_stream serv_data variation_support FT_VALIDATE_DEFAULT ySubscriptYOffset maxMemType1 ySuperscriptXOffset y_ppem_substitute alangTag v_control PS_DriverRec_ ft_raccess_guess_rec FT_Get_TrueType_Engine_Type Lowest_Rec_PPEM FT_Raccess_Get_DataOffsets FT_Stream_GetChar TT_OS2 min_after_BL aname PS_Driver Created FT_ORIENTATION_TRUETYPE __builtin_memcpy FT_New_GlyphSlot FT_SFNT_MAXP level ft_synthesize_vertical_metrics result FT_Outline_New raccess_guess_darwin_ufs_export parameters jump_buffer strings_size ft_frame_uoff3_be encodingID Fail2 hdmx_table TT_Done_Face_Func raccess_guess_darwin_hfsplus TT_Get_Name_Func open_face read_glyph_header FT_Library_Version TT_Load_Table_Func numNameRecords FT_Library_SetLcdFilterWeights is_num FT_Done_Face StrokeWeight TT_Post_25_ FT_Stream_Pos vert_metrics_offset tag_internal sCapHeight filepathname FT_Face_Properties FT_Outline_Funcs_ vert_metrics_size FT_CMap_Done FT_Color_ FT_Stream_ReadULong FT_Orientation_ TT_NameRec get_psname FT_Matrix_Check x_ppem_substitute raccess_guess_vfat FT_Color num_params TT_BDFRec FT_CMap_CharNextFunc ptrdiff_t TTC_HeaderRec TT_ExecContext FT_GlyphLoader_CheckSubGlyphs FT_Outline_LineToFunc FT_CMap_CharIndexFunc sbit_table green FT_RFork_Rule_apple_double FT_Palette_Data_Get nonzero_minval max_before_BL FT_LayerIterator_ ft_glyphslot_clear usLowerOpticalPointSize new_memory_stream stringLength entry_offset FT_F26Dot6 FT_AutoHinter_GlobalResetFunc FT_Stream_GetULong maxStackElements caret_Offset FT_KERNING_UNSCALED FT_PtrDist FT_Get_Glyph_Name have_layers aface TT_HoriHeader FT_List_Add maxCompositeContours caret_Slope_Run FT_Get_Sfnt_Name SymbolSet TT_CMapInfo_ find_variant_selector_charmap sfnt_ps subcnt TT_Load_Strike_Metrics_Func FT_Stream_ReadAt pbytes new_name FormatType TT_Free_Table_Func ft_frame_off3_be TT_Loader_GotoTableFunc kern_table v_cur memory_base pbox akerning usWinAscent TT_PCLT_ FT_Service_KerningRec_ TT_SBIT_TABLE_TYPE_CBLC yStrikeoutSize destroy_size dlen FT_SfntLangTag ft_glyphslot_preset_bitmap FT_Outline_Get_Orientation is_cff2 FT_Load_Char FT_HashnodeRec_ FT_List_Destructor FT_Stream_ReleaseFrame FT_Service_Properties FT_Pixel_Mode_ ft_trig_arctan_table ft_glyphslot_grid_fit_metrics Mac_Style num_names FT_Sfnt_Tag l_anchor TT_CMapInfo TT_SbitTableType FT_Reference_Face map_pos ft_mem_alloc TypeFace apatch FT_RFork_Ref is_darwin_vfs ebdt_size ft_frame_byte FT_Vector_Length base_file_name num_palettes FileName FT_Match_Size ySuperscriptYOffset hdmx_record_sizes TT_SizeRec_ name_table FT_Outline_Translate FT_Stream_ExitFrame yStrikeoutPosition FT_Outline_Embolden FT_SFNT_PCLT gaspFlag FT_Size_RequestRec FT_Sin FT_Tag FT_Tan Fail3 TT_Load_Metrics_Func FT_TRUETYPE_ENGINE_TYPE_NONE y_shift FT_Face_GetCharVariantIsDefault num_properties ft_module_get_service TT_Postscript new_names newpath TT_Loader_ReadGlyphFunc FT_Open_Args_ kern_mode ft_trig_prenorm ft_lookup_glyph_renderer FT_Done_GlyphSlot FT_Frame_Field_ FT_Get_Advances memory_size FT_Outline_Decompose table_end TT_BDFRec_ FT_RFork_Rule_uknown p_transform pfb_pos horz_metrics_size FT_SFNT_MAX FT_Stream_GetUShortLE FT_Stream_ReadFields FT_Kerning_TrackGetFunc face_index_internal max_width sub_index ft_frame_ulong_be numTables TT_Size bsize slash TT_Get_Colr_Layer_Func FT_Hash_LookupFunc serv_id resource_fork_entry_id FT_PsName_GetFunc maxval done_global_hints FT_LCD_FILTER_NONE FT_MulDiv base_file_len _tmp_ TT_Init_Face_Func strlen abitmap FT_Render_Glyph caret_Slope_Rise sxHeight insertion TT_Load_SBit_Image_Func acolor_index FT_Open_Args FT_Service_PsFontName ft_frame_long_be FT_ORIENTATION_FILL_RIGHT FT_LCD_FILTER_LIGHT FT_Select_Metrics FT_Hashkey ySuperscriptYSize sFamilyClass ft_hash_str_free FT_GlyphLoader_Adjust_Subglyphs pstable_index data_offsets FT_Stream_ReadULongLE ft_frame_uoff3_le read_simple_glyph hash_rehash FT_LCD_FILTER_LEGACY1 FT_Get_SubGlyph_Info temp1 psaux CheckSum FT_FloorFix open_face_from_buffer FT_Stream_ReadUShort FT_Service_TTCMaps FT_Get_Sfnt_LangTag usUpperOpticalPointSize TT_Loader TT_HoriHeader_ FT_SFNT_TableLoadFunc maxZones FT_Get_Color_Glyph_Layer Font_Revision FT_List_Remove metric_Data_Format ft_property_do raccess_make_file_name FT_RFork_Rule_linux_netatalk aloader TT_LangTag SFNT_Interface init_data FT_RFork_Rule_apple_single TT_Set_SBit_Strike_Func FT_RFork_Ref_ FT_AutoHinterRec_ value_is_string TT_Post_20Rec FT_Stream_TryRead FT_LCD_FILTER_LEGACY FT_Get_Module interpreter TTC_HeaderRec_ reads scaled_w FT_Int64 func_interface FT_ORIENTATION_FILL_LEFT sfnt FT_List_Up TT_SBit_MetricsRec_ FT_SfntName ft_raccess_guess_func TT_FaceRec_ TT_LangTagRec underlineThickness strcat scaled_h ft_remove_renderer FT_RFork_Rule_darwin_newvfs Do_Conic null_outline FT_HashRec_ open_face_PS_from_sfnt_stream cmap_table mod_name FT_TrueTypeEngineType_ orig_x orig_y before glyf_len load_mac_face aglyph_index in_x FT_List TT_GlyphZoneRec_ FT_Palette_Set_Foreground_Color flag_offset FT_CMap_VariantCharListFunc FT_Palette_Data new_length TypeFamily TT_SBIT_TABLE_TYPE_MAX horz_metrics_offset composites fsType ft_validator_init find_unicode_charmap resource_offset FT_Stream_ReadChar FT_ValidationLevel TT_PCLT TT_Load_Face_Func usLastCharIndex TT_Set_Palette_Func pfb_data ebdt_start ft_glyphslot_set_bitmap left_glyph FT_Stream_Close FT_Sfnt_Table_Info ft_frame_off3_le FT_AutoHinter_GlyphLoadFunc FT_Outline_Funcs ft_corner_orientation FT_KERNING_UNFITTED FT_RFork_Rule_invalid postscript_names usDefaultChar FT_Get_Advance ft_frame_start ft_raccess_guess_table n_curr_contours TT_Gasp_ ft_raccess_guess_rec_ gloader ySubscriptXSize FT_Face_GetCharsOfVariant FT_Orientation offsets_internal apalette_data FT_Reference_Library memmove FT_New_Memory_Face FT_CMap_New IsMacResource n_subs FT_Library_SetLcdGeometry TT_Table raccess_get_rule_type_from_rule_index Success numContours FT_CMap_VariantListFunc FT_Get_Next_Char ucmap min_Top_Side_Bearing min_Bottom_Side_Bearing p_flags dir_tables sbit_table_type maxTwilightPoints FT_CeilFix ft_frame_ulong_le ft_add_renderer FT_Activate_Size filter ft_lcd_padding out_x out_y Units_Per_EM ft_glyphslot_free_bitmap ft_hash_num_lookup FT_Incremental_Interface FT_Pixel_Mode pixel_height FT_LayerIterator base_name FT_Stream_OpenMemory ignore_width item_size gaspRanges FT_Service_PsFontNameRec_ italicAngle FT_Service_TrueTypeEngineRec_ minMemType1 TT_NameTableRec asize FT_List_Iterator colr_blend ft_trig_pseudo_polarize min_Left_Side_Bearing cur_count alpha FT_Outline_Get_Bitmap FT_Service_SFNT_TableRec_ TT_GaspRange destroy_charmaps FT_Angle FT_CMap_InitFunc ft_set_current_renderer hdmx_table_size raccess_guess_darwin_newvfs type_list language_id hinting_engine WidthType FT_Request_Size SerifStyle palette_flags sTypoAscender ft_frame_ushort_be external /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base/ftbase.c area FT_Hash_CompareFunc TT_ExecContextRec_ FT_Library_SetLcdFilter ft_validator_error FT_Matrix_Multiply service_descriptors FT_Outline_Done sign_shift ft_trig_pseudo_rotate ft_mem_qrealloc amajor FT_PIXEL_MODE_BGRA TT_Post_NamesRec_ ft_frame_long_le FT_UInt16 n_of_entries sort_by_res_id FT_Stream_GetULongLE FT_RoundFix load_table FT_Outline_CubicToFunc ft_mem_free ft_trig_downscale ft_hash_str_lookup Exit2 FT_AutoHinter TT_SBit_ScaleRec_ FT_Face_GetVariantsOfChar FT_PIXEL_MODE_MONO strrchr origin TT_LoaderRec_ xstrength FT_Done_Size FT_Vector_Transform_Scaled FT_VALIDATE_TIGHT Glyph_Data_Format GX_Blend FT_Render_Glyph_Internal ft_mem_strcpyn cvt_size FT_VALIDATE_PARANOID FT_Outline_Render read_bytes FT_List_Find FT_Get_X11_Font_Format FT_Validator FT_Kerning_Mode_ TT_VertHeader sbit_table_size ttc_header Reserved have_foreground_color FT_Attach_File ft_frame_short_be FT_SfntLangTag_ new_size load_face_in_embedded_rfork allmatch FT_GlyphLoader_Reset rdata_pos underlinePosition storageOffset Destroy_Driver charvariant_list caret_offset TT_NameRec_ FT_Outline_Check format_tag TT_SBIT_TABLE_TYPE_EBLC FT_Outline_Copy FT_Stream_Skip v_last FT_Lookup_Renderer maxSizeOfInstructions TT_Err_Invalid_Table TT_Err_Invalid_CharMap_Format Ins_SHP TT_Err_Syntax_Error inline_delta tt_face_load_loca nIfs TT_Err_Invalid_Reference is_composite tt_size_reset dualVector GX_HVVarTableRec_ old_range sfnt_id out1 out2 FT_SizeRec TT_Err_Missing_Font_Field codeRangeTable TT_Err_Invalid_Stream_Operation TT_DotFix14_long_long TT_Err_Horiz_Header_Missing TT_Err_Raster_Overflow axisSize Update_Max TT_Err_Too_Many_Function_Defs tt_coderange_font FT_Service_MultiMastersRec_ GX_TC_RESERVED_TUPLE_FLAGS FT_Multi_Master_ GX_TI_RESERVED_TUPLE_FLAG strid avalue cur_range shortDeltaCount delta_cnt storage tt_prepare_zone innerIndex projVector TT_CallRec dummy2 Ins_GETINFO TT_Err_Name_Table_Missing compensations startCoord TT_Project_Func tt_service_properties storage_size cvt_ready tt_size_run_fpgm TT_Err_Glyph_Too_Big TT_Err_Ignore codeSize Compute_Point_Displacement mvar_hlgp_delta FT_F2Dot14 netAdjustment FT_Get_MM_Var_Func TT_CallRec_ all_design_coords Round_None Ins_S45ROUND TT_Err_Invalid_Horiz_Metrics Ins_ODD Ins_SFVTPV Caller_IP tt_size_init y_ratio namedstyle tt_loader_set_pp Ins_MPS Ins_JMPR aIdx1 aIdx2 next_coords_size GX_AVarCorrespondenceRec_ TT_CodeRange_ gv_glyphcnt GX_ItemVarStoreRec_ tt_face_load_prep iupx_called old_point_delta_x old_point_delta_y Ins_GPV start_contour GX_DeltaSetIdxMap tt_get_var_blend Compute_Round Ins_INSTCTRL incr_metrics F_dot_P localpoints tt_driver_done opcode rotated Ins_DEBUG Ins_PUSHB TT_Err_Hmtx_Table_Missing ref2 TT_Process_Simple_Glyph Ins_DIV iupy_called discriminant TT_Err_Invalid_Face_Handle Ins_PUSHW instanceSize TT_Err_Invalid_Stream_Read Ins_SHC control_value_cutin TT_Err_Invalid_Pixel_Size Ins_SHZ psid refp GetShortIns func_write_cvt tt_check_trickyness_sfnt_ids Ins_NPUSHB TT_Err_Missing_Fontboundingbox_Field FT_Set_MM_Design_Func TT_Err_Locations_Missing Ins_CLEAR Ins_NPUSHW grayscale get_mm Ins_FLIPRGOFF GX_TI_INTERMEDIATE_TUPLE instruct_control unrounded GX_VarRegionRec_ Current_Ppem num_axis TT_Init_Glyph_Loading im_start_coords TT_Err_Invalid_Offset TT_Clear_CodeRange Ins_NROUND TT_Process_Composite_Component tt_face_vary_cvt Ins_RTHG TT_Load_Context Ins_DELTAC Ins_FLIPON tt_face_done_loca FT_HAdvance_Adjust_Func cont_limit __builtin_strcmp Exit1 tt_face_load_hdmx TT_Err_Invalid_Library_Handle Round_To_Double_Grid Move_CVT_Stretched incr Ins_UNKNOWN Ins_SCANCTRL Round_Super node2 scan_control dotproduct Ins_SFVTL TT_Err_Invalid_File_Format Ins_RTG cur1 cur2 FT_Get_MM_Blend_Func Round_Down_To_Grid ft_var_to_normalized Normalize TT_GraphicsState_ FT_Var_Axis_ TT_Err_Out_Of_Memory TT_RunIns TT_Err_Invalid_Glyph_Format curs tt_face_free_hdmx Ins_SMD cur_dist vvar_table varData TT_Err_Invalid_Driver_Handle Ins_SANGW table_len GX_TI_PRIVATE_POINT_NUMBERS next_name FT_Service_PropertiesRec axisCoords glyphSize tt_service_gx_multi_masters delta2 TT_CodeRange_Tag_ IUP_Worker end_point Ins_LTEQ ttsize TT_CodeRangeTable hvar_error glyphoffsets FT_Set_MM_Blend_Func FT_Service_TrueTypeEngineRec current_outline header_only mapData Round_Up_To_Grid namedstyle_size new_top mvar_tag LErrorCodeOverflow_ loopcall_counter_max subglyph FT_VAdvance_Adjust_Func round_state ft_var_get_value_pointer TT_Err_Missing_Bitmap GX_DeltaSetIdxMapRec_ Ins_MDRP Ins_ENDF GX_TC_TUPLE_COUNT_MASK TT_Err_Ok Ins_NOT num_axes stackSize subpixel_hinting_lean TT_Err_DEF_In_Glyf_Bytecode Ins_EQ tt_size_ready_bytecode TT_Err_Raster_Uninitialized FT_Set_MM_WeightVector_Func dataSize point_cnt tupleIndex tt_face_load_fpgm coderange TT_Err_Invalid_Version FT_Get_Var_Design_Func has_fpgm outerIndex rsb_adjust tt_get_kerning Ins_IP do_scale Direct_Move_X TT_Set_MM_Blend TT_Err_Table_Missing step_ins p_limit _pbuff Ins_MDAP vertical_lcd_lean TT_GlyphSlot Ins_ABS sharedpoints func_round tt_size_run_prep TT_Set_Var_Design TT_Err_Corrupted_Font_Glyphs Ins_EIF TT_Err_Missing_Encoding_Field tt_interpolate_deltas axisTag tt_size_select TT_Err_Invalid_CodeRange vvar_error Ins_SSW GX_FVar_Head Ins_MSIRP TT_DefRecord_ tt_size_init_bytecode Ins_WCVTF TT_Err_Too_Many_Drivers reexecute Ins_ADD widthMap_offset TT_Err_Missing_Module TT_Err_Invalid_Stream_Skip TT_Load_Simple_Glyph TT_Err_Stack_Underflow regionCount points_out TT_Err_Execution_Too_Long Ins_GT flag_limit Round_To_Grid callStack instanceCount ttslot Ins_SUB Project_x axisCount innerBitCount in_points cvtEntry table_start TT_Err_Unimplemented_Feature tt_driver_init GX_AxisCoords GX_DeltaSetIdxMapRec default_GS func_project Ins_SZP0 Ins_SZP1 Ins_SZP2 TT_Access_Glyph_Frame FT_Service_MetricsVariationsRec _iup_worker_interpolate instruction_trap has_cvt TT_DefArray TT_Err_Lower_Module_Version LNo_Error_ n_ins Ins_FLOOR tt_glyph_load glyphCount vec_limit tt_vadvance_adjust need_init opcode_length single_width_value Ins_AA tt_get_metrics_incr_overrides Ins_IUP TT_Load_Glyph TT_DefRecord max_function_defs num_function_defs tt_glyphzone_new Ins_SWAP Caller_Range phase TT_Err_Invalid_Post_Table Ins_EVEN TT_Err_Invalid_Slot_Handle round_mode Ins_IF numIDefs func_read_cvt tuplecoords TT_Err_Invalid_CharMap_Handle Dual_Project fvaraxis_fields correspondence GX_VarRegion prev_cont func_cur_ppem TT_Forget_Glyph_Frame tt_hvadvance_adjust TT_Err_Bbx_Too_Big Ins_IDEF Ins_CEILING touch Init_Context cvt_deltas TT_Err_Missing_Bbx_Field first_delta TT_Err_ENDF_In_Exec_Stream tupleCount num_coords FExit TT_Size_Metrics fvar_fields TT_Err_Bad_Argument ft_var_load_mvar tt_apply_mvar TT_Err_Corrupted_Font_Header ref1 neg_jump_counter_max SetSuperRound Ins_ISECT manageCvt nump tt_check_trickyness_family TT_Err_Invalid_Opcode TT_Err_Missing_Startfont_Field TT_Err_Stack_Overflow max_ins set_mm_design Fail_Memory tt_services GX_TC_TUPLES_SHARE_POINT_NUMBERS GX_GVar_Head first_touched regionIdxCount tt_property_get scale_valid dummy1 numFDefs FT_VOrg_Adjust_Func Ins_DEPTH TT_Goto_CodeRange sph_fdef_flags glyphIns endCoord ft_var_apply_tuple tt_default_graphics_state Ins_WCVTP tt_sfnt_id_rec_ defaultValue tt_interface vvar_checked avar_segment neg_jump_counter tt_hadvance_adjust subpixel_hinting Ins_Goto_CodeRange Ins_SPVTL Compute_Funcs FT_Set_Instance_Func Ins_RTDG TT_Err_Max func_move_cvt TT_Round_Func Ins_AND period TT_Get_VMetrics inc_stream pedantic_hinting scalar callSize Ins_JROF TT_Set_Named_Instance majorVersion Round_Super_45 /home/computerfido/Desktop/LemonTest/lemon-freetype/src/truetype/truetype.c TT_Err_Cannot_Render_Glyph TT_Err_Could_Not_Find_Context has_delta TT_Err_Too_Many_Hints tt_get_advances tt_size_request mcvt_retain interpreter_version TT_Size_Metrics_ TT_Driver multiplier GX_TupleIndexFlags_ Ins_UTP glyph_data_loaded num_matched_ids tt_synth_sfnt_checksum func_dualproj TT_Err_Invalid_Vert_Metrics orgs Direct_Move minimum_distance Direct_Move_Y Ins_SROUND mapCount ft_var_load_gvar GX_MVarTableRec_ tt_face_get_location Direct_Move_Orig_Y axisList tt_done_blend itemStore maxFunc callrec gep0 gep1 offsetToCoord FT_Set_Var_Design_Func valueCount runcnt tt_face_init FT_StreamRec Ins_SZPS only_height mac_yscale TT_Err_Raster_Negative_Height varRegionList Ins_LT tt_service_metrics_variations sfntd Ins_MIN tt_sfnt_id_rec pairCount num_instances TT_GraphicsState Ins_MD vorg_adjust TT_LoaderRec Fail_Overflow Ins_FLIPOFF TT_Err_Cannot_Open_Stream bsb_adjust FT_UnitVector_ Ins_SRP0 Ins_SRP1 Ins_SRP2 pindex Ins_SxyTCA max_instruction_defs tt_get_interface FT_Get_Var_Blend_Func Ins_NEQ old_stream mvar_table deltaSet TT_Run_Context axis_size Ins_NEG mmvar ft_var_get_item_delta load_truetype_glyph Move_Zp2_Point cur_delta Ins_MPPEM normalized_stylecoords TT_Get_HMetrics num_base_points tt_check_trickyness Ins_GETDATA Ins_MAX use_aw_2 Ins_OR in_twilight FT_Var_Named_Style tt_property_set GX_ItemVarStore opened_frame size_metrics tmp_o TT_Get_CVT_Func TT_Err_Missing_Chars_Field FT_UnitVector FT_MM_Axis_ cvt_dist Direct_Move_Orig_X TT_Err_Too_Many_Caches ft_var_readpackedpoints fvar_start TT_Err_Cannot_Open_Resource maxIns ft_var_load_hvvar spoint_count Ins_RCVT context Ins_CINDEX ft_var_readpackeddeltas axis_rec next_coords num_designs grayscale_cleartype lsb_adjust new_dist tt_cvt_ready_iterator ft_var_load_avar tsb_adjust Ins_POP worker hvar_table vvar_loaded TT_Load_Composite_Glyph TT_Err_CMap_Table_Missing tt_size_done_bytecode TT_CallStack single_width_cutin Ins_ROFF FT_MM_Var peak FT_Service_TTGlyfRec_ num_base_subgs FT_TSB_Adjust_Func TT_Save_Context Ins_RS GX_ItemVarDataRec_ peakCoord innerIndexMask Ins_MIAP set_design_coords _iup_worker_shift SkipCode Ins_SCFS compensation x_ratio Current_Ratio linear_vadvance toCoord TT_Err_Code_Overflow TT_Err_Invalid_Stream_Seek TT_Err_Debug_OpCode TT_Set_CodeRange pedantic tt_loader_done ftsize FT_Int16 ft_var_to_design FT_Metrics_Adjust_Func func_freeProj tt_slot_init TT_Set_CVT_Func Ins_FLIPRGON FT_Done_Blend_Func FT_Service_TTGlyfRec num_records FT_MM_Axis TT_Err_Invalid_Size_Handle fvar_axis_ TT_Err_Invalid_PPem pointSize tmp_r TT_Err_Invalid_Post_Table_Format current_line_gap GX_AVarSegment GX_Value FT_Get_MM_WeightVector_Func Current_Ppem_Stretched named_style tt_delta_interpolate widthp hvar_loaded auto_flip normalizedcoords widthMap FT_Get_MM_Func im_end_coords aRange sbit_metrics minValue num_instruction_defs TT_Err_Missing_Startchar_Field TT_Get_Var_Design gep2 TT_Err_Invalid_Cache_Handle tuplecount TT_Process_Composite_Glyph FT_Service_MetricsVariationsRec_ out_points cur_touched mvar_hasc_delta GX_FVar_Head_ Ins_SFVFS TT_Load_Glyph_Header GX_AVarCorrespondence offsetToData Ins_SPVFS Ins_SSWCI Ins_WS old_cvt_delta GX_ItemVarData FT_MM_Var_ FT_Multi_Master mcvt_load avar_loaded Ins_FLIPPT Ins_ROLL func_move TT_Err_Unknown_File_Format Ins_GETVARIATION GX_HVVarTable new_loca_len curRange maximum Ins_MUL scaledDelta linear_hadvance Ins_SxVTL Ins_CALL TT_CodeRange storeSize LSuiteLabel_ func_move_orig Direct_Move_Orig tt_size_reset_iterator Cur_Count Ins_ALIGNPTS Project_y TT_Get_MM_Var have_diff Read_CVT_Stretched IUP_WorkerRec_ cvtSize TT_Err_Raster_Corrupted region_offset tt_get_sfnt_checksum mac_xscale max_func Ins_SLOOP ft_var_load_item_variation_store GX_TI_TUPLE_INDEX_MASK GX_TupleCountFlags_ axis_flags points_org maxValue gvar_fields delta_base callTop TT_New_Context tt_check_single_notdef axis_flags_size point_deltas_x GX_ItemVarStoreRec point_deltas_y fvar_head mmvar_size Ins_GTEQ Ins_RDTG gvar_head TT_Err_Invalid_Handle here Ins_MINDEX GX_AVarSegmentRec_ orus1 orus2 Ins_LOOPCALL tt_metrics Pop_Push_Count regionIndex stretched Ins_SDPVTL minimum recurse_count tt_get_metrics Ins_SCANTYPE GX_MVarTable TT_Err_Invalid_Composite gvar_start TT_DriverRec_ TT_Err_Invalid_Character_Code delta1 has_prep TT_Err_Nested_Frame_Access cur_base call ttdriver ins_counter TT_Err_Nested_DEFS trick_names regionIndices Ins_FDEF TT_Err_Invalid_Frame_Operation mcvt_modify tt_size_done tt_coderange_glyph tt_face_load_cvt Ins_MIRP ttmetrics Ins_SDB FT_BSB_Adjust_Func Ins_SHPIX Write_CVT TT_Get_MM_Blend TT_Err_Too_Many_Instruction_Defs tt_coderange_cvt tt_face_done Ins_SDS next_name_size fromCoord Round_To_Half_Grid Ins_GC Ins_JROT ft_var_load_delta_set_index_mapping Ins_ELSE TT_Err_Invalid_Stream_Handle freeVector tt_coderange_none TT_Err_Too_Many_Extensions orus_base itemCount maxFDefs tuple_coords bytecode_ready tupleDataSize tt_service_truetype_engine byte_count TT_Err_Post_Table_Missing usePsName Ins_DUP Ins_ALIGNRP tt_delta_shift TT_Err_Missing_Property TT_Err_Array_Too_Large Move_CVT Ins_ROUND Bad_Format have_scale FT_Var_Axis scan_type TT_Move_Func globalCoordCount org_dist GX_FVar_Axis glyf_table_only TT_Err_Divide_By_Zero GX_GVar_Head_ tt_face_get_device_metrics TT_Err_Unlisted_Object tt_loader_init TT_Glyf_GetLocationFunc Ins_RUTG gvar_size tt_glyphzone_done loop TT_Err_Too_Few_Arguments ft_list_get_node_at IUP_WorkerRec entrySize tt_service_truetype_glyf hvar_checked Ins_SCVTCI ft_var_done_item_variation_store TT_Err_Invalid_Frame_Read Fail1 GridPeriod TT_GlyphZone Ins_GFV TT_Err_Invalid_Glyph_Index mmvar_len xy_size TT_Vary_Apply_Glyph_Deltas backward_compatibility tt_set_mm_blend num_twilight_points TT_Err_Invalid_Argument FT_Service_MultiMastersRec Read_CVT GX_ValueRec_ TT_Cur_Ppem_Func dataCount maxIDefs num_points pCrec org1 FT_Var_Named_Style_ org2 FT_LSB_Adjust_Func TT_Err_No_Unicode_Glyph_Name Write_CVT_Stretched loopcall_counter hinted_metrics GX_AxisCoordsRec_ TT_MulFix14_long_long Ins_DELTAP TT_Err_Invalid_Outline unmodified TT_Hint_Glyph old_byte_len GX_TI_EMBEDDED_TUPLE_COORD TT_Err_Missing_Size_Field num_namedstyles FT_RSB_Adjust_Func LErrorLabel_ dataOffsetArray mvar_hdsc_delta TT_Done_Context records_offset compute_glyph_metrics mm_axis_unmap header_string T1_Err_Invalid_File_Format CFF_SubFontRec_ t1_services t1_make_subfont num_other_blues axis_count T1_Err_Ignore PS_GetFontInfoFunc local_subrs_offset t1_cmap_classes cff_decoder_funcs PSH_Globals PS_BlendRec_ PS_DICT_RND_STEM_UP PS_DICT_FONT_NAME sids T1_Err_Invalid_Composite T1_Err_Invalid_Vert_Metrics T1_Token T1_GlyphSlot PS_DICT_BLUE_SHIFT t1glyph top_font CFF_Builder_Add_Contour_Func units_per_em t1_get_name_index PS_DICT_ENCODING_ENTRY num_blue_values T1_FIELD_TYPE_NONE PSH_Globals_Funcs T1_FIELD_LOCATION_FACE T1_ParseState parser CFF_VarRegion num_hints incremental get_glyph_callback design_pos t1_ps_get_font_extra global_subrs_index num_strings AFM_FontInfo PS_Private T1_Driver_Done T1_Load_Glyph max_elems point_tokens T1_Err_Cannot_Open_Resource PS_DICT_OTHER_BLUE T1_Err_Too_Many_Extensions paint_type ps_parser_funcs T1_FontRec adobe_expert_encoding AFM_Parser_FuncsRec_ italic_angle code_last CFF_Size T1_Err_Corrupted_Font_Header T1_Err_DEF_In_Glyf_Bytecode PS_FontExtraRec T1_TokenRec_ T1_Builder_Check_Points_Func PS_DICT_SUBR PS_Parser_FuncsRec_ parse_blend_design_positions T1_Loader T2_HintsRec_ pos_lf CFF_PrivateRec_ CFF_Decoder_FuncsRec CFF_Decoder_ font_offset t1_get_ps_name cid_uid_base global_subrs T1_Parse_Start T1_Err_Divide_By_Zero width_table_length parse_weight_vector FT_CMapRec PS_FontInfoRec_ PS_DICT_NUM_FAMILY_BLUES PS_DICT_WEIGHT parse_private T1_Err_Invalid_Glyph_Index PS_DICT_BLUE_VALUE charset_offset axiscoords single_block blue_scale PSH_Globals_SetScaleFunc T1_Err_Invalid_Stream_Skip T1_Err_Invalid_Offset PS_UniMap T1_Get_MM_WeightVector nominal_width PS_TableRec T1_FIELD_LOCATION_LOADER T1_Get_Var_Design keywords_encountered T1_FIELD_TYPE_MM_BBOX PS_DICT_FAMILY_OTHER_BLUE read_width PS_ParserRec_ PS_FontExtraRec_ T1_FIELD_TYPE_FIXED T1_Err_Invalid_Post_Table_Format the_same PS_Builder_FuncsRec char_string standard_height T1_ParserRec t1_decrypt T1_EncodingRecRec_ CFF_AxisCoords test_cr PS_Dict_Keys cid_count cid_ordering path_begun font_dict_index T1_TokenType t1_get_glyph_name lengths PS_DICT_NUM_OTHER_BLUES usedBV pos_x pos_y PS_DICT_FAMILY_NAME PS_DICT_STD_HW array_size vstore_offset in_memory afm_data charstrings_offset t1_decoder_funcs t1_font PS_DICT_BLUE_FUZZ CFF_Decoder_Get_Glyph_Callback T1_Err_Invalid_Frame_Operation PS_GetGlyphNameFunc T1_FIELD_TYPE_FIXED_1000 private_size T1_Set_MM_Blend PS_GetFontValueFunc T1_Driver_Init token2 t1_ps_get_font_private T1_Err_Table_Missing hints_globals T1_Err_Too_Many_Function_Defs PS_DICT_UNDERLINE_THICKNESS T1_Err_Too_Many_Caches PS_DICT_PASSWORD string_pool private_len CFF_Builder_Start_Point_Func len_buildchar CFF_EncodingRec notdef_glyph parse_subrs T1_Err_ENDF_In_Exec_Stream AFM_ParserRec T1_Err_Too_Many_Hints T1_FIELD_TYPE_STRING cid_font_version T1_FIELD_TYPE_BOOL encoding_table T2_Hints_MaskFunc T1_Done_Metrics private_offset encode start_binary lcoords T1_Err_Invalid_CharMap_Handle t1size PS_DICT_FORCE_BOLD FT_Service_KerningRec t1_builder_funcs swap_table have_integer T1_Err_Raster_Uninitialized T1_Err_Cannot_Render_Glyph T1_FIELD_TYPE_BBOX PS_Decoder_ lenIV vstore PS_UnicodesRec_ T1_DecoderRec ndv_idx strncmp PS_DICT_CHAR_STRING T1_Err_Too_Few_Arguments CFF_IndexRec CFF_SubFontRec T1_EncodingType T1_Err_Bad_Argument CFF_Decoder_FuncsRec_ blue_fuzz T1_Field off_size Again locals_bias FontBBox local_subrs_index T1_TOKEN_TYPE_NONE PS_DICT_NUM_CHAR_STRINGS T1_Face_Done T1_Decoder_Callback CFF_FDSelectRec T1_Set_MM_WeightVector T1_Reset_MM_Blend AFM_Parser T1_ENCODING_TYPE_ISOLATIN1 cid_registry t1_get_index num_locals T1_Field_ParseFunc cid_fd_array_offset glyph_names_block temp_scale T1_Decoder_ZoneRec T1_LoaderRec T1_Finalize_Parser T1_Err_Invalid_Argument is_t1 PSHinter_Service hintmask T1_Err_Invalid_Handle T1_Parse_Have_Width T1_Err_Invalid_CodeRange design_tokens PS_DICT_NOTICE T1_FIELD_LOCATION_BLEND t1_done_loader afont_extra T2_Hints_OpenFunc AFM_Stream globals_bias T1_Err_Missing_Startchar_Field T1_Err_Invalid_Version t1_service_properties force_scaling T1_Hints_SetStem3Func CFF_FDSelectRec_ PS_Table_FuncsRec CFF_FontRecDictRec start_pos PSH_Globals_DestroyFunc builtBV T2_Hints_Funcs initial_random_seed T1_Encoding PS_DICT_NUM_SUBRS T1_Err_Invalid_Stream_Handle lastVsindex n_axis pshinter T1_Compute_Max_Advance T1_Err_Invalid_Library_Handle T1_FIELD_LOCATION_FONT_EXTRA PS_PrivateRec FT_Service_PsCMaps T1_Err_Missing_Fontboundingbox_Field check_type1_format parse_callback parse_state width_only num_flex_vectors T1_EncodingType_ T2_Hints_FuncsRec_ T1_Err_Post_Table_Missing T1_FieldRec embedded_postscript PS_Decoder_Zone CFF_FontRecDictRec_ T1_Err_Invalid_Stream_Operation FT_Service_PsCMapsRec_ unique_id T1_Size T1_Err_Bbx_Too_Big T1_FIELD_TYPE_MAX range_count PS_DICT_PAINT_TYPE FT_Service_PsInfoRec_ charmaprecs t1_service_kerning PS_DICT_IS_FIXED_PITCH T1_FaceRec CFF_CharsetRec_ read_binary_data data_offset PS_Table_FuncsRec_ T1_Hints_ResetFunc CFF_BlendRec_ T1_Builder_Close_Contour_Func T1_FIELD_LOCATION_PRIVATE T1_Decoder_FuncsRec_ T2_Hints max_objects T1_Err_Horiz_Header_Missing no_recurse array_max cache_first blue_shift t1_set_mm_blend t1_parse_font_matrix T1_Err_Syntax_Error notice T1_Err_Stack_Overflow T1_BuilderRec_ synthetic_base T1_Err_Invalid_Frame_Read PS_DICT_ENCODING_TYPE glyph2 ident T1_Get_Kerning PS_DICT_MIN_FEATURE ps_table_funcs T1_Builder_Add_Point_Func flex_state PS_DICT_NUM_BLUE_VALUES T1_Err_Stack_Underflow T1_Err_Invalid_Size_Handle password T1_Hints T1_Read_Metrics T1_Builder_FuncsRec_ cache_fd T1_Decoder_ZoneRec_ notdef_found psdecoder T2_Hints_CloseFunc PS_DICT_NUM_STEM_SNAP_H t1_face PS_DICT_NUM_STEM_SNAP_V T1_Err_Out_Of_Memory T1_ParserRec_ PS_DesignMap_ num_elems T1_Err_Invalid_PPem T1_Err_Invalid_Slot_Handle T1_Err_Missing_Startfont_Field max_ptsize T1_Builder_Start_Point_Func round_stem_up PS_GetFontExtraFunc CFF_Builder_Close_Contour_Func PS_HasGlyphNamesFunc PS_Unicodes_CharIndexFunc T1_FieldLocation_ T1_GlyphSlot_Done custom count_offset T1_FontRec_ full_name T1_Err_Raster_Corrupted T1_Err_Code_Overflow CFF_Decoder T1_Err_Missing_Module T1_Get_MM_Blend CFF_Builder_Check_Points_Func num_snap_heights T1_Size_Request PS_DICT_FONT_BBOX T1_Err_Missing_Font_Field T1_ENCODING_TYPE_EXPERT T1_Font code_table T1_Err_Invalid_Reference subrs_block ps_decoder_init T1_Err_No_Unicode_Glyph_Name blend_top design_points T1_Err_Hmtx_Table_Missing adobe_std_strings T1_FieldLocation index1 index2 encoding_offset PS_Blend pair2 final_blends PS_Builder_FuncsRec_ T1_Err_Invalid_Driver_Handle t1_service_glyph_dict language_group CFF_VarRegion_ min_feature T1_FieldType_ glyph1 T1_Get_Private_Dict old_cursor T1_Err_Cannot_Open_Stream PS_DICT_FS_TYPE T1_Hints_Funcs T1_Decoder_Funcs adobe_std_encoding T1_Decoder_Zone cid_font_type CFF_Builder_ T1_Err_Invalid_Glyph_Format PSHinter_Interface T1_Get_Track_Kerning TrackKerns CFF_VarData_ PS_Macintosh_NameFunc default_weight_vector T1_BuilderRec T1_Hints_OpenFunc T1_Size_Get_Globals_Funcs PS_DesignMap PS_DICT_STEM_SNAP_H point_token T2_Hints_StemsFunc CFF_EncodingRec_ only_immediates CFF_Builder_FuncsRec PS_DICT_STEM_SNAP_V cff_random T1_Set_MM_Design T1_Err_Invalid_Outline /home/computerfido/Desktop/LemonTest/lemon-freetype/src/type1/type1.c T1_TOKEN_TYPE_ARRAY PS_DICT_FAMILY_BLUE PS_Decoder_Zone_ bboxes afont_private T1_Parse_Glyph_And_Get_Char_String num_family_other_blues notdef_index PS_Adobe_Std_StringsFunc T1_Loader_ AFM_TrackKern T1_Err_Lower_Module_Version num_chars base_offset font_infos t1_allocate_blend num_default_design_vector CFF_Builder_Add_Point_Func current_subfont weight T1_TOKEN_TYPE_KEY T1_Decoder cid_supplement NumTrackKern T1_Err_Corrupted_Font_Glyphs CFF_SubFont T1_Get_Advances user_data midi CFF_GlyphSlotRec_ T1_Face_Init IsCIDFont fontdata T1_HintsRec_ CFF_PrivateRec code_first dummy_object T1_Err_Invalid_Table AFM_KernPairRec_ charstrings_block T1_Get_Multi_Master CFF_VarData CFF_Builder PSH_GlobalsRec_ T1_GlyphSlot_Init T1_Builder_Add_Point1_Func base_dict T1_Builder_FuncsRec AFM_StreamRec_ T1_DecoderRec_ cffload atag blend_alloc T1_FIELD_TYPE_INTEGER hdr_size oldcharmap T1_Open_Face PS_FontInfo T2_Hints_ApplyFunc T1_Private charstrings_len T1_Get_MM_Var PSH_Globals_NewFunc T1_Err_Could_Not_Find_Context CFF_SizeRec_ T1_FIELD_LOCATION_CID_INFO PS_Builder T1_Err_Nested_Frame_Access cid_font_revision T1_Err_Nested_DEFS min_kern font_dict stroke_width cid_font_name PSAux_Service T1_ENCODING_TYPE_STANDARD AFM_KernPair T1_Parse_Have_Path T1_New_Parser t1_interface CFF_GlyphSlot subrs_len CFF_CharsetRec PSHinter_Interface_ PS_Table PS_Unicodes_CharNextFunc subrs_hash value_len_ CFF_IndexRec_ PS_TableRec_ __builtin_memcmp axis_token max_kern CFF_VStoreRec_ top_dict_index T1_Err_Ok blend_points PS_FreeGlyphNameFunc default_width T1_Done_Blend full PS_Decoder T1_TOKEN_TYPE_MAX gname T1_Size_Init axismap FT_Service_PsFontNameRec T1_Err_Debug_OpCode PS_DICT_VERSION PSH_Globals_FuncsRec_ T1_Err_Raster_Negative_Height CFF_Decoder_Zone_ PS_BlendRec T1_Hints_ApplyFunc num_snap_widths T1_EncodingRec locals_hash T1_FIELD_LOCATION_MAX p_design parse_blend_axis_types fs_type PS_DICT_LEN_IV T1_Err_Unknown_File_Format num_globals pair1 PS_DICT_LANGUAGE_GROUP char_name CFF_FontRec_ FT_Service_GlyphDictRec capacity T1_Err_Missing_Size_Field KernPairs T1_ParseState_ T1_Err_Invalid_Character_Code PS_FontInfoRec CFF_Font min_ptsize PS_Unicodes_InitFunc T1_ENCODING_TYPE_NONE max_cid T1_Parse_Glyph T1_Err_Invalid_Cache_Handle axis_names parse_buildchar T2_Hints_CounterFunc T1_FaceRec_ T1_Err_Name_Table_Missing AFM_Parser_FuncsRec charstrings_index T1_Err_Invalid_Pixel_Size the_blend T1_FIELD_LOCATION_BBOX FT_GlyphSlotRec T1_Err_Raster_Overflow T1_Err_Missing_Bitmap base_len T1_CMap_Classes hints_funcs blend_bitflags T1_TOKEN_TYPE_ANY copyright t1_keywords T1_Err_Too_Many_Drivers header_length T1_FIELD_TYPE_FIXED_ARRAY T1_Err_Missing_Bbx_Field T1_TOKEN_TYPE_STRING T1_Err_Too_Many_Instruction_Defs CFF_BlendRec read_pfb_tag PS_Unicode_ValueFunc PS_Dict_Keys_ T1_Err_Missing_Chars_Field private_index T1_Read_PFM T1_SizeRec_ lenBV T1_Err_Execution_Too_Long memchr force_bold num_subfonts t1_load_keyword T1_Err_Max T1_FieldRec_ afont_info T1_Size_Done T1_Err_Locations_Missing num_maps mmaster PS_DesignMapRec in_pfb T1_FIELD_LOCATION_FONT_INFO T1_FieldType encoding_type T1_Err_Invalid_Horiz_Metrics CFF_Builder_FuncsRec_ T1_TokenRec T1_Parser min_char num_family_blues PS_DICT_UNDERLINE_POSITION NumKernPair lenNDV PS_Parser_FuncsRec standard_width T1_FIELD_TYPE_INTEGER_ARRAY PS_DICT_MAX cache_count afm_parser_funcs T1_FIELD_TYPE_CALLBACK max_char T1_Err_Invalid_Post_Table old_limit T1_Hints_FuncsRec_ PS_DICT_NUM_FAMILY_OTHER_BLUES T1_Builder PS_ParserRec T1_Parse_Have_Moveto t1_service_ps_name is_fixed_pitch PS_DICT_CHAR_STRING_KEY must_finish_decoder cid_fd_select_offset T1_GlyphSlotRec_ retval PS_Unicodes T1_TokenType_ glyph_width blend_used T1_Err_Glyph_Too_Big force_bold_threshold PS_UniMap_ T1_Err_Invalid_Opcode PS_Builder_ header_size T1_Hints_SetStemFunc T1_Builder_Add_Contour_Func reader PS_PrivateRec_ cf2_instance t1_ps_get_font_info blend_stack T1_Err_Unlisted_Object cdv_idx FT_Service_PsInfoRec AFM_ParserRec_ value_len t1_service_ps_info T1_Decoder_FuncsRec CFF_Decoder_Free_Glyph_Callback PS_DICT_STD_VW T1_Err_Invalid_CharMap_Format T1_Err_Missing_Encoding_Field T1_Err_Unimplemented_Feature privates free_glyph_callback T1_Err_Invalid_Face_Handle PS_DICT_BLUE_SCALE has_font_matrix T1_Err_Invalid_Stream_Read fd_select T1_Err_Invalid_Stream_Seek T1_Err_Missing_Property parse_blend_design_map PS_DICT_UNIQUE_ID top_dict_length PS_GetFontPrivateFunc PS_DICT_FONT_MATRIX data_size CFF_VStoreRec PS_DICT_ITALIC_ANGLE T1_Err_Array_Too_Large CFF_Builder_Add_Point1_Func CFF_AxisCoords_ AFM_FontInfoRec_ locals_len T1_Hints_CloseFunc string_pool_size mm_weights_unmap T1_FIELD_LOCATION_FONT_DICT num_subrs metrics_only dummy T1_Face PSAux_ServiceRec_ PS_DICT_FULL_NAME T1_CMap_ClassesRec_ t1_ps_has_glyph_names local_subrs T1_ENCODING_TYPE_ARRAY lastNDV T1_Set_Var_Design standard axis_tokens t1_service_multi_masters AFM_TrackKernRec_ CFF_Decoder_Zone t1_init_loader PS_Parser t1face T1_FIELD_TYPE_KEY t1_ps_get_font_value T1_Err_CMap_Table_Missing PS_DICT_FONT_TYPE FT_CMap_ClassRec Populate cff_hadvance_adjust CFF_Err_Too_Many_Hints cff_parse_vsindex CFF_Err_Nested_DEFS start_def FT_CID_GetIsInternallyCIDKeyedFunc CFF_Err_Bad_Argument CFF_FDSelect CFF_Err_Invalid_Stream_Operation cff_parse_font_matrix CFF_Err_Invalid_Frame_Operation cff_slot_done axisScalar cff_get_kerning FT_Blend_Build_Vector_Func CFF_Parser CFF_Err_Invalid_Opcode exponent_sign have_overflow CFF_Err_Too_Many_Instruction_Defs start14 cff_parse_fixed cff_service_get_cmap_info num_ranges CFF_InternalRec_ pbyte_len cff_charset_cid_to_gindex cff_get_cid_from_glyph_index FT_CID_GetRegistryOrderingSupplementFunc numOperands CFF_Err_Missing_Property cff_make_private_dict cff_vstore_done CFF_Err_Invalid_CharMap_Handle CFF_Err_Invalid_Reference cff_get_var_design cff_cmap_unicode_class_rec qcount subFont cff_service_ps_info invert Store_Number cff_face_done csindex cff_get_glyph_data CFF_Err_No_Unicode_Glyph_Name cff_sid_to_glyph_name sub_upm sfnt_module CFF_Err_Invalid_Vert_Metrics CFF_Err_Invalid_CharMap_Format CFF_FontRec cff_field_handlers cff_service_cff_load cmaprec next_offset cff_kind_fixed_thousand CFF_Err_Invalid_Frame_Read cff_size_done cff_blend_build_vector FT_Service_TTCMapsRec glyph_sid CFF_Err_Too_Many_Function_Defs cff_set_mm_blend cff_kind_max end14 cff_parse_private_dict CFF_FontRecDict CFF_Err_Unimplemented_Feature CFF_Err_Missing_Size_Field pchar_code CFF_Err_Missing_Bbx_Field CFF_Private CFF_Err_Invalid_Stream_Seek cff_encoding_done CFF_Err_Invalid_Size_Handle cff_load_private_dict CFF_Err_Invalid_Face_Handle cff_get_mm_weightvector cff_fd_select_get FT_Service_MultiMasters org_bytes cff_font_done CFF_VStore CFF_Err_Missing_Font_Field power_ten_limits CFF_Charset cffslot CFF_Err_CMap_Table_Missing CFF_ParserRec cff_cmap_encoding_done cff_size_request cff_get_mm_var FT_Service_CFFLoadRec_ CFF_Err_Debug_OpCode CFF_Err_Name_Table_Missing cff_charset_done cff_get_ps_name CFF_Err_Invalid_File_Format cff_parse_fixed_dynamic cff_cmap_encoding_class_rec cff_get_advances FT_FD_Select_Get_Func cff_service_multi_masters CFF_Internal CFF_Field_Reader FT_Service_CIDRec CFF_Err_Invalid_Library_Handle CFF_ParserRec_ cff_blend_doBlend CFF_Err_Lower_Module_Version remove_style p_end CFF_Err_Hmtx_Table_Missing cff_index_get_pointers topfont poff cff_kind_fixed style_name_length cff_size_get_globals_funcs CFF_Err_Raster_Overflow power_ten CFF_Err_Table_Missing CFF_Err_Too_Few_Arguments cff_parser_run errorp min_scaling cff_service_ps_name CFF_Load_FD_Select cff_get_ros CFF_Err_Invalid_Composite cff_index_get_name CFF_Err_Invalid_Driver_Handle cff_size_init CFF_Err_Cannot_Open_Stream cff_header_fields cff_kind_bool cff_parse_real FT_Service_CFFLoadRec cff_cmap_encoding_init CFF_Err_Invalid_CodeRange CFF_Err_Cannot_Open_Resource cff_service_properties CFF_Err_Array_Too_Large FT_CID_GetCIDFromGlyphIndexFunc CFF_Err_Invalid_Handle sfnt_format new_bytes CFF_Field_Handler_ cff_cmap_unicode_init CFF_Err_Unlisted_Object peak14 cffface cff_parser_done CFF_Index cff_get_mm_blend cff_isoadobe_charset vsOffset cff_services CFF_Err_Missing_Encoding_Field CFF_Err_Missing_Startchar_Field CFF_Field_Handler fullp regionListOffset blend_top_old /home/computerfido/Desktop/LemonTest/lemon-freetype/src/cff/cff.c CFF_Err_Corrupted_Font_Glyphs numBlends family_name_length CFF_Err_Corrupted_Font_Header cff_slot_init cff_blend_clear cff_set_var_design Missing_Table CFF_Err_Invalid_Slot_Handle CFF_Err_Invalid_Outline cur_offset CFF_Err_Locations_Missing CFF_Err_Too_Many_Drivers CFF_Err_Invalid_Post_Table FT_Blend_Check_Vector_Func exponent_add blend_stack_old CFF_Blend cff_get_interface CFF_Err_Ignore cff_index_forget_element CFF_Err_Stack_Underflow cff_size_select CFF_Err_Execution_Too_Long CFF_Err_Invalid_Offset CFF_Err_Horiz_Header_Missing charstring_len CFF_Err_Post_Table_Missing cff_free_glyph_data half_divisor num_args subfont_index CFF_Err_Syntax_Error FT_Load_Private_Dict_Func region cff_get_is_cid max_scaling top_upm glyph_code integer_length cff_kind_num cff_expert_encoding CFF_Encoding cff_index_init string_index CFF_Err_Invalid_Table cff_parse_maxstack CFF_Done_FD_Select cff_get_cmap_info CFF_Err_Invalid_PPem CFF_Err_Ok FT_Get_Standard_Encoding_Func CFF_Face CFF_Err_Raster_Uninitialized cff_service_metrics_variations cff_ps_get_font_info cpriv cff_vstore_load CFF_Err_Missing_Bitmap Skip_Unicode CFF_Err_ENDF_In_Exec_Stream CFF_Err_Invalid_Stream_Read cff_cmap_encoding_char_index varRegion cff_parse_blend cff_ps_has_glyph_names CFF_Err_Invalid_Pixel_Size cff_index_access_element cff_parse_multiple_master do_fixed cff_kind_string CFF_Err_Too_Many_Caches cff_index_done CFF_Err_Code_Overflow CFF_Err_Invalid_Horiz_Metrics CFF_Err_Invalid_Argument cff_get_name_index CFF_Err_Invalid_Cache_Handle continue_search CFF_Err_Raster_Negative_Height CFF_Err_Missing_Chars_Field dict_len cff_driver_done cff_slot_load CFF_Err_DEF_In_Glyf_Bytecode cff_get_var_blend CFF_Err_Invalid_Character_Code cff_get_standard_encoding gids cff_expertsubset_charset CFF_Err_Invalid_Glyph_Format CFF_Err_Out_Of_Memory cff_blend_check_vector CFF_Err_Bbx_Too_Big fdselect CFF_Err_Raster_Corrupted cff_expert_charset cff_set_mm_weightvector scalings CFF_Err_Invalid_Stream_Handle cff_index_get_string cff_metrics_adjust cff_charset_free_cids cff_ps_get_font_extra CFF_Err_Could_Not_Find_Context CFF_Err_Invalid_Version Glyph_Build_Finished cff_parse_integer cff_subfont_load cff_cmap_encoding_char_next exponent cff_cmap_unicode_char_index remove_subset_prefix CFF_Decoder_Funcs pure_cff cff_glyph_load Unlikely kind cff_done_blend cff_subfont_done cff_parser_within_limits CFF_Err_Stack_Overflow has_vertical_info cff_kind_callback CFF_Err_Invalid_Glyph_Index cff_get_glyph_name CFF_Err_Unknown_File_Format absolute_offset object_code cff_encoding_load CFF_Err_Invalid_Stream_Skip nleft cff_index_get_sid_string offsize CFF_Err_Invalid_Post_Table_Format cff_face cff_kind_blend cff_parse_num CFF_Err_Glyph_Too_Big cff_cmap_unicode_done cffsize cff_parser_init fd_index CFF_Err_Divide_By_Zero cff_cmap_unicode_char_next cff_font_load cff_parse_fixed_scaled Load_Data CFF_Err_Missing_Fontboundingbox_Field cff_kind_delta start_fstype cff_index_load_offsets cff_parse_font_bbox cff_charset_compute_cids cff_standard_encoding CFF_Err_Max CFF_CMapStdRec_ new_fraction_length Fail_CID cff_service_cid_info cff_charset_load CFF_Err_Missing_Startfont_Field cff_set_instance CFF_Err_Nested_Frame_Access CFF_Err_Missing_Module cff_strcpy cff_driver_init FT_Service_CFFLoad cff_parse_cid_ros FT_Service_MetricsVariations power_tens cff_index_read_offset FT_Service_CIDRec_ cff_face_init cff_service_glyph_dict CFF_CMapStd CFF_Err_Cannot_Render_Glyph CFF_Err_Too_Many_Extensions cff_kind_none fd_bytes max_offsets cid_face_open CID_Err_ENDF_In_Exec_Stream cid_get_offset gd_bytes CID_Parser CID_Err_Invalid_Frame_Operation CID_Err_Stack_Underflow CID_Err_Invalid_CharMap_Format CID_Err_Invalid_CodeRange CID_Err_Glyph_Too_Big CID_Err_Hmtx_Table_Missing CID_Err_Missing_Chars_Field num_dict CID_Err_Missing_Property cid_size_request CID_Err_Code_Overflow CID_FaceDictRec_ CID_FaceInfoRec_ CID_Err_Raster_Uninitialized upper_nibble CID_Err_Horiz_Header_Missing subrmap_offset CID_Parser_ cid_done_loader CID_Loader CID_FaceDictRec CID_Err_Invalid_Stream_Seek cid_slot_load_glyph CID_Err_Raster_Overflow CID_Err_Missing_Size_Field CID_Err_Invalid_Stream_Operation cid_service_cid_info cid_subrs CID_Err_Invalid_Pixel_Size CID_Err_Missing_Bbx_Field parse_font_name CID_Err_Too_Many_Hints CID_Err_Missing_Fontboundingbox_Field CID_Err_Unknown_File_Format glyph_length CID_Err_Unlisted_Object CID_GlyphSlot CID_Err_Missing_Font_Field cid_driver_done cidface CID_Err_Unimplemented_Feature CID_Err_Table_Missing CID_Err_Invalid_Cache_Handle CID_Err_Invalid_Face_Handle CID_Face cidglyph cid_hex_to_binary CID_Err_Invalid_Outline cid_slot_done cid_version cid_face_done CID_Err_Invalid_Glyph_Format cid_services CID_Size CID_Err_Ignore cid_service_ps_name CID_Err_Invalid_Post_Table CID_Err_Corrupted_Font_Header cid_parse_font_matrix CID_Err_Too_Many_Extensions CID_Err_Could_Not_Find_Context CID_Err_DEF_In_Glyf_Bytecode newlimit cid_interface CID_Err_Post_Table_Missing dlimit CID_Err_Invalid_Handle cid_driver_init CID_Err_Raster_Negative_Height CID_Err_Divide_By_Zero CID_Err_No_Unicode_Glyph_Name CID_Err_Invalid_Stream_Handle font_dicts CID_Err_Invalid_Character_Code CID_Err_Lower_Module_Version binary_length CID_Err_Too_Many_Caches CID_Err_Invalid_Offset CID_Err_Max CID_Err_Ok CID_Err_Invalid_Library_Handle cid_get_interface CID_Err_Invalid_Reference CID_FaceInfo CID_Err_Too_Few_Arguments CID_Err_Too_Many_Drivers CID_SizeRec_ cid_get_ros CID_Err_Invalid_Opcode CID_Err_Stack_Overflow CID_FaceInfoRec CID_Err_Too_Many_Instruction_Defs forcebold_threshold CID_GlyphSlotRec_ CID_Err_Invalid_Composite CID_FaceDict CID_SubrsRec_ cid_ps_get_font_info cid_parser_done CID_Err_Name_Table_Missing CID_Err_Invalid_Version CID_Err_Bbx_Too_Big CID_Err_Missing_Module cid_get_cid_from_glyph_index CID_Loader_ cid_ps_get_font_extra /home/computerfido/Desktop/LemonTest/lemon-freetype/src/cid/type1cid.c CID_Err_Out_Of_Memory cid_service_ps_info cid_load_glyph CID_Err_Debug_OpCode CID_Err_Raster_Corrupted CID_Err_Missing_Startfont_Field cid_load_keyword oldpos CID_Subrs CID_Err_Invalid_File_Format CID_Err_Nested_Frame_Access plimit cidsize CID_Err_Nested_DEFS cid_size_get_globals_funcs CID_Err_Bad_Argument cid_slot_init CID_Err_Invalid_Argument CID_Err_Missing_Encoding_Field CID_Err_Invalid_Size_Handle read_len CID_Err_Cannot_Render_Glyph CID_Err_Invalid_Vert_Metrics CID_Err_Invalid_Horiz_Metrics sd_bytes num_dicts parse_expansion_factor cid_size_done cidmap_offset cid_get_postscript_name CID_Err_Invalid_Stream_Read CID_Err_Invalid_Glyph_Index CID_Err_Corrupted_Font_Glyphs CID_Err_Invalid_Stream_Skip CID_Err_Execution_Too_Long CID_Err_Invalid_Post_Table_Format CID_Err_Invalid_Table postscript_len CID_Err_Syntax_Error CID_Err_Invalid_CharMap_Handle cid_size_init ps_len CID_Err_Invalid_Slot_Handle parse_fd_array cid_field_records cid_get_is_cid CID_Err_Invalid_PPem CID_Err_Invalid_Frame_Read cid_stream stream_len CID_Err_Missing_Bitmap CID_Err_Too_Many_Function_Defs CID_Err_Invalid_Driver_Handle CID_Err_Array_Too_Large CID_Err_Cannot_Open_Resource CID_FaceRec_ CID_Err_Missing_Startchar_Field entry_len cid_service_properties CID_Err_Cannot_Open_Stream CID_Err_Locations_Missing cid_parse_dict cid_init_loader num_xuid CID_Err_CMap_Table_Missing cid_read_subrs cid_face_init cid_parser_new log_font bct_offset PFR_Err_Out_Of_Memory PFR_Err_Cannot_Render_Glyph PFR_Err_Missing_Startchar_Field base_adj num_items PFR_HeaderRec size1 pfr_cmap_done stroke_flags Found_Strike PFR_Err_Raster_Corrupted Failure PFR_Err_Name_Table_Missing phy_font_max_size phy_font_section_offset phys_offset acount PFR_Err_Missing_Property PFR_Err_Missing_Startfont_Field PFR_Err_Invalid_Driver_Handle max_subs pfr_phy_font_load PFR_Err_Invalid_Horiz_Metrics local gps_section_offset kern_items pfr_face_done aformat PFR_Err_Unimplemented_Feature FT_PFR_GetMetricsFunc PFR_LogFontRec num_vert num_log_fonts PFR_ExtraItem_ParseFunc char2 pair_count bct_max_size PFR_Err_Missing_Chars_Field PFR_Err_Too_Few_Arguments prev_code twobytes PFR_Err_Unlisted_Object pdata axsize pfr_get_kerning log_font_section_size PFR_Err_Divide_By_Zero PFR_Err_Ok item_list pfr_metrics_service_rec PFR_Err_Horiz_Header_Missing PFR_Err_Invalid_Cache_Handle item_data char1 pfr_cmap_char_next PFR_Err_Invalid_Reference pfr_extra_item_load_bitmap_info PFR_Err_Invalid_CharMap_Format PFR_Err_Invalid_File_Format log_font_max_size PFR_Err_Invalid_Face_Handle pfr_glyph_curve_to pfr_glyph_end PFR_Err_Max PFR_BitWriter_ PFR_Err_Too_Many_Function_Defs max_horz_stem_snap found_offset chars_offset PFR_SubGlyphRec_ PFR_Err_Invalid_Stream_Skip twobyte_adj stroke_thickness phys PFR_ExtraItem y_count pfr_glyph_load_simple pfr_glyph_close_contour old_points pfr_face_init PFR_DimensionRec_ ametrics_y_scale anadvance PFR_Err_CMap_Table_Missing font_ref_number PFR_Err_Too_Many_Caches log_dir_offset color_flags PFR_DimensionRec item_type PFR_Err_DEF_In_Glyf_Bytecode num_bitmaps PFR_Err_Corrupted_Font_Glyphs pair_size y_ppm PFR_Err_Missing_Fontboundingbox_Field Line1 pfr_extra_items_parse pfr_cmap_init PFR_Err_Missing_Encoding_Field PFR_BitWriter PFR_Err_Hmtx_Table_Missing pfr_get_metrics em_metrics max_xy_control PFR_Glyph FT_Service_PfrMetricsRec pfr_bitwriter_init anoutline_resolution PFR_BitmapCharRec_ pfr_extra_item_load_stem_snaps pfr_glyph_start writer PFR_Err_Invalid_Version phy_font Test_Error PFR_SubGlyphRec y_delta phy_bct_set_max_size PFR_CMapRec_ pfrsize max_y_orus PFR_Err_Lower_Module_Version PFR_Err_Cannot_Open_Stream PFR_Err_Invalid_Table bct_size probe FT_PFR_GetKerningFunc PFR_Err_Invalid_Slot_Handle PFR_BitWriterRec PFR_Err_Unknown_File_Format gps_max_size PFR_Err_Invalid_Stream_Read PFR_Err_Too_Many_Hints PFR_SubGlyph max_vert_stem_snap PFR_ExtraItemRec PFR_Err_Stack_Underflow kern_items_tail pfr_phy_font_done PFR_Err_Debug_OpCode standard_advance PFR_Header em_outline pfrface num_kern_pairs PFR_LogFont PFR_Char pfr_header_load pfr_face_get_kerning phy_font_max_size_high PFR_Err_Missing_Size_Field pfr_header_check pfr_cmap_class_rec Too_Short PFR_PhyFontRec_ pfr_glyph_move_to format_low pfr_glyph_load decreasing PFR_Err_Execution_Too_Long PFR_Err_Invalid_Composite PFR_Err_Invalid_Size_Handle char_len PFR_Err_Table_Missing num_aux FoundPair gps_offset pfr_glyph_done PFR_Err_Raster_Overflow PFR_Err_Invalid_Frame_Operation PFR_Err_Missing_Bbx_Field PFR_Err_Nested_DEFS pfr_get_service PFR_Err_Invalid_Vert_Metrics signature2 PFR_Err_Invalid_PPem PFR_Size PFR_Err_Code_Overflow PFR_Err_Invalid_Post_Table x_ppm PFR_StrikeRec ametrics_x_scale pfr_services miter_limit found_size pfr_phy_font_extra_items avector PFR_Err_Invalid_Post_Table_Format /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pfr/pfr.c control1 control2 PFR_KernItem PFR_Err_Ignore PFR_KernItemRec_ PFR_Err_Invalid_Offset PFR_Err_Raster_Negative_Height Restart power PFR_Err_Invalid_Stream_Operation PFR_Face PFR_Err_No_Unicode_Glyph_Name PFR_SizeRec_ PFR_Err_Invalid_CodeRange PFR_StrikeRec_ PFR_Err_Stack_Overflow pfrslot PFR_Err_Bad_Argument size_increment PFR_Err_Glyph_Too_Big pfr_cmap_char_index PFR_Err_Nested_Frame_Access PFR_Err_Invalid_Outline pfr_extra_items_skip PFR_Strike PFR_Err_Missing_Bitmap PFR_Err_Invalid_Handle PFR_Err_Array_Too_Large flags0 PFR_Err_Too_Many_Extensions PFR_LogFontRec_ FT_PFR_GetAdvanceFunc org_count PFR_ExtraItemRec_ PFR_Err_Corrupted_Font_Header PFR_Err_Syntax_Error Found_It log_font_section_offset PFR_Err_Invalid_Frame_Read scaled_advance pfr_get_advance PFR_Err_Invalid_Opcode PFR_SlotRec_ PFR_Err_Invalid_Glyph_Format pfr_slot_done PFR_BitmapChar ametrics_resolution PFR_Err_Invalid_Glyph_Index PFR_Err_Too_Many_Instruction_Defs pfr_extra_item_load_kerning_pairs axpos PFR_Err_Bbx_Too_Big num_phy_fonts pfr_lookup_bitmap_data PFR_GlyphRec_ aadvance PFR_HeaderRec_ args_format phy_font_section_size astring PFR_CMap PFR_Err_Missing_Module max_x_orus max_blue_values gchar y_pos PFR_Err_Missing_Font_Field PFR_Slot PFR_Err_Locations_Missing PFR_Err_Invalid_Argument phys_size item num_stem_snaps gps_section_size cpair pfr_log_font_count PFR_Err_ENDF_In_Exec_Stream signature pfr_bitwriter_decode_bytes pfr_glyph_line_to num_horz PFR_GlyphRec pfr_load_bitmap_metrics PFR_Err_Invalid_Stream_Seek pfr_slot_load max_strikes counts pfr_log_font_load pfr_slot_load_bitmap PFR_Err_Invalid_Character_Code PFR_FaceRec_ pfr_bitwriter_decode_rle2 PFR_Err_Post_Table_Missing pfr_header_fields aypos pfr_slot_init old_count PFR_Err_Cannot_Open_Resource FT_Service_PfrMetricsRec_ PFR_Err_Invalid_CharMap_Handle PFR_Err_Invalid_Pixel_Size PFR_PhyFont PFR_Err_Invalid_Stream_Handle PFR_PhyFontRec pfr_glyph_load_rec pfr_aux_name_load num_subs pfr_glyph_init PFR_Err_Raster_Uninitialized PFR_Err_Could_Not_Find_Context pfr_glyph_load_compound PFR_Err_Invalid_Library_Handle pfr_bitwriter_decode_rle1 pfr_load_bitmap_bits gps_size bold_thickness aysize log_dir_size PFR_CharRec_ x_control max_chars PFR_Err_Too_Many_Drivers pfr_extra_item_load_font_id t42_get_ps_font_name T42_GlyphSlot real_size T42_Err_DEF_In_Glyf_Bytecode t42_ps_has_glyph_names t42_services T42_Driver_Init T42_Size_Select T42_Err_Nested_DEFS T1_FontInfo T42_Err_Unknown_File_Format T42_Err_Post_Table_Missing T42_Err_Missing_Startchar_Field t42_ps_get_font_private t42_loader_done T42_Err_Invalid_Cache_Handle T42_Err_Unimplemented_Feature T42_Face_Init t42_parse_font_matrix T42_Err_Invalid_Frame_Read T42_Err_Invalid_Glyph_Format T42_Err_Lower_Module_Version T42_Err_Nested_Frame_Access T42_Open_Face T42_Err_Missing_Size_Field T42_Err_Invalid_Version t42_interface T42_Err_Out_Of_Memory t42_service_ps_font_name T42_Err_Cannot_Render_Glyph T42_Err_Missing_Property ttclazz T42_Parser T42_Err_Invalid_Frame_Operation T42_ParserRec t42_service_ps_info T42_Size_Init T42_Load_Status_ T42_Err_Invalid_Stream_Handle T42_Err_Invalid_Handle T42_Err_Name_Table_Missing t42_parse_dict T42_GlyphSlotRec_ ttf_size T42_Err_Invalid_Stream_Skip T42_Err_Missing_Fontboundingbox_Field t42_get_glyph_name status T42_Loader BEFORE_START T42_Size T42_Err_Divide_By_Zero T42_Err_CMap_Table_Missing T42_Err_Hmtx_Table_Missing T42_Err_Ignore T42_Err_Invalid_Vert_Metrics T42_Err_Invalid_CharMap_Handle T42_LoaderRec T42_Err_Invalid_Table unicode_map t42size t42_service_glyph_dict T42_Err_Invalid_Glyph_Index T42_Err_Stack_Underflow ttf_face T42_Err_Raster_Overflow T42_Err_Missing_Module t42_loader_init T42_Loader_ T42_Get_Interface T42_Err_Invalid_Stream_Seek T42_DriverRec_ t42_parse_sfnts T42_Err_Could_Not_Find_Context T42_Err_Invalid_Face_Handle T42_Err_Array_Too_Large T42_Err_No_Unicode_Glyph_Name T42_Err_Unlisted_Object T42_Err_Invalid_Offset T42_Err_Invalid_Post_Table_Format T42_Err_Raster_Negative_Height T42_GlyphSlot_Init T42_Err_Invalid_Reference T42_Err_Invalid_File_Format T42_Err_Execution_Too_Long T42_Err_Table_Missing T42_Err_Invalid_Character_Code T42_Err_Invalid_Horiz_Metrics T42_Err_Invalid_Outline have_literal T42_Err_Debug_OpCode t42face OTHER_TABLES PS_UnicodesRec T42_Err_Missing_Startfont_Field t42_parser_done T42_Err_Invalid_Library_Handle T42_Err_Bbx_Too_Big T42_Err_Invalid_Post_Table T42_Driver t42_ps_get_font_info T42_Err_Missing_Bbx_Field T42_Load_Status T42_Err_Cannot_Open_Resource T42_FaceRec_ T42_GlyphSlot_Done T42_Err_Glyph_Too_Big T42_Err_Too_Many_Drivers T42_Err_Invalid_Stream_Operation T42_Err_Invalid_Pixel_Size T42_Err_Syntax_Error T42_Err_Code_Overflow T42_SizeRec_ t42_load_keyword string_buf t42slot T42_Err_Corrupted_Font_Header t42_is_space T42_Err_Invalid_PPem ttf_data T42_Err_Bad_Argument T42_Err_Invalid_Driver_Handle T42_Err_Too_Many_Caches t42_get_name_index T42_Err_Invalid_Slot_Handle T42_Err_ENDF_In_Exec_Stream ttmodule T42_Err_Raster_Corrupted T42_Err_Ok T42_ParserRec_ T42_Err_Cannot_Open_Stream T42_Err_Invalid_Opcode T42_Err_Too_Few_Arguments T42_Err_Missing_Bitmap t42_parser_init t42_ps_get_font_extra T42_Err_Raster_Uninitialized T42_Err_Corrupted_Font_Glyphs t42_parse_charstrings T42_Err_Invalid_Argument T42_Err_Horiz_Header_Missing T42_Err_Invalid_CodeRange T42_Err_Invalid_Composite T42_Err_Max T42_Err_Too_Many_Extensions n_keywords t42_parse_encoding T42_Face T42_Err_Missing_Encoding_Field T42_Size_Done T42_Driver_Done T42_Err_Locations_Missing T42_Err_Invalid_Stream_Read t42_keywords T42_Face_Done BEFORE_TABLE_DIR T42_Size_Request t42_glyphslot_clear old_string_size T42_GlyphSlot_Load T42_Err_Too_Many_Hints /home/computerfido/Desktop/LemonTest/lemon-freetype/src/type42/type42.c T42_Err_Missing_Chars_Field T42_Err_Stack_Overflow T42_Err_Invalid_CharMap_Format T42_Err_Too_Many_Function_Defs T42_Err_Too_Many_Instruction_Defs T42_Err_Invalid_Size_Handle T42_Err_Missing_Font_Field WinPE_RsrcDirEntryRec WinNE_HeaderRec_ winpe_rsrc_dir_entry_fields fntface bits_offset dir_entry2 dir_entry3 WinMZ_HeaderRec_ WinPE_RsrcDirEntryRec_ root_dir FNT_Face_Done ne_header first_char A_space aheader FNT_Size_Select pitch_and_family size_shift pe32_header WinMZ_HeaderRec bytes_per_row rsrc_virtual_address last_char winne_header_fields WinPE32_HeaderRec_ column new_format FT_Service_WinFntRec FNT_Face_Init winpe32_header_fields WinPE32_SectionRec FT_WinFNT_HeaderRec nominal_point_size face_instance_index fnt_font_done italic B_space fnt_font_load FNT_CMap magic32 winpe32_section_fields winmz_header_fields FT_WinFnt_GetHeaderFunc strike_out fnt_cmap_char_next Found_rsrc_section /home/computerfido/Desktop/LemonTest/lemon-freetype/src/winfonts/winfnt.c x_res lang_dir_offset root_dir_offset characteristics WinPE32_SectionRec_ rname_tab_offset winpe_rsrc_dir_fields WinPE_RsrcDirRec number_of_named_entries winpe_rsrc_data_entry_fields FT_Service_WinFntRec_ time_date_stamp name_dir_offset C_space FT_WinFNT_HeaderRec_ name_dir color_table_offset WinPE32_HeaderRec FNT_Size_Request default_char winfnt_service_rec resource_tab_offset number_of_id_entries avg_width fnt_frame WinPE_RsrcDirRec_ WinPE_RsrcDataEntryRec internal_leading size_of_optional_header FNT_FontRec_ code_page horizontal_resolution pe32_section dir_entry1 type_id winfnt_services device_offset offset_to_data FNT_CMapRec_ mz_header WinNE_HeaderRec fnt_cmap_init WinPE_RsrcDataEntryRec_ FNT_FaceRec_ file_type major_version rsrc_size fnt_cmap_char_index winfnt_get_service external_leading fnt_face_get_dll_font bits_pointer fnt_cmap_class_rec res_offset family_size minor_version winfnt_header_fields fnt_cmap_class pointer_to_raw_data reserved1 fnt_size size_of_raw_data number_of_sections FNT_Load_Glyph data_entry break_char winfnt_get_header FT_WinFNT_Header vertical_resolution lfanew FNT_Font FNT_Face machine underline lang_dir y_res face_name_offset PCF_Err_Horiz_Header_Missing drawDirection pcfcmap FT_Stream_OpenLZW PCF_Err_Invalid_Stream_Read pcf_enc_header PCF_ParseProperty pcf_table_header PCF_ParsePropertyRec BDF_PropertyRec_ PCF_Err_Glyph_Too_Big fontDescent pcf_read_TOC charcodeCol PCF_Err_Invalid_Library_Handle PCF_Face_Done orig_nprops charcodeRow PCF_Err_Unimplemented_Feature PCF_Err_Invalid_Stream_Operation pcf_load_font pcf_service_bdf PCF_Err_Code_Overflow PCF_Enc pcf_cmap_char_index PCF_Err_Missing_Chars_Field PCF_Err_Invalid_CharMap_Format PCF_Err_Invalid_Reference acharset_registry ink_maxbounds PCF_Err_Invalid_Frame_Operation pcfface PCF_Err_Missing_Startchar_Field PCF_Err_Missing_Fontboundingbox_Field PCF_Toc pcf_seek_to_table_type ntables PCF_Err_Invalid_Character_Code PCF_TableRec_ PCF_Err_Ok PCF_Err_Stack_Overflow PCF_CMap pcf_driver_done constantWidth nbytes PCF_Err_Invalid_Slot_Handle PCF_Err_Out_Of_Memory PCF_EncRec_ BDF_PROPERTY_TYPE_ATOM PCF_ParsePropertyRec_ PCF_Err_Invalid_Stream_Skip pcf_metric_header TwoByteSwap FourByteSwap PCF_EncRec PCF_Err_CMap_Table_Missing pcf_cmap_init PCF_Err_Divide_By_Zero PCF_Err_Invalid_Vert_Metrics hasBDFAccelerators PCF_Err_Invalid_Frame_Read sizebitmaps inkInside PCF_Err_Post_Table_Missing PCF_Err_ENDF_In_Exec_Stream isString PCF_Err_Invalid_Version PCF_Err_Invalid_CodeRange PCF_Err_Too_Many_Caches pcf_get_metrics PCF_Size_Request PCF_Err_Invalid_Size_Handle PCF_Err_Syntax_Error PCF_Err_Cannot_Open_Resource PCF_Size_Select pcf_property_msb_header pcf_property_header PCF_Err_Bad_Argument PCF_Err_Invalid_Table pcf_driver_requester PCF_Err_Too_Many_Function_Defs pcf_service_properties pcf_driver_init terminalFont PCF_TocRec_ PCF_Err_Stack_Underflow PCF_Err_Debug_OpCode pcf_find_property PCF_Err_Unlisted_Object PCF_Err_Invalid_Driver_Handle PCF_Err_Missing_Size_Field defaultChar PCF_AccelRec_ PCF_Err_Locations_Missing pcf_cmap_done firstCol PCF_Compressed_MetricRec PCF_Err_Invalid_Outline pcf_accel_header Bail PCF_Err_Name_Table_Missing PCF_Err_DEF_In_Glyf_Bytecode PCF_Err_Too_Many_Instruction_Defs PCF_Err_Nested_Frame_Access PCF_Err_Too_Few_Arguments firstRow PCF_Err_Invalid_Pixel_Size PCF_Err_Missing_Startfont_Field PCF_Face fontAscent PCF_TocRec PCF_Err_Raster_Overflow inkMetrics resolution_y PCF_FaceRec_ error3 PCF_TableRec PCF_Err_No_Unicode_Glyph_Name PCF_Err_Ignore PCF_Err_Missing_Font_Field PCF_Err_Bbx_Too_Big PCF_Err_Raster_Corrupted PCF_Err_Execution_Too_Long PCF_Err_Cannot_Open_Stream PCF_Err_Invalid_Glyph_Index FT_BDF_GetPropertyFunc bitmapSizes PCF_Err_Raster_Negative_Height PCF_Property BitOrderInvert pcf_get_properties defaultCharEncodingOffset acharset_encoding PCF_Err_Table_Missing pcf_toc_header ink_minbounds PCF_Err_Invalid_Glyph_Format PCF_Face_Init PCF_Err_Array_Too_Large pcf_get_encodings pcf_get_accel pcf_compressed_metric_header PCF_MetricRec_ PCF_Err_Missing_Encoding_Field PCF_CMapRec_ PCF_Err_Corrupted_Font_Glyphs PCF_Err_Invalid_Face_Handle PCF_Err_Invalid_Post_Table_Format PCF_Err_Invalid_Stream_Seek BDF_PROPERTY_TYPE_CARDINAL acharcode rightSideBearing PCF_Err_Invalid_PPem prop_name bitmapsFormat PCF_Err_Lower_Module_Version PCF_Err_Missing_Property PCF_Err_Missing_Bbx_Field nencoding PCF_Err_Corrupted_Font_Header have_change aproperty BDF_PropertyType PCF_Compressed_MetricRec_ BDF_PropertyRec pcf_interpret_style PCF_Err_Hmtx_Table_Missing pcf_enc_msb_header BDF_PropertyType_ pcf_get_metric characterWidth BDF_PROPERTY_TYPE_NONE PCF_Err_Invalid_Offset leftSideBearing pcf_cmap_char_next cardinal orig_nmetrics PCF_Glyph_Load FT_BDF_GetCharsetIdFunc PCF_Err_Invalid_Horiz_Metrics resolution_x PCF_Err_Cannot_Render_Glyph attributes pcf_has_table_type pcf_services PCF_Accel lastCol PCF_Err_Invalid_Handle BDF_PROPERTY_TYPE_INTEGER PCF_Err_Max comp_source defaultCharCol /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pcf/pcf.c pcf_get_bitmaps PCF_Err_Invalid_Composite FT_Stream_OpenGzip maxOverlap lastRow PCF_Err_Nested_DEFS PCF_Err_Invalid_Opcode FT_Service_BDFRec_ PCF_Err_Too_Many_Extensions pcf_metric_msb_header PCF_Err_Raster_Uninitialized pcf_accel_msb_header PCF_Err_Invalid_Argument PCF_Table encodingOffset PCF_Err_Invalid_CharMap_Handle PCF_PropertyRec_ PCF_AccelRec pcf_get_charset_id PCF_Err_Unknown_File_Format PCF_Err_Too_Many_Hints PCF_Err_Missing_Bitmap PCF_Err_Could_Not_Find_Context pcf_get_bdf_property PCF_Metric comp_stream defaultCharRow PCF_Err_Invalid_Stream_Handle PCF_Err_Missing_Module constantMetrics pcf_cmap_class noOverlap PCF_Err_Invalid_File_Format PCF_MetricRec PCF_Err_Too_Many_Drivers FT_Service_BDFRec PCF_Err_Invalid_Post_Table PCF_Err_Invalid_Cache_Handle pcf_property_set pcf_property_get orig_nbitmaps compr BDF_Err_Missing_Fontboundingbox_Field _bdf_readstream bdf_property_t bdf_driver_requester _bdf_list_shift BDF_Err_Table_Missing BDF_Err_Too_Many_Instruction_Defs bdf_options_t_ BDF_CMap _bdf_atol BDF_Err_Missing_Encoding_Field _bdf_atos BDF_Err_Invalid_Offset bdf_free_font BDF_Err_Raster_Uninitialized buf_size bdf_load_font BDF_Err_Invalid_Driver_Handle num_encodings /home/computerfido/Desktop/LemonTest/lemon-freetype/src/bdf/bdf.c BDF_Err_Raster_Overflow keep_comments client_data BDF_Err_Raster_Negative_Height BDF_Err_Corrupted_Font_Header bdf_bbx_t_ _bdf_parse_glyphs BDF_Err_Bad_Argument glyphs_size maxas BDF_Err_Horiz_Header_Missing BDF_Err_No_Unicode_Glyph_Name BDF_Err_Invalid_Face_Handle BDF_Err_Invalid_Post_Table BDF_Err_Invalid_Stream_Operation vlen BDF_Err_Locations_Missing props_used BDF_Err_Invalid_Outline BDF_Err_Invalid_Table BDF_Err_Too_Many_Drivers nibble_mask _bdf_list_split bdf_cmap_init BDF_Err_Invalid_Stream_Skip separators nuser_props extmemory x_offset BDF_Err_Invalid_Stream_Read bdf_glyph_t_ BDF_Err_Invalid_CharMap_Format _bdf_set_default_spacing BDF_Glyph_Load BDF_Err_Nested_DEFS BDF_encoding_el _bdf_add_comment _num_bdf_properties call_data alen BDF_Err_Array_Too_Large BDF_Err_Invalid_Handle maxds bdf_get_property nbuf BDF_Err_Invalid_Version BDF_Err_Invalid_Post_Table_Format BDF_Err_Invalid_CodeRange correct_metrics BDF_Err_Divide_By_Zero BDF_Size_Request bdf_cmap_char_next _bdf_opts oldsize _bdf_atous bigsize BDF_Err_Ok BDF_Err_Nested_Frame_Access BDF_Err_Code_Overflow _bdf_list_t_ BDF_Err_Corrupted_Font_Glyphs bdf_cmap_class default_glyph bdf_service_bdf _bdf_parse_start Missing_Encoding monowidth BDF_Err_Max BDF_Err_Could_Not_Find_Context BDF_Err_Missing_Chars_Field BDF_Err_Unlisted_Object bdf_font_t keep_unencoded BDF_Err_Invalid_PPem BDF_Err_Bbx_Too_Big BDF_Err_Glyph_Too_Big BDF_Err_Too_Many_Extensions BDF_FaceRec_ BDF_Err_Cannot_Open_Resource BDF_Err_Too_Many_Hints ddigits bdf_property_t_ comments_len _bdf_is_atom BDF_Err_Invalid_File_Format propid BDF_Err_Unknown_File_Format font_ascent BDF_Err_Invalid_Frame_Read bdf_get_charset_id BDF_Err_Invalid_Vert_Metrics bdf_glyph_t BDF_Err_Invalid_Cache_Handle BDF_Err_Invalid_Composite BDF_Err_Invalid_Argument BDF_Err_Invalid_Size_Handle BDF_Err_CMap_Table_Missing props_size proptbl minlb font_descent slen _bdf_list_ensure _bdf_list_done BDF_Err_Hmtx_Table_Missing linelen BDF_Size_Select BDF_CMapRec_ BDF_Err_Too_Many_Function_Defs BDF_Err_Missing_Bbx_Field BDF_Err_Missing_Size_Field lineno _bdf_add_property BDF_Face_Init seps _bdf_list_t bdf_interpret_style BDF_Err_Invalid_Character_Code BDF_Err_Invalid_Stream_Handle BDF_Err_Name_Table_Missing hdigits BDF_Err_Cannot_Open_Stream BDF_Err_DEF_In_Glyf_Bytecode BDF_Err_Stack_Overflow BDF_Err_Invalid_Pixel_Size BDF_Face_Done BDF_Err_Invalid_CharMap_Handle by_encoding BDF_Err_Stack_Underflow BDF_Face _bdf_parse_properties BDF_Err_Invalid_Frame_Operation maxrb BDF_Err_Missing_Font_Field _bdf_atoul BDF_Err_Invalid_Library_Handle final_empty BDF_Err_Invalid_Opcode BDF_Err_Invalid_Glyph_Index _bdf_parse_t BDF_Err_Invalid_Slot_Handle BDF_Err_Missing_Module BDF_Err_ENDF_In_Exec_Stream BDF_Err_Too_Few_Arguments BDF_Err_Too_Many_Caches bdf_services BDF_Err_Out_Of_Memory BDF_Err_Raster_Corrupted BDF_Err_Missing_Bitmap bdf_get_bdf_property bdf_options_t swidth BDF_Err_Unimplemented_Feature BDF_Err_Invalid_Glyph_Format bdf_bbx_t BDF_Err_Missing_Property bdfface BDF_Err_Post_Table_Missing builtin bdf_create_property FT_HashRec BDF_Err_Invalid_Horiz_Metrics sprintf unencoded_used _bdf_list_join BDF_Err_Debug_OpCode BDF_Err_Invalid_Stream_Seek en_table BDF_Err_Execution_Too_Long bdf_font_t_ _bdf_parse_end BDF_Err_Missing_Startfont_Field mask_index glyph_enc BDF_Err_Syntax_Error nibbles BDF_Err_Lower_Module_Version glyphs_used dwidth font_spacing bitmap_size unencoded_size bdfcmap BDF_Err_Missing_Startchar_Field to_skip _bdf_line_func_t bdf_cmap_char_index BDF_Err_Ignore maxlb _bdf_parse_t_ BDF_Err_Cannot_Render_Glyph BDF_encoding_el_ bdffont BDF_Err_Invalid_Reference bdf_get_font_property avail bdf_cmap_done newsize rbearing _bdf_list_init SFNT_Err_Invalid_Library_Handle lastVarSel SFNT_Err_Debug_OpCode tt_face_load_kern NoCpal FT_Bitmap_Done tt_cmap14_char_var_index tt_cmap6_class_rec sfnt_get_name_id sfnt_interface NoBitmap table1 table2 sfnt_header woff_offset min_after_bl SFNT_Err_Invalid_Argument cur_gindex type_offset char_type SFNT_Err_Invalid_Slot_Handle TT_SBitDecoderRec_ strike_idx instance_values TT_CMap srcSlot tt_cmap12_validate instance_offset char_lo TT_CMapRec_ SFNT_Err_Invalid_Reference tt_face_palette_set base_glyph_offset tt_cmap8_validate numVar tt_face_free_cpal last_end keys count2 SFNT_Err_Bbx_Too_Big get_win_string SFNT_Err_Too_Many_Function_Defs SFNT_Err_Unimplemented_Feature num_segs metaLength SFNT_Err_Invalid_Handle tt_face_load_head num_pairs has_head SFNT_Err_Missing_Encoding_Field tt_cmap8_char_next tt_cmap0_class_rec max_before_bl SFNT_Err_Invalid_CharMap_Handle old_pair TT_Name_ConvertFunc tt_face_colr_blend_layer post_len tt_get_cmap_info tt_cmap14_class_rec tt_cmap10_get_info tt_face_free_name wval SFNT_Err_Invalid_Post_Table storage_start load_post_names maxProfile tt_cmap2_get_info cur_group tt_cmap14_get_nondef_chars sfnt_find_encoding tt_cmap2_char_next bitmap_allocated num_components variantCode SFNT_Err_Nested_DEFS tt_face_load_sbit TT_CMap_ClassRec_ tt_face_load_strike_metrics tt_cmap14_char_index SFNT_Err_Missing_Startchar_Field SFNT_Err_Invalid_Stream_Read tt_get_glyph_name entrySelector TT_CMap_ClassRec SFNT_Err_Glyph_Too_Big tt_face_get_colr_layer originOffsetX originOffsetY subfamily_name tt_face_load_hmtx SFNT_Err_Invalid_Outline NoColr SFNT_Err_Ok TT_CMap4 SFNT_Err_Stack_Overflow get_apple_string_error found_unicode tt_cmap14_init SFNT_Err_Post_Table_Missing SFNT_Err_Code_Overflow woff_header_fields property_len TT_CMap12 max_gid recurse_depth tt_face_get_kerning ignore_typographic_family post_limit SFNT_Err_Missing_Chars_Field sfnt_get_var_ps_name privOffset TT_CMapRec SFNT_Err_Corrupted_Font_Header image_format sfnt_service_sfnt_table TT_CMap13 TT_CMap14 TT_CMap4Rec_ PSname tt_cmap10_char_next tt_cmap12_init sfnt_is_alphanumeric pwrite report_invalid_characters tt_cmap12_next glyph_id graphicType charCode tt_face_load_font_dir entry_label_offset num_groups tt_name_ascii_from_utf16 sfnt_stream_close get_sfnt_table tt_cmap14_def_char_count SFNT_Err_Stack_Underflow rangeShift totalSfntSize num_base_glyphs SFNT_Err_Corrupted_Font_Glyphs FT_Bitmap_Init sfnt_table_info TEncoding_ SFNT_Err_Missing_Module psnames_error sfnt_init_face NoData TT_CMap13Rec_ SFNT_Err_Invalid_Table tt_face_load_gasp tt_cmap_unicode_char_next load_format_25 TT_SBitDecoder_LoadFunc found_win SFNT_Err_Invalid_Frame_Operation duplicate tt_cmap14_validate tt_sbit_decoder_load_bitmap SFNT_Err_Cannot_Open_Resource prev_end sfnt_services varSel default_values TT_SBitDecoderRec y_min image_size FoundStrike aprop NextTable cmap4 tt_cmap14_char_map_nondef_binary SFNT_Err_Invalid_Stream_Seek eblc_base tt_face_free_ps_names tt_cmap2_class_rec check_table_dir tt_sbit_decoder_init SFNT_Err_CMap_Table_Missing SFNT_Err_Invalid_Offset tt_face_get_metrics new_map tt_cmap4_validate Next_Segment byte_size starts SFNT_Err_Invalid_Stream_Skip default_value_offset glyph_ids fixed2float tt_cmap0_validate last_start FT_Gzip_Uncompress tt_cmap0_get_info tt_cmap13_char_index tt_cmap4_char_map_binary SFNT_Err_Invalid_Driver_Handle offset1 offset2 cur_end SFNT_Err_Raster_Negative_Height range_index found_apple_roman sfnt_ps_map tt_cmap13_char_map_binary valid_entries SFNT_Err_Raster_Corrupted tt_cmap13_validate metaOffset tt_face_load_sbix_image WOFF_HeaderRec TEncoding sfnt_offset SFNT_Err_Invalid_Character_Code tt_face_free_colr nblocks bit_depth tt_cmap14_char_next has_CBDT found_apple post_fields SFNT_Err_Nested_Frame_Access tt_cmap4_class_rec image_offset ptable_offset SFNT_Err_ENDF_In_Exec_Stream /home/computerfido/Desktop/LemonTest/lemon-freetype/src/sfnt/sfnt.c tt_face_load_hhea privLength has_unicode tt_face_get_ps_name tt_cmap2_char_index tt_cmap14_variant_chars tt_face_load_cmap find_base_glyph_record cur_start tt_face_goto_table p_next SFNT_Err_Horiz_Header_Missing nuni cur_charcode tt_cmap13_class_rec SFNT_Err_Missing_Fontboundingbox_Field SFNT_Err_Cannot_Render_Glyph ptable_size SFNT_Err_Table_Missing avgwidth first_code tt_cmap10_char_index tt_cmap12_get_info tt_face_load_maxp sfnt_open_font tt_cmap14_char_map_def_binary ttcmap numMappings maxp_fields metrics_loaded has_CBLC base_glyph_begin SFNT_HeaderRec convert validator tt_sbit_decoder_alloc_bitmap tt_module tt_cmap_unicode_char_index TT_Validator instance_size ignore_typographic_subfamily TT_NameTable BaseGlyphRecord_ woff tt_cmap12_class_rec is_apple_sbit char_type_func table_dir_entry_fields is_apple_sbix tt_cmap12_char_next TT_TableRec SFNT_Err_Ignore SFNT_Err_Array_Too_Large tt_encodings ppem_ tt_face_load_any tt_cmap6_char_index tt_face_load_bhed SFNT_Err_Locations_Missing code_count tt_cmap0_char_next tt_cmap4_get_info get_win_string_error tt_cmap_unicode_init tt_sbit_decoder_load_compound tt_cmap14_get_def_chars InvalidTable found_apple_english sfnt_get_ps_name FoundRange tt_cmap_unicode_done BadTable sfnt_is_postscript TT_CMap_ValidateFunc SFNT_Err_Invalid_Glyph_Index SFNT_Err_Invalid_Stream_Operation tt_cmap4_set_range woff_open_font tt_cmap12_char_index tt_name_ascii_from_other Cpal_ SFNT_Header bit_height get_apple_string tt_face_load_colr SFNT_Err_Bad_Argument SFNT_Err_Invalid_Glyph_Format tt_cmap4_char_next is_english SFNT_Err_Invalid_Opcode start_id SFNT_Err_Invalid_CodeRange sfnt_get_interface name_table_fields pclazz bsize_idx SFNT_Err_Execution_Too_Long Next_SubHeader sfnt_load_face key0 tt_sbit_decoder_load_metrics duni offset_table_fields SFNT_Err_Invalid_Cache_Handle upem sfnt_service_bdf old_tag tt_cmap4_char_map_linear retry SFNT_Err_Divide_By_Zero tt_cmap8_char_index strike_index_array pcharcode has_outline murmur_hash_3_128 entry_selector searchRange SFNT_Err_Too_Few_Arguments tt_cmap13_get_info SFNT_Err_Too_Many_Instruction_Defs nbits tt_cmap12_char_map_binary tt_face_load_bdf_props flavor minorVersion tt_sbit_decoder_done sfnt_get_glyph_name pclt_fields SFNT_Err_Invalid_Face_Handle maxp_fields_extra tt_cmap14_ensure tt_cmap4_init WOFF_TableRec_ nondefOff SFNT_Err_Raster_Uninitialized tt_cmap10_class_rec tt_cmap6_validate tt_sbit_decoder_load_image table_pos SFNT_Err_Invalid_Size_Handle rval tt_cmap4_next SFNT_Err_Missing_Size_Field hexdigits tt_cmap14_char_variants tt_cmap6_char_next SFNT_Err_Out_Of_Memory bit_width Colr_ dstSlot lastUni ttc_header_fields tt_sbit_decoder_load_bit_aligned tt_cmap0_char_index tt_face_build_cmaps search_range tt_face_load_cpal frac_part tt_face_load_generic_header SFNT_Err_DEF_In_Glyf_Bytecode tt_cmap8_get_info bit_size FT_Bitmap_Convert SFNT_Err_Invalid_Pixel_Size range_shift SFNT_Err_Missing_Font_Field strike_offset SFNT_Err_Syntax_Error tt_cmap14_char_var_isdefault load_format_20 num_segs2 SFNT_Err_Max storage_limit next_end tt_cmap8_class_rec SFNT_Err_Invalid_Stream_Handle lastBase abearing langTag_record_fields SFNT_Err_Invalid_File_Format tt_cmap_unicode_class_rec SFNT_Err_Unknown_File_Format check_length TT_Post_Names WOFF_Table SFNT_Err_Name_Table_Missing image_start tt_face_load_name os2_fields_extra5 line_bits os2_fields image_end SFNT_HeaderRec_ gaspranges TT_SBit_Metrics name_record_fields compare_offsets name_strings SFNT_Err_Raster_Overflow SFNT_Err_Could_Not_Find_Context SFNT_Err_Too_Many_Caches SFNT_Err_Invalid_PPem has_meta tt_face_lookup_table SFNT_Err_Invalid_Composite cur_values layer_offset sfnt_get_name_index astrike_index SFNT_Err_Too_Many_Drivers colors_offset tt_cmap14_get_info next_start tt_face_done_kern tt_cmap6_get_info metaOrigLength metrics_header_fields TT_ValidatorRec tt_face_free_sbit SFNT_Err_Hmtx_Table_Missing tt_sbit_decoder_load_byte_aligned cur_pair SFNT_Err_Missing_Property max_results os2_fields_extra1 os2_fields_extra2 SFNT_Err_No_Unicode_Glyph_Name tt_cmap_classes tt_face_set_sbit_strike tt_service_get_cmap_info SFNT_Err_Missing_Startfont_Field SFNT_Err_Unlisted_Object output_len sfnt_service_ps_name array_start is32 SFNT_Err_Cannot_Open_Stream tt_face_get_name CompLength TT_Post_20 TT_Post_25 TT_CMap14Rec_ cmap12 cmap13 cmap14 dcnt tt_cmap14_find_variant FT_Service_SFNT_TableRec tt_cmap2_validate SFNT_Err_Too_Many_Extensions TT_ValidatorRec_ strike_index_count tt_face_find_bdf_prop sfnt_get_charset_id num_colors SFNT_Err_Invalid_Version sfnt_service_glyph_dict BaseGlyphRecord setjmp offset_table index_format SFNT_Err_Invalid_Frame_Read tt_cmap2_get_subheader WOFF_HeaderRec_ SFNT_Err_Lower_Module_Version sfnt_done_face tt_face_load_pclt num_base_glyph color_indices nameid SFNT_Err_Missing_Bbx_Field construct_instance_name OrigOffset fvar_len TT_CMap12Rec_ int_part SFNT_Err_Invalid_Post_Table_Format tt_cmap14_done old_p fmix32 tt_face_free_bdf_props defp tt_cmap_init tt_cmap14_variants tt_face_load_os2 tt_face_load_sbit_image num_selectors eblc_limit p_start FT_ValidatorRec first_layer_index tt_cmap13_char_next tt_cmap10_validate SFNT_Err_Invalid_Horiz_Metrics SFNT_Err_Too_Many_Hints char_hi tt_cmap13_next tt_face_load_post SFNT_Err_Missing_Bitmap TT_CMap_Class tt_cmap13_init has_sing tt_cmap4_char_index TT_BDF num_cmaps num_results TT_SBitDecoder SFNT_Err_Invalid_CharMap_Format SFNT_Err_Invalid_Vert_Metrics af_warper_compute af_latn_titl_style_class AF_BLUE_STRING_LATIN_SUBS_SMALL_DESCENDER af_telu_dflt_style_class AF_COVERAGE_ORDINALS style_metrics_size AF_BLUE_STRING_MYANMAR_TOP shaper_buf AF_CJKMetrics af_iup_shift AF_BLUE_STRING_TAI_VIET_BOTTOM AF_BLUE_STRING_MAX AF_AxisHintsRec_ AF_ScriptClass axhints af_lao_script_class height_threshold af_latn_c2cp_style_class AF_BLUE_STRINGSET_TFNG p_last AF_Err_Raster_Corrupted af_none_script_class AF_STYLE_LATB_DFLT af_grek_sups_style_class pp1x_uh af_face_globals_new AF_BLUE_STRING_GEORGIAN_MKHEDRULI_ASCENDER AF_Err_Raster_Uninitialized has_last_stem af_cjk_writing_system_class AF_BLUE_STRING_ETHIOPIC_TOP is_top_right_blue AF_Err_Ok af_osge_dflt_style_class AF_BLUE_STRING_TAMIL_BOTTOM AF_SCRIPT_KALI AF_STYLE_LATN_C2CP af_kali_uniranges AF_Err_Corrupted_Font_Glyphs AF_BLUE_STRING_LAO_BOTTOM AF_WritingSystemClassRec_ af_limb_script_class af_gujr_dflt_style_class AF_SCRIPT_SAUR AF_Err_Invalid_Reference af_dsrt_uniranges af_cari_uniranges AF_STYLE_VAII_DFLT AF_Err_Missing_Fontboundingbox_Field af_thai_uniranges AF_BLUE_STRING_GLAGOLITIC_SMALL_BOTTOM af_nkoo_script_class AF_BLUE_STRING_MYANMAR_DESCENDER prev_min_pos AF_Err_Unknown_File_Format AF_Err_Raster_Negative_Height af_axis_hints_new_segment AF_BLUE_STRING_GURMUKHI_BASE AF_BLUE_STRING_ARABIC_TOP af_cjk_hints_detect_features AF_BLUE_STRING_LAO_TOP AF_BLUE_STRING_SINHALA_BOTTOM af_nkoo_dflt_style_class AF_STYLE_SUND_DFLT AF_COVERAGE_PETITE_CAPITALS_FROM_CAPITALS AF_BLUE_STRING_ADLAM_SMALL_BOTTOM AF_BLUE_STRING_GUJARATI_BOTTOM AF_WRITING_SYSTEM_LATIN Is_Weak_Point points_limit prev_min_coord AF_AxisHints af_goth_script_class af_gujr_uniranges last_touched af_guru_nonbase_uniranges AF_BLUE_STRING_KHMER_SYMBOLS_WANING_BOTTOM AF_BLUE_STRINGSET_SUND AF_BLUE_STRING_LATIN_SUBS_CAPITAL_BOTTOM af_beng_uniranges af_cjk_hints_link_segments af_avst_dflt_style_class org_len AF_Warper af_sund_dflt_style_class af_cjk_hints_init af_bamu_uniranges af_cjk_metrics_scale_dim seg_delta AF_BLUE_STRING_OLD_TURKIC_TOP AF_BLUE_STRINGSET_NONE AF_COVERAGE_SMALL_CAPITALS_FROM_CAPITALS AF_Err_Invalid_Character_Code AF_Err_Invalid_Size_Handle af_ethi_uniranges AF_BLUE_STRINGSET_THAI AF_STYLE_ETHI_DFLT AF_BLUE_STRINGSET_ARMN AF_COVERAGE_PETITE_CAPITALS AF_STYLE_ORKH_DFLT AF_SCRIPT_OSMA AF_BLUE_STRINGSET_OLCK AF_Err_Raster_Overflow style_metrics_scale style_metrics dist_score FT_Prop_GlyphToScriptMap AF_BLUE_STRING_SHAVIAN_SMALL_TOP af_loader_init af_latn_sups_style_class inverse af_avst_nonbase_uniranges af_geok_uniranges af_deva_dflt_style_class af_mong_uniranges af_beng_nonbase_uniranges script_uni_nonbase_ranges af_cyrl_pcap_style_class af_blue_stringsets AF_Err_Bbx_Too_Big af_cans_dflt_style_class AF_SCRIPT_BENG AF_StyleMetricsRec af_osge_nonbase_uniranges AF_STYLE_CYRL_SUBS AF_BLUE_STRINGSET_BUHD af_glyph_hints_done AF_CJKAxisRec_ AF_SCRIPT_ETHI af_tfng_dflt_style_class AF_BLUE_STRING_GEORGIAN_NUSKHURI_DESCENDER af_shaw_uniranges best_distort AF_STYLE_LATN_SUBS AF_Dimension_ af_orkh_nonbase_uniranges AF_BLUE_STRING_DEVANAGARI_HEAD AF_Err_Invalid_Post_Table_Format xx1max AF_BLUE_STRINGSET_ETHI AF_BLUE_STRING_MONGOLIAN_TOP_BASE AF_WRITING_SYSTEM_INDIC AF_Err_Invalid_Driver_Handle AF_Err_Invalid_CodeRange AF_Err_Invalid_Composite af_mymr_uniranges af_latn_script_class af_grek_c2sc_style_class AF_Module fpos is_round AF_BLUE_STRING_DEVANAGARI_BASE AF_BLUE_STRING_KAYAH_LI_TOP AF_SCRIPT_GURU AF_COVERAGE_SCIENTIFIC_INFERIORS AF_STYLE_CHER_DFLT AF_Err_Nested_Frame_Access AF_BLUE_STRING_LATIN_SUPS_CAPITAL_BOTTOM AF_STYLE_CYRL_SINF prev_max_coord af_warper_compute_line_best d_off1 darken_by_font_units_x AF_LatinAxisRec AF_BLUE_STRING_COPTIC_SMALL_TOP AF_STYLE_LATN_SINF old_rsb best_round af_saur_nonbase_uniranges af_cyrl_script_class AF_StyleClassRec AF_Err_Invalid_Table AF_BLUE_STRING_GEORGIAN_MKHEDRULI_TOP AF_WRITING_SYSTEM_DUMMY AF_SCRIPT_KNDA scale_down_matrix AF_SCRIPT_CAKM AF_BLUE_STRING_OSAGE_CAPITAL_DESCENDER num_segments af_avst_uniranges style_metrics_done edge_distance_threshold warper af_cari_nonbase_uniranges af_orkh_script_class best_score trans_delta AF_WritingSystem_ x2max idx_max AF_CJKMetricsRec AF_BLUE_STRING_CYPRIOT_TOP af_cjk_hints_compute_segments AF_ModuleRec_ AF_BLUE_STRING_TAI_VIET_TOP af_limb_nonbase_uniranges AF_ScriptClassRec_ af_orkh_dflt_style_class AF_BLUE_STRING_NKO_SMALL_TOP af_hint_normal_stem AF_Err_Too_Many_Extensions AF_LatinMetricsRec_ AF_Err_Missing_Startchar_Field AF_STYLE_NKOO_DFLT AF_DIR_DOWN prev_min_on_coord AF_BLUE_STRING_GURMUKHI_DIGIT_TOP af_tfng_nonbase_uniranges AF_LatinMetricsRec af_glag_uniranges af_buhd_script_class oldmap af_style_classes af_cans_script_class scaler af_grek_sinf_style_class reference stdHW AF_BLUE_STRING_ARMENIAN_SMALL_ASCENDER af_glyph_hints_rescale af_none_dflt_style_class AF_BLUE_STRINGSET_GLAG max_segments AF_BLUE_STRING_KANNADA_BOTTOM af_knda_uniranges AF_SCRIPT_CANS AF_STYLE_SAUR_DFLT AF_Style AF_COVERAGE_DEFAULT AF_SCRIPT_SYLO af_blue_strings AF_STYLE_GEOK_DFLT AF_Err_Invalid_Frame_Operation af_armn_dflt_style_class AF_BLUE_STRING_MALAYALAM_BOTTOM AF_BLUE_STRINGSET_COPT AF_Err_Invalid_Version AF_Err_Missing_Font_Field AF_BLUE_STRINGSET_GUJR curr af_face_globals_is_digit AF_Err_Corrupted_Font_Header best_contour_last next_u af_geor_nonbase_uniranges AF_BLUE_STRING_MALAYALAM_TOP AF_STYLE_MAX AF_BLUE_STRING_CHEROKEE_SMALL_DESCENDER AF_Err_Invalid_Outline AF_LatinBlueRec AF_STYLE_CAKM_DFLT extra_light af_vaii_nonbase_uniranges af_bamu_dflt_style_class AF_Err_Missing_Property AF_Err_Too_Many_Drivers af_dsrt_script_class af_cjk_metrics_init_blues af_indic_get_standard_widths af_property_get FT_Prop_GlyphToScriptMap_ best_x af_latn_subs_style_class af_cher_uniranges af_osge_script_class AF_BLUE_STRINGSET_KALI AF_LoaderRec af_cjk_get_standard_widths AF_LatinAxis AF_BLUE_STRING_LAO_DESCENDER AF_STYLE_GREK_C2CP AF_BLUE_STRING_LATIN_SUPS_SMALL best_on_point_last af_geok_nonbase_uniranges AF_BLUE_STRINGSET_SAUR Try_x3 Try_x4 AF_STYLE_GURU_DFLT is_serif AF_Width AF_Script_UniRange AF_WarpScore AF_LatinBlueRec_ blue_stringset AF_BLUE_STRING_GEORGIAN_ASOMTAVRULI_TOP prev_max_pos AF_BLUE_STRING_GUJARATI_TOP af_deva_nonbase_uniranges AF_BLUE_STRING_SINHALA_TOP FT_Prop_IncreaseXHeight af_autofitter_init AF_SCRIPT_LAO AF_BLUE_STRING_VAI_BOTTOM prev_segment af_lisu_dflt_style_class AF_BLUE_STRING_LATIN_SUBS_SMALL af_lisu_script_class neutral2 AF_SCRIPT_CARI AF_BLUE_STRING_GURMUKHI_HEAD AF_SCRIPT_MLYM af_loader_reset af_loader_load_glyph af_cans_nonbase_uniranges near_limit2 AF_AxisHintsRec af_hani_dflt_style_class AF_Err_Invalid_Frame_Read latin af_hani_nonbase_uniranges AF_CJKBlueRec_ AF_Err_Too_Many_Instruction_Defs AF_STYLE_TAML_DFLT AF_BLUE_STRING_GEORGIAN_ASOMTAVRULI_BOTTOM AF_BLUE_STRING_LATIN_SMALL_BOTTOM AF_COVERAGE_SUBSCRIPT org_delta AF_BLUE_STRING_ARMENIAN_SMALL_DESCENDER af_cyrl_sups_style_class af_mymr_dflt_style_class AF_BLUE_STRING_DESERET_SMALL_TOP AF_SCRIPT_VAII AF_STYLE_GUJR_DFLT af_latp_script_class af_shaper_get_elem AF_BLUE_STRING_KAYAH_LI_DESCENDER af_hebr_script_class AF_WritingSystem_DoneMetricsFunc AF_BLUE_STRING_KAYAH_LI_LARGE_DESCENDER AF_BLUE_STRING_GUJARATI_ASCENDER af_sinh_uniranges AF_BLUE_STRING_CARIAN_BOTTOM AF_Err_Divide_By_Zero af_sund_uniranges AF_Err_Stack_Underflow AF_Direction_ AF_LatinAxisRec_ x2min af_latb_nonbase_uniranges idx_min af_grek_dflt_style_class AF_STYLE_MONG_DFLT AF_SCRIPT_LIMB AF_STYLE_TELU_DFLT AF_BLUE_STRING_ETHIOPIC_BOTTOM af_latn_sinf_style_class AF_CJKAxis scaler_flags af_vaii_script_class first_v near_limit blue_sorted af_latn_smcp_style_class AF_STYLE_CYRL_C2CP AF_BLUE_STRING_KHMER_TOP af_latin_snap_width AF_STYLE_SYLO_DFLT prev_v af_hebr_uniranges af_tibt_nonbase_uniranges started AF_STYLE_TIBT_DFLT af_tavt_script_class AF_ScalerRec AF_Err_Invalid_Stream_Read af_buhd_nonbase_uniranges af_face_globals_free AF_BLUE_STRING_SHAVIAN_BOTTOM AF_BLUE_STRING_GREEK_SMALL_DESCENDER AF_Err_Missing_Size_Field af_blue_1_2 AF_BLUE_STRINGSET_BENG AF_BLUE_STRING_SUNDANESE_BOTTOM AF_DIMENSION_VERT script_uni_ranges af_osma_dflt_style_class best_dist0 af_buhd_uniranges af_none_nonbase_uniranges AF_BLUE_STRING_BENGALI_TOP af_latin_hint_edges AF_BLUE_STRINGSET_CAKM AF_SCRIPT_GLAG org_scale AF_STYLE_GREK_SUBS AF_SCRIPT_MYMR warping af_latin_hints_compute_blue_edges af_arab_uniranges af_indic_writing_system_class touch_flag AF_STYLE_CYRL_SUPS stem_flags af_limb_uniranges AF_SCRIPT_MONG af_dsrt_dflt_style_class af_sund_script_class AF_Point /home/computerfido/Desktop/LemonTest/lemon-freetype/src/autofit/autofit.c af_glyph_hints_init AF_BLUE_STRING_KAYAH_LI_ASCENDER AF_SCRIPT_TELU best_blue dist_threshold AF_BLUE_STRING_THAI_TOP AF_STYLE_CYRL_SMCP asegment AF_BLUE_STRING_BUHID_SMALL AF_BLUE_STRING_MYANMAR_ASCENDER AF_BLUE_STRING_GURMUKHI_TOP AF_STYLE_CARI_DFLT AF_BLUE_STRING_BENGALI_HEAD stem_width_per_1000 cur_pos1 cur_pos2 AF_STYLE_LATN_SMCP skipped af_latin_sort_blue increase_x_height edge1 edge2 ft_module AF_SCRIPT_MAX AF_STYLE_MLYM_DFLT edge3 af_armn_uniranges FT_AutoHinter_InterfaceRec AF_STYLE_GREK_SINF AF_Err_Invalid_Face_Handle af_autofitter_load_glyph af_cher_nonbase_uniranges AF_BLUE_STRINGSET_KNDA AF_BLUE_STRING_BENGALI_BASE AF_BLUE_STRING_CYPRIOT_SMALL af_glyph_hints_reload prev_max_on_coord AF_BLUE_STRING_AVESTAN_BOTTOM best_scale stdVW AF_BLUE_STRING_GEORGIAN_NUSKHURI_BOTTOM AF_BLUE_STRING_HEBREW_DESCENDER AF_SCRIPT_AVST AF_Err_Lower_Module_Version AF_STYLE_GREK_SUPS AF_BLUE_STRING_BUHID_TOP AF_BLUE_STRINGSET_LAO wmin AF_Err_CMap_Table_Missing af_cyrl_ordn_style_class af_mlym_script_class Hint_Metrics af_loader_compute_darkening AF_Err_Invalid_Stream_Operation AF_LoaderRec_ af_latin_align_linked_edge AF_BLUE_STRING_LAO_LARGE_ASCENDER af_saur_script_class af_guru_uniranges AF_SCRIPT_TAML af_face_globals_get_metrics af_dummy_writing_system_class af_saur_uniranges AF_SCRIPT_SHAW af_khms_uniranges af_cans_uniranges AF_BLUE_STRING_KHMER_DESCENDER old_advance AF_STYLE_GREK_PCAP AF_Err_Name_Table_Missing AF_STYLE_OSMA_DFLT AF_BLUE_STRING_MYANMAR_BOTTOM best_delta style_metrics_init af_tfng_script_class af_vaii_dflt_style_class af_indic_hints_apply af_lao_nonbase_uniranges AF_STYLE_GREK_SMCP AF_STYLE_GREK_ORDN af_property_set AF_STYLE_COPT_DFLT af_taml_uniranges AF_BLUE_STRING_TELUGU_TOP AF_BLUE_STRINGSET_BAMU em_ratio af_cjk_metrics_check_digits AF_FaceGlobalsRec_ AF_SCRIPT_LISU af_goth_uniranges af_cher_script_class best_on_point_first AF_BLUE_STRING_GEORGIAN_NUSKHURI_ASCENDER AF_Err_Too_Many_Hints AF_BLUE_STRING_COPTIC_CAPITAL_TOP af_lisu_nonbase_uniranges size_internal af_grek_ordn_style_class AF_BLUE_STRING_KAYAH_LI_BOTTOM Use_y4 af_cjk_align_serif_edge AF_Err_Invalid_Vert_Metrics AF_BLUE_STRING_CYRILLIC_CAPITAL_BOTTOM af_blue_2_1 af_blue_2_2 AF_BLUE_STRINGSET_CANS af_ethi_script_class AF_BLUE_STRING_SHAVIAN_TOP AF_ScalerRec_ FT_Prop_IncreaseXHeight_ AF_Err_Invalid_Argument af_nkoo_nonbase_uniranges AF_WarperRec_ af_latb_script_class xx1min af_shaper_buf_destroy AF_COVERAGE_TITLING af_thai_dflt_style_class af_osma_nonbase_uniranges AF_BLUE_STRING_OSAGE_SMALL_ASCENDER AF_STYLE_ORYA_DFLT AF_BLUE_STRING_ARMENIAN_CAPITAL_BOTTOM best_segment_last dist2 af_sinh_nonbase_uniranges d_off af_beng_script_class AF_BLUE_STRING_CANADIAN_SYLLABICS_SUPS_TOP contour_limit style_hints_init AF_STYLE_LATN_SUPS new_scale AF_SegmentRec AF_BLUE_STRINGSET_GURU AF_StyleClassRec_ af_cyrl_smcp_style_class af_olck_uniranges af_cakm_dflt_style_class is_under_ref AF_Err_Nested_DEFS AF_STYLE_CPRT_DFLT AF_BLUE_STRING_CHEROKEE_SMALL_ASCENDER af_thai_script_class AF_WritingSystem_ApplyHintsFunc af_grek_subs_style_class AF_CJKMetricsRec_ AF_Err_Invalid_CharMap_Handle af_axis_hints_new_edge AF_BLUE_STRING_LATIN_SMALL_F_TOP AF_BLUE_STRING_OLD_TURKIC_BOTTOM af_tavt_uniranges AF_BLUE_STRING_CANADIAN_SYLLABICS_SMALL_TOP AF_Err_Hmtx_Table_Missing anedge num_rounds af_cjk_hint_edges AF_BLUE_STRINGSET_DEVA af_deva_uniranges segment_limit base_delta ydelta af_khms_nonbase_uniranges AF_BLUE_STRING_ARMENIAN_SMALL_TOP AF_BLUE_STRING_OL_CHIKI AF_STYLE_SHAW_DFLT af_latin_writing_system_class AF_Blue_String_ AF_Blue_StringRec_ af_goth_nonbase_uniranges af_telu_script_class AF_STYLE_MYMR_DFLT opos af_get_interface AF_BLUE_STRINGSET_CPRT is_straight link af_latn_c2sc_style_class AF_BLUE_STRING_SUNDANESE_DESCENDER AF_BLUE_STRINGSET_MAX af_cyrl_nonbase_uniranges other_flags xdelta has_serifs old_best_point AF_BLUE_STRINGSET_CARI AF_Err_Invalid_File_Format AF_BLUE_STRINGSET_MLYM af_cyrl_sinf_style_class AF_STYLE_AVST_DFLT af_geok_dflt_style_class AF_COVERAGE_SUPERSCRIPT af_cher_dflt_style_class stem_darkening_for_ppem af_shaper_buf_create AF_BLUE_STRING_CHAKMA_TOP AF_SCRIPT_NKOO AF_CJKBlue AF_STYLE_OSGE_DFLT AF_Coverage AF_Err_Invalid_CharMap_Format AF_SCRIPT_DSRT AF_SCRIPT_ADLM a_delta control_overshoot AF_BLUE_STRINGSET_VAII af_arab_dflt_style_class big_max af_telu_uniranges AF_Err_Ignore AF_BLUE_STRING_ARMENIAN_SMALL_BOTTOM af_limb_dflt_style_class AF_STYLE_HANI_DFLT AF_STYLE_GREK_C2SC AF_STYLE_ADLM_DFLT af_glag_dflt_style_class af_latin_hints_detect_features af_lao_uniranges AF_DIR_UP af_khmr_uniranges AF_GlyphHintsRec AF_BLUE_STRING_HEBREW_BOTTOM af_glyph_hints_align_edge_points scaled_stem AF_BLUE_STRING_BAMUM_TOP EndContour num_flats AF_BLUE_STRING_NKO_BOTTOM af_latin_hints_init AF_Err_Unimplemented_Feature u_off1 u_off2 AF_Err_Too_Many_Function_Defs AF_STYLE_LAO_DFLT AF_Err_Locations_Missing AF_Err_Code_Overflow af_latin_hints_compute_segments scores AF_BLUE_STRING_COPTIC_CAPITAL_BOTTOM AF_STYLE_DEVA_DFLT passed AF_BLUE_STRING_KANNADA_TOP style_options AF_BLUE_STRING_KHMER_BOTTOM AF_BLUE_STRING_LATIN_SMALL_TOP AF_BLUE_STRING_THAI_LARGE_ASCENDER edge_next AF_WritingSystem_InitMetricsFunc new_lsb left2right AF_BLUE_STRING_CHAKMA_BOTTOM AF_SCRIPT_TAVT AF_SCRIPT_GEOK AF_BLUE_STRING_LATIN_CAPITAL_TOP AF_SCRIPT_GEOR AF_Err_Invalid_Offset AF_BLUE_STRING_CHAKMA_DESCENDER len_score out_dir best_contour_first af_taml_script_class AF_DIMENSION_HORZ af_mlym_nonbase_uniranges gstyles AF_STYLE_GOTH_DFLT AF_BLUE_STRINGSET_MYMR af_sort_pos idx0 u_off AF_BLUE_STRING_GUJARATI_DIGIT_TOP af_cprt_nonbase_uniranges af_geok_script_class embedded af_nkoo_uniranges AF_Err_Syntax_Error last_v AF_SCRIPT_BUHD AF_BLUE_STRING_OSAGE_SMALL_DESCENDER af_loader_done af_beng_dflt_style_class af_ethi_nonbase_uniranges AF_BLUE_STRING_GEORGIAN_MTAVRULI_BOTTOM AF_BLUE_STRING_ADLAM_SMALL_TOP standard_vertical_width AF_BLUE_STRING_LATIN_CAPITAL_BOTTOM af_latn_nonbase_uniranges af_sund_nonbase_uniranges af_buhd_dflt_style_class blue_ref af_grek_script_class AF_STYLE_LATP_DFLT AF_BLUE_STRING_KHMER_LARGE_DESCENDER AF_BLUE_STRING_LISU_BOTTOM af_lisu_uniranges AF_BLUE_STRINGSET_AVST AF_STYLE_GLAG_DFLT af_grek_pcap_style_class af_loader_embolden_glyph_in_slot AF_BLUE_STRING_OSAGE_CAPITAL_TOP AF_WritingSystem_ScaleMetricsFunc af_adlm_nonbase_uniranges af_cjk_metrics_init af_bamu_script_class AF_BLUE_STRING_OSAGE_SMALL_BOTTOM AF_FaceGlobals AF_STYLE_BAMU_DFLT AF_Err_Out_Of_Memory AF_SCRIPT_GOTH AF_SCRIPT_ORKH af_telu_nonbase_uniranges AF_STYLE_CYRL_DFLT margin af_dummy_hints_apply af_glyph_hints_align_weak_points prev_min_flags AF_Err_Array_Too_Large AF_SCRIPT_CYRL AF_BLUE_STRING_OSMANYA_TOP AF_Err_Invalid_Slot_Handle AF_SCRIPT_COPT fitted_width AF_BLUE_STRING_HEBREW_TOP AF_BLUE_STRINGSET_MONG AF_STYLE_LATN_DFLT af_armn_nonbase_uniranges AF_Err_Horiz_Header_Missing AF_EdgeRec AF_SCRIPT_TFNG af_copt_uniranges af_taml_dflt_style_class AF_BLUE_STRINGSET_TAML AF_BLUE_STRING_SAURASHTRA_TOP af_indic_metrics_scale AF_BLUE_STRINGSET_SHAW AF_BLUE_STRING_CYPRIOT_BOTTOM af_lao_dflt_style_class AF_GlyphHintsRec_ AF_Segment AF_Err_Invalid_Glyph_Index AF_CJKAxisRec AF_Err_Invalid_PPem af_knda_script_class af_autofitter_done af_latp_dflt_style_class AF_Err_Unlisted_Object cur_idx AF_SCRIPT_HANI af_hebr_dflt_style_class af_orkh_uniranges best_pos AF_SCRIPT_OSGE af_ethi_dflt_style_class AF_BLUE_STRINGSET_LISU af_kali_script_class AF_Err_Invalid_Stream_Skip org_pos AF_BLUE_STRING_GUJARATI_DESCENDER af_latin_metrics_init_blues AF_STYLE_KHMS_DFLT af_geor_dflt_style_class af_saur_dflt_style_class af_mymr_script_class AF_Style_ AF_BLUE_STRING_LATIN_SUPS_SMALL_F_TOP af_tibt_dflt_style_class seg0 top_to_bottom_hinting seg2 AF_SCRIPT_GREK AF_BLUE_STRING_LISU_TOP af_sylo_script_class af_hebr_nonbase_uniranges AF_PointRec_ af_sylo_dflt_style_class af_latin_get_standard_widths AF_Err_Too_Few_Arguments AF_STYLE_KHMR_DFLT AF_SCRIPT_LATB best_blue_is_neutral af_cakm_nonbase_uniranges new_delta AF_SCRIPT_LATN AF_SCRIPT_LATP AF_COVERAGE_SMALL_CAPITALS AF_BLUE_STRING_GEORGIAN_MKHEDRULI_DESCENDER darken_amount AF_BLUE_STRING_NKO_TOP AF_Err_Missing_Startfont_Field AF_STYLE_KALI_DFLT af_blue_1_1_1 af_blue_1_1_2 len_threshold af_property_get_face_globals AF_EdgeRec_ AF_BLUE_STRING_OSAGE_SMALL_TOP AF_BLUE_STRING_AVESTAN_TOP AF_SCRIPT_DEVA AF_STYLE_CANS_DFLT af_grek_titl_style_class af_cyrl_c2sc_style_class af_khms_script_class AF_Blue_Stringset_ glyph_styles af_cjk_align_edge_points af_cprt_script_class best_y_extremum AF_SCRIPT_ARAB af_grek_c2cp_style_class segment_dir blue_count AF_BLUE_STRING_OSAGE_CAPITAL_BOTTOM AF_Err_Execution_Too_Long af_latin_metrics_init_widths af_knda_nonbase_uniranges AF_BLUE_STRING_TAMIL_TOP AF_Err_Invalid_Library_Handle af_latin_metrics_scale_dim AF_STYLE_TFNG_DFLT trans_matrix AF_BLUE_STRING_KHMER_SYMBOLS_WAXING_TOP endpoint num_edges af_mong_script_class AF_Blue_StringRec AF_Coverage_ af_orya_script_class af_latp_nonbase_uniranges AF_BLUE_STRING_ARABIC_BOTTOM AF_DIMENSION_MAX AF_CJKBlueRec size_changed AF_STYLE_KNDA_DFLT AF_BLUE_STRING_THAI_BOTTOM af_warper_weights AF_BLUE_STRING_SINHALA_DESCENDER AF_Err_Invalid_Handle AF_WritingSystem_GetStdWidthsFunc af_sylo_uniranges af_autofitter_interface AF_SCRIPT_SINH AF_BLUE_STRING_LAO_ASCENDER max_edges af_latin_hints_compute_edges af_cjk_align_linked_edge scale_down_factor AF_BLUE_STRINGSET_TAVT AF_BLUE_STRING_GOTHIC_TOP AF_BLUE_STRING_LATIN_SUPS_CAPITAL_TOP af_script_classes AF_Script_UniRangeRec AF_SCRIPT_BAMU AF_BLUE_STRING_CANADIAN_SYLLABICS_BOTTOM AF_BLUE_STRINGSET_NKOO AF_STYLE_LIMB_DFLT AF_BLUE_STRINGSET_DSRT AF_Err_Table_Missing wmax AF_BLUE_STRINGSET_ADLM af_hani_uniranges AF_BLUE_STRING_NKO_SMALL_BOTTOM af_khmr_dflt_style_class af_sylo_nonbase_uniranges af_armn_script_class af_glyph_hints_scale_dim af_osge_uniranges segment_width_threshold AF_Script_UniRangeRec_ AF_BLUE_STRING_GLAGOLITIC_SMALL_TOP af_cyrl_c2cp_style_class AF_SCRIPT_CPRT AF_BLUE_STRING_ADLAM_CAPITAL_BOTTOM AF_STYLE_CYRL_TITL AF_SCRIPT_KHMR AF_SCRIPT_KHMS p_first AF_WritingSystemClassRec AF_BLUE_STRING_COPTIC_SMALL_BOTTOM AF_STYLE_SINH_DFLT darken_x darken_y AF_Err_Missing_Bbx_Field AF_Err_Invalid_Post_Table AF_STYLE_LATN_TITL AF_STYLE_BUHD_DFLT base_edge AF_Scaler AF_BLUE_STRING_CYRILLIC_CAPITAL_TOP writing_system AF_SCRIPT_CHER AF_COVERAGE_RUBY AF_BLUE_STRING_LATIN_SMALL_DESCENDER AF_STYLE_LATN_C2SC best_y bdelta pp2x_uh af_guru_dflt_style_class link1 af_knda_dflt_style_class AF_BLUE_STRING_VAI_TOP af_mong_nonbase_uniranges af_tavt_nonbase_uniranges af_copt_script_class AF_BLUE_STRING_GEORGIAN_MTAVRULI_TOP AF_BLUE_STRINGSET_GEOK AF_BLUE_STRING_CHEROKEE_CAPITAL AF_BLUE_STRINGSET_GEOR af_khmr_nonbase_uniranges AF_BLUE_STRING_GURMUKHI_BOTTOM af_latn_ordn_style_class AF_BLUE_STRING_TIFINAGH AF_WRITING_SYSTEM_MAX segment_length_threshold af_latn_uniranges style_metrics_getstdw AF_STYLE_ARAB_DFLT ametrics AF_BLUE_STRING_GLAGOLITIC_CAPITAL_BOTTOM af_cjk_hints_apply seg1 af_cakm_script_class af_latin_hints_apply AF_BLUE_STRING_THAI_DIGIT_TOP AF_BLUE_STRING_BUHID_BOTTOM AF_BLUE_STRING_ARMENIAN_CAPITAL_TOP AF_STYLE_LISU_DFLT af_glag_script_class AF_ScriptClassRec AF_BLUE_STRING_SHAVIAN_DESCENDER AF_BLUE_STRING_LATIN_SUPS_SMALL_DESCENDER af_orya_nonbase_uniranges old_charmap AF_BLUE_STRING_DESERET_CAPITAL_TOP AF_STYLE_HEBR_DFLT af_grek_uniranges af_geor_uniranges af_latin_align_serif_edge AF_BLUE_STRING_CJK_BOTTOM AF_Err_Invalid_Stream_Handle AF_StyleMetrics af_cjk_hints_compute_blue_edges standard_horizontal_width af_dummy_hints_init AF_LatinBlue AF_Err_Invalid_Pixel_Size AF_Direction af_indic_hints_init num_idx af_goth_dflt_style_class af_mlym_dflt_style_class af_taml_nonbase_uniranges AF_Err_Post_Table_Missing af_cjk_metrics_scale af_tibt_uniranges is_neutral_blue AF_DIR_LEFT xmax_delta AF_BLUE_STRINGSET_GOTH in_dir AF_BLUE_STRINGSET_ORKH AF_BLUE_STRING_CARIAN_TOP af_khmr_script_class af_olck_script_class AF_BLUE_STRING_GEORGIAN_MKHEDRULI_BOTTOM old_lsb NextContour af_shaw_nonbase_uniranges af_service_properties AF_BLUE_STRINGSET_CYRL AF_Err_Missing_Encoding_Field AF_SCRIPT_HEBR AF_WidthRec_ af_face_globals_compute_style_coverage af_hani_script_class af_osma_script_class AF_WarperRec af_mlym_uniranges af_arab_script_class AF_Err_Debug_OpCode AF_STYLE_GREK_DFLT AF_BLUE_STRING_KHMER_SUBSCRIPT_TOP AF_SCRIPT_ORYA af_olck_dflt_style_class af_gujr_nonbase_uniranges af_copt_nonbase_uniranges af_shaw_script_class AF_Err_Invalid_Opcode edge_limit AF_Err_Stack_Overflow AF_BLUE_STRINGSET_HEBR af_adlm_dflt_style_class AF_Script af_direction_compute fallback_script d_off2 AF_BLUE_STRING_GREEK_SMALL_BETA_TOP AF_STYLE_CYRL_C2SC AF_BLUE_STRING_GOTHIC_BOTTOM af_kali_nonbase_uniranges Skip_Loop default_script af_cyrl_dflt_style_class style_hints_apply dflt AF_BLUE_STRINGSET_HANI width_count AF_STYLE_TAVT_DFLT AF_BLUE_STRINGSET_OSGE AF_Err_Cannot_Render_Glyph laxis num_widths af_avst_script_class is_top_blue AF_STYLE_OLCK_DFLT stem_edge AF_Err_Glyph_Too_Big af_shaper_get_cluster AF_BLUE_STRING_THAI_DESCENDER af_shaw_dflt_style_class af_latb_dflt_style_class af_cyrl_subs_style_class AF_BLUE_STRING_DEVANAGARI_BOTTOM af_guru_script_class blue_edge AF_Err_DEF_In_Glyf_Bytecode point_limit AF_BLUE_STRINGSET_GREK AF_STYLE_DSRT_DFLT segments_end Done_Width AF_BLUE_STRING_LATIN_SUBS_CAPITAL_TOP AF_BLUE_STRING_SAURASHTRA_BOTTOM af_latp_uniranges AF_BLUE_STRING_GREEK_SMALL AF_Err_Too_Many_Caches AF_SCRIPT_SUND AF_BLUE_STRINGSET_LATB af_tavt_dflt_style_class AF_DIR_NONE AF_BLUE_STRINGSET_LATN AF_BLUE_STRINGSET_LATP AF_BLUE_STRING_DESERET_SMALL_BOTTOM is_major_dir af_cprt_dflt_style_class AF_SCRIPT_NONE AF_BLUE_STRING_GREEK_CAPITAL_BOTTOM af_cjk_compute_stem_width fitted af_vaii_uniranges dist1 AF_WritingSystemClass darken_by_font_units_y af_cari_script_class AF_SCRIPT_THAI af_latb_uniranges AF_Edge AF_SCRIPT_ARMN AF_BLUE_STRING_OSMANYA_BOTTOM AF_StyleMetricsRec_ AF_Script_ af_cjk_hints_compute_edges AF_Err_No_Unicode_Glyph_Name dist_demerit AF_SCRIPT_OLCK AF_BLUE_STRING_GREEK_CAPITAL_TOP AF_Blue_Stringset best_dist pp2x af_tibt_script_class AF_Err_Invalid_Horiz_Metrics af_dsrt_nonbase_uniranges AF_BLUE_STRING_CHEROKEE_SMALL AF_BLUE_STRINGSET_ARAB AF_Dimension AF_BLUE_STRING_CANADIAN_SYLLABICS_SUPS_BOTTOM AF_BLUE_STRING_BAMUM_BOTTOM AF_BLUE_STRING_CANADIAN_SYLLABICS_SMALL_BOTTOM AF_BLUE_STRING_SUNDANESE_TOP AF_BLUE_STRING_DESERET_CAPITAL_BOTTOM af_sinh_script_class af_sinh_dflt_style_class AF_Err_Missing_Module AF_STYLE_NONE_DFLT AF_STYLE_ARMN_DFLT AF_Err_Invalid_Cache_Handle af_latin_hints_link_segments Store_Point af_glyph_hints_align_strong_points on_edge af_services AF_BLUE_STRING_THAI_LARGE_DESCENDER xmin_delta AF_STYLE_CYRL_PCAP AF_Err_Max af_tfng_uniranges AF_Blue_String AF_BLUE_STRINGSET_SINH AF_Err_Missing_Chars_Field AF_BLUE_STRING_ARABIC_JOIN AF_StyleClass aglobals AF_STYLE_LATN_PCAP AF_BLUE_STRING_SHAVIAN_SMALL_BOTTOM fallback_style AF_Err_Missing_Bitmap af_bamu_nonbase_uniranges AF_GlyphHints af_indic_metrics_init AF_WritingSystem cur_len best_segment_first AF_BLUE_STRING_LATIN_SUBS_SMALL_F_TOP AF_DIR_RIGHT af_latn_pcap_style_class AF_Err_Cannot_Open_Stream base_distort AF_STYLE_CYRL_ORDN log_base_2 standard_charstring num_contours AF_STYLE_THAI_DFLT af_cjk_metrics_init_widths n_edges AF_BLUE_STRINGSET_OSMA af_cari_dflt_style_class digits_have_same_width AF_STYLE_LATN_ORDN edge_delta af_glag_nonbase_uniranges AF_BLUE_STRING_BUHID_LARGE af_cyrl_uniranges AF_SegmentRec_ AF_WRITING_SYSTEM_CJK AF_BLUE_STRING_THAI_ASCENDER af_cprt_uniranges AF_BLUE_STRINGSET_KHMR AF_BLUE_STRINGSET_KHMS AF_BLUE_STRING_CYRILLIC_SMALL af_none_uniranges pp1x AF_Loader slot_internal af_glyph_hints_save AF_WritingSystem_InitHintsFunc AF_STYLE_BENG_DFLT AF_STYLE_GREK_TITL AF_BLUE_STRING_TELUGU_BOTTOM af_latin_metrics_scale AF_BLUE_STRING_MONGOLIAN_BOTTOM_BASE AF_BLUE_STRINGSET_CHER af_blue_1_1 af_deva_script_class AF_LatinMetrics af_kali_dflt_style_class AF_BLUE_STRING_CANADIAN_SYLLABICS_TOP AF_BLUE_STRING_CJK_TOP af_latin_metrics_init af_orya_dflt_style_class af_gujr_script_class af_adlm_uniranges blue_shoot af_grek_smcp_style_class AF_Err_Invalid_Glyph_Format af_mong_dflt_style_class shaper_buf_ last_stem_pos af_blue_2_1_1 af_blue_2_1_2 AF_PointRec AF_BLUE_STRING_GLAGOLITIC_CAPITAL_TOP AF_Err_Cannot_Open_Resource cur_val af_mymr_nonbase_uniranges AF_BLUE_STRING_DEVANAGARI_TOP AF_BLUE_STRING_ADLAM_CAPITAL_TOP af_orya_uniranges af_latin_compute_stem_width AF_Err_Invalid_Stream_Seek a_scale af_sort_and_quantize_widths AF_BLUE_STRINGSET_TELU flat_threshold AF_Err_Bad_Argument af_latin_metrics_check_digits af_cakm_uniranges link2 AF_BLUE_STRING_CYRILLIC_SMALL_DESCENDER af_cyrl_titl_style_class over_ref contour_index af_shaper_get_coverage af_khms_dflt_style_class AF_SCRIPT_TIBT AF_BLUE_STRING_GEORGIAN_NUSKHURI_TOP af_copt_dflt_style_class base_flags AF_STYLE_GEOR_DFLT af_osma_uniranges prev_max_flags AF_Err_ENDF_In_Exec_Stream af_arab_nonbase_uniranges vvector af_grek_nonbase_uniranges af_latn_dflt_style_class af_geor_script_class af_writing_system_classes af_adlm_script_class af_olck_nonbase_uniranges glyph_count AF_Err_Could_Not_Find_Context num_fills af_cjk_snap_width af_iup_interp AF_SCRIPT_GUJR af_thai_nonbase_uniranges AF_WidthRec cur_ab PS_Hint_TableRec t2_hints_stems PS_Mask_TableRec_ align_top PSH_Err_Code_Overflow PSH_Err_Stack_Underflow psh_hint_snap_stem_side_delta /home/computerfido/Desktop/LemonTest/lemon-freetype/src/pshinter/pshinter.c PS_DimensionRec PSH_Err_Invalid_Stream_Skip PSH_Err_Invalid_PPem alignment strongs_0 pshinter_interface glyphrec PSH_ZoneRec PSH_Err_Missing_Property PSH_DIR_UP PSH_Err_Invalid_Composite cur_top PSH_Hint_TableRec_ ps_dimension_done PSH_AlignmentRec_ PSH_Err_Missing_Chars_Field PS_Mask_TableRec org_ab ps_hint_table_ensure PS_Hint_Table ps_hints_init direction psh_globals_scale_widths psh_glyph_find_strong_points ps_dimension_add_counter PSH_Err_Invalid_Character_Code ps_hints_t1reset psh_glyph_interpolate_other_points PS_HINT_TYPE_1 PSH_Alignment PSH_Err_Raster_Uninitialized hint_tables ps_dimension_init T1_Hints_FuncsRec old_y_scale PSH_Err_Unlisted_Object PSH_Err_Raster_Overflow PSH_Err_Invalid_CharMap_Handle psh_globals_new PS_HintsRec psh_glyph_find_blue_points PSH_Err_Table_Missing bit_pos PSH_Err_Cannot_Render_Glyph cur_height fit_count dimension PSH_Hint_TableRec PSH_Err_Too_Many_Hints PSH_Blue_TableRec_ PSH_Glyph finished PSH_Err_Invalid_Argument ps_dimension_add_t1stem PSH_Err_Bad_Argument PSH_DIR_LEFT PSH_Width PSH_Err_Too_Many_Caches PSH_Err_Nested_DEFS scale_ab scale_delta PSH_Err_Too_Many_Extensions org_bottom PSH_Err_Invalid_Outline psh_glyph_compute_extrema cur_max PSH_Err_Nested_Frame_Access ps_hints_stem PSH_Err_Invalid_Cache_Handle PSH_Err_Missing_Encoding_Field PS_Hint_Type read_count PSH_Contour t1_hints_stem PS_HintRec_ PSH_Blue_TableRec PSH_Err_Array_Too_Large max_bits PS_Hinter_Module dir_in psh_glyph_compute_inflections PSH_Err_Corrupted_Font_Glyphs par_cur_center cur_pos PSH_Err_Syntax_Error num_zones dim_x dim_y psh_hint_table_record_mask PSH_Err_Invalid_Version scale_mult fit_len PSH_ContourRec_ do_horz_hints bit_count PS_Hinter_Module_Rec_ PSH_Err_Horiz_Header_Missing ps_hints no_overshoots PSH_Err_Too_Many_Function_Defs PSH_Err_Too_Few_Arguments PSH_Err_Corrupted_Font_Header PS_Dimension PSH_DimensionRec sort_global do_horz_snapping no_shoots PSH_Err_Invalid_CharMap_Format n_prev is_others ps_mask_set_bit psh_hint_table_find_strong_points psh_blues_set_zones PSH_Hint_Table PS_Hints PSH_GlyphRec PSH_Err_DEF_In_Glyf_Bytecode PSH_Err_Invalid_Frame_Read min_flag max_masks PSH_Err_No_Unicode_Glyph_Name PSH_Err_Stack_Overflow psh_dimension_quantize_len PSH_Dimension PS_Hint ahint psh_blues_set_zones_0 wmask left_nearest ps_hints_apply t1_hints_funcs_init psh_globals_destroy mask1 align_bot PSH_Err_Invalid_Handle PSH_Err_Lower_Module_Version PSH_Blue_Zone num_masks rmask PSH_Widths PSH_Err_Invalid_Opcode PSH_BluesRec right_disp orient_prev PS_Mask PS_DimensionRec_ PSH_Err_Raster_Corrupted blue_threshold PSH_Err_Invalid_Glyph_Format PSH_Err_Out_Of_Memory ps_mask_table_merge pshinter_get_globals_funcs psh_globals_set_scale PSH_Err_Invalid_Reference org_ac cur_a PSH_Err_Invalid_Glyph_Index cur_c PSH_HintRec_ ps_mask_table_ensure PSH_Err_Invalid_Face_Handle PSH_Err_Invalid_Slot_Handle cur_u PSH_Hint old_x_scale t2_hints_funcs_init PSH_DimensionRec_ PSH_Err_Missing_Size_Field hint2 ps_mask_table_done ps_mask_test_bit PSH_Err_Invalid_Vert_Metrics ps_hints_close PS_HINT_TYPE_2 PSH_Err_Missing_Module org_top psh_calc_max_height PSH_Err_Unknown_File_Format do_vert_snapping PSH_Err_Invalid_CodeRange PSH_ZoneRec_ PSH_Err_Too_Many_Instruction_Defs ps_hints_t2mask psh_blues_snap_stem count_top stem_bot T2_Hints_FuncsRec hint_masks PSH_Err_Execution_Too_Long ps_hinter_done PSH_Err_Invalid_Stream_Handle ps_dimension_set_mask_bits ps_hints_open psh_hint_table_activate_mask psh_glyph_load_points count1 PSH_Err_ENDF_In_Exec_Stream max_hints ps_hint_table_alloc zone2 count_bot point_dir psh_compute_dir pshinter_get_t2_funcs PSH_Globals_FuncsRec left_disp ps_mask_table_alloc psh_glyph_interpolate_strong_points n_next PSH_Err_Invalid_Stream_Seek stand PSH_Err_Glyph_Too_Big psh_hint_table_align_hints PSH_Err_CMap_Table_Missing PSH_Err_Name_Table_Missing PSH_WidthsRec ps_dimension_end_mask normal_top PSH_Err_Invalid_Table Next_Contour family_top PSH_Err_Cannot_Open_Stream PSH_DIR_NONE ps_mask_table_merge_all PSH_Err_Invalid_Pixel_Size counter_masks org_v hint1 hint3 flags2 PSH_Err_Cannot_Open_Resource PSH_Err_Invalid_Size_Handle points_end family_bottom cur_bottom PSH_GlyphRec_ PSH_Err_Max PSH_Err_Missing_Startfont_Field ps_hints_t2counter aindex PSH_Err_Hmtx_Table_Missing PSH_Err_Missing_Font_Field PSH_Err_Ignore psh_blues_scale_zones PSH_Err_Invalid_Frame_Operation psh_hint_align PSH_Err_Unimplemented_Feature PSH_WidthRec_ ps_hinter_init cur_org_center source_bits psh_hint_table_record PSH_Err_Raster_Negative_Height orient_cur psh_glyph_interpolate_normal_points counters PSH_WidthsRec_ top_table psh_hint_overlap cur_ref delta0 par_org_center PSH_Blues Extremum org_ref right_nearest PSH_Err_Too_Many_Drivers PSH_Zone PSH_Blue_ZoneRec PSH_Err_Post_Table_Missing psh_hint_table_done psh_hint_table_init PS_Hint_Type_ PSH_PointRec_ PSH_Blue_Table PSH_Err_Invalid_Stream_Operation PS_Hint_TableRec_ PS_MaskRec_ ps_mask_table_set_bits mask2 PSH_DIR_RIGHT stem_top PS_Mask_Table t2_hints_open normal_bottom PSH_Err_Could_Not_Find_Context PSH_Err_Invalid_Library_Handle psh_glyph_done PS_MaskRec source_pos pshinter_get_t1_funcs PSH_Err_Divide_By_Zero ps_mask_table_test_intersect t1_hints_open PS_HintsRec_ do_stem_adjust org_c PSH_Err_Invalid_Stream_Read PSH_AlignmentRec PSH_Err_Invalid_Post_Table_Format minor_dir ps_mask_clear_bit psh_glyph_save_points PSH_Err_Bbx_Too_Big PSH_DIR_DOWN org_a PSH_Err_Invalid_Post_Table num_bits num_strongs do_vert_hints org_u PSH_WidthRec max_scale dir_out ps_mask_table_last PSH_Err_Invalid_File_Format PSH_Err_Missing_Bbx_Field PSH_Err_Invalid_Horiz_Metrics PSH_Err_Debug_OpCode hint_mask ps_mask_done PSH_BluesRec_ PSH_Err_Missing_Bitmap psh_globals_funcs_init ps_hints_done hint_type ps_dimension_end do_snapping ps_hint_table_done max_flag PSH_Err_Locations_Missing ps_dimension_reset_mask zone1 psh_hint_table_deactivate ps_hints_t1stem3 PSH_Err_Missing_Startchar_Field amask PSH_Err_Invalid_Offset ps_mask_ensure PSH_Err_Ok count_others psh_glyph_init PSH_Point PSH_Blue_ZoneRec_ bot_table PSH_Err_Missing_Fontboundingbox_Field PSH_Err_Invalid_Driver_Handle Line_Up Raster_Err_Missing_Chars_Field Raster_Err_Nested_DEFS High max_Y Raster_Err_Out_Of_Memory Raster_Err_Could_Not_Find_Context Raster_Err_Unlisted_Object y_turns Decompose_Curve ft_raster1_init lastY Cubic_To joint Raster_Err_Missing_Startfont_Field min_Y Raster_Err_Invalid_File_Format ymin2 Raster_Err_Locations_Missing TStates Raster_Err_Stack_Underflow TProfileList Horizontal_Sweep_Init Raster_Err_Invalid_CharMap_Format black_TBand_ start_arc Raster_Err_Missing_Fontboundingbox_Field Bezier_Down band_stack Raster_Err_Ok precision Sort Bezier_Up ft_raster1_set_mode Raster_Err_Invalid_Table Raster_Err_Invalid_Size_Handle Raster_Err_Invalid_CodeRange P_Right Function_Sweep_Span Raster_Err_Too_Many_Function_Defs draw_left Raster_Err_Invalid_Driver_Handle Raster_Err_CMap_Table_Missing Raster_Err_Raster_Overflow New_Profile target_map ymax1 black_PRaster Raster_Err_Unimplemented_Feature Proc_Sweep_Span Skip_To_Next Raster_Err_Invalid_Character_Code Raster_Err_Raster_Uninitialized InsNew araster Vertical_Sweep_Span Raster_Err_Too_Many_Caches Raster_Err_ENDF_In_Exec_Stream Raster_Err_Invalid_Outline End_Profile ft_black_done Next_Line Raster_Err_Invalid_Post_Table_Format Raster_Err_Divide_By_Zero Raster_Err_Table_Missing /home/computerfido/Desktop/LemonTest/lemon-freetype/src/raster/raster.c Raster_Err_Too_Many_Extensions Proc_Sweep_Drop Flat_State pool_base Raster_Err_Array_Too_Large Conic_To Raster_Err_Invalid_Reference TPoint Raster_Err_Invalid_Glyph_Index countL precision_bits y_change ymin Unknown_State Horizontal_Sweep_Step PProfileList cProfile band_top Raster_Err_Debug_OpCode Raster_Err_Invalid_Frame_Operation traceOfs Raster_Err_Missing_Size_Field Raster_Err_Corrupted_Font_Glyphs ft_standard_raster Line_Down Raster_Err_Missing_Encoding_Field Raster_Err_Invalid_Stream_Seek Raster_Err_DEF_In_Glyf_Bytecode ft_black_init P_Left Raster_Err_Cannot_Open_Stream Raster_Err_Corrupted_Font_Header Raster_Err_Invalid_Pixel_Size Raster_Err_Missing_Bbx_Field precision_half Scan_DropOuts ft_raster1_render ft_raster1_get_cbox Raster_Err_Missing_Font_Field Raster_Err_Too_Many_Drivers gProfile numTurns Raster_Err_Invalid_PPem arcs num_Profs traceIncr Raster_Err_Horiz_Header_Missing Raster_Err_Invalid_Argument Raster_Err_Invalid_Cache_Handle Convert_Glyph flipped ft_black_reset Raster_Err_Max Raster_Err_Cannot_Open_Resource TProfile Raster_Err_Too_Many_Hints Horizontal_Sweep_Drop Raster_Err_Nested_Frame_Access Raster_Err_Invalid_Stream_Operation mode_tag Raster_Err_Invalid_Composite Raster_Err_Cannot_Render_Glyph Raster_Err_Invalid_Vert_Metrics Raster_Err_Code_Overflow black_TBand black_TWorker Raster_Err_Post_Table_Missing Vertical_Sweep_Drop bWidth TSplitter Raster_Err_Too_Few_Arguments sizeBuff maxBuff Raster_Err_Name_Table_Missing dropouts oldProfile lastProfile precision_step Horizontal_Sweep_Span fProfile maxY Raster_Err_Invalid_Stream_Handle Raster_Err_Invalid_CharMap_Handle Raster_Err_Missing_Startchar_Field maxy ft_black_set_mode Raster_Err_Execution_Too_Long bOrigin Raster_Err_Ignore splitter Raster_Err_Glyph_Too_Big Ascending_State aState dropOutControl black_TWorker_ ft_black_new precision_jitter ymax ymax2 fresh Raster_Err_Hmtx_Table_Missing Vertical_Sweep_Init Raster_Err_Invalid_Offset Raster_Err_Raster_Corrupted Insert_Y_Turn DelOld black_TRaster_ second_pass PByte state_bez Raster_Err_Stack_Overflow PLong Raster_Err_Invalid_Stream_Skip TPoint_ Raster_Err_Invalid_Slot_Handle Proc_Sweep_Init Descending_State ft_black_render Render_Single_Pass Raster_Err_Invalid_Handle Raster_Err_Invalid_Stream_Read Split_Conic black_PWorker Raster_Err_Invalid_Opcode Raster_Err_Missing_Property Split_Cubic Function_Sweep_Init Finalize_Profile_Table Raster_Err_No_Unicode_Glyph_Name Init_Linked ft_raster1_transform precision_scale Vertical_Sweep_Step Raster_Err_Invalid_Frame_Read lastX waiting Raster_Err_Lower_Module_Version Raster_Err_Invalid_Horiz_Metrics Raster_Err_Bbx_Too_Big Set_High_Precision Raster_Err_Missing_Bitmap Raster_Err_Invalid_Glyph_Format Raster_Err_Missing_Module Raster_Err_Too_Many_Instruction_Defs TStates_ Raster_Err_Raster_Negative_Height Line_To minY Draw_Sweep Raster_Err_Invalid_Library_Handle Function_Sweep_Step Raster_Err_Bad_Argument miny Raster_Err_Invalid_Post_Table Proc_Sweep_Step Raster_Err_Invalid_Face_Handle Raster_Err_Syntax_Error Raster_Err_Invalid_Version TProfile_ PProfile draw_right ymin1 Raster_Err_Unknown_File_Format Smooth_Err_Missing_Startchar_Field Smooth_Err_Hmtx_Table_Missing Smooth_Err_Too_Many_Extensions FT_Trace_Enable Smooth_Err_Glyph_Too_Big ft_smooth_render Smooth_Err_Too_Many_Instruction_Defs ft_smooth_set_mode gray_render_conic Smooth_Err_Invalid_File_Format bands gray_raster_reset gray_raster_render gray_move_to Smooth_Err_Invalid_Offset Smooth_Err_Invalid_Horiz_Metrics gray_sweep ft_smooth_render_lcd_v gray_render_line Smooth_Err_Missing_Chars_Field Smooth_Err_Stack_Overflow Smooth_Err_Cannot_Open_Resource Smooth_Err_Missing_Font_Field Smooth_Err_Missing_Fontboundingbox_Field dx_r Smooth_Err_Invalid_Handle TPixmap_ Smooth_Err_Raster_Overflow Smooth_Err_Missing_Size_Field gray_split_conic Smooth_Err_Too_Few_Arguments Smooth_Err_Invalid_Opcode PCell Smooth_Err_Invalid_Outline Smooth_Err_Invalid_Post_Table ft_smooth_render_generic TArea Smooth_Err_Invalid_CodeRange gray_PRaster gray_hline Smooth_Err_Bad_Argument Smooth_Err_Missing_Encoding_Field Smooth_Err_Array_Too_Large gray_raster_new Smooth_Err_Invalid_Table prod pcell Smooth_Err_Invalid_Slot_Handle Smooth_Err_Raster_Negative_Height Smooth_Err_Too_Many_Drivers ft_smooth_transform Smooth_Err_Missing_Bitmap TCell gray_convert_glyph Smooth_Err_Invalid_Glyph_Format Smooth_Err_Locations_Missing Smooth_Err_Unimplemented_Feature gray_raster_done Smooth_Err_Invalid_Size_Handle Smooth_Err_Bbx_Too_Big Smooth_Err_Invalid_Stream_Seek Smooth_Err_Max Smooth_Err_Invalid_Driver_Handle Smooth_Err_Code_Overflow /home/computerfido/Desktop/LemonTest/lemon-freetype/src/smooth/smooth.c cover Smooth_Err_Lower_Module_Version continued Smooth_Err_ENDF_In_Exec_Stream Smooth_Err_Missing_Startfont_Field TPixmap Smooth_Err_Invalid_Frame_Operation min_ex gray_PWorker ycells gray_convert_glyph_inner num_spans to_x to_y Smooth_Err_Invalid_Stream_Handle ft_smooth_render_lcd Smooth_Err_Invalid_CharMap_Handle max_cells Smooth_Err_Nested_DEFS Split Smooth_Err_Table_Missing Smooth_Err_Invalid_Frame_Read gray_set_cell Smooth_Err_Could_Not_Find_Context Smooth_Err_Invalid_Library_Handle num_cells min_ey FT_Trace_Disable gray_raster_set_mode Smooth_Err_Divide_By_Zero Smooth_Err_DEF_In_Glyf_Bytecode Smooth_Err_Syntax_Error Smooth_Err_Ignore Smooth_Err_Invalid_CharMap_Format Smooth_Err_Invalid_Glyph_Index gray_conic_to gray_TRaster_ Smooth_Err_Missing_Bbx_Field TCoord gray_render_cubic render_span_data bez_stack gray_cubic_to Smooth_Err_Debug_OpCode Smooth_Err_Invalid_Stream_Operation Smooth_Err_No_Unicode_Glyph_Name Smooth_Err_Too_Many_Function_Defs gray_TWorker Smooth_Err_CMap_Table_Missing Smooth_Err_Name_Table_Missing Smooth_Err_Raster_Corrupted Smooth_Err_Cannot_Open_Stream ft_smooth_init required_mode Smooth_Err_Stack_Underflow Smooth_Err_Invalid_Pixel_Size Smooth_Err_Invalid_Face_Handle hmul gray_TWorker_ Smooth_Err_Invalid_Stream_Skip Smooth_Err_Raster_Uninitialized gray_record_cell Smooth_Err_Invalid_Stream_Read draw TCell_ Smooth_Err_Invalid_Composite ft_grays_raster Smooth_Err_Invalid_Argument Smooth_Err_Invalid_PPem Smooth_Err_Nested_Frame_Access Smooth_Err_Unlisted_Object Smooth_Err_Invalid_Character_Code ft_smooth_get_cbox vmul Smooth_Err_Invalid_Vert_Metrics gray_split_cubic Smooth_Err_Invalid_Cache_Handle Smooth_Err_Out_Of_Memory TPos Smooth_Err_Too_Many_Caches max_ex max_ey Smooth_Err_Post_Table_Missing Smooth_Err_Horiz_Header_Missing Smooth_Err_Cannot_Render_Glyph Smooth_Err_Invalid_Post_Table_Format band Smooth_Err_Too_Many_Hints gray_line_to Smooth_Err_Invalid_Reference Smooth_Err_Corrupted_Font_Glyphs Smooth_Err_Missing_Property Smooth_Err_Missing_Module Smooth_Err_Ok Smooth_Err_Execution_Too_Long dy_r render_span Smooth_Err_Invalid_Version Smooth_Err_Corrupted_Font_Header Smooth_Err_Unknown_File_Format WASH ft_gzip_file_skip_output ft_gzip_alloc voidpf Gzip_Err_Invalid_Vert_Metrics nowrap Gzip_Err_Post_Table_Missing inflate_codes_new Gzip_Err_Invalid_Table CHECK1 Gzip_Err_Invalid_Cache_Handle total_in Gzip_Err_Missing_Size_Field Gzip_Err_Ok window Gzip_Err_Invalid_Slot_Handle zalloc fixed_bd Gzip_Err_Array_Too_Large fixed_bl Gzip_Err_Missing_Fontboundingbox_Field Gzip_Err_Execution_Too_Long Gzip_Err_Invalid_Offset zstream Gzip_Err_Max z_stream CODES inflate_block_mode Gzip_Err_Invalid_Horiz_Metrics ft_gzip_file_fill_output Gzip_Err_Hmtx_Table_Missing inflate_codes_free check_func inflate_mask inflate total_out cpdext Gzip_Err_Invalid_Size_Handle __mlibc_errno checkfn Gzip_Err_Invalid_Opcode Gzip_Err_Corrupted_Font_Glyphs Gzip_Err_Code_Overflow uLong Gzip_Err_Missing_Property Gzip_Err_DEF_In_Glyf_Bytecode adler DICT1 DICT2 DICT3 DICT4 inflate_codes_state inflateReset FT_GZipFileRec_ Bytef Gzip_Err_Ignore TABLE marker trees BLOCKS inflateEnd inflate_trees_bits Gzip_Err_Missing_Bitmap Gzip_Err_Invalid_Stream_Operation DISTEXT Gzip_Err_Debug_OpCode inflate_huft_s zip_buff Gzip_Err_Too_Many_Drivers DTREE Gzip_Err_Invalid_PPem Gzip_Err_Table_Missing next_out Gzip_Err_Nested_Frame_Access Gzip_Err_Missing_Bbx_Field INFLATE_DONE inflate_blocks_reset decode Gzip_Err_Invalid_Argument BADCODE inflate_flush Gzip_Err_Missing_Encoding_Field avail_out lbits Gzip_Err_Invalid_Post_Table Gzip_Err_Invalid_Glyph_Index program_invocation_name method Gzip_Err_Raster_Negative_Height Gzip_Err_Too_Many_Function_Defs Gzip_Err_No_Unicode_Glyph_Name CHECK2 CHECK3 CHECK4 zcalloc Gzip_Err_Unimplemented_Feature inflate_blocks_free ft_gzip_file_reset Gzip_Err_Syntax_Error Bits inflate_blocks_statef inflateInit2_ inflate_codes need Gzip_Err_Missing_Chars_Field inflate_huft dtree ft_gzip_file_done Gzip_Err_ENDF_In_Exec_Stream Gzip_Err_Invalid_Composite inflate_trees_fixed COPY z_stream_s ft_gzip_get_uncompressed_size Gzip_Err_Invalid_Stream_Seek FT_GZipFile alloc_func free_func Gzip_Err_Stack_Underflow Gzip_Err_Stack_Overflow avail_in Gzip_Err_Glyph_Too_Big Gzip_Err_Raster_Corrupted uLongf z_streamp bitb Gzip_Err_Invalid_Post_Table_Format bitk inflate_blocks_state Gzip_Err_Invalid_Reference BTREE Gzip_Err_Divide_By_Zero dbits zcfree Gzip_Err_Out_Of_Memory Gzip_Err_Raster_Uninitialized Gzip_Err_Lower_Module_Version Gzip_Err_Unlisted_Object Gzip_Err_Raster_Overflow ft_gzip_file_init ft_gzip_stream_close Gzip_Err_Could_Not_Find_Context opaque Gzip_Err_Cannot_Render_Glyph uIntf Gzip_Err_Invalid_Face_Handle ft_gzip_file_io inflate_trees_dynamic fixed_td fixed_tl Gzip_Err_Locations_Missing Gzip_Err_Too_Many_Caches Gzip_Err_Invalid_CharMap_Format Gzip_Err_Corrupted_Font_Header Gzip_Err_Invalid_Frame_Read what /home/computerfido/Desktop/LemonTest/lemon-freetype/src/gzip/ftgzip.c Gzip_Err_Invalid_Outline inflate_mode Gzip_Err_Too_Many_Instruction_Defs next_in program_invocation_short_name METHOD adler32 INFLATE_BAD Gzip_Err_Unknown_File_Format Gzip_Err_Bad_Argument Gzip_Err_Too_Few_Arguments Gzip_Err_Too_Many_Extensions LENEXT ltree inflate_blocks_new input_len DICT0 Gzip_Err_Missing_Startchar_Field Gzip_Err_Invalid_Version Gzip_Err_Nested_DEFS ft_gzip_free Exop Gzip_Err_Invalid_File_Format Gzip_Err_Missing_Startfont_Field cpdist ft_gzip_stream_io Gzip_Err_Invalid_Frame_Operation Gzip_Err_Invalid_Handle Gzip_Err_Invalid_Driver_Handle inflate_blocks ft_gzip_check_header old_pos Gzip_Err_CMap_Table_Missing ft_gzip_file_fill_input Gzip_Err_Invalid_Stream_Skip Gzip_Err_Invalid_Glyph_Format Gzip_Err_Name_Table_Missing zfree data_type uInt Gzip_Err_Invalid_Stream_Read Gzip_Err_Horiz_Header_Missing Gzip_Err_Cannot_Open_Stream Gzip_Err_Invalid_Pixel_Size zip_size huft_build cplens DIST STORED Gzip_Err_Invalid_Character_Code Gzip_Err_Too_Many_Hints Gzip_Err_Missing_Font_Field Gzip_Err_Invalid_Stream_Handle stream_size Gzip_Err_Invalid_CharMap_Handle Gzip_Err_Invalid_CodeRange inflate_codes_mode Gzip_Err_Missing_Module internal_state border LENS blens Gzip_Err_Invalid_Library_Handle cplext inflate_codes_statef Gzip_Err_Cannot_Open_Resource hufts Gzip_Err_Bbx_Too_Big wbits ft_lzw_file_done LZW_Err_Invalid_Glyph_Index LZW_Err_Missing_Size_Field LZW_Err_Out_Of_Memory LZW_Err_Could_Not_Find_Context LZW_Err_Invalid_Library_Handle stack_top LZW_Err_Invalid_Frame_Read LZW_Err_Invalid_CharMap_Format LZW_Err_Stack_Overflow LZW_Err_Missing_Bbx_Field NextCode LZW_Err_Invalid_Horiz_Metrics LZW_Err_Invalid_Face_Handle ft_lzw_stream_close LZW_Err_Invalid_Opcode LZW_Err_Locations_Missing LZW_Err_Syntax_Error LZW_Err_Invalid_Stream_Skip LZW_Err_Cannot_Open_Resource LZW_Err_Too_Few_Arguments /home/computerfido/Desktop/LemonTest/lemon-freetype/src/lzw/ftlzw.c LZW_Err_Invalid_Stream_Read ft_lzw_file_reset LZW_Err_Missing_Bitmap LZW_Err_Invalid_Vert_Metrics LZW_Err_Nested_DEFS LZW_Err_Debug_OpCode LZW_Err_Missing_Module ft_lzwstate_refill old_char LZW_Err_Max LZW_Err_Horiz_Header_Missing ft_lzw_stream_io LZW_Err_Invalid_Composite LZW_Err_Invalid_Stream_Operation FT_LzwStateRec LZW_Err_Invalid_Post_Table_Format prefix_size LZW_Err_Array_Too_Large buf_total LZW_Err_Invalid_Stream_Handle FT_LZW_PHASE_START ft_lzw_check_header LZW_Err_Cannot_Render_Glyph LZW_Err_Invalid_Argument LZW_Err_Post_Table_Missing FT_LZW_PHASE_CODE free_bits out_size ft_lzw_file_fill_output LZW_Err_Invalid_CharMap_Handle LZW_Err_Ignore old_size LZW_Err_Invalid_Offset LZW_Err_Invalid_PPem ft_lzw_file_skip_output buf_clear ft_lzw_file_io LZW_Err_Invalid_Reference LZW_Err_DEF_In_Glyf_Bytecode LZW_Err_Too_Many_Instruction_Defs LZW_Err_Missing_Chars_Field LZW_Err_Invalid_Driver_Handle buf_tab LZW_Err_Bbx_Too_Big LZW_Err_No_Unicode_Glyph_Name ft_lzwstate_get_code LZW_Err_Unimplemented_Feature LZW_Err_Too_Many_Hints FT_LzwStateRec_ LZW_Err_Invalid_Table LZW_Err_Invalid_File_Format LZW_Err_CMap_Table_Missing LZW_Err_Name_Table_Missing LZW_Err_Too_Many_Function_Defs LZW_Err_Cannot_Open_Stream LZW_Err_Invalid_Pixel_Size LZW_Err_Lower_Module_Version FT_LZWFile FT_LZW_PHASE_STACK LZW_Err_Invalid_Handle LZW_Err_Raster_Corrupted LZW_Err_Missing_Font_Field FT_LzwPhase_ ft_lzwstate_reset LZW_Err_Invalid_Glyph_Format stack_0 LZW_Err_Missing_Property FT_LzwState LZW_Err_Raster_Negative_Height LZW_Err_Divide_By_Zero LZW_Err_Too_Many_Extensions LZW_Err_Code_Overflow suffix FT_LZW_PHASE_EOF LZW_Err_Missing_Fontboundingbox_Field ft_lzwstate_prefix_grow LZW_Err_Corrupted_Font_Glyphs LZW_Err_Glyph_Too_Big FT_LZWFileRec_ LZW_Err_Execution_Too_Long LZW_Err_Invalid_CodeRange LZW_Err_Invalid_Slot_Handle LZW_Err_Table_Missing LZW_Err_Corrupted_Font_Header LZW_Err_Stack_Underflow ft_lzwstate_done LZW_Err_Missing_Encoding_Field LZW_Err_Hmtx_Table_Missing ft_lzw_file_init old_code ft_lzwstate_stack_grow LZW_Err_ENDF_In_Exec_Stream LZW_Err_Bad_Argument LZW_Err_Ok LZW_Err_Invalid_Size_Handle LZW_Err_Raster_Overflow LZW_Err_Raster_Uninitialized numread LZW_Err_Invalid_Stream_Seek LZW_Err_Invalid_Character_Code LZW_Err_Missing_Startchar_Field LZW_Err_Missing_Startfont_Field LZW_Err_Too_Many_Caches LZW_Err_Invalid_Frame_Operation LZW_Err_Invalid_Outline ft_lzwstate_init LZW_Err_Too_Many_Drivers FT_LzwPhase LZW_Err_Unknown_File_Format LZW_Err_Nested_Frame_Access ft_lzwstate_io LZW_Err_Invalid_Cache_Handle LZW_Err_Unlisted_Object LZW_Err_Invalid_Version LZW_Err_Invalid_Post_Table buf_offset free_ent in_eof max_free in_code cf2_builder_lineTo FieldArray CF2_Err_Missing_Startchar_Field bitCount PSaux_Err_Syntax_Error moveUp op_endchar cf2_hint_isPair AFM_VALUE_TYPE_STRING haveWidth ps_table_new needWinding PSaux_Err_Missing_Startchar_Field aint CF2_Matrix_ cf2_cmdRLINETO cf2_stack_pushFixed vStemHintArray summand1 cf2_escRANDOM AFM_TOKEN_CAPHEIGHT CF2_Err_Too_Many_Instruction_Defs AFM_TOKEN_XHEIGHT cf2_hintmask_setCounts charstring_base PSaux_Err_Invalid_Post_Table_Format cff_builder_start_point PSaux_Err_Table_Missing in_offset darkenX darkenY afm_key_table T1_CMapStd t1_cmap_custom_init PSaux_Err_Invalid_Glyph_Index currentCS PSaux_Err_Unknown_File_Format PSaux_Err_Bad_Argument cf2_cmdCALLGSUBR cf2_arrstack_init CF2_PathOpQuadTo topHintEdge initialHintMap csFlatEdge CF2_Err_Invalid_Version CF2_BluesRec charstringIndex AFM_TOKEN_STARTKERNDATA otherBlues PSaux_Err_Name_Table_Missing PSaux_Err_Invalid_PPem CF2_StackNumber_ ps_builder_done cf2_hint_isPairTop op_hlineto flatFamilyEdge CF2_MAX_HINTS curp familyBlues cff_decoder cff_builder_funcs ps_tobool captured currentDS ps_table_release PSaux_Err_Invalid_Reference cf2_escGET CF2_Err_Corrupted_Font_Glyphs PSaux_Err_Corrupted_Font_Header cf2_buf_isEnd PSaux_Err_Too_Many_Instruction_Defs logBase2 AFM_TOKEN_VVECTOR t1_builder_add_contour CF2_Err_Corrupted_Font_Header CF2_BufferRec AFM_TOKEN_W1X CF2_Err_Invalid_CharMap_Format normalizedV t1_cmap_expert_init emBoxTop emBoxBottomEdge psaux_get_glyph_name cf2_cmdRESERVED_17 PSaux_Err_Missing_Chars_Field renderingFlags upMoveDown CF2_Err_Too_Many_Extensions PSaux_Err_Missing_Bitmap cf2_escFLEX1 PSaux_Err_Raster_Corrupted cf2_cmdBLEND afm_stream_read_one intersection cf2_glyphpath_computeIntersection hintOffset t1_cmap_std_init PSaux_Err_Missing_Module CF2_HintRec PSaux_Err_Cannot_Open_Resource CF2_Err_Invalid_Handle cf2_cmdCNTRMASK emRatio FT_Fast op_hsbw cf2_stack_popInt dsCoord AFM_VALUE_TYPE_INTEGER PSAux_Interface sizeItem t1_lookup_glyph_by_stdcharcode_ps AFM_TOKEN_STARTCOMPOSITES AFM_TOKEN_W0X AFM_TOKEN_W0Y AFM_TOKEN_AXISTYPE CF2_Outline factor2 cf2_getNominalWidthX AFM_VALUE_TYPE_FIXED PSaux_Err_Invalid_Slot_Handle CF2_Err_Bbx_Too_Big blueFuzz cf2_cmdHMOVETO cf2_getT1SeacComponent CF2_Err_Debug_OpCode cf2_cmdVSINDEX PSaux_Err_ENDF_In_Exec_Stream AFM_TOKEN_STARTKERNPAIRS1 cf2_stack_clear PSaux_Err_Lower_Module_Version op_vhcurveto CF2_Err_Invalid_Face_Handle cf2_hint_isValid flatEdge CF2_Err_Invalid_Stream_Read get_callback cf2_getOtherBlues AFM_TOKEN_CC AFM_TOKEN_CH ps_parser_skip_spaces cf2_hintmask_init CF2_StackNumber cf2_glyphpath_curveTo PSaux_Err_Glyph_Too_Big AFM_Token cf2_hintmap_dump CF2_Err_Code_Overflow cf2_cmdVSTEMHM t1_cmap_std_char_index have_underflow hStemHintArray cf2_hintmap_build ps_table_add CF2_Err_Glyph_Too_Big PSaux_Err_Invalid_Argument chunk PSaux_Err_Missing_Bbx_Field PSaux_Err_Cannot_Render_Glyph AFM_TOKEN_FONTNAME pflags cff_builder_add_point known_othersubr_result_cnt op_hstem cf2_escDUP AFM_TOKEN_NOTICE scaleX scaleY snapThreshold cf2_escMUL cf2_escNOT darkenAmount CF2_GhostTop fracUp PSaux_Err_Execution_Too_Long pathIsClosing glyphWidth ps_builder_add_contour afm_parse_kern_pairs bottomHintEdge doConditionalLastRead cf2_escPUT ps_parser_load_field_table end_section CF2_NumberType_ CF2_Err_Missing_Chars_Field emBoxBottom CF2_Err_Missing_Module skip_procedure CF2_PairBottom CF2_Err_Missing_Font_Field cf2_hint_lock curX curY skip_literal_string op_div CF2_Callback_Type t1_cmap_standard_init cf2_getScaleAndHintFlag afm_stream_read_string CF2_NumberFrac cf2_cmdVHCURVETO ps_parser_to_fixed_array ps_parser_to_int lsb_x lsb_y subtrahend CF2_Err_Invalid_Opcode CF2_Err_Cannot_Open_Resource doEmBoxHints instructionLimit afm_parse_kern_data CF2_HintMaskRec_ dsMove ps_table_done CF2_HintMove cf2_builder_cubeTo cf2_getBlueValues cf2_arrstack_finalize CF2_HintMoveRec PSaux_Err_Invalid_Stream_Seek CF2_NumberInt op_rrcurveto PSaux_Err_Raster_Overflow cf2_cmdHHCURVETO CF2_GlyphPathRec_ CF2_Err_Missing_Startfont_Field AFM_TOKEN_ITALICANGLE AFM_TOKEN_C CF2_Err_Post_Table_Missing CF2_Blues AFM_TOKEN_L cond2 AFM_TOKEN_N PSaux_Err_Invalid_Post_Table PSaux_Err_Stack_Underflow arrstack AFM_TOKEN_STARTAXIS cf2_arrstack_push t1_cmap_unicode_char_index PSaux_Err_Debug_OpCode AFM_TOKEN_ENDCOMPOSITES AFM_TOKEN_METRICSSETS cf2_glyphpath_closeOpenPath cf2_escRESERVED_8 CF2_HintMask shared_vals cf2_free_instance dummyWidth cf2_escSETCURRENTPT prevP0 cff_decoder_init xOffset1 xOffset3 ps_parser_to_fixed afm_parser_read_int elemIsQueued Unexpected_OtherSubr cf2_outline_init PSaux_Err_Missing_Fontboundingbox_Field AFM_TOKEN_ENDAXIS ps_builder_funcs PS_Conv_EexecDecode CF2_Err_Stack_Underflow PSaux_Err_DEF_In_Glyf_Bytecode afm_compare_kern_pairs secondHintEdge AFM_STREAM_STATUS_EOL stemWidthPer1000 bchar_index cf2_cmdHLINETO CF2_Locked cf2_cmdHINTMASK CF2_Err_Invalid_Stream_Handle outerTransform AFM_TOKEN_CHARACTERSET cf2_setError AFM_TOKEN_BLENDDESIGNMAP in_charstring_type CF2_ArrStackRec_ ps_builder_init PSaux_Err_Could_Not_Find_Context AFM_TOKEN_ENCODINGSCHEME yOffset3 CF2_Err_Invalid_Horiz_Metrics t1_builder_done glyphpath boost cf2_hintmap_isValid PSaux_Err_Too_Many_Caches hintmap cf2_stack_pop maskByte CF2_Err_Invalid_Post_Table_Format CF2_BufferRec_ CF2_GlyphPath op_callothersubr reverseWinding PSaux_Err_Invalid_Pixel_Size cf2_cmdHSBW hintOriginY AFM_TOKEN_ISFIXEDPITCH windingMomentum AFM_TOKEN_ENDKERNPAIRS decimal iSrc AFM_TOKEN_ENDKERNDATA cff_builder_done cf2_computeDarkening downMoveUp cf2_hintmap_init cf2_blues_init CF2_Err_Invalid_Glyph_Index reallocate_t1_table CF2_RenderingFlags PSaux_Err_Too_Few_Arguments op_dotsection CF2_Err_Invalid_Library_Handle psaux_driver_class upMinCounter AFM_TOKEN_WEIGHTVECTOR CF2_Err_Unknown_File_Format innerTransform maskPtr cf2_getBlueMetrics AFM_VALUE_TYPE_BOOL op_setcurrentpoint PSaux_Err_Raster_Negative_Height PS_Conv_Strtol cf2_hint_isBottom PS_Conv_ASCIIHexDecode cf2_stack_count AFM_TOKEN_ISBASEFONT doingSeac cf2_doBlend ps_parser_to_bytes cf2_getUnitsPerEm cf2_builder_moveTo CF2_StackRec_ isCFF2 AFM_TOKEN_STARTFONTMETRICS cf2_getPpemY opIdx PSaux_Err_Invalid_Stream_Operation cf2_initGlobalRegionBuffer CF2_Err_Too_Many_Hints CF2_OutlineCallbacksRec_ cff_builder_close_contour iDst stemHint cf2_hint_isSynthetic ps_builder_check_points CF2_Err_Invalid_Frame_Read PSaux_Err_Invalid_CodeRange t1_cmap_custom_class_rec PSaux_Err_Nested_Frame_Access CF2_Err_Unimplemented_Feature blueValues cf2_hintmask_getMaskPtr cf2_glyphpath_lineTo prevElemP0 prevElemP3 cf2_escDROP code_to_sid cf2_cmdVVCURVETO CF2_ICF_Top t1_cmap_unicode_done CF2_NumberType FT_UFast CF2_Err_Invalid_CodeRange CF2_Err_Raster_Uninitialized CF2_PathOp_ numElements embed PSaux_Err_Invalid_Size_Handle minDS indexStemHint cf2_cmdCLOSEPATH CF2_Err_Locations_Missing CF2_Font cf2_freeT1SeacComponent PSaux_Err_Too_Many_Drivers PSaux_Err_Too_Many_Hints opStack CF2_Err_Invalid_Outline cf2_cmdVSTEM cf2_getVStore CF2_ArrStack /home/computerfido/Desktop/LemonTest/lemon-freetype/src/psaux/psaux.c op_rmoveto PSaux_Err_Invalid_Library_Handle CF2_Err_Nested_Frame_Access CF2_Err_Missing_Size_Field CF2_Err_Table_Missing csBottomEdge ps_builder_add_point AFM_TOKEN_STARTKERNPAIRS0 cf2_escVSTEM3 CF2_Err_Divide_By_Zero initial_map_ready csFuzz CF2_Stack PSaux_Err_Cannot_Open_Stream cf2_glyphpath_hintPoint csUnitsPerPixel stemHintArray cf2_arrstack_getPointer cf2_glyphpath_moveTo t1builder T1_CMap_ClassesRec cf2_escHSTEM3 T1_CMapCustomRec_ cf2_arrstack_size CF2_Err_CMap_Table_Missing is_expert CF2_Err_Invalid_Character_Code CF2_OutlineCallbacks metrics_sets cf2_initLocalRegionBuffer op_pop cf2_stack_getReal t1_builder_start_point no_stem_darkening_driver cf2_cmdHSTEM cf2_cmdEXTENDEDNMBR AFM_Token_ PSaux_Err_Invalid_Character_Code numOtherBlues CF2_Err_Syntax_Error cf2_hintmask_read AFM_TOKEN_BLENDDESIGNPOSITIONS AFM_TOKEN_ENDCHARMETRICS PSaux_Err_Invalid_Table num_elements start_idx callbacks AFM_TOKEN_KPH AFM_TOKEN_KPX AFM_TOKEN_KPY afm_parse_track_kern PSaux_Err_Invalid_Version CF2_Err_Stack_Overflow lastVal CF2_Err_Invalid_CharMap_Handle ps_parser_skip_PS_token PS_Conv_ToFixed op_hstem3 CF2_Err_Missing_Encoding_Field prevElemOp AFM_TOKEN_ENDDIRECTION CF2_Err_Bad_Argument cff_decoder_prepare CF2_Err_Name_Table_Missing t1_decoder cf2_getStdHW t1_cmap_custom_char_index ps_parser_to_coord_array cf2_getFamilyBlues PSaux_Err_Missing_Font_Field cf2_getFamilyOtherBlues CF2_Err_Could_Not_Find_Context PSaux_Err_Invalid_Cache_Handle cf2_cmdRLINECURVE fractionalTranslation counterHintMap CF2_HintMoveRec_ initialMap t1_decoder_init op_sbw CF2_OutlineRec_ prevP1 CF2_MAX_HINT_EDGES old_cur PSaux_Err_Max cf2_interpT2CharString cf2_cmdVLINETO CF2_OutlineRec N_AFM_TOKENS ft_char_table syntheticEmboldeningAmountX syntheticEmboldeningAmountY CF2_Err_Invalid_Slot_Handle PSaux_Err_Invalid_Stream_Skip acur AFM_TOKEN_UNDERLINEPOSITION old_base factor1 t1_builder_init AFM_TOKEN_FULLNAME cff_builder_add_contour useIntersection op_hmoveto AFM_TOKEN_CHARWIDTH AFM_ValueRec PSaux_Err_Ok CF2_Err_Missing_Bbx_Field psaux_interface cf2_cmdVMOVETO cf2_cmdCALLSUBR op_vlineto cf2_hint_isLocked cf2_escRESERVED_38 AFM_TOKEN_TRACKKERN counterMask flexStore scaledStem PSaux_Err_Out_Of_Memory AFM_TOKEN_ISFIXEDV hintMap ps_builder_add_point1 newSize downMoveDown CF2_Err_Invalid_Cache_Handle AFM_VALUE_TYPE_NAME CF2_CallbackParamsRec CF2_Err_Hmtx_Table_Missing cf2_escPOP cf2_cmdRETURN PSaux_Err_Missing_Property CF2_PathOpMoveTo cf2_escRESERVED_13 readFromStack AFM_TOKEN_ENDFONTMETRICS PSaux_Err_Invalid_Driver_Handle cf2_cmdRMOVETO PS_Conv_ToInt T1_Operator_ csTopEdge gr_idx cf2_escSQRT CF2_Err_Missing_Bitmap op_callsubr PSaux_Err_Ignore newHintMap t1_cmap_custom_char_next cf2_outline_close CF2_Err_Missing_Property newPtr miterLimit cf2_getMaxstack cf2_escDOTSECTION AFM_TOKEN_KP cf2_escINDEX CF2_Err_Too_Many_Drivers prevElemP1 cf2_cmdHSTEMHM scaleC CF2_Err_Raster_Corrupted PSaux_Err_Array_Too_Large CF2_HintMapRec_ op_rlineto cf2_stack_init free_callback CF2_Err_Raster_Overflow cf2_escRESERVED_25 byteCount CF2_Err_Invalid_Glyph_Format PSaux_Err_Too_Many_Extensions max_bytes achar cf2_escFLEX AFM_TOKEN_ESCCHAR CF2_CallbackParamsRec_ afm_parser_init CF2_StemHintRec cf2_escSUB summand2 cf2_arrstack_setCount cf2_doFlex CF2_Err_Invalid_Frame_Operation t1_decoder_parse_metrics cff_compute_bias PSaux_Err_Invalid_Handle cf2_glyphpath_init afm_parser_skip_section CF2_Matrix CF2_HintMap cf2_buf_readByte cf2_stack_pushInt CF2_StemHint PSaux_Err_Corrupted_Font_Glyphs moveIsPending numFamilyOtherBlues CF2_Err_Cannot_Render_Glyph cf2_escRESERVED_31 CF2_PathOpCubeTo translation isHFlex PSaux_Err_CMap_Table_Missing CF2_Err_Nested_DEFS PSaux_Err_Horiz_Header_Missing PSaux_Err_Invalid_Stream_Handle cf2_getDefaultWidthX quadTo sid_to_string ps_parser_done PSaux_Err_Unlisted_Object delimiters CF2_BlueRec afm_parser_done t1_cmap_expert_class_rec cf2_glyphpath_finalize hintOrigin hasVariations CF2_HintRec_ AFM_TOKEN_BLENDAXISTYPES boldenX CF2_Err_DEF_In_Glyf_Bytecode nextP0 midpoint cf2_glyphpath_pushMove AFM_TOKEN_STDHW fieldrec CF2_Err_Array_Too_Large AFM_TOKEN_CHARACTERS dividend PSaux_Err_Invalid_Glyph_Format cf2_getWindingMomentum AFM_TOKEN_FONTBBOX pnum_bytes pnum_tokens zoneHeight PSaux_Err_Invalid_File_Format savedMove CF2_Err_Invalid_Composite ps_builder_close_contour CF2_Err_Horiz_Header_Missing cff_check_points max_values stemhint CF2_Err_Unlisted_Object cond1 ps_tocoordarray afm_stream_skip_spaces Store_Integer cf2_hintmap_insertHint CF2_Err_Out_Of_Memory cf2_hintmask_isNew cf2_checkTransform cf2_escHFLEX1 AFM_TOKEN_STDVW CF2_Err_Invalid_Stream_Seek AFM_TOKEN_UNKNOWN cff_builder_add_point1 cf2_cmdHVCURVETO CF2_Err_Invalid_Size_Handle AFM_TOKEN_B needExtraSetup cf2_escOR CF2_ArrStackRec advWidth boldenAmount t1_args_count CF2_Err_Too_Few_Arguments stemDarkened CF2_OutlineCallbacksRec subrStack firstHintEdge integral cf2_arrstack_getBuffer bchar ps_parser_to_token maxScale hintMoves PSaux_Err_Raster_Uninitialized ps_decoder AFM_TOKEN_AXISLABEL minuend AFM_TOKEN_ENDTRACKKERN AFM_TOKEN_UNDERLINETHICKNESS CF2_FontRec_ cf2_escRESERVED_32 cff_lookup_glyph_by_stdcharcode cf2_escSBW cf2_getStdVW cf2_cmdENDCHAR PSaux_Err_Invalid_Opcode lenNormalizedV PSaux_Err_Stack_Overflow afm_tokenize PSaux_Err_No_Unicode_Glyph_Name PSaux_Err_Missing_Startfont_Field cf2_stack_setReal suppressOvershoot op_vstem AFM_STREAM_STATUS_EOF CF2_Err_Raster_Negative_Height CF2_Err_No_Unicode_Glyph_Name CF2_HintMapRec AFM_TOKEN_DESCENDER AFM_ValueRec_ CF2_CallbackParams upMoveUp PSaux_Err_Post_Table_Missing ps_parser_init pathIsOpen PSaux_Err_Invalid_CharMap_Handle PSaux_Err_Code_Overflow T1_Operator AFM_VALUE_TYPE_INDEX CF2_Err_Invalid_Driver_Handle byte2 cf2_escHFLEX numFamilyBlues cf2_setGlyphWidth darken PSaux_Err_Divide_By_Zero lastIndex cf2_escAND indexInsert isT1 op_return op_vstem3 byte4 CF2_Err_Invalid_File_Format CF2_Err_Too_Many_Function_Defs AFM_Value CF2_Err_Execution_Too_Long CF2_Frac CF2_F16Dot16 CF2_Err_Cannot_Open_Stream AFM_TOKEN_VV byte3 AFM_TOKEN_W0 AFM_TOKEN_W1 AFM_TOKEN_ASCENDER CF2_Err_Invalid_Argument ps_parser_load_field t1_cmap_unicode_init PSaux_Err_Invalid_CharMap_Format cf2_glyphpath_pushPrevElem cf2_hintmap_adjustHints hasWidthArg PSaux_Err_Invalid_Frame_Read subr_no idx2 T1_CMapCustom AFM_TOKEN_WX AFM_TOKEN_WY byte1 CF2_HintMaskRec cf2_freeSeacComponent PSAux_ServiceRec CF2_Err_Missing_Fontboundingbox_Field cf2_cmdRCURVELINE t1_cmap_custom_done cf2_cmdRESERVED_2 t1_cmap_standard_class_rec firstHintMap prevElemP2 t1_cmap_std_done numBlueValues CF2_BluesRec_ PSaux_Err_Missing_Encoding_Field PSaux_Err_Invalid_Outline CF2_GlyphPathRec cf2_getLanguageGroup no_stem_darkening_font op_none cf2_escNEG PSaux_Err_Too_Many_Function_Defs skip_comment afm_parser_next_key PSaux_Err_Invalid_Composite saveEdge skip_string emBoxTopEdge t1_builder_add_point AFM_STREAM_STATUS_EOC AFM_ValueType_ max_tokens alternate op_vmoveto CF2_Synthetic cf2_hintmask_setAll AFM_TOKEN_FAMILYNAME AFM_TOKEN_STARTCHARMETRICS PSaux_Err_Invalid_Offset cf2_getSubfont CF2_Err_Invalid_Post_Table cf2_decoder_parse_charstrings offsetStart0 cf2_stack_roll PSaux_Err_Missing_Size_Field No_Width CF2_ICF_Bottom cf2_doStems dsFlatEdge achar_index op_seac divider CF2_Hint lastSubfont PSaux_Err_Bbx_Too_Big cf2_hintmask_isValid moveDown CF2_PathOpLineTo maxDS PSaux_Err_Invalid_Horiz_Metrics AFM_TOKEN_STARTDIRECTION minDiff PSaux_Err_Invalid_Face_Handle PSaux_Err_Invalid_Stream_Read cf2_hintmask_setNew ps_tofixedarray AFM_TOKEN_MAPPINGSCHEME cffbuilder cf2_cmdRRCURVETO cf2_escSEAC cf2_glyphpath_computeOffset cf2_hint_initZero cf2_escEQ t1_builder_add_point1 AFM_STREAM_STATUS_NORMAL max_coords cf2_escEXCH CF2_Err_Max yOffset1 AFM_TOKEN_PCC cf2_cmdESC AFM_TOKEN_STARTTRACKKERN halfWidth dsNew bottomZone CF2_Err_Invalid_Stream_Skip AFM_TOKEN_VERSION CF2_NumberFixed PSaux_Err_Invalid_Vert_Metrics cf2_font_setup afm_parser_read_vals cf2_arrstack_setNumElements hintMask op_hvcurveto t1_cmap_unicode_class_rec subrNum T1_CMapStdRec_ CF2_Err_Invalid_Table darkenParams lastIsX cf2_hint_isTop t1_builder_close_contour cf2_escABS lastError cf2_escROLL CF2_Err_Invalid_Pixel_Size ps_builder_start_point cf2_stack_free blueScale glyphPath boldenY new_root hintMove cf2_escIFELSE CF2_Err_Ok maxZoneHeight t1_builder_check_points currentTransform cf2_hintmap_map cf2_cmdRESERVED_0 cf2_escRESERVED_19 CF2_StemHintRec_ ps_builder PSaux_Err_Nested_DEFS arg_cnt num_limit AFM_TOKEN_STARTKERNPAIRS CF2_Err_Invalid_Stream_Operation CF2_Err_Invalid_Reference downMinCounter cf2_outline_reset CF2_Err_Invalid_Vert_Metrics cf2_getNormalizedVector afm_parser_parse large_int CF2_Err_Too_Many_Caches nominalWidthX shift_elements cf2_escCALLOTHERSUBR cf2_getSeacComponent AFM_TOKEN_W1Y CF2_Err_Invalid_Offset CF2_BlueRec_ CF2_Err_ENDF_In_Exec_Stream AFM_TOKEN_ISCIDFONT unitsPerEm PSaux_Err_Unimplemented_Feature op_max darkened fracDown op_unknown15 cf2_hint_init CF2_Err_Lower_Module_Version cf2_stack_popFixed hinted nextP1 cf2_getGlyphOutline CF2_PairTop CF2_GhostBottom offsetStart1 t1_cmap_std_char_next tempHintMask PSaux_Err_Invalid_Frame_Operation totalSize CF2_Err_Ignore CF2_Err_Invalid_PPem familyOtherBlues CF2_Buffer AFM_TOKEN_WEIGHT cf2_blues_capture op_closepath component cff_builder_init cf2_escADD PSaux_Err_Hmtx_Table_Missing cf2_escDIV AFM_TOKEN_W t1_decoder_done PSaux_Err_Locations_Missing ps_parser_to_token_array cf2_arrstack_clear stemWidth blueShift csCoord t1_cmap_unicode_char_next PSnames_Err_Invalid_CodeRange pscmaps_services NextIter PSnames_Err_Unknown_File_Format PSnames_Err_Unimplemented_Feature pscmaps_interface PSnames_Err_Too_Many_Extensions compare_uni_maps PSnames_Err_Invalid_PPem ft_adobe_glyph_list PSnames_Err_Syntax_Error PSnames_Err_Invalid_Post_Table ps_get_macintosh_name PSnames_Err_Too_Many_Function_Defs t1_standard_encoding PSnames_Err_Name_Table_Missing /home/computerfido/Desktop/LemonTest/lemon-freetype/src/psnames/psnames.c PSnames_Err_Nested_DEFS PSnames_Err_Invalid_Slot_Handle PSnames_Err_Glyph_Too_Big PSnames_Err_Ignore PSnames_Err_Corrupted_Font_Glyphs PSnames_Err_Invalid_Composite ft_extra_glyph_names ft_sid_names ft_standard_glyph_names PSnames_Err_Missing_Chars_Field PSnames_Err_No_Unicode_Glyph_Name PSnames_Err_Corrupted_Font_Header PSnames_Err_Code_Overflow PSnames_Err_Invalid_Post_Table_Format PSnames_Err_Too_Many_Hints PSnames_Err_Missing_Bbx_Field PSnames_Err_Bbx_Too_Big PSnames_Err_Cannot_Open_Resource PSnames_Err_Missing_Module map1 map2 ft_extra_glyph_unicodes PSnames_Err_Invalid_Version PSnames_Err_Invalid_Argument PSnames_Err_Invalid_Vert_Metrics PSnames_Err_Invalid_Frame_Read PSnames_Err_Invalid_Reference PSnames_Err_Missing_Encoding_Field PSnames_Err_Out_Of_Memory free_glyph_name PSnames_Err_Too_Many_Instruction_Defs PSnames_Err_Invalid_Stream_Seek PSnames_Err_Raster_Negative_Height PSnames_Err_Post_Table_Missing ft_mac_names PSnames_Err_Missing_Startchar_Field PSnames_Err_Max PSnames_Err_Invalid_Offset PSnames_Err_Missing_Startfont_Field PSnames_Err_Ok PSnames_Err_Stack_Overflow NotFound PSnames_Err_Bad_Argument PSnames_Err_Invalid_Stream_Operation PSnames_Err_CMap_Table_Missing PSnames_Err_Unlisted_Object PSnames_Err_Invalid_Handle PSnames_Err_Invalid_File_Format PSnames_Err_Invalid_Library_Handle PSnames_Err_Nested_Frame_Access PSnames_Err_Invalid_Pixel_Size PSnames_Err_Missing_Bitmap PSnames_Err_Invalid_Opcode FT_Service_PsCMapsRec PSnames_Err_Invalid_Size_Handle unicode1 PSnames_Err_Raster_Corrupted PSnames_Err_Missing_Font_Field PSnames_Err_DEF_In_Glyf_Bytecode PSnames_Err_Invalid_Glyph_Index PSnames_Err_Invalid_Table PSnames_Err_Lower_Module_Version PSnames_Err_Invalid_CharMap_Handle ft_extra_glyph_name_offsets psnames_get_service ps_unicodes_char_index PSnames_Err_Divide_By_Zero ps_unicode_value PSnames_Err_Array_Too_Large PSnames_Err_Invalid_Glyph_Format PSnames_Err_Could_Not_Find_Context unicode2 PSnames_Err_Invalid_Horiz_Metrics PSnames_Err_Invalid_Character_Code PSnames_Err_Too_Many_Drivers PSnames_Err_Invalid_Frame_Operation PSnames_Err_Cannot_Open_Stream PSnames_Err_Table_Missing PSnames_Err_Invalid_CharMap_Format PSnames_Err_Invalid_Face_Handle PSnames_Err_Missing_Fontboundingbox_Field ps_check_extra_glyph_unicode ft_get_adobe_glyph_index PSnames_Err_Horiz_Header_Missing extra_glyphs PSnames_Err_Invalid_Stream_Skip PSnames_Err_Stack_Underflow PSnames_Err_Execution_Too_Long PSnames_Err_Missing_Property PSnames_Err_Invalid_Stream_Read PSnames_Err_Missing_Size_Field PSnames_Err_Hmtx_Table_Missing PSnames_Err_Locations_Missing PSnames_Err_Invalid_Stream_Handle ps_unicodes_char_next uni_char PSnames_Err_Raster_Overflow PSnames_Err_Too_Few_Arguments ps_unicodes_init ps_get_standard_strings PSnames_Err_Debug_OpCode extra_glyph_list_states PSnames_Err_Cannot_Render_Glyph PSnames_Err_Invalid_Cache_Handle t1_expert_encoding PSnames_Err_Too_Many_Caches PSnames_Err_Invalid_Outline PSnames_Err_ENDF_In_Exec_Stream PSnames_Err_Invalid_Driver_Handle PSnames_Err_Raster_Uninitialized ps_check_extra_glyph_name malloc ft_ansi_stream_close fseek /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base/ftsystem.c ft_realloc fopen ft_alloc fread fclose ft_free ftell ft_ansi_stream_io ft_debug_init /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base/ftdebug.c FT_Trace_Get_Count FT_Trace_Get_Name source_lly source_ury ft_bitmap_assure_buffer source_offset_ target_pitch_sign xstr source_llx bit_last source_urx source_ /home/computerfido/Desktop/LemonTest/lemon-freetype/src/base/ftbitmap.c atarget_offset target_llx target_lly target_ury xStrength limit_r final_llx final_rows yStrength target_size FT_Bitmap_Copy final_width FT_Bitmap_Embolden source_pitch_sign final_lly final_urx final_ury null_bitmap limit_p ft_gray_for_premultiplied_srgb_bgra free_source_bitmap FT_Bitmap_Blend target_urx FT_GlyphSlot_Own_Bitmap FT_Bitmap_New new_pitch ypixels xpixels old_target_pitch ystr free_target_bitmap_on_error                       �      �       U�      �       �U��      �       U                  �      �       S                          �      �       U�      H       \H      K       �U�K      q       \q      t       �U�                                     P      J       ]J      W       PW      Z       ]                        �             P             SK      Z       SZ      n       P                        4       V                                 
 ��F     �      '       S'      ,       sx�,      4       S                        @       J        UJ       �       S�      �       �U��      �       S                  V       j        P                                  _       �        P�       �        T�       /       R/      �       V�      �       P�      �       P�      �       T�      �       R�      �       V                        �       (       T(      }       R�      �       T�      �       R                                    �       �        Q�       �        U�       �        Q�       �        0��       �        P�       �        U      
       P(      /       0�/      @       P@      D       TW      \       P                                      U       2        V2       3        �U�                                    
 ��F     �               S       $        sx�$       1        S                      `�      w�       Uw�      ��       �U���      ��       U                            `�      ~�       T~�      ��       V��      ��       �T���      ��       V��      ��       �T���      ��       T                            `�      ~�       Q~�      ��       \��      ��       �Q���      ��       \��      ��       �Q���      ��       Q                        w�      ~�       U~�      ��       S��      ��       U��      ��       U                     `�      ��       0���      ��       P��      ��       0�                    ~�      ��       S��      ��       S                    ��      Ӷ       PԶ      ޶       P                      �      3�       U3�      7�       u�7�      _�       U                    �      7�       T7�      _�       T                    �      "�       Q"�      K�       �Q�                        е      �       U�      ��       V��      �       U�      �       �U�                        е      �       T�      ��       S��      �       T�      �       �T�                        е      ׵       Q׵      ��       \��      �       R�      �       �Q�                  �      �       Q                        P�      m�       Um�      ��       �U���      ��       U��      ǵ       �U�                            P�      k�       Tk�      }�       ]}�      ��       �T���      ��       ]��      ��       T��      ǵ       ]                            P�      m�       Qm�      ��       V��      ��       �Q���      ��       V��      ��       Q��      ǵ       V                            P�      m�       Rm�      ��       \��      ��       �R���      ��       \��      ��       R��      ǵ       \                 P�      ǵ       ��                              P�      m�       Qm�      ��       V��      ��       �Q���      ��       V��      ��       Q��      ǵ       V                       P�      m�       Um�      ��       �U���      ��       U��      ǵ       �U�                         P�      q�       0�q�      }�       P��      ��       P��      ��       0���      ǵ       P                                  ��      ��       U��      �       Z�      %�       �U�%�      a�       Za�      t�       �U�t�      ��       Z��      ��       �U���      ��       Z��      Ս       �U�                                ��      �       T�      %�       �T�%�      Y�       TY�      t�       �T�t�      ��       T��      ��       �T���      ��       T��      Ս       �T�                                  ��      ��       Q��      �       U�      %�       �Q�%�      \�       U\�      t�       �Q�t�      ��       U��      ��       �Q���      ��       U��      Ս       �Q�                            ��      �       R�      %�       �R�%�      J�       RJ�      t�       �R�t�      ��       R��      Ս       �R�                                    ��      �       X�      a�       Xa�      l�       �X�l�      t�       Pt�      ��       X��      ��       �X���      ��       S��      ��       P��      ��       X��      Ս       w                                   ��      �       Y�      %�       �Y�%�      a�       Ya�      t�       w t�      ��       Y��      ��       w ��      ��       �`��      ��       Y��      Ս       �h                             ��      �       0��      $�       S$�      %�       y %�      ��       0���      ��       S��      ��       y ��      Ս       0�                  ��      Ս       P                   t�      ��       X��      ��       �X�                   t�      ��       Z��      ��       �U�                    ��      	�       U	�      X�       �U�                          ��      	�       T	�      �       V�      3�       �T�3�      H�       VH�      X�       �T�                        ��      	�       Q	�      2�       ^2�      3�       �Q�3�      X�       ^                          ��      	�       R	�      �       S�      3�       �R�3�      ;�       S;�      X�       �R�                            ��      	�       X	�      �       �X��      �       P�      0�       ]0�      3�       P3�      X�       ]                        ��      ��       Y��      .�       \.�      3�       �Y�3�      X�       \                        �n      �n       U�n      �n       �U��n      �n       U�n      �n       �U�                            �n      �n       T�n      �n       S�n      �n       �T��n      �n       S�n      �n       T�n      �n       S                          �n      �n       Q�n      �n       V�n      �n       �Q��n      �n       Q�n      �n       V                 �n      �n       ���                              �n      �n       T�n      �n       S�n      �n       �T��n      �n       S�n      �n       T�n      �n       S                       �n      �n       U�n      �n       �U��n      �n       U�n      �n       �U�                         �n      �n       0��n      �n       P�n      �n       0��n      �n       P�n      �n       R                  fn      �n       P                      0n      Gn       UGn      Hn       �U�Hn      Qn       U                        0n      ;n       T;n      Gn       u Gn      Hn       �T�Hn      Qn       T                      0n      Gn       QGn      Hn       �Q�Hn      Qn       Q                        Pm      |m       U|m      �m       �U��m      �m       U�m      "n       �U�                          Pm      �m       T�m      �m       S�m      �m       �T��m      �m       T�m      "n       S                          Pm      �m       Q�m      �m       V�m      �m       �Q��m      �m       Q�m      "n       V                      �m      �m       P�m      �m       \�m      "n       \                           �m      �m       U�m      �m       w �m      �m       U�m      �m       U�m      �m       u ��m      n       u �ɚ�r@J$" %�n      n       w �ɚ�r@J$" %�n      n       U                  �m      �m       1��m      �m       1��m      n       	��                          0l      xl       Uxl      �l       �U��l      �l       U�l      m       �U�m      #m       U                          �l      �l       P�l      �l       S�l      �l       s ��l      �l       r ��l      m       S                           �l      �l       Q�l      �l       u �l      �l       Q�l      �l       Q�l      �l       q ��l      �l       q �ɚ�r@J$" %��l      �l       u �ɚ�r@J$" %��l      �l       Q                  �l      �l       1��l      �l       1��l      �l       	��                            �j      k       Uk      �k       S�k      �k       �U��k      l       Sl      l       �U�l      !l       U                        �j      k       Tk      &k       Z&k      l       �T�l      !l       T                        "k      &k       P&k      �k       V�k      l       Vl      l       R                 rk      �k       1v$�                           +k      =k       Q=k      Mk       u Mk      Mk       T�k      �k       Q�k      �k       q ��k      �k       q �ɚ�r@J$" %��k      �k       u �ɚ�r@J$" %��k      �k       T                  +k      Mk       1��k      �k       1��k      �k       	��                         Mk      _k       Q_k      jk       �`jk      jk       Q�k      �k       Q�k      �k       q ��k      �k       q �ɚ�r@J$" %��k      �k       �`�ɚ�r@J$" %��k      �k       Q                 Mk      jk       1��k      �k       1��k      �k       	��                      pj      �j       U�j      �j       u �j      �j       �U�                      pj      �j       T�j      �j       t �j      �j       �T�                      �i      �i       U�i      j       Qj      nj       �U�                      j      ;j       P;j      @j       R@j      ij       u                      j      .j       1�.j      3j       	��3j      =j       T=j      @j       t �@j      ij       T                 j      Qj       Q                        &j      ;j       P;j      @j       R@j      Ej       PEj      ij       R                    \j      ij       Pij      nj       q �                 \j      ij       P                      �i      �i       U�i      �i       T�i      �i       �U�                      �i      �i       U�i      �i       T�i      �i       �U�                  �i      �i       W                      �i      �i       U�i      �i       T�i      �i       �U�                      �i      �i       U�i      �i       T�i      �i       �U�                  �i      �i       W                            �f      g       Ug      |g       V|g      �g       �U��g      i       Vi      6i       U6i      �i       V                          �f      �f       T�f      g       s|��g      �g       s|��h      �h       Si      i       Si      6i       T                            �f      g       Qg      ~g       \~g      �g       �Q��g      i       \i      6i       Q6i      �i       \                              g      7g       0�7g      Yg       PYg      ^g       �L�g      �g       0��g      �h       0��h      �h       P�h      i       0�6i      �i       0�                          �f      g       0�g      �g       ]�g      �g       ]�g      �h       ]�h      �h       1��h      i       ]i      6i       0�6i      �i       ]                                           g      7g       Q�g      �g       Q�g      �g       q��g      h       Qh      h       q�h      0h       Q0h      8h       q�8h      =h       Q=h      Hh       q�Hh      Qh       QQh      `h       q�`h      xh       Qxh      �h       q��h      �h       Q�h      �h       q��h      �h       Q�h      i       Qi      i       X6i      [i       Qbi      �i       Q�i      �i       Q                                 �g      �g       P�g      �g       P)h      0h       P2h      =h       PLh      Qh       Psh      xh       P�h      �h       P�h      �h       P�h      i       P                         �g      �g       8��g      �g       R)h      0h       8�2h      =h       0�Lh      Qh       0�sh      xh       @��h      �h       @��h      �h       H�                        �g      �g       R�h      i       R6i      Pi       s~�
��| "�bi      ni       s~�
��| "��i      �i       s~�
��| "�                          g      7g       s}���i      i       s}���6i      Pi       s}���bi      ni       s}����i      �i       s}���                 <g      vg       V                 Cg      Yg       v8                  Gg      Yg       T                  Gg      Yg       v8                        Pf      �f       U�f      �f       S�f      �f       �U��f      �f       S                            Pf      cf       Tcf      �f       V�f      �f       �T��f      �f       V�f      �f       �T��f      �f       V                       Pf      �f       0��f      �f       Q�f      �f       q��f      �f       0��f      �f       s t "��f      �f       Q                     Pf      �f       0��f      �f       P�f      �f       0�                        �c      $d       U$d      Gd       SGd      `d       �U�`d      ld       S                            �c      d       Td      Hd       VHd      Id       �T�Id      _d       V_d      `d       �T�`d      ld       V                       �c      4d       0�4d      4d       Q4d      :d       q�Id      `d       0�`d      hd       s t "�hd      ld       Q                     �c      :d       0�:d      Id       PId      ld       0�                        `c      �c       U�c      �c       S�c      �c       �U��c      �c       S                            `c      sc       Tsc      �c       V�c      �c       �T��c      �c       V�c      �c       �T��c      �c       V                       `c      �c       0��c      �c       Q�c      �c       q��c      �c       0��c      �c       s t "��c      �c       Q                     `c      �c       0��c      �c       P�c      �c       0�                        �b      c       Uc      /c       S/c      Hc       �U�Hc      \c       S                            �b      �b       T�b      0c       V0c      1c       �T�1c      Gc       VGc      Hc       �T�Hc      \c       V                       �b      c       0�c      c       Qc      "c       q�1c      Hc       0�Hc      Xc       s t "�Xc      \c       Q                     �b      "c       0�"c      1c       P1c      \c       0�                        _      D_       UD_      o_       So_      �_       �U��_      �_       S                            _      #_       T#_      p_       Vp_      q_       �T�q_      �_       V�_      �_       �T��_      �_       V                       _      T_       0�T_      T_       QT_      b_       q�q_      �_       0��_      �_       s t "��_      �_       Q                     _      b_       0�b_      q_       Pq_      �_       0�                            �^      �^       U�^      �^       S�^      �^       �U��^      �^       S�^      �^       �U��^      _       S                            �^      �^       T�^      �^       V�^      �^       �T��^      �^       V�^      �^       �T��^      _       V                  _      _       P                    t^      �^       Q�^      �^       q��^      �^       Q                   p^      �^       0��^      �^       P                    T^      `^       Q`^      f^       q�f^      o^       Q                   P^      j^       0�j^      o^       P                    $^      0^       Q0^      ;^       q�;^      N^       Q                    ^      I^       0�I^      N^       P                    �]       ^       Q ^      ^       q�^      ^       Q                   �]      ^       0�^      ^       P                    �]      �]       Q�]      �]       q��]      �]       Q                   �]      �]       0��]      �]       P                 �]      �]       0�                              �[      \       U\      v\       Sv\      |\       �U�|\      �\       S�\      �\       �U��\      �\       U�\      ]       S                                    �[      \       T\      w\       Vw\      |\       �T�|\      �\       T�\      �\       V�\      �\       �T��\      �\       T�\      �\       �T��\      �\       T�\      ]       V                      �[      m\       0�m\      q\       P|\      �\       0��\      �\       P�\      �\       0��\      ]       @�                       B\      S\       PS\      q\       ]�\      �\       P�\      �\       ]                 �[      \       u8                  \      )\       �Y  |\      �\       �Y  �\      �\       �Y                      \      \       T\      )\       V|\      �\       T�\      �\       V                  \      )\       0�|\      �\       0��\      �\       0��\      �\       @�                    \       \       0� \      )\       P|\      �\       0��\      �\       P�\      �\       0�                 G\      S\       T                    �[      �[       U�[      �[       �U�                      �[      �[       T�[      �[       S�[      �[       �T�                   �[      �[       u8�[      �[       P                  �[      �[       T                    �[      �[       u8�[      �[       P                       ]      0]       U0]      R]       SR]      T]       �U�                     ]      0]       T0]      T]       �T�                       ]      0]       Q0]      S]       VS]      T]       �Q�                  1]      T]       P                        @[      o[       Uo[      w[       Sw[      �[       �U��[      �[       S                            @[      m[       Tm[      o[       Qo[      �[       �T��[      �[       T�[      �[       X�[      �[       �T�                            @[      j[       Qj[      o[       Ro[      �[       �Q��[      �[       Q�[      �[       R�[      �[       �Q�                               @[      s[       0�s[      w[       V�[      �[       0��[      �[       Y�[      �[       sp ��[      �[       ss��[      �[       Q�[      �[       V                          �Z      �Z       U�Z      �Z       V�Z      [       �U�[      [       U[      -[       V                        �Z      �Z       T�Z      �Z       S�Z      [       �T�[      -[       S                        �Z      �Z       Q�Z      [       �Q�[      *[       P*[      -[       �Q�                          �Z      �Z       R�Z      �Z       ]�Z      [       �R�[      *[       R*[      -[       ]                   �Z       [       0� [      [       U�[      -[       0�                    �Z      �Z       \[      -[       \                        `�      ޳       U޳      ��       �U���      �       U�      ô       �U�                    `�      ��       T��      ô       �T�                      `�      ó       Qó      �       S�      ��       �Q���      ô       S                      ��      ޳       U޳      �       �U���      �       U�      ô       �U�                   ǳ      �       V��      ô       V                  ��      ô       \                  �      ô       ]                   1�      L�       _��      ��       _��      ��       _                   1�      L�       ]��      ��       ]��      ��       ]                  1�      L�       0���      ��       0���      ��       0�                  b�      f�      	 v �
���                  b�      f�       Q                    b�      f�       Uf�      g�       ]                 s�      ��       v                 s�      ��       \                        �      @�       U@�      w�       �U�w�      ��       U��      Q�       �U�                    �      (�       T(�      Q�       �T�                        �      $�       Q$�      h�       Vh�      w�       �Q�w�      Q�       V                 f�      h�       0�                       �      @�       U@�      h�       �U�w�      ��       U��      Q�       �U�                    +�      h�       Sw�      Q�       S                  ��      Q�       \                  ��      Q�       ]                   ��      ۲       _
�      �       _C�      C�       _                   ��      ۲       ]
�      �       ]C�      C�       ]                  ��      ۲       0�
�      �       0�C�      C�       0�                  �      ��       R                  �      ��       s                    �      ��       U��      ��       ]                 �      '�       s                 �      (�       \                          @o      To       UTo      �o       S�o      �o       �U��o      �o       S�o      
p       �U�                            @o      do       Tdo      �o       V�o      �o       T�o      �o       �T��o      p       Vp      
p       �T�                          @o      do       Qdo      �o       \�o      �o       �Q��o      p       \p      
p       �Q�                           @o      �o       0��o      �o       P�o      �o       S�o      �o       P�o      �o       S�o      p       P                      �o      �o       P�o      �o       ]�o      �o       P                  �o      �o       V�o      �o       V                  po      �o       } p "�                    �s      �s       U�s      Pt       �U�                      �s      �s       T�s      �s       ���s      Pt       �T�                          �s      �s       Q�s      	t       V	t      8t       �Q�8t      Mt       VMt      Pt       �Q�                 �s      It       0�                          �s      t       Pt      t       St      t       Pt      4t       S4t      Kt       P                        �s      	t       V	t      t       �Q�8t      Mt       VMt      Pt       �Q�                    �s      t       ��  8t      Pt       ��                      �s      t       �T�8t      Pt       �T�                    �s      t       U8t      Pt       U                    �s      t       �U�8t      Pt       �U�                  �s      -t        �8t      Pt        �                t      -t       0�                t      -t       V                 t      -t       \                 t      "t       V                 "t      -t       V                 "t      -t       \                              Pt      st       Ust      �t       V�t      �t       �U��t      �t       V�t      �t       �U��t      �t       V�t      �t       �U�                    Pt      Ut       TUt      �t       �T�                      Pt      Zt       QZt      wt       Twt      �t       �Q�                              Pt      wt       Rwt      �t       ]�t      �t       �R��t      �t       ]�t      �t       �R��t      �t       ]�t      �t       �R�                              Pt      wt       Xwt      �t       ^�t      �t       �X��t      �t       ^�t      �t       �X��t      �t       ^�t      �t       �X�                            xt      �t       P�t      �t       S�t      �t       0��t      �t       S�t      �t       } �t      �t       �R�t      �t       P                      �t      �t       P�t      �t       �L�t      �t       P                      pt      �t       \�t      �t       \�t      �t       \                 �t      �t       S                 �t      �t       \                              �t      u       Uu      Ku       VKu      Ru       �U�Ru      bu       Vbu      iu       �U�iu      {u       V{u      �u       �U�                    �t      �t       T�t      �u       �T�                      �t      �t       Q�t      u       Tu      �u       �Q�                              �t      u       Ru      Ou       ]Ou      Ru       �R�Ru      fu       ]fu      iu       �R�iu      u       ]u      �u       �R�                              �t      u       Xu      Qu       ^Qu      Ru       �X�Ru      hu       ^hu      iu       �X�iu      �u       ^�u      �u       �X�                            u      -u       P-u      Au       SAu      Ru       0�Ru      au       Sau      fu       } fu      iu       �Riu      yu       P                      .u      @u       P@u      Ru       �LRu      iu       P                      u      Mu       \Ru      du       \iu      }u       \                 6u      Au       S                 6u      Au       \                    p      'p       U'p      Tp       �U�                    p      p       Tp      Tp       �T�                      p      p       Qp      +p       T+p      Tp       �Q�                          p      +p       R+p      Dp       VDp      Ep       �R�Ep      Sp       VSp      Tp       �R�                          p      +p       X+p      Cp       SCp      Ep       �X�Ep      Rp       SRp      Tp       �X�                        ,p      7p       P7p      Dp       v Dp      Ep       �REp      Qp       P                 p      p       u                     `p      wp       Uwp      �p       �U�                    `p      dp       Tdp      �p       �T�                      `p      ip       Qip      {p       T{p      �p       �Q�                          `p      {p       R{p      �p       V�p      �p       �R��p      �p       V�p      �p       �R�                          `p      {p       X{p      �p       S�p      �p       �X��p      �p       S�p      �p       �X�                        |p      �p       P�p      �p       v �p      �p       �R�p      �p       P                 `p      ap       u                         @q      Hq       UHq      �q       _�q      �q       �U��q      �q       _                    @q      fq       Tfq      �q       �T�                        @q      fq       Qfq      �q       \�q      �q       �Q��q      �q       \                        @q      fq       Rfq      �q       ^�q      �q       �R��q      �q       ^                        @q      fq       Xfq      �q       ]�q      �q       �X��q      �q       ]                     @q      �q       0��q      �q       P�q      �q       P                 gq      �q                              gq      �q       P�q      �q       S�q      �q       S                        �p      �p       U�p      q       _q      q       �U�q      @q       _                    �p      �p       T�p      @q       �T�                        �p      �p       Q�p      q       \q      q       �Q�q      @q       \                        �p      �p       R�p      	q       ^	q      q       �R�q      @q       ^                        �p      �p       X�p      q       ]q      q       �X�q      @q       ]                     �p      �p       0��p      �p       Pq      q       P                 �p      �p                              �p      �p       P�p      �p       Sq      !q       S                              �u      �u       U�u      �u       V�u      �u       �U��u      v       Vv      	v       �U�	v      v       Vv      "v       �U�                    �u      �u       T�u      "v       �T�                      �u      �u       Q�u      �u       T�u      "v       �Q�                              �u      �u       R�u      �u       ]�u      �u       �R��u      v       ]v      	v       �R�	v      v       ]v      "v       �R�                              �u      �u       X�u      �u       ^�u      �u       �X��u      v       ^v      	v       �X�	v      !v       ^!v      "v       �X�                            �u      �u       P�u      �u       S�u      �u       0��u      v       Sv      v       } v      	v       �R	v      v       P                      �u      �u       P�u      �u       �L�u      	v       P                      �u      �u       \�u      v       \	v      v       \                 �u      �u       S                 �u      �u       \                    �e      �e       U�e      f       �U�                        �e      f       Tf      f       Uf      f       �T�f      f       T                      �e      f       Qf      f       �Q�f      f       Q                      �e      f       Rf      f       �R�f      f       R                      �e      f       Xf      f       �X�f      f       X                      �X      �X       U�X      |Y       _|Y      }Y       �U�                      �X      �X       T�X      zY       ^zY      }Y       �T�                    �X      �X       Q�X      }Y       ��                    �X      �X       R�X      }Y       �R�                      �X      �X       X�X      xY       ]xY      }Y       �X�                      �X      �X       Y�X      vY       \vY      }Y       �Y�                       �X      �X       0��X      1Y       S1Y      5Y       s�;Y      `Y       S`Y      dY       s�                 �X      Y       0�RY      RY       0�                 �X      Y       ^RY      RY       ^                 �X      Y       0�RY      RY       0�                        @�      ��       U��      5�       �U�5�      B�       UB�      ��       �U�                        @�      }�       T}�      +�       S+�      5�       �T�5�      ��       S                              @�      z�       Qz�      $�       _$�      5�       �Q�5�      B�       QB�      W�       �Q�W�      ��       _��      ��       �Q�                        @�      x�       Rx�      5�       ��5�      B�       RB�      ��       ��                                @�      ��       X��      $�       ^$�      5�       �X�5�      B�       XB�      �       ^�      �       �X��      �       ^�      ��       �X�                        @�      ��       Y��      5�       �Y�5�      B�       YB�      ��       �Y�                        ��      ʗ       0�ʗ      $�       Vg�      �       V�      �       V                                 �      �       0��      ��       \��      �       \�      �       \O�      \�       0�\�      v�       Qv�      z�       q���      ��       \��      ��       0�                        ��      ��      	 p 0$0&���      $�       \I�      �       \�      �       \                      �      ��      	 p 0$0&���      �       ���0$0&�g�      ��       ���0$0&�                          ʗ      ܗ       Pܗ      �       ] �      $�       Pg�      �       ]�      �       ]                      ��      �      	 p 0$0&�g�      ��      	 p 0$0&���      �       _�      �       _                          d�      h�       Ph�      ��       u ��      5�       ��5�      B�       u B�      ��       ��                        E�      Q�       PQ�      ��       _�      �       _��      ��       _                         d�      $�       0�5�      �       0��      G�       0�G�      ��       P��      ��       0�                             d�      $�       0�5�      �       0��      ��       P��      ��       ]��      �       0��      �       ]�      �       0��      ��       ]                    d�      z�       Qz�      ��       _5�      B�       Q                    d�      }�       T}�      ��       S5�      B�       S                  d�      ��       0�5�      B�       0�                  ��      ��       _�      �       _                  ��      ��       S�      �       S                  ��      ��       0��      �       0�                   �      )�       2���      ��       2�                   �      )�       S��      ��       S                    �      U�       ^ə      ��       ^                        �      ��       Sə      �       S�      �       S��      ��       S                       �      ��       0�ə      �       0��      �       0���      ��       0�                   M�      w�       4��      �       4�                   M�      w�       S�      �       S                      U�      ��       ^�      �       ^��      ��       ^                      U�      ��       S�      �       S��      ��       S                     U�      ��       0��      �       0���      ��       0�                 �      ��       ]                 �      ��       ��                        �_      �_       U�_      �b       �U��b      �b       U�b      �b       �U�                                �_      �_       T�_      Db       SDb      Lb       �T�Lb      db       Sdb      nb       �T�nb      �b       S�b      �b       �T��b      �b       S                              �_      �_       Q�_      a       \a      nb       �Q�nb      b       \b      �b       �Q��b      �b       Q�b      �b       �Q�                                  �_      �_       R�_      Kb       ^Kb      Lb       �R�Lb      mb       ^mb      nb       �R�nb      �b       ^�b      �b       �R��b      �b       R�b      �b       ^                                  �_      �_       X�_      Ib       ]Ib      Lb       �X�Lb      kb       ]kb      nb       �X�nb      �b       ]�b      �b       �X��b      �b       X�b      �b       ]                :b      =b       0�                        }`      .a       U.a      b       \Lb      Zb       \nb      b       U�b      �b       \                    �`      a       Qnb      b       Q                    �`      a       Pnb      b       P                  �a      �a       T                    �a      �a       R�b      �b       R                    �a      �a       P�a      �a       p�                  b      b      	 p 0$0&�                    �_      �_       Q�_      �_       \�b      �b       Q                    �_      �_       T�_      �_       S�b      �b       S                
  �_      �_       0��b      �b       0�                 �_      �_       @�                   �_      �_       Q�_      �_       ���                   �_      �_       U�_      �_       S                  .a      Va       \Lb      Zb       \                  .a      Va       SLb      Zb       S                  .a      Va       0�Lb      Zb       0�                 wa      ~a       @�                   wa      {a       Q{a      ~a       �@�                   wa      {a       U{a      ~a       S                   �a      �a       8��b      �b       8�                   �a      �a       S�b      �b       S                    �a      b       V�b      �b       V                   �a      =b       S�b      �b       S                  �a      =b       0��b      �b       0�                   b      :b       \�b      �b       \                   b      :b       S�b      �b       S                  b      :b       0��b      �b       0�                    �W      �W       U�W      �X       X                  �W      X       T                    �W      �W       U�W      �X       X                 WX      �X       x� �                 WX      �X       Q                  TX      WX       R                 TX      WX       Q                  IX      LX       R                 IX      LX       Q                            0U      KU       UKU      �V       \�V      �V       �U��V      �V       \�V      �V       �U��V      �W       \                  0U      SU       T                              0U      7U       Q7U      qU       ^qU      �U       �Q��U      �U       ^�U      �V       �Q��V      �V       ^�V      �W       ^                    0U      <U       R<U      �W       �R�                            FU      KU       UKU      �V       \�V      �V       �U��V      �V       \�V      �V       �U��V      �W       \                     �U      �U       }d��U      �U       ^�U      yV       ^                  �U      yV       Q                   �U      TV       ~TV      yV       X                  �U      yV       P                   �U      TV       ~TV      yV       Z                   �U      TV       ~TV      yV       R                   �U      TV       ~TV      yV       Y                   �U      TV       ~TV      yV       T                 �U      TV       ~                  qU      �U       ^                   �V      �V       ^�V      �V       �Q�                   rW      �W       ^�W      �W       ^                 �W      �W       ^                  �W      �W       P                 dW      rW       ^                    CW      CW       PCW      MW       p  $0 $+( ��W      �W       P                 �W      �W       ^                      @O      �O       U�O      P       [P      �P       �U�                    �O      �O       y p ��O      �P       Z                    �O      �O       y p ��O      �P       Y                 �O      �P       V                         ;P      AP       T��AP      �P       T�^��P      �P       �^��P      �P       Q�R��P      �P       T�^�                    yP      �P       Q���P      �P       Q�R�                 �O      P       0�                 AP      bP       Q                     �O      P       0�P      bP       Q�P      �P       Q                     qO      P       0�P      �P       U�P      �P       U                  *P      �P       S                 �O      �O       T                   �O      �O       U�O      �O       [                          �P      3Q       U3Q      DQ       �U�DQ      QQ       UQQ      U       ��U      U       U                      �P      Q       TQ      ,Q       �T�U      U       T                            �P      1Q       Q1Q      3Q       P3Q      DQ       ��DQ      QQ       PQQ      U       ��U      U       Q                          lQ      �Q       ^�Q      �Q       _�Q      rT       ^rT      �T       _�T       U       ^                     lQ      �Q       0��Q      kT       ���T       U       ��                           lQ      �Q       0��Q      �Q       ^�Q      �Q       V�Q      rT       \rT      �T       ^�T       U       \                  �Q      �Q       Y                        VQ      dQ       PdQ       U       �� U      
U       P
U      U       ��                  �Q      �Q       0��0��1R      ;R      	 ����@�                           �Q      �Q       0��0���Q      GR      
 ��~���~�GR      �R      
 ��~���~��R      �R       ���~��R      rT      
 ��~���~��T       U      
 ��~���~�                                     -S      -S       U��-S      0S       U�P�0S      jS       U���~�jS      nS       U���~�nS      �S       U���S      T       P��'T      .T       �P��T      �T       U���~��T      �T       U���T      �T       �P��T      �T       U���T       U       P��                        �Q      �Q       0��Q      1R       ]1R      ;R       Z;R      �S       ]`T      �T       ]                       R      GR       Z|R      �R       ��~�R      `T       Z�T       U       Z                   �Q      �Q       0��Q       U       ��~                    �S      .T       ]�T       U       ]                       jS      nS      N w � $ &{ w � $ &{ ?&"#��@& $ &��������?&"#��@& $ &�nS      "T       w �T      �T       R�T       U       w                               �R      �S       X�S      �S       ���S      &T       X&T      .T       ���T      �T       X�T      �T       X�T       U       ��                       �Q      �Q       Y�Q      IT       SIT      MT       q�MT       U       S                  �Q       U       V                     �Q      �Q       	���Q      �R       ���R       U       ��                �R      �R       ��                �R      �R       P                 �R      �R       T�R      �R       t ��~"#���                �R      �R       t ?&�                �R      �R       �@                �R      �R       U                   �R      �R       X�R      �R      
 q x "#���                  �R      �R       x ?&��R      �R       Q                �S      �S       w                 �S      �S       ��                �S      �S       w                 �S      �S       ��                   �S      �S       P�S      �S      
 p r "#���                  �S      �S       p ?&��S      �S       R                 �S      �S       X                 �S      �S       ]                 �S      �S       X                 �S      �S       ]                �S      �S       w                 �S      �S       ��                �S      �S       w                 �S      �S       ��                   �S      �S       R�S      �S      
 q r "#���                  �S      �S       r ?&��S      �S       Q                     U      'U       U'U      (U       �U�                     U      'U       T'U      (U       �T�                      �N      �N       U�N      �N       �U��N      �N       U                      �N      �N       T�N      �N       �T��N      �N       T                          �N      �N       Q�N      �N       w �N      �N       �Q��N      �N       Q�N      �N       w                      �N      �N       W�N      �N       w���N      �N       W                     �N      �N       T�N      �N       �T��N      �N       T                     �N      �N       U�N      �N       �U��N      �N       U                        yM      �M       0��M      N       Y%N      <N       Y=N      BN       0�                        yM      �M       0��M      �M       R%N      <N       R=N      BN       0�                  �M      <N       Z                   �M      �M       Q�M      �M       qp��M      �M       Q                    �M      �M       P�M      �M       p��M      �M       P                    �M      �M       S���M      �M       S�[�                    �M      
N       P
N      N       p�N      !N       P                    �M      N       QN      N       q�N      )N       Q                  N      N       R                      PL      �L       U�L      �L       �U��L      M       U                      PL      �L       T�L      �L       S�L      �L       �T��L      M       T                    kL      �L       VM      M       V                  �L      �L       T                  �L      �L       V                 �L      �L       T                 �L      �L       V                 �L      �L       T                 �L      �L       V                          �K      �K       U�K      �K       S�K      �K       �U��K      	L       U	L      ML       S                              �K      �K       T�K      �K       V�K      �K       �T��K      	L       T	L      "L       V"L      0L       T0L      ML       V                   �K      �K       v �1��K      �K       Q                    0K      TK       UTK      �K       �U�                    9K      zK      	 t 0$0&�zK      �K      	 t0$0&�                  =K      �K      	 x 0$0&�                    `K      lK       RlK      �K       Q�K      �K       R                      `K      dK       RdK      �K       Q�K      �K       R                  `K      lK       PlK      pK       p�                            ��      �       U�      i�       Vi�      x�       �U�x�      ��       U��      ͕       V͕      ֕       U                              ��      �       T�      #�       R#�      i�       _i�      x�       �T�x�      ��       T��      ͕       _͕      ֕       T                            ��      �       Q�      i�       \i�      x�       �Q�x�      ��       Q��      ͕       \͕      ֕       Q                            ��      �       R�      i�       Si�      x�       �R�x�      ��       R��      ͕       S͕      ֕       R                        ��      s�       ]x�      ��       ]��      ��       u ��      ͕       ]                                    F      vF       UvF      �G       ��~�G      �G       �U��G      �J       ��~�J      �J       �U��J      �J       ��~�J      �J       U�J      �J       �U��J      �J       U�J      )K       ��~                                    F      vF       TvF      �G       w �G      �G       �T��G      �J       w �J      �J       �T��J      �J       w �J      �J       T�J      �J       �T��J      �J       T�J      )K       w                                     F      vF       QvF      �G       ��~�G      �G       �Q��G      �J       ��~�J      �J       �Q��J      �J       ��~�J      �J       Q�J      �J       �Q��J      �J       Q�J      )K       ��~                        �F      �F       U���F      �F       U�T��F      �F       u s ����$ ��T��F      G      " u s ����$ ��t s ����$ ���G      �G      " u s ����$ ��t s ����$ ���G      �G       �t s ����$ ��                                         �F      2G       ^2G      ;G       U;G      �G       _�G      �G       ^�G      �G       _�G      H       UH      #J       _�J      �J       ^�J      �J       _�J      K       _K      K       u�K      K       _K      "K       u0�                          �F      �G       V�G      �J       V�J      �J       V�J      �J       v��J      �J       V�J      )K       V                                            �F      G       [G      2G       ��~2G      ;G       ^;G      �G       ~��G      �G       [�G      �G       ~��G      H       ^H      GH       ~�GH      �H       ~��H      �H       ^�H      #I       ~�#I      #J       \�J      �J       [�J      �J       \�J      K       ~�K      )K       ~�                                    G      7G       P}G      �G       P�G      H       PH      H       P�H      �H       PZI      eI       P
J      J       P7J      DJ       P�J      �J       P$K      )K       P                               >F      vF       0�vF      �G       ��~�G      UJ       ��~UJ      XJ       p�XJ      jJ       PjJ      wJ       ��~�#��J      �J       ��~�J      )K       ��~                     >F      vF       0�vF      �F       [UJ      �J       [                                   �F      G      	 r 8$8&�;G      >G       p 38$8&�>G      bG       ~�38$8&��G      �G      	 r 8$8&�H      RH       ~�38$8&��H      �H       ~�38$8&�3I      ZI      	 z 8$8&�ZI      �I       0��I      �I      	 q 8$8&��I      #J       0�                        :F      �G       S�G      �J       S�J      �J       S�J      )K       S                                    >F      vF       ^vF      2G       _2G      �G       ]�G      �G       _�G      H       ]H      H       _H      7J       ]7J      �J       _�J      �J       _�J      �J       ]�J      )K       ]                            PF      vF      	 p 0$0&�vF      �G       ��~�0$0&��G      �J       ��~�0$0&��J      �J      	 u 0$0&��J      �J       ��~�0$0&��J      )K       ��~�0$0&�                      @E      E       TE      �E       �T��E      �E       T                      @E      �E       Q�E      �E       �Q��E      �E       Q                      @E      �E       R�E      �E       �R��E      �E       R                   @E      �E       6��E      �E       0��E      �E       6�                    }E      �E       P�E      �E       �T����34$z "�                      �D      E       UE      /E       �U�/E      3E       U                     �D      E       0�E      #E       P#E      3E       0�                  E      E       P                  E      E       P                          pC      �C       U�C      �D       \�D      �D       0��D      �D       U�D      �D       \�D      �D       U                      �C      �C       P�C      �D       ���D      �D       ��                 �C      �C       0�                          �C      �C       0��C      �C       v��C      7D       V7D      ;D       v��D      �D       0�                    �C      �C       S�C      CD       S                  �C      D       ~                 yD      �D       \                 yD      �D       ��                     0C      9C       0�9C      XC       YXC      jC       0�                     0C      =C       0�=C      XC       XXC      jC       0�                     0C      @C       0�@C      XC       PXC      jC       0�                        �q      r       Ur      Kr       SKr      Mr       �U�Mr      Vr       U                        �q      r       Tr      Lr       VLr      Mr       �T�Mr      Vr       T                       �q      r       0�r      r       Pr      Mr       QMr      Vr       0�                    �B       C       U C      C       �U�                    �B       C       T C      C       �T�                    �B       C       Q C      C       �Q�                    �B       C       R C      C       �R�                    �B      �B       U�B      �B       �U�                    �B      �B       T�B      �B       �T�                    �B      �B       Q�B      �B       �Q�                    �B      �B       R�B      �B       �R�                    �B      �B       U�B      �B       �U�                    �B      �B       T�B      �B       �T�                    �B      �B       Q�B      �B       �Q�                    �B      �B       R�B      �B       �R�                         A      `A       U`A      �B       �U��B      �B       U�B      �B       �U�                             A      �A       T�A      �A       S�A      �A       �T��A      �B       S�B      �B       T�B      �B       S                      A      >A       PDA      pA       PpA      tA       px�tA      �A       P                              A      >A       QDA      `A       Q`A      �A       U�A      0B       U�B      �B       U�B      �B       U�B      �B       qx�                     �A      �A       S�A      �A       0��A      �B       S�B      �B       S                      �A      �A       ]�A      �B       ]�B      �B       ]                     �A      �A       ^�A      �B       ^�B      �B       ^                     �A      �A       \�A      �B       \�B      �B       \                 �A      �A       S                 �A      �A       ]                 �A      �A       S                  �A      �A       S                  �A      �A       Q                  �A      �A      
 pl@     �                      �A      �A       s ��A      �A       U�A      �A       s �                    �A      �B       S�B      �B       S                    �A      �B       \�B      �B       \                   �A      0B       | �B      �B       |                       'B      GB       VGB      �B       0��B      �B       V�B      �B       0�                 �A      'B       S                 �A      'B       |��                  B      'B       V                   'B      �B       S�B      �B       S                 0B      @B       V                 0B      @B       |��                   GB      �B       \�B      �B       \                  GB      vB       0��B      �B       0�                  GB      vB       ltuo��B      �B       ltuo�                  GB      vB       \�B      �B       \                   OB      vB       P�B      �B       P                	   GB      vB       0��B      �B       0�                    VB      iB       QmB      vB       Q                    0@      8@       U8@      W@       �U�                    0@      8@       T8@      W@       �T�                    9@      A@       PJ@      R@       P                    �?      �?       U�?      0@       �U�                      �?      �?       T�?      @       \@      0@       �T�                 �?      @       S                  �?      @       ]                              Љ      +�       U+�      �       V�      �       �U��      6�       U6�      �       V�      ��       U��      ��       V                              Љ      +�       T+�      �       w �      �       ���      6�       T6�      �       w �      ��       T��      ��       w                       ��      �       ]6�      �       ]��      ��       ]                                   Љ      +�       0�+�      9�       _<�      ��       _��      ��       P��      �       S�      6�       0�6�      m�       Sm�      v�       0�v�      �       S�      ��       0���      ��       S                    �      +�       0��      ��       0�                 Ԋ      ؊       S                 A�      c�       S                   6�      �       S)�      5�       S��      ��       S                   6�      �       V)�      5�       V��      ��       V                    :�      �       \)�      5�       \��      ��       \                             :�      O�       0�O�      S�       PS�      Ջ       _Ջ      �       T�      �       _)�      5�       _��      ��       T��      ��       _                   [�      5�       S��      ��       S                      ^�      ��       Q��      ��       ��)�      5�       ��                 ��      ɋ       _                   ��      ��       v����      ɋ       U                   ɋ      �       V��      ��       V                  ɋ      ��       0���      ��       0�                  ɋ      ��       ltuo���      ��       ltuo�                  ɋ      ��       V��      ��       V                   Ћ      ��       P��      ��       P                   ɋ      ��       0���      ��       0�                    ڋ      �       Q�      ��       Q                      �      �       T�      )�       _)�      5�       _��      ��       _                    �      )�       \)�      5�       \��      ��       \                 c�      m�       S                 c�      m�       ]                          �{      �{       U�{      �{       P�{      �{       �U��{      �{       P�{      �{       U                        �{      �{       T�{      �{       Q�{      �{       �T��{      �{       T                 �{      �{       r�#                          �y      �y       U�y      �y       V�y      z       �U�z      ;z       U;z      �{       V                        �y      �y       T�y      �y       S�y      z       �T�z      �{       S                        �y      �y       Q�y      �y       \�y      z       �Q�z      �{       \                                     �y      �y       0�z      Rz       0�Rz      az       Phz      mz       P�z      �z       P�z      �z       _�z      �z       P�z      {       7�{      8{       P8{      l{       _l{      �{       0�                 �y      �y       t                       �z      {       XK{      ]{       X]{      g{       pg{      l{       X                   z      �z       ^l{      �{       ^                    @z      Qz       Pl{      r{       P                     fz      hz       Phz      �z       ���{      �{       ��                    �z      �z       Q�z      �z       q 4!��z      �z       Q                       �y      �y       0��z      �z       0��z      g{       ]g{      l{       Pr{      �{       0�                 �y      �y       �Q                   �y      �y       P                 �y      �y       V                  �y      �y       ]                 �y      �y       0�                    �y      �y       X�y      �y       }�y      �y       X                  ({      l{       �Q                    ({      l{       Q                  ({      l{       V                  8{      l{       P                 ({      l{       0�                      K{      ]{       Xa{      g{       pg{      l{       X                          P�      ��       U��      ۷       X۷      (�       �U�(�      F�       XF�      V�       U                                  P�      ��       T��       �       V �      �       �T��      �       V�      �       �T��      #�       V#�      (�       �T�(�      F�       VF�      V�       T                          P�      ��       Q��      ۷       Y�      (�       Q(�      F�       YF�      V�       Q                        P�      ۷       R۷      ��       S�      �       S�      V�       R                    ��      ۷       T(�      F�       T                             P�      ۷       0�۷      �       P�      ��       0���      ��       P�      �       0��      (�       6�(�      V�       0�                      ŷ      ��       ]�      �       ]?�      F�       ]                  ��      ��       V                  ��      ��       U                 ��      ��       T                  �?      �?       0��?      �?       0�                  �?      �?       T�?      �?       T                  �?      �?       U�?      �?       U                    �?      �?       Q�?      �?       Q                  �?      �?       0��?      �?       0�                      �?      �?       P�?      �?       q�?      �?       P�?      �?       P                        �>      �>       P�>      �>       u �>      �>       P�>      �>       u                           �;      �;       U�;      �;       S�;      �;       �U��;      	<       S	<      <       U                 �;      �;       P                   �;      �;       Q�;      �;       s                   �;      �;       U                   �;      �;       0��;      �;       P                            @;      l;       Ul;      �;       S�;      �;       �U��;      �;       S�;      �;       �U��;      �;       U                 r;      ~;       P                   M;      W;       PW;      a;       u                   T;      q;       Q                   T;      r;       0�r;      ~;       P                            �:      �:       U�:      ;       S;      ;       �U�;      ";       S";      (;       �U�(;      >;       U                            �:      �:       T�:      ;       V;      ;       �T�;      #;       V#;      (;       �T�(;      >;       T                            �:      �:       Q�:      ;       \;      ;       �Q�;      %;       \%;      (;       �Q�(;      >;       Q                            �:      �:       R�:      ;       ];      ;       �R�;      ';       ]';      (;       �R�(;      >;       R                   �:      	;       P;      !;       P                    �:      �:       Y1;      =;       Y                       �:      �:       0��:      	;       P;      !;       P1;      =;       0�                                 :      ]:       U]:      w:       Sw:      :       U:      �:       �U��:      �:       U�:      �:       S�:      �:       �U��:      �:       U                                 :      V:       TV:      x:       Vx:      :       T:      �:       �T��:      �:       T�:      �:       V�:      �:       �T��:      �:       T                                 :      ^:       Q^:      z:       \z:      :       Q:      �:       �Q��:      �:       Q�:      �:       \�:      �:       �Q��:      �:       Q                                 :      ^:       R^:      |:       ]|:      :       R:      �:       �R��:      �:       R�:      �:       ]�:      �:       �R��:      �:       R                                 :      ^:       X^:      ~:       ^~:      :       X:      �:       �X��:      �:       X�:      �:       ^�:      �:       �X��:      �:       X                   _:      v:       P�:      �:       P                    2:      ^:       Y�:      �:       Y                       2:      _:       0�_:      v:       P�:      �:       P�:      �:       0�                              �9      �9       U�9      �9       S�9      �9       U�9      �9       �U��9      :       S:      	:       �U�	:      :       U                              �9      �9       T�9      �9       V�9      �9       T�9      �9       �T��9      :       V:      	:       �T�	:      :       T                   �9      �9       P�9      :       P                  �9      �9       Q                     �9      �9       0��9      �9       P�9      :       P                                   9      ?9       U?9      K9       SK9      L9       UL9      M9       �U�M9      n9       Sn9      o9       �U�o9      �9       S�9      �9       U�9      �9       S                   ?9      B9       Pk9      k9       0��9      �9       P                         09      B9       PM9      Z9       Pk9      k9       0�w9      �9       P�9      �9       P                   W9      k9       Uo9      v9       U                      W9      k9       0�o9      w9       0�w9      �9       P�9      �9       P                                 8      d8       Ud8      v8       Sv8      x8       Ux8      y8       �U�y8      �8       S�8      �8       �U��8      �8       U�8      9       S                                   8      d8       Td8      w8       Vw8      x8       Tx8      y8       �T�y8      �8       T�8      �8       V�8      �8       �T��8      �8       T�8      9       V                             8      d8       Qd8      y8       �Q�y8      �8       Q�8      �8       �Q��8      �8       Q�8      9       w                              8      d8       Rd8      y8       �R�y8      �8       R�8      �8       �R��8      �8       R�8      9       �\                    d8      g8       P�8      �8       0��8      �8       P                        N8      g8       P�8      �8       0��8      �8       P�8      9       P                    y8      �8       U�8      �8       U                     y8      �8       0��8      �8       0��8      9       P                                `7      �7       U�7      �7       S�7      �7       U�7      �7       �U��7      �7       U�7      �7       S�7      �7       �U��7      8       S                                `7      �7       T�7      �7       V�7      �7       T�7      �7       �T��7      �7       T�7      �7       V�7      �7       �T��7      �7       T�7      8       V                   �7      �7       P�7      �7       0��7      �7       P                       {7      �7       P�7      �7       P�7      �7       0��7      8       P                   �7      �7       U�7      �7       U                    �7      �7       0��7      �7       0��7      8       P                            p>      �>       U�>      �>       S�>      �>       �U��>      �>       S�>      �>       �U��>      �>       U                            p>      �>       T�>      �>       V�>      �>       �T��>      �>       V�>      �>       �T��>      �>       T                    �>      �>       P�>      �>       P                 �>      �>       P                   �>      �>       s��>      �>       T                            >      (>       U(>      K>       SK>      N>       �U�N>      W>       SW>      Y>       �U�Y>      c>       U                            >      %>       T%>      L>       VL>      N>       �T�N>      X>       VX>      Y>       �T�Y>      c>       T                    ->      M>       PN>      V>       P                 2>      M>       P                   2>      K>       s�K>      M>       T                            �=      �=       U�=      �=       S�=      �=       �U��=      >       S>      >       �U�>      >       U                    �=      �=       P�=      >       P                 �=      �=       P                   �=      �=       s��=      �=       T                      �=      �=       U�=      �=       �U��=      �=       U                            �=      �=       T�=      �=       S�=      �=       �T��=      �=       S�=      �=       �T��=      �=       T                            �=      �=       Q�=      �=       V�=      �=       �Q��=      �=       V�=      �=       �Q��=      �=       Q                    �=      �=       P�=      �=       P                 �=      �=       P                          =      D=       UD=      `=       S`=      l=       �U�l=      q=       Sq=      w=       �U�                          =      A=       TA=      g=       Vg=      l=       �T�l=      t=       Vt=      w=       �T�                          =      H=       QH=      i=       \i=      l=       �Q�l=      v=       \v=      w=       �Q�                    I=      k=       Pl=      s=       P                       I=      `=       s�`=      k=       Tl=      q=       s�q=      w=       �U#�                 N=      k=       P                  �6      �6       T                    �6      �6       Q�6      V7       Q                   �6      P7       0�P7      V7       7�                        �5      �5       U�5      �5       V�5      �5       U�5      	6       �U�                        �5      �5       T�5      �5       �T��5      �5       T�5      	6       �T�                          �5      �5       Q�5      �5       \�5      �5       Q�5      6       \6      	6       �Q�                   �5      �5       0��5      	6       Q                       �5      �5       0��5      �5       P�5      �5       0��5      6       P                  �5      �5       S                      6      06       U06      p6       Sp6      �6       �U�                      6      B6       TB6      �6       V�6      �6       �T�                       6      a6       0�a6      c6       Pc6      r6       0�r6      �6       P                 <6      J6       0�c6      c6       0�                 <6      J6       Sc6      c6       S                   <6      E6       0�E6      J6       PJ6      J6       0�c6      c6       P                 <6      D6       U                            P�      ��       U��      %�       S%�      8�       �U�8�      T�       UT�      b�       Sb�      ��       �U�                        P�      ��       T��      8�       ��8�      T�       TT�      ��       ��                          P�      ��       Q��      /�       V/�      8�       �Q�8�      T�       QT�      ��       V                          P�      ��       R��      1�       \1�      8�       �R�8�      T�       RT�      ��       \                   ��      3�       ]T�      ��       ]                   ��      7�       _T�      ��       _                            f�      ��       0���      ��       P��      5�       ^8�      T�       0�T�      }�       ^}�      �       T��      ��       0���      ��       ^                   T�      }�       ^}�      �       T                 T�      s�       ~                 T�      s�       ~                  b�      ��       S                   t�      }�       ^}�      �       T                 t�      ��       S                              �      b�       Ub�      m�       �U�m�      ��       U��      *�       V*�      /�       �U�/�      1�       U1�      F�       V                      &�      j�       \m�      ,�       \1�      F�       \                   &�      b�       |�m�      ��       |�                           &�      I�       0�I�      T�       PT�      [�       S[�      ]�       p�]�      b�       Pm�      r�       0�                    ��      �       Q1�      F�       Q                    ��      .�       ]1�      F�       ]                 ��      $�       V$�      /�       0�                 ��      �       v                 ��      �       v                   	�      )�       S                 �      $�       V                 �      $�       S                          5      +5       0�+5      ;5       P;5      =5       q�=5      C5       QC5      J5       0�                        <      F<       UF<      �<       ]�<      �<       �U��<      �<       U                        <      F<       TF<      �<       V�<      �<       �T��<      �<       T                      '<      �<       S�<      �<       S�<      �<       u�                   ?<      �<       \                      p4      �4       T�4      �4       �T��4      �4       T                        �4      �4       P�4      �4       P�4      �4       P�4      �4       u�                     �4      �4       R�4      �4       R                              �3      4       U4      $4       S$4      *4       U*4      +4       �U�+4      :4       S:4      @4       �U�@4      f4       U                              �3      �3       T�3      )4       ])4      *4       T*4      +4       �T�+4      ?4       ]?4      @4       �T�@4      f4       T                              �3      4       Q4      %4       V%4      *4       Q*4      +4       �Q�+4      ;4       V;4      @4       �Q�@4      f4       Q                              �3      4       R4      '4       \'4      *4       R*4      +4       �R�+4      =4       \=4      @4       �R�@4      f4       R                   4      4       P+4      94       P                    �3      4       XV4      f4       X                       �3      4       0�4      4       P+4      94       PV4      f4       0�                              �1      -2       U-2      /3       S/3      53       �U�53      ;3       S;3      A3       �U�A3      g3       Ug3      �3       S                                �1      -2       T-2      A3       �T�A3      J3       TJ3      M3       �T�M3      U3       TU3      X3       �T�X3      e3       Te3      �3       �T�                        �1      -2       Q-2      A3       �Q�A3      g3       Qg3      �3       �Q�                              �1      $2       R$2      43       \43      53       �R�53      @3       \@3      A3       �R�A3      g3       Rg3      �3       \                              �1      -2       X-2      23       V23      53       �X�53      <3       V<3      A3       �X�A3      g3       Xg3      �3       V                         �1      02       0�02      M2       PM2      :3       TA3      g3       0�g3      �3       T                      �1      2       P2      2       u�A3      J3       u�                       �2      �2       R�2      �2       v �3      �3       R�3      �3       v                        �2      �2       U�2      3       X3      .3       vg3      �3       U                  �2      �2       I��3      �3       I�                    �2      �2       p 
����2      �2      	 y�
����3      �3      	 y�
���                      �2      �2       R�2      �2       v �3      �3       R�3      �3       v                   �2      �2       1��3      �3       1��3      �3       	��                    �2      �2       p 
����2      �2      	 y�
����3      �3      	 y�
���                  �2      �2       I��3      �3       I�                       �2      �2       p�-I�-� ��2      �2       p �-I�-� ��2      �2       z �-I�-� ��3      �3       <p �-I�-� ��3      �3       <y�
��v �-I�-� �                 	   �2      �2       R�3      �3       <p �-I�-� ��3      �3       <y�
��v �-I�-� �                  �2      3       I�g3      �3       I�                    �2      �2       p 
����2      3      	 y�
���g3      �3      	 y�
���                      �2      �2       U�2      3       X3      3       vg3      �3       U                  �2      3       1�g3      g3       1�g3      �3       	��                    �2      �2       p 
����2      3      	 y�
���g3      �3      	 y�
���                  �2      3       I�g3      �3       I�                       �2      3       p�-I�-� �3      3       p �-I�-� �3      3       u �-I�-� �g3      �3       <p �-I�-� ��3      �3       <y�
��u �-I�-� �                    3      3       Xg3      �3       <p �-I�-� ��3      �3       <y�
��u �-I�-� �                  I2      r2       y                   I2      r2       v                  I2      k2       y                  I2      k2       v                       U2      W2       PW2      _2      
 p q "#���_2      k2       R                       U2      W2       p ?&�W2      c2       Qc2      g2       p ?&�g2      k2       v � $ &y � $ &?&�                 v2      �2       y(                 v2      �2       v                 v2      �2       y(                 v2      �2       v                     v2      x2       Px2      �2      
 p q "#����2      �2       U                   v2      x2       p ?&�x2      �2       Q                      p1      �1       U�1      �1       �U��1      �1       U                        p1      �1       T�1      �1       Q�1      �1       �Q��1      �1       Q                          p1      }1       Q}1      �1       �Q��1      �1       Q�1      �1       �Q��1      �1       Q                      �0      11       U11      71       �U�71      b1       U                      �0      �0       TR1      [1       T[1      ]1       �T�                          �0      �0       Q�0      1       �Q�71      71       �Q�71      R1       �Q@+( �R1      ]1       Q]1      b1       �Q@+( �                            �0      1       R1      11       R71      K1       XK1      R1       �X�R1      ]1       R]1      b1       X                          �0      1       X1      11       X71      K1       XK1      R1       �X�R1      b1       X                           0      30       U30      ]0       S]0      ^0       �U�^0      v0       Uv0      �0       S                             0      W0       TW0      ^0       �T�^0      �0       T�0      �0       �T��0      �0       T�0      �0       �T�                         0      X0       0�X0      X0       P^0      �0       0��0      �0       P�0      �0       0�                     ?0      W0       s�#v0      �0       s�#�0      �0       s�#                     �0      �0       �h��0      �0       R�0      �0       �h�                   �0      �0       0��0      �0       0�                     �0      �0       T�0      �0       �T��0      �0       T                   �0      �0       S�0      �0       S                              �+      �+       U�+      �+       V�+      ,       U,      =,       �U�=,      �-       V�-      �-       U�-      �/       V                                    �+      =,       T=,      �,       R�,      O-       �T�O-      h-       Rh-      �-       �T��-      (.       R(.       /       �T� /      5/       R5/      |/       �T�|/      �/       R                          �+      ,       \,      7,       s�=,      �-       \�-      �-       T�-      �/       \                                        �+      �+       0�=,      W,       0�W,      g,       Tw,      w,       TO-      h-       0��-      �-       0��-      �-       T�-      .       0�.      .       T.      .       0�.      (.       T /      5/       0�|/      �/       0�                                              �+      �+       0�=,      ],       0�],      t,       Yw,      =-       YO-      h-       0��-      �-       0��-      �-       T�-      .       0�.      .       T.      #.       0�#.      f.       Yo.      �.       Y�.       /       Y /      5/       0�5/      |/       Y|/      �/       0�                                         �+      �+       0�=,      �,       0��,      O-       [O-      h-       0��-      �-       [�-      �-       {`��-      (.       0�(.      j.       [j.      o.       Po.       /       [ /      5/       0�5/      |/       [|/      �/       0�                                         �+      �+       0�=,      �,       0��,      O-       ZO-      h-       0��-      �-       Z�-      �-       z`��-      (.       0�(.      �.       Z�.      �.       P�.       /       Z /      5/       0�5/      |/       Z|/      �/       0�                   �,      -       T�.      �.       T                   �,      -       [�.      �.       [                   �,      -       1��.      �.       1��.      �.       	��                   �,      -       [�.      �.       [�.      �.       { �                   �,      -       T�.      �.       T                      �,      -       t 1%{ @$"�-t �-� �-      -       P�.      �.       { @$t 1%"�-t �-� �                    �,      -       t 1%{ @$"�-t �-� �-      -       P�.      �.       { @$t 1%"�-t �-� �                     -      /-       Y�.       /       Y5/      U/       Y                     -      /-       Z�.       /       Z5/      U/       Z                     -      /-       1��.      �.       1��.       /       	��5/      U/       1�                     -      /-       Z�.      �.       Z�.       /       z �5/      U/       Z                     -      /-       Y�.       /       Y5/      U/       Y                       /       /       z @$y 1%"�-y �-� �5/      M/       y 1%z @$"�-y �-� �M/      U/       P                     /       /       z @$y 1%"�-y �-� �5/      M/       y 1%z @$"�-y �-� �M/      U/       P                  w-      �-       s                     w-      �-       P�-      �-      
 v��
���                 w-      �-       U                 w-      �-      
 v��
���                      �-      �-       U�-      �-      
 q u "#����-      �-       [                   �-      �-       u ?&��-      �-       Q                 �-      �-       s(                 �-      �-      
 v��
���                		 �-      �-       X�-      �-       Z                 �-      �-       P                   (.      T.       Y�.      �.       Y                   (.      T.       Z�.      �.       Z                   (.      T.       1��.      �.       1��.      �.       	��                   (.      T.       Z�.      �.       Z�.      �.       z �                   (.      T.       Y�.      �.       Y                    ?.      T.       y 1%z @$"�-y �-� ��.      �.       z @$y 1%"�-y �-� �                  ?.      T.       y 1%z @$"�-y �-� ��.      �.       z @$y 1%"�-y �-� �                    `*      d*       Td*      �+       �T�                            o*      �*       r��*      �*       T�*      �+       r��+      �+       T�+      �+       r��+      �+       T                           o*      �*       T�*      �*       �T5$u� "��*      &+       �T5$u� "�&+      ]+       T]+      �+       �T5$u� "��+      �+       �T5$u� "�                    �*      �*      
 u��
����*      �*       T�*      +       T                    �*      �*       Q�*      +       Q+      +       �T5$u� "#                  �*      �*       1��*      �*       1��*      +       	��                    �*      �*       Q�*      �*       Q�*      +       q �+      +       �T5$u� "#�                   �*      �*       T�*      +       T                          �*      �*       t 1%q @$"�-t �-� ��*      �*       t 1%�T5$u� "#@$"�-t �-� ��*      �*       P�*      +       q @$t 1%"�-t �-� �+      +       �T5$u� "#@$t 1%"�-t �-� �                   �*      �*       t 1%q @$"�-t �-� ��*      +       q @$t 1%"�-t �-� �+      +       �T5$u� "#@$t 1%"�-t �-� �                      �*      �*       T+      &+       Tk+      �+       T�+      �+       T�+      �+      
 u��
���                          �*      �*       Y�*      �*       �T5$u� "#+      &+       Yk+      y+       Py+      �+       Y�+      �+       Y�+      �+       �T5$u� "#                    �*      �*       1�+      &+       1�k+      �+       1��+      �+       1��+      �+       	��                           �*      �*       Y�*      �*       �T5$u� "#+      +       Yk+      y+       Py+      �+       Y�+      �+       Y�+      �+       y ��+      �+       �T5$u� "#�                      �*      �*       T+      &+       Tk+      �+       0��+      �+       T�+      �+      
 u��
���                            �*      �*       t 1%y @$"�-t �-� ��*      �*       t 1%�T5$u� "#@$"�-t �-� ��*      �*       P�+      �+       y @$t 1%"�-t �-� ��+      �+       �T5$u� "#@$t 1%"�-t �-� ��+      �+      - �T5$u� "#@$u��
��1%"�-u��
���-� �                      �*      �*       P�+      �+       y @$t 1%"�-t �-� ��+      �+       �T5$u� "#@$t 1%"�-t �-� ��+      �+      - �T5$u� "#@$u��
��1%"�-u��
���-� �                       7       t                           (       u��0$0&�(      0       Q0      7       u��0$0&�                       7       t                       7       u��0$0&�                   0      7       Q7      7      
 p q "#���                  0      7       q ?&�7      7       P                [      b       t                [      b       u��0$0&�                [      b       t                [      b       u��0$0&�                  [      b       Qb      b      
 p q "#���                  [      b       q ?&�b      b       P                w      �       t                    w             u��0$0&�      �       P�      �       u��0$0&�                w      �       t                w      �       u��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       t                    �      �       u��0$0&��      �       P�      �       u��0$0&�                �      �       t                �      �       u��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                      �)      !*       T!*      (*       �T�(*      `*       T                      �)      �)       Q�)      �)       u�)      `*       X                            �(      )       U)      6)       S6)      A)       �U�A)      X)       UX)      �)       S�)      �)       U                   �(      6)       0�A)      �)       0�                          �(      6)       \A)      U)       \U)      X)       u #�X)      �)       \�)      �)       \                     �(      )       |A)      U)       |U)      X)      	 u #�#                          �(      <)       VA)      S)       VS)      X)       u X)      �)       V�)      �)       V                     )      )       R)      6)       0�X)      �)       0�                   �(      )       UA)      X)       U                     �(      )       v��A)      S)       v��S)      X)       u #��                    �(      )       RA)      X)       R                 )      )       R                 )      )       v��                          ��      �       U�      �       S�      �       �U��      ��       S��      Ɖ       U                          ��      �       T�      �       \�      �       �T��      ��       \��      Ɖ       T                    ؈      �       V�      ��       V                 ш      �       P                   ш      �       ^�      ��       ^                           ��      ��       0���      �       P�      �       ]�      )�       P)�      ��       ]��      Ɖ       0�                               ��      �       0��      �       0��      1�       0�1�      5�       P5�      E�       _E�      ]�       P]�      ��       _��      ��       T��      Ɖ       0�                           ��      �       0��      5�       0�E�      ^�       0�^�      n�       Pn�      w�       }� ��      Ɖ       0�                �      �       ]                �      �       V                 5�      E�       _                 5�      E�       V                 ��      ��       T                 ��      ��       U                         (      e(       Ue(      �(       S�(      �(       �U��(      �(       U                    (      �(       #��(      �(       0��(      �(       #�                 8(      �(       V                 8(      i(       v                   [(      q(       Rr(      �(       0�                 8(      [(       U                 8(      [(       v �                  <(      [(       R                 [(      j(       R                 [(      j(       v �                        0v      Yv       UYv      �v       V�v      �v       �U��v      w       U                        0v      ev       Tev      �v       S�v      �v       �T��v      w       T                      fv      jv       Pjv      �v       7��v      �v       P�v      �v       �L                      Hv      tv       \�v      �v       \�v      �v       u�                   jv      tv       |tv      �v       P                  �v      �v       v  $0.��                   �v      �v       �X�v      �v       0�                  �v      �v       S                 �v      �v       �X                 �v      �v       S                      w      5w       U5w      ;w       �U�;w      Fw       U                        w      !w       T!w      5w       �H5w      ;w       �T�;w      Fw       T                                                                    ��      �       U�      ��       S��      ��       �U���      �       S�      #�       ��|#�      |�       �U�|�      ��       ��|��      ��       �U���      ��       S��      y�       ��|y�      ��       U��      ��       �U���      H�       ��|H�      z�       �U�z�      ��       ��|��      ��       S��      ��       �U���      ��       ��|��      Ȩ       SȨ      @�       ��|@�      C�       �U�C�      n�       ��|n�      ��       �U���      �       ��|�      ��       �U���      ӫ       ��|                                                        ��      �       T�      #�       V#�      |�       �T�|�      ��       V��      ��       �T���      y�       Vy�      ��       T��      ��       �T���      H�       VH�      z�       �T�z�      ;�       V;�      C�       _C�      �       V�      ��       _��      �       V�      )�       _)�      t�       �T�t�      ~�       _~�      ��       V��      ӫ       �T�                              ��      ��       Q��      :�       ��|:�      |�       �Q�|�      y�       ��|y�      ��       Q��      ��       �Q���      ӫ       ��|                          ��      �       R�      y�       ��|y�      ��       R��      ��       �R���      ӫ       ��|                                                  ��      �       X�      #�       ^#�      |�       �X�|�      ��       ^��      ��       �X���      y�       ^y�      ��       X��      ��       �X���      H�       ^H�      z�       �X�z�      ��       ^��      C�       �X�C�      �       ^�      ��       �X���      �       ^�      ~�       �X�~�      ӫ       ^                                                      ��      =�       0�=�      |�       [|�      ��       ��|��      ��       _��      �       0��      #�       [W�      \�       ��||�      ��       [��      ɥ       0�ɥ      L�       _L�      d�       [d�      y�       _y�      ��       0���      �       _�      >�       [>�      M�       ��|z�      ��       [��      Ȩ       [�      �       _~�      ��       _��      ��       0���      ӫ       _                                                 ��      %�       0�%�      (�       P(�      |�       s |�      ��       ��|��      �       0��      s�       ��||�      ��       ��|��      ��       s ��      ɥ       ��|ɥ      y�       ��|y�      ��       0���      ��       ��|��      ��       s ��      ��       ��|��      Ȩ       s Ȩ      n�       ��|�      ӫ       ��|                                 Ģ      ��       0���      ѣ       Pѣ      ף       T��      \�       0�|�      ��       0���      n�       0�٪      �       P�      ~�       0���      ӫ       0�                                �      #�       ]|�      ��       ]��      y�       ]��      H�       ]z�      0�       ]C�      �       ]��      �       ]~�      ӫ       ]                            ��      y�       S��      �       Sz�      ��       S��      ��       S��      ��       ��|#���      ��       S                        ��      y�       \��      �       \z�      ��       \��      ӫ       \                     I�      U�       0�U�      |�       X��      Ȩ       0�                     I�      Y�       0�Y�      |�       Y��      Ȩ       0�                     ɥ      ԥ       0�ԥ      إ       Xd�      y�       0�                   ɥ      إ       0�d�      y�       0�                  ��      զ       0��      �       0�                       ��      ��       X��      ͦ       ��|�      �       X�      �       ��|                 ��      զ       0��      �       0�                  ��      Ϋ       ]                  ��      ʫ       Sʫ      Ϋ       0�                  ��      Ϋ       V                 ��      ��       S                 ��      ʫ       S                 ��      ʫ       V                  b�      ��       0�                   ��      ��       P��      ��       P                    ��      Ѫ       P~�      ��       P                   ģ      ѣ       Pѣ      ף       T                 ģ      ѣ       x�# �                  #�      (�       ��|W�      \�       0�                  0�      \�       V                 N�      W�       V                                �      7�       V��      ��       VȨ      ;�       V;�      C�       _C�      n�       V�      ��       _��      �       V�      )�       _)�      b�       �T�t�      ~�       _                      �      7�       ��|��      ��       ��|Ȩ      n�       ��|�      b�       ��|t�      ~�       ��|                      �      7�       ��|��      ��       ��|Ȩ      n�       ��|�      b�       ��|t�      ~�       ��|                 �      >�       ��|                       �      7�       ��|��      ��       ��|Ȩ      @�       ��|C�      n�       ��|��      �       ��|                        �      7�       P��      ��       U�Ȩ      ը       U�a�      n�       P��      �       Pb�      b�       0�                 �      �       ��|                 �      �       ��|                 �      >�       ��|                 �      �       ��|                   d�      y�       0�y�      ��       P                         �      �      	 q  $ &��      �       Q�      �       q���      �      , ���H0H%�$!0)( 8/�� $ &�                        �      �       q  $ &#	�#���      �       q� $ &#	�#���      �      4 ���H0H%�$!0)( 8/�� $ &#	�#���      �       Q                &�      d�       0�                 &�      >�       ��|                &�      d�       0�                 d�      y�       ��                     d�      l�       ��~�l�      x�       Px�      y�       ��|                           �      ;�       V;�      C�       _�      ��       _�      )�       _)�      t�       �T�t�      ~�       _                      �      C�       ��|�      ��       ��|�      b�       ��|t�      ~�       ��|                      �      C�       ��|�      ��       ��|�      b�       ��|t�      ~�       ��|                           �      �       P�      @�       S@�      C�       ^�      ��       ^�      "�       ^t�      ~�       ^                         ��      6�       ^6�      C�       ��|�      ��       ��|�      b�       ��|t�      ~�       ��|                                  ��      @�       2�@�      V�       P��      ��       P��      ܩ       Pܩ      �       ��|�      C�       P�      )�       P)�      b�       \b�      b�       0�t�      ~�       P                            �      @�       0�@�      �       \�      �       |�&�      C�       \�      ��       \�      )�       0�t�      ~�       \                        @�      �       S4�      C�       1��      ��       St�      ~�       S                         ��      @�       0�@�      C�       V�      ��       V�      �       Vt�      y�       V                 ��      ��       0�                    ��      ܩ       Tܩ      �       ��|                    ũ      ܩ       Qܩ      �       ��|                   ũ      ܩ       Tܩ      �       ��|                 �      ��       T                 �      ��       Q                         @�      &�       ^&�      C�       ^�      ��       ^�      "�       ^t�      ~�       ^                 &�      4�       \                 9�      ?�       T                 9�      @�       ^                 H�      b�       ��|                 Y�      u�       V                 Y�      b�       ��|                 l�      u�       V                  ��      ��       } ��                  ��      ��       S                    б      ڱ       Uڱ      ۱       �U�                    б      ڱ       Tڱ      ۱       �T�                    б      ڱ       Qڱ      ۱       �Q�                    б      ڱ       Rڱ      ۱       �R�                                                    ��      ��       U��      ��       V��      �       �U��      ��       V��      =�       ��~=�      v�       �U�v�      ��       V��      ?�       ��~?�      �       �U��      :�       V:�      E�       ��~E�      [�       �U�[�      {�       V{�      ��       �U���      ��       V��      +�       �U�+�      V�       VV�      ��       �U�                                          ��      ��       T��      ��       S��      �       �T��      =�       S=�      v�       �T�v�      Ġ       SĠ      �       �T��      {�       S{�      ��       �T���      ��       S��      +�       �T�+�      _�       S_�      ��       �T�                    ��      ��       Q��      ��       �Q�                                ��      �       R�      ��       \��      �       �R��      ��       \��      b�       �R�b�      l�       \l�      ��       |���      ��       �R�                    ��      �       X�      ��       ��~                                �      ��       P��      �       w �      �       ��~�      +�       w +�      K�       ��~K�      U�       w U�      z�       ��~z�      ��       w                                            ��      ��       P�      F�       PG�      t�       Px�      y�       Py�      қ       Zқ      �       ��~$�      .�       ��b�      ��       P=�      B�       Zv�      ��       Z��      ��       ���      �       1��      �       Z�      �       ^��      ��       0�                        ��      ˛       Q˛      қ       �R~ �v�      ��       Q�      �       Q                           ��      $�       ��~v�      ��       ��~�      �       ��~�      :�       ��~[�      {�       ��~��      ��       ��~+�      V�       ��~                            ��      ��       Q��      ��       \v�      ��       \�      �       \�      0�       \[�      {�       \��      ��       \                       ��      ɛ       Rɛ      қ       ~ v�      ��       R�      �       R                       ��      Λ       TΛ      қ       ��v�      ��       T�      �       T                           ��      $�       Sv�      ��       S�      �       S�      :�       S[�      {�       S��      ��       S+�      V�       S                           ��      $�       Vv�      ��       V�      �       V�      :�       V[�      {�       V��      ��       V+�      V�       V                             ��      қ       v қ      $�       ��~v�      ��       v �      �       v �      :�       ��~[�      {�       ��~��      ��       ��~+�      V�       ��~                               ��      ��       0���      М       PМ      $�       \v�      ��       0��      �       0��      0�       0�[�      {�       0���      ��       0�+�      V�       \                           ��      ^�       ]^�      $�       }|�v�      ��       ]�      �       }|�[�      {�       ]��      ��       ]+�      V�       }|�                            �      A�       PA�      $�       _�      �       _0�      :�       _[�      {�       P��      ��       _+�      V�       _                	           ��      b�       0�v�      ��       0��      :�       0�[�      {�       0���      ��       0�+�      V�       0�                  ��      �       ]v�      ��       ]                  ��      �       Sv�      ��       S                  ��      �       0�v�      ��       0�                   ^�      ��       ]�      �       ]                   ^�      ��       S�      �       S                  ^�      ��       0��      �       0�                 ̜      ۜ       _                   ̜      М       PМ      ۜ       \                   ̜      М       UМ      ۜ       S                 +�      V�       \                 +�      V�       ��~                      )�      .�       T��      ��       ���      �       } ��      ��       T                      )�      D�       w ��      ��       w �      �       w ��      ��       w                             v�      =�       ��~��      �       ��~:�      [�       ��~{�      ��       ��~��      +�       ��~V�      ��       ��~                      v�      =�       _��      �       _:�      P�       _                                  v�      7�       ^��      ��       ^��      "�       ^"�      ߠ       ��~:�      E�       ^P�      [�       ��~{�      ��       ��~��      +�       ��~V�      ��       ��~                                  v�      =�       S��      Ġ       SĠ      �       �T�:�      [�       S{�      ��       �T���      ��       S��      +�       �T�V�      _�       S_�      ��       �T�                                  v�      ��       V��      =�       ��~��      ?�       ��~?�      �       �U�:�      E�       ��~E�      [�       �U�{�      ��       �U���      +�       �U�V�      ��       �U�                               ~�      ��       v ��      =�       ��~��      �       ��~:�      E�       ��~P�      [�       ��~{�      ��       ��~��      +�       ��~V�      ��       ��~                                 ~�      =�       0���      �       0��      �       P�      ڠ       _ڠ      ߠ       0�:�      P�       0�P�      [�       _{�      ��       _��      +�       _V�      ��       _                                          ��      ��       0���      �       ]�      �       }��      =�       ]��      ��       ]��      �       }��      ?�       0�?�      ��       \��      ��       |���      Ġ       \:�      E�       }�P�      [�       \��      ߡ       |�V�      ��       \                             �      ?�       1�?�      7�       ��~7�      _�       P_�      ߠ       ��~P�      [�       ��~{�      ��       ��~��      +�       ��~V�      ��       ��~                  ��      ��       P                                   �      ?�       0�?�      7�       ^7�      _�       R_�      ߠ       ^P�      [�       ^{�      ��       ^��      ˡ       ^ˡ      �       R�      #�       ^V�      ~�       ^~�      ��       R                                  ��      ��       0���      =�       \��      �       \�      ߠ       ��:�      E�       \P�      [�       ��{�      ��       ����      +�       ��V�      ��       ��                                 �      ?�       6�?�      2�       V2�      ;�       v�;�      C�       ]C�      I�       v�I�      O�       v�O�      U�       v�U�      ��       Q��      Ġ       VP�      [�       V��      ��       V��      ˡ       Pˡ      ԡ       p�ԡ      �       QV�      g�       Vg�      ~�       P~�      ��       p���      ��       Q                                 �      ?�       2�?�      ;�       ];�      C�       t}�C�      ߠ       ]P�      [�       ]{�      ��       ]��      ˡ       ]ˡ      +�       SV�      ~�       ]~�      ��       S                              x�      ��       P��      ؟       ��~؟      ��       R��      ��      ( ��~20��~#������������������+( �P�      [�       RV�      b�       Rb�      ��      ( ��~20��~#������������������+( �                    ڝ      �       P��      ��       P                  ��      ŝ       V'�      2�       V                  ��      ŝ       S'�      2�       S                 ��      ŝ       0�'�      2�       0�                      ?�      P�       XP�      _�       ��~��      Ġ       X                   ?�      c�       S��      Ġ       S                  ?�      c�       0���      Ġ       0�                   z�      ��       R��      ��      ( ��~20��~#������������������+( �                   z�      ��        q "���      ��       Q                 z�      ��       S                 ̠      ڠ       _                 ̠      ڠ       ��~                  =�      B�       ���      �       ^                  =�      Y�       w �      �       w                                  �      X�       UX�      ��       ]��      ��       �U���      .�       ].�      3�       �U�3�      R�       ]R�      W�       �U�W�      f�       U                                 �      C�       TC�      �       V�      ��       �T���      *�       V*�      3�       �T�3�      N�       VN�      W�       �T�W�      f�       T                                 �      P�       QP�      ��       ^��      ��       �Q���      0�       ^0�      3�       �Q�3�      T�       ^T�      W�       �Q�W�      f�       Q                                 �      `�       R`�      �       w �      ��       ��~��      �       w �      3�       �R�3�      ;�       w ;�      W�       �R�W�      f�       R                       �      `�       X`�      W�       ��~W�      f�       X                                 �      `�       Y`�      ��       \��      ��       �Y���      ,�       \,�      3�       �Y�3�      P�       \P�      W�       �Y�W�      f�       Y                           ��      ݬ       0�ݬ      �       P�      �       w ;�      L�       w L�      W�       ��~W�      f�       6�                      �      ��       0���      �       S��      )�       S3�      f�       0�                    �      +�       u W�      f�       u                    �      ��      
 `H@     �3�      ;�      
 `H@     �                   �      ��       �ܝ  3�      ;�       �ܝ                       �      P�       QP�      ��       ^3�      ;�       ^                     �      C�       TC�      ��       V3�      ;�       V                     �      X�       UX�      ��       ]3�      ;�       ]                
       �      d�       0�d�      h�       Ph�      ��       S3�      ;�       S                p�      ��       ^                p�      ��       V                p�      ��       S                 ��      �       S                 �      )�       S                    ;�      N�       VN�      W�       �T�W�      f�       0�                 W�      f�       u                       �             U             S             �U�                 �      �       u8                  �             T                      ��      ��       U��      ��       �U���      Ʊ       U                        ��      ��       T��      ��       ����      ��       �T���      Ʊ       T                        ��      ��       Q��      ��       �@��      ��       �Q���      Ʊ       Q                        ��      ��       R��      ��       P��      ��       �R���      Ʊ       R                        ��      ��       X��      ��       R��      ��       �X���      Ʊ       X                      �      �       U�      �       �U��      �       U                        �      ��       T��      �       �H�      �       �T��      �       T                      �      �       Q�      �       �Q��      �       Q                      �      �       R�      �       �R��      �       R                            ��      ��       U��      �       _�      ��       �U���      �       _�      u�       �U�u�      ��       _                        ��      ��       T��      ��       \��      ��       �T���      ��       \                    ��      ��       Q��      ��       �Q�                    ��      ��       R��      ��       ��                        ��      ��       X��      ��       ]��      ��       �X���      ��       ]                    ��      ��       Y��      ��       ��                    ��      �       S��      ��       S                    ��      ��       V��      ��       V                                ��      Ȇ       0�Ȇ      �       P�      ߇       ^߇      �       0���      �       P�      7�       ^7�      ^�       U^�      u�       ^u�      |�       P|�      ��       ^                           ��      �       0��      �       P�      ��       _ч      �       0���      �       0��      u�       _u�      ��       0�                  3�      M�       P                 (�      B�       0�                    ��      ��       S��      �       SX�      c�       S                        ��      ��       ^��      �       P�      �       ^X�      b�       Ub�      c�       ^                  Ç      ч       _��      ��       0�                  Ç      ч       S��      ��       S                 ч      ߇       ^                 ч      ߇       S                  t      �       T                        �      �       R�      �       P�      �       R�      �       R                           &      (&       U(&      �&       V�&      �&       U�&      �&       �U��&      '       V                           &      )&       T)&      �&       S�&      �&       T�&      �&       �T��&      '       S                       &      )&       Q)&      �&       ]�&      '       �Q�                  &      �&       \                 A&      ]&       ]                 A&      ]&       V                 A&      ]&      
 �G@     �                     A&      M&       s��M&      \&       U\&      ]&       s��                 v&      �&       V                 v&      �&       S                      �&      �&       s
 0.���&      �&       } 
 0.���&      '       } 
 0.��                    �&      �&       \�&      
'       \
'      '       0�                    �&      �&       ^�&      '       ^                 �&      �&       \                 �&      
'       \                 �&      
'       ^                 �&      �&       T                 �&      �&       V                     �&      �&       S�&      �&       T�&      �&       �T�                     �&      �&       V�&      �&       U�&      �&       �U�                              )       U)      d       Vd      g       Ug      h       �U�                              *       T*      c       Sc      g       Tg      h       �T�                            *       Q*      f       \f      h       �Q�                  B      O       T                  B      T       V                     \      c       Sc      g       Tg      h       �T�                     \      d       Vd      g       Ug      h       �U�                          0�      G�       UG�      j�       Sj�      o�       Uo�      p�       �U�p�      v�       U                      0�      R�       TR�      p�       �T�p�      v�       T                          0�      R�       QR�      k�       Vk�      o�       Qo�      p�       �Q�p�      v�       Q                     <�      R�       TR�      `�       �T�`�      o�       T                   L�      R�       TR�      `�       �T�                 L�      `�       S                     L�      X�       0�X�      ]�       P]�      `�       T                 L�      R�       U                                      �{      |       U|      P~       \P~      Q       �U�Q      _       U_      d�       \d�      p�       Up�      ��       \��      �       �U��      N�       \N�      i�       �U�i�      p�       \                                    �{      +|       T+|      '       ^'      -       u-      .       �T�.      @       ^@      Q       �T�Q      _       T_      d�       ^d�      p�       Tp�      p�       ^                                        �{      +|       Q+|      �|       V�|      .}       �Q�.}      4}       V4}      7}       v :!�7}      :}       p �Q�Q
  $0.( :!�:}             V              s�#H       -       u�#H.      <       s�#HQ      _       Q_      d�       Vd�      p�       Qp�      p�       V                                                �}      �}       P�}      �~       R�~      �~       R�~      �~       w �~      -       R.      <       R<      @       w _      {       R��      ��       P��      ��       P��      d�       RɁ      �       P.�      1�       P1�      ��       R�      [�       R[�      i�       w                          .}      i}       Q{      �       Q�      �       w �      �       Qi�      p�       Q                         |              S       -       U.      @       S_      d�       Sp�      p�       S                       .}      i}       q{      �       q�      �       qi�      p�       q                         .}      �}       _{      ؀       _p�      ?�       _�      �       _i�      p�       _                                     �{      |       U|      P~       \P~      Q       �U�Q      _       U_      d�       \d�      p�       Up�      ��       \��      �       �U��      N�       \N�      i�       �U�i�      p�       \                        �      �       R�      ��       ��p�      �       ��i�      p�       R                    )�      4�       0�p�      �       0�                  �      �       \i�      p�       \                    �      �       0��      �       Ui�      p�       0�                     �      �       Q�      �       w i�      p�       Q                   �      �       0�i�      p�       0�                 �      !�       u #(                   ��      !�       Z!�      ?�       ��                 ��      �       w                         �}      *~       q�*~      ?~       |�#�?�      o�       q�o�      ��       |�#�                   �}      ~       @�?�      d�       @�                   �}      ~       U?�      d�       U                       �}      �}       P�}      ~       s� ?�      D�       PD�      d�       s�                    �}      ~       1�~      ~       1�?�      ?�       1�?�      d�       	��                       �}      �}       P�}      ~       s� ?�      ?�       P?�      D�       p �D�      P�       s� �                  �}      ~       U~      ~       u �?�      d�       U                  �}      ~       @�?�      d�       @�                      ~      ~       t 6%�~      ~       P\�      _�       P_�      d�       p �                    ~      ~       P\�      _�       P_�      d�       p �                   ~      ;~       @�d�      ��       @�                   ~      ;~       Td�      ��       T                       ~      '~       P'~      ;~       s� d�      l�       Pl�      ��       s�                     ~      3~       1�3~      ;~       1�d�      d�       1�d�      x�       	��x�      ��       	��                       ~      '~       P'~      3~       s� d�      d�       Pd�      l�       p �l�      x�       s� �                  ~      3~       T3~      ;~       t �d�      x�       Tx�      ��       t �                  ~      ;~       @�d�      ��       @�                      3~      ;~       q 6%�;~      ;~       P��      ��       P��      ��       p �                    ;~      ;~       P��      ��       P��      ��       p �                      P~      �~       \��      �       \N�      i�       \                    �~      �~       U��      �       0�N�      i�       0�                     c~      �~       S��      �       SN�      i�       S                   c~      j~       Pj~      �~       s��      ��       s                    n~      �~       P�~      �~      	 s#�#��      ��      	 s#�#                    u~      �~       U�~      �~       p�~      �~       U��      ��       0�                     ~      �~       0���      �       0�N�      i�       0�                     ~      �~       Q��      ��       QN�      [�       Q                       ~      �~       P�~      �~      	 s#�#��      ��      	 s#�#N�      [�      	 s#�#                   �~      �~       P��      ��       P                     ~      �~       0���      �       0�N�      i�       0�                    �~      �~       U�~      �~       p                 �~      �~       \                 �~      �~       U                  ��      �       X                  ��      �       Y                  ��      �       s��                     ǂ      т       0�т      ۂ       Q�      �       Q                  ǂ      �       P                 W�      i�       \                   W�      [�       U[�      i�       ]                                        t ?�             T             v @&?�      -       T.      <       T                 |      .}       S                   ��      d�       y  $0.��      N�       y  $0.�                   ��      d�       S�      N�       S                   ��      d�       s0��      N�       s0�                          �      �       p x "#?	���      $�       x ��"#?	��$�      +�       P+�      ?�       x ��"#?	��)�      :�       t ��"#?	��B�      E�       T                     �      8�       ��u "#?	��8�      ;�       P;�      ?�       ��u "#?	��                      '      c'       Uc'      y'       �U�y'      �'       U                      '      _'       Ty'      �'       T�'      �'       �T��'      �'       T                   '      k'       Qy'      �'       Q                    '      x'       Py'      �'       P                          `%      �%       U�%      �%       S�%      �%       T�%      �%       �U��%      �%       U                        s%      �%       q��%      �%       u#��%      �%       s#��%      �%       q�                          �%      �%       V�%      �%      	 u#�#�%      �%       V�%      �%       U�%      �%       V                        �%      �%       0��%      �%       R�%      �%       R�%      �%       R�%      �%       0�                         �%      �%       R�%      �%       r�%      �%       R�%      �%       r�%      �%       r�%      �%       R                     �%      �%       S�%      �%       T�%      �%       �U�                   �%      �%       V�%      �%       U                              �w      x       Ux      3x       S3x      =x       �U�=x      �x       S�x      �x       �U��x      y       Uy      yy       S                              �w      x       Tx      4x       V4x      =x       �T�=x      �x       V�x      �x       �T��x      y       Ty      yy       V                 �w      x       P                 �w      x       p                      x      8x       ]=x      �x       ]y      yy       ]                              �w      x       0�x      x       Px      .x       \=x      �x       \�x      �x       �T�x      y       0�y      Ey       \Ey      Ny       0�Ny      yy       \                   Ex      �x       \y      /y       \Ny      ty       \                    Vx      �x       _y      /y       _Ny      ty       _                      jx      nx       Pnx      �x       w y      /y       w Ny      ty       w                    jx      �x       ^y      /y       ^Ny      ty       ^                           jx      �x       0��x      �x       P�x      �x       Xy      &y       X&y      /y       ��Ny      hy       ��                  "y      /y       ��Ny      [y       ��                    "y      &y       U&y      /y       ^Ny      [y       ^                    "y      'y       0�'y      /y       PNy      [y       P                 ;y      Ey       \                 ;y      Ey       ]                        �!      �!       U�!      �!       S�!      �!       �U��!      �!       S                    �!      �!       V�!      �!       V                 �!      �!       v                    �!      �!       \�!      �!       \                 �!      �!       s�                 �!      �!       \                  �!      �!       U                        Pw      �w       U�w      �w       S�w      �w       �U��w      �w       S                        Pw      ~w       T~w      �w       \�w      �w       �T��w      �w       T                    pw      �w       V�w      �w       V                  ~w      �w       T                  ~w      �w       V                      @%      P%       UP%      ]%       S]%      _%       �U�                      @%      P%       TP%      ^%       V^%      _%       �U#�                         "      U"       UU"      �#       [�#      �#       U�#      7%       [                           "      Z"       TZ"      �#       ^�#      �#       �T��#      �#       T�#      7%       ^                         "      ."       Q."      �#       �Q��#      �#       Q�#      7%       �Q�                        "      U"       u��U"      �#       {���#      �#       u���#      7%       {��                        "      U"       u��U"      �#       {���#      �#       u���#      7%       {��                         �"      D#       Z�#      �#       Z�#      1$       5�1$      �$       1��$      �$       6��$      7%       1�                                                                    �"      �"       P���"      �"       P�\���"      �"      	 w �\���"      �"       w �\�S���"      #       w �\�S�Y�#      #       X�\�S�Y�#      #       X�R�S�Y�#      #       X�R�P�Y�#      $#       X�R�P�Q�$#      m#       X�R�T�Q�m#      �#       X�R��Q��#      �#       X��Q��#      �#       X���#      �#       X�R�T�Q��#      R$       w �\�S�Y�R$      U$       X�\�S�Y�U$      y$       X�\�T�Y�y$      |$       X�R�T�Y�|$      �$       X�R�T�Q��$      �$       X�R�T�Q��$      �$       w �\�S�Y��$      �$       X�\�T�Y��$      �$       X�\�T�Y��$      %       X�R�T�Q�%      %       X�r��T�Q�%      %       X�\�T�Y�%      !%       X�\�T�Y�!%      ,%       X�R�T�Q�,%      7%       X�R�T�Q�                          "      *"       0�*"      7"       P7"      >"       S>"      H"       �Q�#      �#       0�                          "      ."       0�."      :"       Q:"      B"       ]B"      H"       �Q#�#      �#       0�                     #      �#       X�#      �#       X�$      �$       X,%      7%       X                     #      �#       Q�#      �#       Q�$      �$       Q,%      7%       Q                     $#      U#       P�#      �#       P�$      �$       t x �,%      7%       t x �                       '#      �#       Y�#      �#       Y�$      �$       Y2%      7%       1�                      D#      �#       U�#      �#       U�$      �$       U                   K"      Z"       ���Z"      _"       T                   K"      U"       u��U"      _"       {��                        `r      �r       U�r      ts       �U�ts      �s       U�s      �s       �U�                            `r      �r       T�r      �r       S�r      �r       �T��r      ts       Sts      �s       T�s      �s       S                            `r      �r       Q�r      �r       \�r      �r       �Q��r      ts       \ts      �s       Q�s      �s       \                     �r      �r       ^�r      ts       ^�s      �s       ^                               `r      �r       0��r      �r       P�r      �r       V�r      #s       V#s      +s       0�+s      hs       Vhs      is       Tts      �s       0��s      �s       V                 �r      �r       P                 �r      �r       s                 �r      �r       V                 s      #s       V                 s      #s       ^                     /s      9s       V`s      hs       Vhs      is       T                   /s      9s       ^`s      ts       ^                    �       �        U�       �        �U�                      �       �        T�       �        u� �       �        �T�                   �       �        U�       �        �U�                               )        U)       0        S0       a        �U�a       k        U                                   0        T0       R        VR       S        �T�S       `        V`       a        �T�a       k        T                            L        0�L       S        PS       k        0�                            )        U)       Q        Sa       k        U                        p      �       T�              �T�              T      x       �T�                        p      �       Q�              �Q�              Q      x       �Q�                        s      �       p���              �T#��       P       p��P      x       �T#��                    @      J       UJ      c       �U�                    @      J       TJ      c       �T�                   @      J       U��J      c       �U���                    F      J       TJ      c       �T�                  K      U       P                                 U      1       �U�                                 T      1       �T�                                U�      1       �U��                                T      1       �T�                        #       P                    0�      6�       U6�      7�       �U�                    0�      6�       T6�      7�       �T�                    0�      6�       Q6�      7�       �Q�                    0�      6�       R6�      7�       �R�                     �      $�       U$�      %�       �U�                     �      $�       T$�      %�       �T�                     �      $�       Q$�      %�       �Q�                     �      $�       R$�      %�       �R�                     ��      �       U�      %�       \M�      l�       \                                ��      �       T�      �       ]�      ,�       �T�,�      [�       ][�      c�       �T�c�      ��       ]��      �       �T��      �       ]                        ��      �       Q�      "�       S"�      ,�       �Q�,�      �       S                        ��      �       R�      )�       ^)�      ,�       �R�,�      �       ^                          �      �       P,�      A�       PB�      W�       PW�      [�        c�      ��                                �      �       P�      �       _,�      [�       _c�      ��       _                 �      �       P                   c�      ��       ^�      �       ^                   c�      ��       S�      �       S                    ��      ��       _�      �       _                      ��      ��       _��      �       \�      �       _                  ܖ      �       P                    ��      ��       0��      �       0�                   ��      ��       \�      �       \                  �      �       _�      �       _                  �      �       ^�      �       ^                        �      �       U�             ]             �U�      	       U                        �      �       T�      �       V�             �T�      	       T                    �      �       P�      �       u                  �      �       S                 �      �       0�                  �      �       T                  �      �       V                 �      �       }                  �      �       V                      ��      ��       U��      �       S�      �       �U�                      ��      Ƒ       TƑ      ��       U��      �       �T�                     ��      Ƒ       TƑ      ��       U��      ��       �T�                 ��      ��       1�                   ��      ��       U��      ��       S                      д      ڴ       Uڴ      %�       S%�      &�       �U�                      д      �       T�      �       U�      &�       �T�                     ڴ      �       T�      �       U�      �       �T�                 Դ      �       0�                   Դ      ڴ       Uڴ      �       S                      �       �        T�              V             �T�                   �       �        0��       �        P                  �       
       \                    �              S             P                    �      �       U�             �U�                    �      �       T�             �T�                      C       j        Qj       n        Rn       �        u � $ &�                              F       S        PS       V        q ��V       c        Pc       j        q �5$q 	�$"q ��j       n        r �5$r 	�$"r ��n       t        u ��Ou � $ &	�$"�t       �        R                         1        T                                    0�       +        P+       1        0�                 5      �       u�                 5      �       u� �                    A      d      	 p 0$0&�d      j       u� �0$0&�                 A      �      	 r 0$0&�                 T      j       0�                 �      '       u� �                 �             U                 �      '       u�                 �      '       u� �                       &       U                       '       u�                       '       u� �                          0�      U�       UU�      \�       �U�\�      z�       Uz�      ��       V��      ��       �U�                    0�      O�       TO�      ��       �T�                    E�      U�       Z\�      ��       Z                          O�      U�       T\�      r�       Tr�      ��       S��      ��       v��      ��       �U#                   O�      U�       Q\�      ��       Q                         M�      U�       u�U�      \�       �U#�\�      z�       u�z�      ��       v���      ��       �U#�                         M�      U�       u� �U�      \�       �U#`�\�      z�       u� �z�      ��       v� ���      ��       �U#`�                   ��      ��       V��      ��       �U�                   ��      ��       v���      ��       �U#�                   ��      ��       v� ���      ��       �U#`�                                ��      ?�       U?�      D�       SD�      N�       �U�N�      ��       S��      ��       �U���      ��       S��      Đ       �U�Đ      )�       S                    ��      �       T�      )�       �T�                            ��      �       Q�      4�       \4�      N�       �Q�N�      �       \�      Ր       �Q�Ր      )�       \                        �      I�       ]N�      ��       ]��      ��       ]Đ      )�       ]                               �      ?�       u�?�      D�       s�D�      N�       �U#�N�      ��       s���      ��       �U#���      ��       s���      Đ       �U#�Đ      )�       s�                               �      ?�       u� �?�      D�       s� �D�      N�       �U#`�N�      ��       s� ���      ��       �U#`���      ��       s� ���      Đ       �U#`�Đ      )�       s� �                        �      ?�       0�N�      я       0�я      �       1�5�      ��       1�Đ      Ր       1�Ր      )�       0�                                  �      4�       T4�      G�       \N�      V�       TV�      �       V�      ��       \��       �       |}� �      ��       \Đ      Ր       \Ր      )�       V                           �      /�       _/�      ?�       QN�      ��       _��      %�       QĐ      Ր       QՐ      )�       _                 >�      ��       S                 >�      ��       s�                 >�      ��       s� �                      `�      x�       Ux�      �       S�      ��       �U�                 `�      a�       u                 ю      �       S                ю      �       s�                ю      �       s� �                      P      h       Uh      P       SP      R       �U�                  `      Q       V                 `      j       T                 `      k       V                 w      �       T                 w      �       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                 �      �       T                 �      �       V                       D       S                         P       s�P      R       �U#�                         P       s� �P      R       �U#`�                 m      {       U                              �      �       U�             S             �U�      /       U/      1       S1      7       �U�7      S       U                          �      �       T�             �T�      /       T/      7       �T�7      S       T                              �      �       Q�             V             �Q�      /       Q/      4       V4      7       �Q�7      S       Q                    �             P/      3       P                         �      �       U�             S             �U�/      1       S1      7       �U�                 �      �       u�                            `      r       Ur      u       �U�u      �       U�             �U?&�U'�U?&�             U      -       �U?&�U'�U?&�                              `             T      �       �T��      �       T�      �      
 �Ty 'y ��             �T?&�T'�T?&�             T      -      
 �Ty 'y �                            `      �       Q�      �       �Q��      �       Q�             �Q?&�Q'�Q?&�      $       Q$      -       �Q?&�Q'�Q?&�                            `      �       R�      �       �R��      �       R�            
 �Ru 'u �      +       R+      -      
 �Ru 'u �                        g      �       P�      �       �U�Q"��             Y      -       P                      k      �       X�      �       �T�R"��      -       X                      �      �       T�             T       -       T                  �             R                  �      �       P                    @      J       TJ      Z       �T�                    @      D       RD      Z       �R�                    M      W       RW      Z      
 �Ru t �                     S      �       R�      �       Y�             R                      W      �       Q�      �       P�      �       Q                  �      j       R                         H       x x t t " ��H      g       q @<$�                      `      i       Ri      �       Y�      (       Y                        b      �       Q�      �       P�      �       P�      (       P                        �       X                          �       T(      =       T                                  �      �       Q�      �       X�      �       Q�      �       P�      �       P      
       Q
             X      (       Q(      =       P                     W      i       1�i      o       	��o      �       Z�      =       Z                   W      �       1��      �       [�      =       [                      �      �       S�      �       \      :       \                        �      �       U�      5       S5      =       �U�=      A       U                      �      �       T�      =       [=      A       T                      �      �       Q�      =       �Q�=      A       Q                                   | p "�      8       \8      =       �U                      *      0       v p "�0      6       V6      =       �U#                       �      �       q @$��      �       Q�      =       Z=      A       q @$�                        P      x       Ux      7       �U�7      C       UC      �       �U�                                       X�Y�Z�[�      %       X�Y�Z�S�%      -       X�Y�Z��-      4      
 �Y�Z��4      ;       �Z��                     �      �      
 ���������             Ut      �       U      $       U                   �      �       0��             Tt      |       T                  N      i       R                    R      \       P\      i       z { "�                   �      7       RC      �       R                t      �       
�Z�                 t      |       T                t      �       1�                 t      |       T                t      �       
�Z�                    �      7       RC      �       R                �      �       R                  �      �       R      7       R                   �      �       U      $       U                  �      �       1�             1�      7       	��                	   �      �       U             U      $       u �                
  �      �       R      7       R                  �      �       P      $       u @$t "�-r �-� �                 �      �       P      $       u @$t "�-r �-� �                   �      �       R�      �       R                       �      �       X�      �       �U�      �       X�      �       �U                  �      �       1��      �       1��      �       	��                      �      �       X�      �       �U�      �       X�      �       x ��      �       �U�                   �      �       R�      �       R                    �      �       P�      �       x @$t "�-r �-� ��      �       �U@$t "�-r �-� �                   �      �       P�      �       x @$t "�-r �-� ��      �       �U@$t "�-r �-� �                   �      �       R|      �       R                       �      �       Y�      �       �U#|      �       Y�      �       �U#                  �      �       1�|      |       1�|      �       	��                      �      �       Y�      �       �U#|      |       Y|      �       y ��      �       �U#�                   �      �       R|      �       R                    �      �       P|      �       y @$t "�-r �-� ��      �       �U#@$t "�-r �-� �                   �      �       P|      �       y @$t "�-r �-� ��      �       �U#@$t "�-r �-� �                   �      �       Rb      |       R                       �      �       Z�      �       �U#b      l       Zl      |       �U#                  �      �       1�b      b       1�b      |       	��                      �      �       Z�      �       �U#b      b       Zb      l       z �l      |       �U#�                   �      �       Rb      |       R                    �      �       Pb      l       z @$t "�-r �-� �l      |       �U#@$t "�-r �-� �                   �      �       Pb      l       z @$t "�-r �-� �l      |       �U#@$t "�-r �-� �                   �             RC      b       R                       �             [             �U#C      L       [L      b       �U#                   �             1�C      C       1�C      b       	��                       �             [             �U#C      C       [C      L       { �L      b       �U#�                   �             RC      b       R                                     { @$t "�-r �-� �             �U#@$t "�-r �-� �             PC      L       { @$t "�-r �-� �L      b       �U#@$t "�-r �-� �                                  PC      L       { @$t "�-r �-� �L      b       �U#@$t "�-r �-� �                               Y       UY      �       S�      9       �U�9      A       U                             V       TV      9       [9      A       T                             ;       Q;      9       �Q�9      A       Q                  }      �      	 w ��"�                  �      �       v ��"�                  �      �      	 ���@"�                                    ~ p "�      6       ^6      9       {                              ;       q @$�;      b       Qb      9       Z9      A       q @$�                    �      �       r z ��             R                               4       T�      �       T�             TY      d       Tq      �       T�      �       T                                                X      A       u�      �       X�      �       u�      �       X�             uY      q       uq      |       X|      �       u�      �       X�             u                 `      �       X                 `      �       T                `      �       X                `      �       T                   r      �       R�      �      
 r { "#���                  r      �       r ?&��      �       [                �      �       Y                �      �       Q                �      �       Y                �      �       Q                  �      �       P�      �      
 p z "#���                  �      �       p ?&��      �       Z                    �      �       RI      o       R       )       R�      �       R                        �      �       Q�      �       uI      S       QS      o       u       )       u�      �       u                    �      �       1�I      I       1�I      o       	��       #       	��#      )       1��      �       1��      �       	��                          �      �       Q�      �       uI      I       QI      S       q �S      W       QW      o       u�       )       u��      �       u                       �      �       RI      o       R               R       )       r ��      �       R�      �       r ��      �       Z                              �      �       q { "�-r �-� ��      �       u@${ "�-r �-� �o      �       P�      �       u)      /       q { "�-r �-� �/      9       u@${ "�-r �-� ��      �       P                 �      �       q { "�-r �-� �o      o       P)      )       q { "�-r �-� ��      �       P                   �             Rs      �       R�      �       R9      Y       R                           �      �       Y�             us      �       Y�      �       u�      �       Y�      �       u9      F       YF      Y       u                   �             1�s      |       1�|      �       	���      �       1��      �       1��      �       	��9      B       1�B      Y       	��                            �      �       Y�             us      |       Y|      �       y ��      �       u��      �       Y�      �       y ��      �       u�9      B       YB      F       y �F      Y       u�                    �      �       R�      �       R9      Y       r �                             P�      �       Y                           $       R�      �       R�      �       Rq      �       R�      �       R                                            X      $       u�      �       X�      �       u�      �       X�      �       uq      |       X|      �       u�      �       X�      �       u                           $       1��      �       1��      �       	���      �       1�q      q       1�q      �       	���      �       1��      �       	���      �       1�                                              X      $       u�      �       X�      �       x ��      �       u��      �       X�      �       uq      q       Xq      |       x �|      �       u��      �       X�      �       x ��      �       u�                $      $       P�      �       P                       '      =       R�             RY      q       R�      �       R�             R                       '      4       T�             TY      d       T�      �       T�      �       T                       '      =       1��             1�Y      Y       1�Y      q       	���      �       1��      �       	���      �       1��             	��                       '      4       T�             TY      Y       TY      d       t ��      �       T�      �       t ��      �       T�      �       t �                      �      �       U�      9       �U�9      A       U                     q      |      $ s  "#��@& $ &{ ~ "#��@& $ &"�|      �       s @& $ &{ ~ "#��@& $ &"��      �       s @& $ &{ @& $ &"�                     �      �      $ s x "#��@& $ &r u "#��@& $ &"��      �       x @& $ &r u "#��@& $ &"��             x @& $ &r @& $ &"�                              t                               u                                 t       C       X                              u                    8      f       Sf      f      
 s  "#���                  8      f       s ?&�f      f       _                f      q       t                f      q       u                f      q       t                f      q       u                  f      q       [q      q      
 { ~ "#���                  f      q       { ?&�q      q       ^                q      q       t                q      q       t                q      q       t                q      q       u                q      q       t                q      q       u                q      q       Yq      q      
 p y "#���                q      q       P                q      q       u                q      q       t                 q      q       u                q      q       Xq      q       x w "#���                q      q       x ?&�                �      �       t                �      �       �U#                �      �       t                �      �       �U#                q      �       t                  q      �       u�      �       �U#                !q      �       t                !  q      �       u�      �       �U#                   �      �       R�      �      
 r u "#���                  �      �       r ?&��      �       U                �      �       t                �      �       �U#                �      �       t                �      �       �U#                  �      �       P�      �      
 p v "#���                  �      �       p ?&��      �       V                             3       U3      8       u �8      v       �U�                             @       T@      E       YE      E       t �E      v       �T�                             M       QM      R       XR      R       q �R      v       �Q�                              3       1�3      8       	��8      B       RB      E       r �E      O       RO      R       r �R      v       R                        v       U                      #      @       T@      E       YE      v       T                        &      M       QM      R       XR      a       Qa      v       X                    h      u       Pu      v       q �                   h      u       Pu      v       q �                      0m      ;m       U;m      Dm       u Dm      Jm       �U�                    0m      Dm       TDm      Jm       �T�                                    0�      ��       U��      ��       S��      ��       �U���      ȅ       Sȅ      х       Uх      ҅       �U�҅      ޅ       Uޅ      ��       S��      �       �U��      &�       U                                      0�      ��       T��      ��       ]��      ��       �T���      ��       T��      ͅ       ]ͅ      х       Tх      ҅       �T�҅      ޅ       Tޅ      �       ]�      �       �T��      &�       T                                        0�      |�       Q|�      ��       V��      ��       �Q���      ��       Q��      Ʌ       VɅ      х       Rх      ҅       �Q�҅      ޅ       Qޅ      ��       V��      �       R�      �       �Q��      &�       Q                                        0�      ��       R��      ��       \��      ��       �R���      ��       R��      ˅       \˅      х       Xх      ҅       �R�҅      ޅ       Rޅ      ��       \��      �       T�      �       �R��      &�       R                    r�      ��       P��      ��       P                    ��      ��       Pޅ      �       P                     ޅ      ��       S��      �       u�~��      �       �U�                     ޅ      ��       V��      �       R�      �       �Q�                 ޅ      �       1�                     ޅ      ��       \��      �       T�      �       �R�                             M       QM      P       q���}�P      �       Q�      �       q�����      �       Q                    n      �       R�      �       R                                        #      6       R6      C       PC      F       RF      P       r �P      _       P_      w       Sz      �       S�      �       S�      �       u �      �       R�      �       S�      �       R�      �       P�      �       S�      �       R                                &      6       P6      C       [C      P       PP      S       RS      �       [�      �       P�      �       p ��      �       R�      �       P                               6      C       PC      _       Pw      �       S�      �       S�      �       u �      �       S�      �       P�      �       S                    n      �       X�      �       X                        n      t       p 3$ �F     "�t      z       p3$ �F     "�z      �       p3$(�F     "��      �       p 3$ �F     "��      �       p3$ �F     "��      �       p3$(�F     "�                                 :      ^       Sa      �       S�      �       sx��      �       S�      �       t �      �       ���}��      �       S�      �       S�      �       t                     :      P       Ra      �       R                                                  [       +       Q:      :       [:      G       { z "�G      ^       [a      t       [t      {       { z �{      �       [�      �       P�      �       [�      �       p ��      �       P�      �       { ��      �       [                                  +       Q:      ^       Qa      �       Q�      �       P�      �       p ��      �       [�      �       P�      �       Q                        G      ^       [{      �       [�      �       P�      �       [                      :      ^       Xa      �       X�      �       X                        :      D       p 3$ �F     "�D      J       p3$ �F     "�J      V       p3$(�F     "�a      x       p 3$ �F     "�x      ~       p3$ �F     "�~      �       p3$(�F     "�                              :       Y:      @       u D      R       YR      X       u                               =       X=      @       t D      U       XU      X       t                       +      5       Oq �5      D       q~�D      O       Oq �O      [       R[      \       P                            `      �       U�      .       �U�.      6       U6      |       �U�|      �       U�      �       �U�                                    `      �       T�              S       .       �T�.      6       T6      W       SW      b       �T�b      r       Sr      |       �T�|      �       T�      �       S                                        `      �       Q�      &       \&      -       T-      .       �Q�.      6       Q6      Z       \Z      a       Ta      b       �Q�b      u       \u      |       �Q�|      �       Q�      �       \                                        `      �       R�      (       ](      -       Q-      .       �R�.      6       R6      \       ]\      a       Qa      b       �R�b      w       ]w      |       �R�|      �       R�      �       ]                            `      �       X�      .       �X�.      6       X6      |       �X�|      �       X�      �       �X�                            `      �       Y�      .       �Y�.      6       Y6      |       �Y�|      �       Y�      �       �Y�                  �      �       ��                        �      ,       _6      `       _b      {       _�      �       _                                    �      �       R�      (       ](      -       Q-      .       �R�6      \       ]\      a       Qa      b       �R�b      w       ]w      |       �R��      �       ]                                    �      �       Q�      &       \&      -       T-      .       �Q�6      Z       \Z      a       Ta      b       �Q�b      u       \u      |       �Q��      �       \                                �      �       T�              S       .       �T�6      W       SW      b       �T�b      r       Sr      |       �T��      �       S                        �      �       U�      .       �U�6      |       �U��      �       �U�                       �      *       ^6      ^       ^b      y       ^�      �       ^                        �      $       V6      X       Vb      s       V�      �       V                    �             P6      D       P                                P6      D       P                      �      �       T�      /       �T�/      6       T                      �      �       Q�      /       �Q�/      6       Q                      �      �       R�      /       �R�/      6       R                  �      /       U                 �      �       0�                     �      �       @��             @�      /       @�                     �      �       U�             U      /       U                           �      �       P�      �       t �      �       tx�      �       P�             t       /       t                      �      �       1��      �       1��      �       1��             	��             1�      /       	��                        �      �       P�      �       t �      �       P�      �       p ��             t �      /       t                    �      �       U�      �       u ��             U             U      /       u �                    �      �       @��             @�      /       @�                           �      �       p 6%��      �       p 6%��      �       P             P             p �-      /       P                   �      �       P             P-      /       P                        @      �       U�      %       �U�%      1       U1      D       �U�                    @      �       T�      D       �T�                    @      \       Q\      D       Z                          �      �       0��      �       u��             U             u�1      D       U                      x      �       Y�      �       y 	���      D       Y                        �      �       X�      �       x`��      /       X1      D       X                       �      �       tP��             tp�             tP�1      D       tp�                        P      f       Uf      �       �U��      �       U�      �       �U�                   m      �       U�      �       R                   m      �       R�      �       R                     m      |       U|      �       Y�      �       R                     m      |       R|      �       X�      �       R                  _      �       P                  m      �       Z                      �      �       Q�      �       p �      �       pp                  �      �       Q                        �      �       U�      �	       \�	      �	       �U��	      �	       \                          �      �       T�      �       U�      �	       [�	      �	       �T��	      �	       [                        �      �       Q�      �	       V�	      �	       �Q��	      �	       V                          �	      �	       C��	      �	       P�	      �	       C��	      �	       P�	      �	       C�                         S	      �	       R�	      �	       R�	      �	       q�	      �	       R�	      �	       R                        [	      �	       S�	      �	       Q�	      �	       S�	      �	       S                  �      �       W                      �      �       T�      �       U�      �       [                 �	      �	       ��                   �	      �	       ltuo�                 �	      �	       \                    �	      �	       Q�	      �	       S                 �	      �	       0�                      �	      �	       R�	      �	       q�	      �	       R                     
      W
       TW
      �
       �T�                         _
      o
      $ x z "#��@& $ &r t "#��@& $ &"�o
      s
       p @& $ &r t "#��@& $ &"�s
      ~
      $ x z "#��@& $ &r t "#��@& $ &"�~
      �
       x z "#��@& $ &p @& $ &"��
      �
      $ x z "#��@& $ &r t "#��@& $ &"�                  
      
       t                   
      
       u                   
      
       t                     
      
       u 
      #
       R                   
      *
       P*
      *
      
 p s "#���                  
      *
       p ?&�*
      *
       S                *
      =
       t                *
      =
       u                *
      =
       t                *
      =
       u                  *
      =
       Y=
      =
      
 y { "#���                  *
      =
       y ?&�=
      =
       [                =
      I
       t                =
      I
       t                  =
      I
       XI
      I
      
 x z "#���                	  =
      I
       x ?&�I
      I
       Z                  I
      W
       tW
      _
       �T#                I
      _
       u                  I
      W
       tW
      _
       �T#                I
      _
       u                  I
      _
       R_
      _
      
 r t "#���                  I
      _
       r ?&�_
      _
       T                    �
      �
       U�
      �
       �U�                      �
      �
       T�
      �
       \�
      �
       �T�                  �
      �
       S                  �
      �
       V                 �
      �
       \                 �
      �
       S                      �
      �
       T�
      �
       Q�
             �T�                            1       U1      �       \�      �       �U�                            +       T+      �       ^�      �       �T�                         1       0�1      k       S                  <      �       V                <      o       V                 <      `       v                 <      `       v                  O      o       _                 a      o       V                 a      o       _                 �      �       |�                  �      �       ^                  �      �       P                  �             P                  �             Q                            2       U2      |       _|      }       �U�                            2       T2      _       ]_      }       �T�                            2       Q2      _       V_      }       �Q�                            2       R2      _       ^_      }       �R�                     $      W       SW      Y       TZ      Z       0�Z      s       S                  <      _       \                 <      M       s                   N      W       SW      Y       T                 N      Z       V                      �      �       U�      �       u ��             �U�                      �      �       T�      �       Y�      �       t ��             �T�                      �      �       Q�      �       X�      �       q ��             �Q�                       �      �       1��      �       	���      �       R�      �       r ��      �       R�      �       r ��             R                 �              U                      �      �       T�      �       Y�             T                          �      �       Q�      �       X�             Q             P             X                                 P             q �                                P             q �                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  �      �       T�      �       �T�                �      �       U                   �      �       T�      �      
 p t "#���                  �      �       t ?&��      �       P                      �      �       U�      �       u ��      �       �U�                     �      �       1��      �       	���      �       X�      �       x ��      �       X                 �      �       U                    �      �       T�      �       R                    �      �       P�      �       q �                   �      �       P�      �       q �                    �      �       U�      �       �U�                  �      �       U                 �      �       0�                 �      F       u�                 �      F       u� �                        `      p       Up      �       S�      �       T�      �       �U�                    l      �       V�      �       U                     q      �       S�      �       T�      �       �U�                   q      �       V�      �       U                      �      �       U�      �       �U��      �       U                              �       �        U�       �        S�       �        T�       �        �U��       �        S�       �        �U��       !       U                            �       �        T�       �        V�       �        �T��       �        V�       �        �T��       !       T                      �       �        \�       �        U�       �        \                   �       �        U�       �        S                     �       �        S�       �        T�       �        �U�                   �       �        \�       �        U                        !      B!       UB!      a!       Sa!      b!       �U�b!      t!       U                   /!      B!       u#�B!      D!       s#�                 /!      D!       T                   /!      B!       u#�B!      D!       s#�                    O!      a!       Sa!      b!       �U�                      �)      �)       U�)      �)       �U��)      �)       U                      �)      �)       T�)      �)       �T��)      �)       T                      �)      �)       Q�)      �)       �Q��)      �)       Q                      �/      �/       U�/      �/       �U��/       0       U                        �/      �/       T�/      �/       �T��/      �/       T�/       0       �T�                        �/      �/       T�/      �/       �T��/      �/       T�/       0       �T�                      �/      �/       U�/      �/       �U��/       0       U                     �/      �/       u�#�/      �/      	 �U#�#�/      �/       u�#                        `5      |5       U|5      �5       S�5      �5       �U��5      �5       U                      `5      ~5       T~5      �5       �T��5      �5       T                     `5      5       0�5      �5       P�5      �5       0�                 y5      ~5       P                   �<      �<       T	=      =       T                   �<      �<       V�<      =       V                     �<      �<       T�<      �<       S�<      =       S                    ?      Z?       R]?      q?       R                      =?      H?       PH?      Q?       rQ?      Z?       P]?      q?       P                        `@      �@       U�@      �@       V�@      �@       �U��@      �@       U                        `@      �@       T�@      �@       \�@      �@       �T��@      �@       T                          `@      �@       Q�@      �@       �Q��@      �@       Q�@      �@       �Q��@      �@       Q                     `@      �@       0��@      �@       P�@      �@       0�                  �@      �@       �Q�                  �@      �@       \                  �@      �@       V                     �@      �@       0��@      �@       P�@      �@       0�                    �@      �@       P�@      �@       v                  �@      �@       S                  �@      �@       ]                      �E      F       UF      F       �U�F      F       U                      �E      F       TF      F       �T�F      F       T                      �E      F       QF      F       �Q�F      F       Q                      �E      F       RF      F       �R�F      F       R                      �E      F       XF      F       �X�F      F       X                    �E      F       XF      F       �X�                    �E      F       RF      F       �R�                    �E      F       QF      F       �Q�                    �E      F       TF      F       �T�                    �E      F       UF      F       �U�                   �E      F       UF      F       �U�                 �E      F       u�                       M      .M       U.M      /M       �U�/M      1M       U                    @M      UM       UUM      oM       �U�                     NM      UM       0�UM      [M       RiM      nM       R                  NM      nM       P                      PN      cN       UcN      dN       �U�dN      �N       U                      PN      cN       TcN      dN       �T�dN      �N       T                      PN      cN       QcN      dN       �Q�dN      �N       Q                       O      O       TO      O       �T�O      O       T                       O      .O       U.O      /O       �U�/O      1O       U                       O      .O       T.O      /O       �T�/O      1O       T                      �Y      �Y       U�Y      �Y       �U��Y      �Y       U                          �Y      
Z       U
Z      Z       SZ      Z       �U�Z      0Z       S0Z      2Z       �U�                            �Y      
Z       T
Z      Z       VZ      Z       �U#Z      &Z       T&Z      1Z       V1Z      2Z       �T�                              @Z      fZ       UfZ      xZ       VxZ      yZ       �U�yZ      �Z       U�Z      �Z       V�Z      �Z       �U��Z      �Z       U                          @Z      eZ       TeZ      yZ       �T�yZ      �Z       T�Z      �Z       �T��Z      �Z       T                        YZ      wZ       SwZ      xZ       vxZ      yZ       �U#yZ      �Z       S                            YZ      fZ       UfZ      xZ       VxZ      yZ       �U�yZ      �Z       U�Z      �Z       V�Z      �Z       �U�                 YZ      �Z       0�                    0[      >[       U>[      ?[       �U�                      0[      :[       T:[      >[       Q>[      ?[       �T�                      0[      6[       Q6[      >[       R>[      ?[       �Q�                      `]      z]       Uz]      �]       S�]      �]       �U�                   k]      z]       u8z]      |]       P                  n]      |]       T                    n]      z]       u8z]      |]       P                            pd      �d       U�d      �d       S�d      �d       �U��d      �e       S�e      �e       �U��e      �e       S                          pd      �d       T�d      �d       V�d      �d       �T��d      �d       V�d      �e       �T�                            pd      �d       Q�d      �d       \�d      �d       �Q��d      �e       \�e      �e       �Q��e      �e       \                 pd      �e       �Av  �                 pd      �e       �'v  �                    �d      �d       P�d      �d       P                   pd      �d       0��d      �d       0�                      e      e       Pe      e       ^�e      �e       ^                      e      e       0�e      e       ]�e      �e       ]                    We      le       P�e      �e       P                  �e      �e       V                     pd      �d       0��d      e       0��e      �e       0�                   �d      �d       @��e      �e       @�                   �d      �d       S�e      �e       S                    �d      e       V�e      �e       V                      �d      �e       S�e      �e       �U��e      �e       S                   e      5e       8�he      e       8�                   e      5e       She      e       S                   e      =e       Vpe      e       V                   e      =e       Spe      e       S                  e      =e       0�pe      e       0�                     f      #f       U#f      Ff       �U�                         f      7f       T7f      ;f       U;f      <f       �T�<f      Ff       T                       f      2f       Q2f      <f       �Q�<f      Ff       Q                       f      ;f       R;f      <f       �R�<f      Ff       R                       f      ;f       X;f      <f       �X�<f      Ff       X                      �j      �j       T�j      �j       �T��j      �j       T                       o      o       Uo      1o       S1o      3o       �U�                       o      	o       T	o      2o       V2o      3o       �T�                    o      o       0�o      0o       P                                    p�       �       U �      ��       \��      ��       U��      ��       �U���      ��       \��      ��       �U���      ��       U��      �       \�      #�       u�~�#�      $�       �U�                                      p�      ��       T��      <�       S<�      ��       �T���      ��       S��      ��       �T���      ��       S��      ��       �T���      ׄ       Sׄ      ��       T��      �       S�      $�       �T�                                        p�      ��       Q��      /�       _/�      ��       �Q���      ��       _��      ��       �Q���      ��       _��      ��       �Q���      ׄ       _ׄ      ��       Q��      �       _�      #�       Q#�      $�       �Q�                                        p�      ��       R��      '�       ]'�      ��       �R���      ��       ]��      ��       �R���      ��       ]��      ��       �R���      ׄ       ]ׄ      ��       R��      �       ]�      #�       R#�      $�       �R�                                        p�      ��       X��      <�       V<�      ��       �X���      ��       V��      ��       �X���      ��       V��      ��       �X���      ׄ       Vׄ      �       X�      �       V�      #�       T#�      $�       �X�                         ��      ��       P��       �       u  �      �       | ��      ��       u ��      ׄ       u                                 ��      ��       ^��      ��       ^��      ��       �T�Q"���      ׄ       ^��      �       ^�      �       �T "��      #�       �Tq "�#�      $�       �T�Q"�                                у      ��       X��      <�       V<�      ��       �X���      ��       V��      ׄ       V��      �       V�      #�       T#�      $�       �X�                            у      ��       ]��      ��       ]��      ׄ       ]��      �       ]�      #�       R#�      $�       �R�                              у      /�       _/�      ��       �Q���      ��       _��      ׄ       _��      �       _�      #�       Q#�      $�       �Q�                              у      ��       T��      <�       S<�      ��       �T���      ��       S��      ׄ       S��      �       S�      $�       �T�                              у       �       U �      ��       \��      ��       \��      ׄ       U��      �       \�      #�       u�~�#�      $�       �U�                           �      �       P�      <�       0�U�      k�       0�k�      w�       P��      ��       P��      #�       P                    �      �       P��      ׄ       P                     7�      U�       0�U�      ^�       1�^�      ��       0�                  7�      ��       _                       ��      ��       \��      �       \�      #�       u�~�#�      $�       �U�                       ��      ��       ]��      �       ]�      #�       R#�      $�       �R�                       ��      ��       _��      �       _�      #�       Q#�      $�       �Q�                       ��      ��       V��      �       V�      #�       T#�      $�       �X�                      ��      ��       U��      ˌ       �U�ˌ      �       U                      ��      ��       T��      ˌ       �T�ˌ      �       T                        ��      ��       Q��      ʌ       Sʌ      ˌ       �Q�ˌ      �       Q                       ��      ǌ       0�ǌ      ˌ       Rˌ      ݌       0�݌      �       R                       ��      ��       0���      ˌ       Pˌ      ݌       0�݌      �       P                                  p�      ��       U��      ˭       ]˭      �       �U��      ��       ]��      ��       ����      ��       �U���      ��       ]��      ��       ����      
�       �U�
�      s�       ��                          p�      ��       T��      ��       U��      
�       _
�      �       �T��      s�       _                        p�      ��       Q��      �       S�      �       �Q
���Q�Q0+( ��      s�       S                    p�      ��       R��      s�       ��                 p�      s�       �S �                 p�      s�       �F �                      ��      ��       P��      ��       } ��      s�       ��                	                    ��      ˭       0��      ��       0���      Ү       ^8�      L�       PL�      j�       ^j�      n�       ~�n�      ��       ^��      ��       0�ԯ      ܯ       ^ܯ      �       ~��      ��       ^
�      N�       ^O�      s�       ^                
                        ��      ˭       0��      ��       0���      Ү       PM�      n�       Pn�      r�       pj�r�      ��       P��      ��       0�ԯ      �       P�      �       ph��      ��       P
�      �       P�      h�       [h�      w�       ���      &�       [O�      s�       P                        ��      ��       P��      ��       w ��      �       ���      s�       w                           ��      ˭       0��      ��       0�r�      ��       1���      ��       0��      ��       0�O�      a�       1�a�      s�       0�                               ��      ˭       0��      �       0��      ��       0���      ��       0���      ��       P��      �       V�      &�       0�&�      O�       VO�      s�       0�                          ��      í       �  �      �       �  �      ��       �  ��      ��       �  
�      �       �  O�      s�       �                            ��      í       �  �      �       �  �      ��       �  ��      ��       �  
�      �       �  O�      s�       �                            ��      í       �  �      �       �  �      ��       �  ��      ��       �  
�      �       �  O�      s�       �                            ��      í       S�      �       S�      ��       S��      ��       S
�      �       SO�      s�       S                            ��      ��       U��      í       _�      �       _�      ��       _��      ��       _
�      �       _O�      s�       _                              4�      <�       P<�      ��       \��      ��       ����      ��       \��      ��       ��
�      �       ��O�      s�       ��                            r�      ��       	����      ��       ]��      ��       ]
�      �       ]O�      W�       ]a�      i�       ]                                ��      í       P�      ,�       P��      Ү       \�      �       P�      ��       \��      ��       \
�      �       \O�      s�       \                          r�      ��       0���      ��       V��      ��       V
�      �       VO�      s�       V                   8�      j�       6���      ��       6�                   8�      j�       _��      ��       _                      @�      ��       V��      ��       ��      ��       V                    @�      ��       _��      s�       _                   @�      ��       0���      s�       0�                    �      �       4���      ԯ       4�                    �      �       _��      ԯ       _                    ��      8�       ^��      ԯ       ^                        ��      Ү       _��      ��       _��      ��       _
�      s�       _                       ��      Ү       0���      ��       0���      ��       0�
�      s�       0�                   ��      ��       T��      ��       U                ��      ��       0�                  ˭      ��       w ��      ��       w                   ˭      ��       _��      ��       _                  ˭      ��       0���      ��       0�                   N�      {�       ^�      &�       ^                   N�      {�       _�      &�       _                  N�      {�       0��      &�       0�                 ��      ̰       V                 ��      ̰       _                 &�      O�       V                 &�      O�       ��                      0�      7�       U7�      8�       �U�8�      A�       U                      0�      7�       T7�      8�       �T�8�      A�       T                    h�      ��       P��      ��       P                    �      %�       P7�      F�       P                     �      �       t�      6�       Q7�      F�       Q                  "�      6�       T                  "�      6�       U                      ��      θ       Uθ      ϸ       �U�ϸ      Ѹ       U                      ��      θ       Tθ      ϸ       �T�ϸ      Ѹ       T                      ��      θ       Qθ      ϸ       �Q�ϸ      Ѹ       Q                      ��      θ       Rθ      ϸ       �R�ϸ      Ѹ       R                        @E      fE       UfE      �E       S�E      �E       �U��E      BF       S                          @E      \E       T\E      fE       QfE      �E       V�E      �E       �T��E      BF       V                  �E      �E       0�=F      BF       P                   WE      �E       \�E      �E       \                      �E      F       ]F      F       }|�F      BF       ]                  �E      BF       \                            �      �       T�      )       Y)      2       T2      �       Y�      �       T�      �       Y                           �             0�      (       P)      P       0�P      �       P�      �       0��      �       P                               �             0�             P      )       X)      P       0�P      p       Pp      �       X�      �       0��      �       X�      �       P�      �       X                        �      �       T�             t�5      5       T5      X       t�X      p       t��      �       t��      �       t��      �       [                        �              Z5      M       r 1$x "�M      `       Z`      �      
 r 1$u�	"��      �       Z                    p:      z:       Uz:      :       �U�                 �      �       U                      �      �       U�      �       �U��      �       S                            �      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T�                    �      �       V�      �       V                   �      �       u� ��      �       s� �                I      _       u�                 I      _       v��0$0&�                   X      _       P_      _      
 p r "#���                  X      _       p ?&�_      _       R                w      �       u�                 w      �       v��0$0&�                   �      �       P�      �      
 p r "#���                  �      �       p ?&��      �       R                �      �       u�                    �      �       v��0$0&��      �      	 p 0$0&�                   �      �       X�      �      
 p x "#���                  �      �       x ?&��      �       P                �      �       s�                 �      �       v��0$0&�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                      p       x        Ux       �        S�       �        �U�                     p       x        Ux       �        S�       �        �U�                 �      �       U                      �      �       U�      h        Sh       j        �U�                     �      �       U�      h        Sh       j        �U�                 �      �       u                   �      i        V                         )      9)       U9)      �+       V�+      �+       �U��+      �+       V                     )      \)       T\)      �+       �T�                    2)      �+       ]�+      �+       ]                    �)      �+       \�+      �+       \                    �)      �+       P�+      �+       P                     =)      \)       0�\)      �)       R�)      �)       Q                    =)      Q)       UQ)      \)       v�6&�                \)      o)       q 2$y "                   h)      o)       Po)      o)      
 p t "#���                  h)      o)       p ?&�o)      o)       T                 �)      �)       Q                 �)      �)       R                 �)      �)       2�                 �)      �)       \                 �)      	*       3�                 �)      	*       \                 +      �+       V                 +      �+       \                 �+      �+       0��+      �+       1��+      �+       2�                 �+      �+       0�                 �+      �+       2�                 �+      �+       \                 �+      �+       |��                        �:      �:       U�:      �;       S�;      �;       �U��;      �;       U                       �:      �:       U�:      �;       S�;      �;       �U��;      �;       U                  �:      �;       ]                  �:      �;       V                  �:      �:       \                 �:      �:       S                 �:      �:       s�                 �:      ;       S                 �:      ;       \                 �:      ;       |8                        `�      ��       U��      ̥       ^̥      ;�       s���      ��       ^ի      �       s�                                  `�      ��       T��      B�       SB�      V�       �T�V�      �       S�      ի       �T�ի      �       S�      ܭ       �T�ܭ      �       S�      կ       �T�                    `�      ��       Q��      կ       ��~                                  `�      ��       R��      B�       \B�      V�       �R�V�      d�       \d�      ��       �R���      ��       \��      ի       �R�ի      �       \�      կ       �R�                                  `�      ��       X��      B�       ]B�      V�       �X�V�      u�       ]u�      ��       �X���      ��       ]��      ի       �X�ի      �       ]�      կ       �X�                                                             ��      ɥ       Pɥ      ̥       V̥      ץ       Pץ      >�       V>�      B�       PV�      w�       Pw�      ��       V��      �       V�      m�       ��~ܧ      X�       ��~��      �       P�      �       V�      �       0�:�      :�       0�P�      ��       V��      ��       ��~ƫ      Ϋ       PΫ      ի       Pի      ݫ       V�      ��       P��      �       ��~�      �       V�       �       P �      E�       VE�      Z�       P��      ��       Pܭ      �       V                 `�      b�       t�#                              ��      ��       P��      B�       _V�      ��       _��      ��       P��      �       _ի      �       _ܭ      �       _                                 `�      ��       T��      B�       SB�      V�       �T�V�      �       S�      ի       �T�ի      �       S�      ܭ       �T�ܭ      �       S�      կ       �T�                        W�      d�       Td�      ��       ��~�@%��      �       T�      &�       ��~�@%�                           V�      ��       S��      �       S�      ի       �T��      ܭ       �T�ܭ      �       S�      կ       �T�                         ��      �       S�      X�       �T���      ��       �T���      �       �T�ܭ      �       S                           �      Q�       0�ܧ      �       0��      X�       V��      ��       Vt�      ��       0���      �       V                             �      �       0��      m�       ��~ܧ      X�       ��~��      ��       ��~��      ��       ��~��      �       ��~ܭ      �       0�                           �      �       0��      m�       ��~ܧ      X�       ��~��      ��       ��~��      �       ��~ܭ      �       0�                             �      �       0��      m�       ��~ܧ      �       ��~�      X�       ��~��      ��       ��~��      �       ��~ܭ      �       0�                             �      �       0��      W�       ��~\�      m�       Pܧ      X�       ��~��      ��       ��~��      �       ��~ܭ      �       0�                 �      �       0�                  �      ��       X                   ��      t�       ��~��      �       ��~                     ��      6�       S6�      `�       ��~��      �       S                            ۩      �       \�      �       |��      �       \�      4�       ��~4�      ;�       P��      �       \                   ֩      h�       ]��      �       ]                    �      ��       P��      �       P                       ۩      ��       0���      ;�       V;�      `�       S��      �       0�                        �      ;�       3�;�      M�       VM�      T�       v�T�      [�       V                       `�      ��       S��      ƫ       S�      
�       SZ�      ��       S                        v�      ��       \��      ƫ       \�      
�       \Z�      ��       \                        m�      ��       0���      ��       T��      ��       Q��      ��       T                         �      �       p 
����      G�       ZG�      ��       ��~�      �       p 
���Z�      r�       Z                        �      ��      , ��H$��@$!��8$!��!�������      �      	 ~ ������      «       ^�      �      � �H0H%�$!0)( 8/��
���H0H%�$!0)( 8/���H0H%�$!0)( 8/����������+( �����Z�      ��       ^                          ͪ      ͪ       _ͪ      ͪ       �ͪ      �       ��      ��       ���      ��       x r "���      ��        r "#���      ��       x r "��      
�       �Z�      ��       �                      ͪ      G�      	  ��~"�G�      ��        ��~"��      �      	  ��~"�Z�      r�      	  ��~"�                 ̨      �       S&�      E�       S                    �      �       P�      �       0�&�      B�       PE�      E�       P                	 �      :�       S��      ��       S                    �      :�       P:�      :�       0���      ��       P��      ��       P                 L�      L�       0�                      +�      B�       0�B�      ��       ^��      կ       ^                        +�      B�       0�B�      m�       ]s�      ��       ]��      կ       ]                          +�      B�       0�B�      `�       \`�      s�       |�s�      ��       \��      ��       1���      կ       1�                  ��      ǯ       P                 d�      ��       S                      
�      �       S��      ܭ       S�      �       S��      ��       S                           ,�      C�       PC�      q�       Vq�      ��       P�      �       P��      ܭ       PJ�      `�       V                          ��      ��       2���      ì       R�      �       1���      ��       2���      ʮ       1�ʮ      �       R                      �      �       T�      J�       ]`�      ��       ]                   �      J�       V`�      ��       V                    �      J�       \`�      ��       \                    �      5�       P`�      �       P                       �      �       �����      �       R�      J�       Rt�      ��       R                   �      �       0��      ,�       T                  �      ,�       Q                      �             U      t       St      {       �U�                  �      z       V                                                                    ж      *�       U*�      *�       _*�      V�       UV�      4�       _4�      5�       �U�5�      ��       _��      1�       U1�      A�       _A�      ��       U��      ��       _��      ��       U��      ��       _��      �       U�      ��       _��      ��       U��      P�       _P�      w�       Uw�      ��       _��      ��       U��      ��       _��      �       U�      ��       _��      ��       U��      �       _�      (�       U(�      ��       _                             ж      _�       0�_�      0�       ]5�      ��       ]��      1�       0�1�      A�       ]A�      ��       0���      ��       ]                  8�      M�       T                      F�      P�       0�P�      X�       QX�      d�       q�                                                                                            �      =�       Vù      ι       Vι      Թ      
 83$0"���      ̻       V��      ̼       V�      b�       V^�      v�       V�      �       V�      <�       q 3$x "�<�      E�      	 83$x "���      ��       V��      ,�       V��      q�       V��      �       Vi�      ��       Vq�      �       V2�      ��       R��      ��       V��      ��      	 83$x "�N�      ��       V��      ��       q 3$x "���      ��      	 83$x "��      |�       V|�      ��      
 83$0"���      ��       V��      �       V&�      ��       V��      ��       V��      ��       V�      �       V8�      9�       VV�      o�      	 83$x "�u�      ��       V��      �       VQ�      {�       R{�      ��       Vp�      ��       V��      ��      	 83$x "�                                                                                                                                                                                                                      �      =�       �ù      Թ       ���      ǻ       ���      ��       ���      ̼       ��      /�       �9�      B�       �P�      O�       �^�      n�       ��      ��       ���      ��       �ѿ      �       �+�      7�       �L�      c�       �t�      ��       ���      #�       �7�      M�       �[�      q�       ���      ��       ���      ��       ��      
�       ��      E�       ���      ��       ���      �       �5�      O�       �]�      b�       �s�      ��       ���      ��       ���      ��       ���      ,�       ���      %�       ���      ��       ���      ��       ���      /�       ���      �       ���      ��       ��      <�       ���      �       �i�      y�       ���      ��       �q�      ��       ���      P�       ���      ��       ��      9�       ���      ��       ���      ��       ���      �       �'�      ��       �2�      2�       �2�      ��       	����      ��       �N�      ��       ���      �       ��      ��       ���      ��       ���      �       �)�      :�       �w�      ��       ���      ��       ���      ��       ���      ��       ��      &�       �7�      K�       �\�      {�       ���      ��       ��      ��       �N�      `�       �q�      ��       ��      L�       �]�      ��       ���      ��       ��      .�       �@�      O�       �j�      ��       ���      ��       ���      t�       ���      �       �&�      ;�       �@�      j�       �~�      ��       ���      ��       ���      ��       ��      �       �8�      \�       ���      ��       ���      ��       ���      V�       �y�      ��       ���      ��       ���      U�       ���      �       �(�      3�       �V�      o�       �u�      ��       ���      �       �Q�      {�       	����      @�       �~�      ��       ���      ��       �}�      ��       ���      ��       �                 ��      ��       V                         ��      q�       _��      ��       _��      �       _�      8�       _��      ��       _                         ��      q�       V��      ��       V��      �       V�      8�       V��      ��       V                       ��      ��       1���      ��       S��      q�       S��      ��       S                      ��      ��       T��      g�       T��      ��       T                      �      ,�       P,�      7�       ��
��p "�7�      I�       P��      ��       P                            ��      ��       P��      q�       \��      ��       \��      �       \�      8�       \��      ��       \                                 ��      ��       r 3$p "��      �       r 3$p "�      ?�       r 3$0"?�      B�       q 3$0"B�      M�       ux�M�      S�       US�      W�       QW�      a�       q 6��
������$�a�      g�        p pp0*( 6��
������$���      ��       r 3$0"                   �      '�       Vy�      ��       V                   �      '�       _y�      ��       _                      �      '�       Py�      ��       P��      ��       v                        ��      �       V��      M�       V��      ��       V}�      ��       V                       ��      �       _��      M�       _��      ��       _}�      ��       _                       ��      �       v��      @�       v��      ��       v}�      ��       v                          ��      ��       P��      �       v ��      @�       v ��      ��       v }�      ��       v                                       5�      =�       0���      ��       Q
�      �       P�      �       Q.�      @�       0�D�      H�       PH�      M�       Q��      ��       P��      ��       Q��      ��       P��      ��       Q                      ��      ��       P��      @�       v �
��4$� "�}�      ��       P                      ��      ��       Q��      @�       v�
��4$�"�}�      ��       v�
��4$�"�                ��      �       Y                      ��       �       t z � �      �       P�      �       t z ��      �       v �
��4$� "�z �                   �      �       P�      �      
 p t "#���                  �      �       p ?&��      �       T                  �       �       Q �       �      
 q r "#���                  �       �       q ?&� �       �       R                ��      ��       �                 ��      ��       P                   ��      ��       P��      ��      
 p q "#���                  ��      ��       p ?&���      ��       Q                  ��      ��       P                  ��      ��       R                 ǹ      ι       _                 ǹ      ι       V                   ;�      ��       RQ�      {�       R                   ;�      ��       _Q�      {�       _                    >�      ��       XQ�      {�       X                     >�      l�       ql�      ��       TQ�      {�       T                          [�      l�       0�l�      o�       p�o�      {�       P{�      ��       p�Q�      f�       0�                     ��      ��       V8�      ��       VM�      ~�       V                     ��      ��       _8�      ��       _M�      ~�       _                    ~�      ��       Zy�      ~�       Z                       ~�      ��       0���      ��       Y��      ��       y���      ��       Y                 �      %�       V                 �      %�       _                 y�      ��       V                 y�      ��       _                 P�      b�       V                   P�      ^�       _��      p�       _                	 P�      O�       v                 
 P�      O�       v                 P�      O�       v                    ]�      ��       X��      O�       v                   ]�      ��       Q��      O�       v                     y�      ^�       V��      p�       V                          ��      ��       ��~p "���      ޾       ��~u "�޾      �       P�       �       ��~u "���      ��       ��~u "�                 4�      9�       r ��~�                     4�      O�       | �s "#�O�      K�       | ��~���      �       | ��~�                      4�      O�       UO�      ^�       ��~��      p�       ��~                 4�      K�       ��~                 ��      �       ��}                      �      O�       y | �O�      K�       ��~| ���      ��       ��~| �                  #�      p�       \                 ^�      n�       _                 ��      ��       _                  ��      ��       V                 ��      ѿ       _                  ��      ѿ       V                 ѿ      �       _                 ѿ      �       V                ѿ      �       �                ѿ      �       v                    �      �       Q�      �      
 q r "#���                  �      �       q ?&��      �       R                 �      �       _                 �      �       V                 �      +�       _                  �      +�       V                 +�      L�       V                    /�      ?�       P?�      L�       v                 L�      [�       _                 [�      t�       V                 t�      ��       _                  �      ��       P                  ��      ��       R                 t�      ��       �                 ��      ��       V                 ��      ��       _                  ��      ��       T��      ��       P                   ��      ��      	 p 0$0&���      ��       U                   ��      ��      	 t 0$0&���      ��       T                     ��      ��       ����      ��       Q��      ��       ��                   ��      ��      	 t 0$0&���      ��       T                   ��      ��      	 p 0$0&���      ��       U                 ��      7�       V                 ��      7�       _                  �      �       T�      #�       P                   �      �      	 p 0$0&��      #�       U                   �      �      	 t 0$0&��      #�       T                     �      �       ���      #�       Q#�      7�       ��                   �      �      	 t 0$0&��      #�       T                   �      �      	 p 0$0&��      #�       U                 7�      [�       V                 7�      [�       _                 [�      ��       V                 [�      ��       _                 ��      ��       V                 ��      ��       _                    ��      ��       P��      ��       v                  ��      �       V                 ��      �       _                  ��      �       Q                   �      <�       q 3$x "�<�      E�      	 83$x "�                  �      ��       _                 �      ��       V                    S�      \�       P\�      c�       S                  c�      s�       R                     ��      ��       _V�      y�       _��      �       _                          ��      ��       Q��      ��       �� $ &5$�"���      ��       r $ &5$�"�V�      h�       Qh�      o�       �� $ &5$�"�                    X�      h�       qh�      y�       Q                  X�      y�       T                  X�      y�       _                   ��      �       V��      ��       V                   ��      �       _��      ��       _                       �      �       Q�      �       r� $ &3$ "#���      ��       Q��      ��       r� $ &3$ "#�                       �      �       P�      �       v ��      ��       P��      ��       v                    �      �       _��      ��       _                     
�      �       q p "��      �       P��      ��       p q ���      ��       P                 s�      ��       V                  w�      ��       Q                  �      ��       P                 �      ��       v                  5�      ]�       V                 5�      ]�       _                 ]�      s�       V                 ��      ��       V                 ��      ��       _                 ��      ��       _                 ��      R�       V                 ��      R�       _                  ��      R�       T                 ��      #�       v                            �      �      	 q  $ &��      �       R�      �      	 q  $ &��      �      
 q   $ &��      R�       1t�$ $ &�                 R�      s�       _                 s�      ��       V                 s�      ��       _                 ��      ��       V                 ��      ��       _                 ��      ��       _                 ��      ��       V                 ��      ��       _                 ��      ��       _                    ,�      ]�       Vi�      ��       V                    ��      ��       P��      ��       p �                   ��      ��       V-�      ��       V                   ��      ��       _-�      ��       _                     ��      ��       0���      ��       S-�      ��       S                  A�      ^�       P                   ��      ��       V��      ��       V                   ��      ��       _��      ��       _                    �      ��       [��      ��       [                    �      ��       Y��      ��       Y                      �      .�       PY�      ��       P��      ��       P                    ��      ��       z  $0.���      ��       z  $0.�                   ��      ��       V{�      ��       V                    ��      ��       _{�      ��       _                   ��      s�       S{�      ��       S                    \�      ��       P{�      ��       P                    s�      ��       Z��      ��       Z                       s�      ��       P��      ��       Y��      ��       y���      ��       Y                 ��      ��       _                    #�      6�       Pa�      ��       P                   ��      �       V~�      ��       V                   ��      �       _~�      ��       _                      ��      ��       x ����      �       U~�      ��       U                        ��      ��       1���      ��       P��      ��       p�~�      ��       1�                       �      q�       V��      ��       V��      ��       V��      ��       V                       �      ��       _��      ��       _��      ��       _��      ��       _                
     �      <�       v��      ��       v��      ��       v                            �      .�       P.�      ��       S��      ��       P��      ��       P��      ��       S��      ��       S                          G�      Z�       PZ�      ��       \��      ��       P��      ��       P��      ��       \                    q�      ��       P��      ��       V                	         �      <�       �<�      ��       ��}��      ��       ���      ��       ���      ��       ��}                     ~�      ��       | p ���      ��       | v ���      ��       R                 ��      �       V                 ��      i�       _                      ��      ��       x ����      �       U�      i�       x ��                 �      �       0�                   �      +�       _+�      U�       _                 i�      ��       V                 i�      ��       _                  u�      ��       V��      ��       V                   u�      ��       _��      ��       _                 ��      ��       V                       ��      ��       VC�      V�       V��      �       Vp�      }�       V                       ��      ��       _C�      V�       _��      �       _p�      }�       _                        ��      =�       T=�      _�       vC�      V�       T��      �       T                      N�      w�       Pw�      ��       r $ &5$�"�p�      }�       r $ &5$�"�                            ��      ��      	 t (q "���      ��       Q��      ��       r $ &5$�"#C�      V�       Q��      ��      	 t (q "���      �       t (�"�p�      }�       Q                    ��      �       UC�      V�       U                     t�      ��       q��      ��       Qp�      }�       q                   t�      ��       Tp�      }�       T                   t�      ��       _p�      }�       _                 ��      �       V                  ��      �       _                 ��      �       Q                   ��      ��       	����      �       R                 �      ��       V                 �      ��       _                  :�      T�       P                  	�      ��       S                   ��      ��       V��      ��       V                   ��      ��       _��      ��       _                      ��      ��       P��      ��       v ��      ��       v                       ��      ��       P��      ��       P��      ��       Q                 ��      ��       V                 ��      ��       _                  ��      ��       T                 ��      '�       V                 ��      '�       _                  �      �       T                     '�      �       V��      ��       V�      (�       V                       '�      ��       _��      �       U��      ��       _�      (�       U                      E�      �       Y��      ��       Y�      (�       Y                    P�      ��       R��      ��       R                     �      ��       V��      ��       V�      �       V                       �      ��       _��      ��       U��      ��       _�      �       U                   @�      ��       Q��      ��       Q                      1�      ��       Y��      ��       Y�      �       Y                    @�      ��       R��      ��       R                 ��      h�       V                 ��      h�       _                   ��      ��       0���      h�       P                  ��      h�       t�                       h�      ��       V��      ��      	 83$x "�V�      o�      	 83$x "���      ��      	 83$x "�                     h�      N�       _9�      u�       _��      ��       _                                        ��      ��       P��      ��       U�      1�       P1�      =�       U9�      >�       P>�      P�       UV�      ]�       P]�      o�       U��      ��       U��      ��       P��      ��       U��      ��       P                                    ��      ��       Q��      ��       P�      .�       Q.�      =�       P9�      >�       Q>�      P�       TV�      ]�       Q]�      o�       T��      ��       P��      ��       Q��      ��       P��      ��       Q                      ��      ��       Q.�      =�       Q��      ��       Q��      ��       Q                       h�      ��       v��      ��      
 83$x "#V�      o�      
 83$x "#��      ��      
 83$x "#                          t�      ��       Q��      ��       v ��      ��       83$x "V�      o�       83$x "��      ��       83$x "                       h�      ��       �%�      (�       SV�      o�       ���      ��       �                        ��      ��       T��      ��       �| "�V�      o�       �| "���      ��       �| "�                        ��      ��       Q��      ��       �v "�V�      o�       �v "���      ��       �v "�                            ��      ��       ��1�      =�       ��>�      V�       ��]�      u�       ����      ��       ����      ��       ����      ��       ����      ��       ��                      ��      ��       P]�      o�       T��      ��       P��      ��       Q                      ��      ��       U]�      o�       U��      ��       U��      ��       P                      ��      N�       \9�      V�       \��      ��       \                      �      N�       V9�      V�       V��      ��       V                      1�      =�       ��>�      V�       ����      ��       ����      ��       ��                      1�      =�       P>�      P�       T��      ��       P��      ��       Q                      1�      =�       U>�      P�       U��      ��       U��      ��       P                 R�      ^�       _                 R�      ^�       V                 ^�      y�       _                     ��      ��       V�      -�       V��      ��       V                     ��      ��       _�      -�       _��      ��       _                      �      k�       Rk�      ��       v �      -�       R                      ��      ��       Q��      ��       r $ &5$�"���      ��       r $ &5$�"�                          �      '�      	 r (p "�'�      ��       P�      (�      	 r (p "�(�      -�       r (�"���      ��       P��      ��       r $ &5$�"#                  1�      Z�       T                    ��      ��       p��      ��       Q��      ��       p                  ��      ��       T��      ��       T                  ��      ��       _��      ��       _                 ��      ��       V                 ��      ��       V                 �      )�       V                   )�      w�       V��      ��       V                     )�      P�       _P�      w�       U��      ��       U                      :�      w�       Y��      ��       Y��      ��       y���      ��       Y                    :�      w�       0���      ��       0�                 w�      ��       V                 ��      ��       V                 ��      ��       V                 ��      �       V                 �      �       _                 �      "�       _                 "�      7�       V                 7�      \�       V                 \�      i�       V                 i�      q�       V                 '�      1�       V                 ��      ��       _                 ��      ��       V                 ��      ��       _                 ��      ��       V                 ��      ��       _                 ��      ��       V                      ��      ��       Y��      ��       y p ���      �       Y                   �      ��       V��      �       V                    �      ��       _��      �       _                   ��      �       V��      K�       V                    ��      �       _��      K�       _                   �      ��       V��      p�       V                    �      ��       _��      p�       _                 ��      ��       _                 ��      ��       _                     ��      N�       _@�      j�       _p�      ��       _                      ��      �       P1�      E�       PE�      H�       q 3$x "                 N�      \�       V                     q�      ��       V��      ��       q 3$x "���      ��      	 83$x "�                 q�      �       _                  u�      �       \                     u�      ��       v��      ��      	 q 3$x "#��      ��      
 83$x "#                      ��      ��       S��      ��       R��      �       s �                 �      ]�       V                 �      ]�       _                  �      ]�       Q                �      :�       �                �      :�       v                   ,�      :�       P:�      :�      
 p t "#���                  ,�      :�       p ?&�:�      :�       T                   ]�      '�       V��      ��       V                   ]�      '�       _��      ��       _                    d�      '�       R��      ��       R                 +�      F�       _                 +�      F�       V                   F�      ��       V�      C�       V                   F�      ��       _�      C�       _                  ��      ��       Q                  l�      ��       R                    n�      ��       Q��      ��       U                   ��      �       VK�      z�       V                   ��      �       _K�      z�       _                  ��      �       Q                  ��      �       R                    ��      ��       Q��      �       T                 �      �       _                 �      �       V                 �      @�       V                 �      @�       _                 @�      j�       V                 @�      j�       _                   n�      |�       Vu�      ��       V                    n�      |�       _u�      ��       _                   n�      |�       Ru�      ��       R                  ��      ��       S                 ��      ��       V                 ��      ��       V                   ��      �       _z�      ��       _                   ��      �       Vz�      ��       V                 �      �       V                 �      '�       _                 �      '�       V                 U�      ��       V                 U�      ��       _                  d�      ��       R                    t�      ��       P��      ��       p�                 ��      �       V                 ��      Q�       _                   ��      �       s�~��      Q�       s�                 �      �       0�                   �      �       _�      Q�       _                    �      }�       Q}�      ��       �� $ &5$�"#                    ��      C�       RC�      ��       ������53$�"�                    U�      p�       Pp�      ��       �� $ &5$�"�                   m�      }�       q}�      ��       Q                 m�      ��       T                 m�      ��       _                     �      V�       u�V�      _�       �A�      ��       u�                                                             �      V�       UV�      4�       _4�      5�       �U�5�      ��       _1�      A�       _A�      ��       U��      ��       _��      ��       U��      ��       _��      �       U�      ��       _��      ��       U��      P�       _P�      w�       Uw�      ��       _��      ��       U��      ��       _��      �       U�      ��       _��      ��       U��      �       _�      (�       U(�      ��       _                    MQ      �Q       P�Q      	R       P                        UQ      �Q       Q�Q      �Q       u������53$u�"��Q      �Q       Q�Q      	R       u������53$u�"�                  �Q      �Q       Q                     �Q      �Q       p�Q      �Q       Q R      	R       p                   �Q      �Q       T R      	R       T                     �Q      �Q       X�Q      �Q       U R      	R       U                            �      �       U�      |       S|      �       �U��             S             �U�      s       S                        �      �       T�      �       V�      j       �T�j      s       V                      �      �       ]�             ]      s       ]                           �      �       1��      :       \D      w       \�      �       \      j       \j      s       1�                          �      1       QU      w       Q�      �       Q�      �       Q      j       Q                                     T      )       s��
��t "�)      1       P�      �       P�      �       T                          �      �       P�      w       ^�             ^      j       ^j      s       P                                     �             u 3$p "      1       u 3$s0"U      w       u 3$p "�      �       t 3$s0"�      �       rx��      �       R�      �       T�      �      / u 3$s0"?7u 3$s0"?8u 3$s0"?80*( ��      �       R�      �       u 3$s0"      j       R                              0�      ��       U��      .�       ^.�      m�       Um�      |�       �U�|�      ��       U��      9�       ^9�      N�       U                      m�      ��       @���      .�       ]|�      ��       8���      9�       ]                   ق      �       Z��             Z                    ق      .�       V��      9�       V                 ��      9�       S                       ��             S      �       _�      ��       R�      9�       _                            ��      ��       Z��      �       S�      .�       Z��      ��       S��             P      9�       \                       ��      ��       0���      �       Y�      .�       Y��             Y                            �       \1�      <�       \<�      A�       _                              �       _�      ��       R1�      8�       _8�      A�       t�                            ��       Q��      �       |�1�      A�       Q                          ��       T1�      A�       T                              �       ����      ��       U��      �       ���1�      A�       ���                  M�      ��       S                  M�      ��       _                  M�      ��       V                    M�      y�       Ty�      ��       
���                      M�      p�       ���p�      y�       Uy�      ��       ���                  ��             S                  ��             _                    ��      ��       Q��             s�                  ��      ��       Z                      ��      ��       �����      ��       U��             ���                   Ǆ      ܄       ����      9�       ���                    Ǆ      ܄       S�      9�       S                    Ǆ      ܄       V�      9�       V                      Ǆ      ܄       Z�      ��       Z��       �       z  �                          �      ��       Z��      
�       z  ��      %�       P%�      -�       p�-�      9�       P                      ք      ڄ      
 r u q "�ڄ      ܄       R�      9�       R                            @      �       U�      =       S=      G       �U�G      �       S�      �       �U��      P       S                          �             ���      �       ��"      �       ��0      5       PK      P       P                                   P�      �       ��"      �       ��                      �             \�      �       \      P       \                      �             V�      �       V      P       V                        {      �       1�l      �       0�      "       1��      P       0�                                    t u "#��@& $ &���            ( t u "#��@& $ &��q r "#��@& $ &��            M s��
��4$s�"�y  $ &s�� $ &u "#��@& $ &��q r "#��@& $ &��            u s��
��4$s�"�y  $ &s�� $ &s��
��4$s�"�y  $ &s�� $ &?&"#��@& $ &��q r "#��@& $ &��      *      � s��
��4$s�"�y  $ &s�� $ &s��
��4$s�"�y  $ &s�� $ &?&"#��@& $ &��s��
��4$s�"#�x  $ &s�� $ &r "#��@& $ &��                  �      �       U�             s�                    �      �       t y ��      �       T�             s��
��4$s�"�y �                   �             T            
 t u "#���                  �             t ?&�             U                               Q            
 q r "#���                               q ?&�             R                      �      �       _�      �       p 3$�U#0""      �       _                          r      �       P�      �       ^d      i       Px      �       R�      �       ^                      �      �       Px      �       P�      �       ��                       4      8       p t "#��@& $ &���8      @      ( p t "#��@& $ &��q u "#��@& $ &��@      H      + p ?&p "#��@& $ &��q u "#��@& $ &��H      O      I p ?&p "#��@& $ &��s�r "#�z  $ &s�� $ &u "#��@& $ &��O      [      j p ?&p "#��@& $ &��s�r "#�z  $ &s�� $ &s�r "#�z  $ &s�� $ &?&"#��@& $ &��                      4       [                                t p �      -       T                   &      4       P4      4      
 p t "#���                  &      4       p ?&�4      4       T                  4      8       Q8      8      
 q u "#���                  4      8       q ?&�8      8       U                        �      P       UP      (       S(      2       �U�2      �       S                    �             T      �       �T�                      �      /       ^/      2       �U#�2      �       ^                       �             t#�      P       t�2      Z      	 �T##�Z      j       t�                              [      �       ]�             ]j      x       ]x      {       P{      �       ]�      �       P�      �       ]                    �      �       P�      �       P                          V      [       P[      �       R�      �       ��j      �       R�      �       R                      &      -       P-             _j      �       _                 �      �       u�                 �      �       u�                       b      k       p r �k      {       P�      �       }  ��      �       P                   j      �       t 3�#<3$s "#�      �       t 3�#<3$s "#                         j      x       ]x      {       P{      �       ]�      �       P�      �       ]                   j      �       S�      �       S                        p      O       UO      �       S�      �       �U��      7       U                      p      C       TC      �       ���      7       T                            p      �       Q�      �       V�      �       �Q��      �       Q�      .       V.      7       �Q�                      p      O       RO      �       �R��      7       R                      p      O       XO      �       �X��      7       X                                                    �      �       Q��8�      �       Q�_��6�      �       Q�_�^�[��2�      �       Q�_�^�[�S�Y��(�      �       Q�_�^�[�u� �Y��(�      �       Q�_�^�[�u� �Y�Z�� �      �       Q�_�^�[����Y�Z�� �      -       r �_�^�[����Y�Z�� -      4       �_�^�[����Y�Z�� 4      O       �_�^�[����Y��(O      �       �_�^������0�      �       Q��8�      �       Q�_��6�      �       Q�_�^�[�����0�      �       Q�_�^�[����Y��(�      4       Q�_�^�[����Y�Z�� 4      6       Q�_��[����Y�Z�� 6      7       Q��[����Y�Z��                     �      1       P1      O       x              P                    e      i       Pi      �       ]                     
      3
       T3
      X
       �T�                     
      6
       Q6
      X
       �Q�                 
      I
       u��0$0&�                 
      I
       u��0$0&�                   
      B
       QB
      I
       �Q�                 
      I
       T                     >
      B
       RB
      I
       QI
      I
      	 p q "#�@�                  B
      I
       q ?&�I
      I
       P                    �	      �	       T�	      
       �T�                    �	      �	       Q�	      
       �Q�                �	      	
       u��0$0&�                �	      	
       u��0$0&�                  �	      
       Q
      	
       �Q�                �	      	
       T                     �	      
       R
      	
       Q	
      	
      	 p q "#�@�                  
      	
       q ?&�	
      	
       P                                    �      �       T�      �       R�      &	       �T�&	      2	       R2	      H	       �T�H	      w	       Rw	      �	       �T��	      �	       R�	      �	       �T��	      �	       R                                  �      �       Q�      &	       �Q�&	      D	       QD	      H	       �Q�H	      �	       Q�	      �	       �Q��	      �	       Q�	      �	       �Q��	      �	       Q                    @      G       QG      P       �Q�                    0      7       Q7      ?       �Q�                    �             Q      -       �Q�                    �      �       Q�      �       �Q�                            �      �       U�      �       V�      �       �U��      �       U�      1       V1      :       �U�                          �      �       T�      �       \�      �       �T��      3       \3      :       �T�                            �      �       Q�      �       S�      �       �Q��      �       Q�      
       S
      :       �Q�                            �      �       R�      �       ]�      �       �R��      �       R�      5       ]5      :       �R�                   �      �       T�             T                          @      �       U�      �       V�             �U�      '       U'      k       V                        @      _       T_      �       \�             �T�      k       \                          @      �       Q�      �       S�             �Q�      $       Q$      k       S                          @      �       R�             �R�      8       R8      O       ��O      k       �R�                        _      �       T�      �       T      8       TO      k       T                      �4      �4       U�4      �4       S�4      �4       �U�                      �4      �4       T�4      �4       V�4      �4       �T�                      �4      �4       Q�4      �4       ]�4      �4       �Q�                       5      5       U5      #5       S#5      05       �U�                       5      5       T5      /5       \/5      05       �T�                       5      5       Q5      -5       V-5      05       �Q�                      05      @5       U@5      S5       SS5      i5       �U�                      05      @5       T@5      T5       VT5      i5       �T�                  A5      X5       P                     A5      S5       v 3$s�"�S5      T5       v 3$�U#�"�T5      Z5       �T3$�U#�"�                   X5      Z5       PZ5      Z5      
 p q "#���                  X5      Z5       p ?&�Z5      Z5       Q                      p5      x5       Ux5      �5       S�5      �5       �U�                  y5      �5       P                     y5      �5      
 s��
����5      �5       q 
����5      �5       �U#��
���                   �5      �5       P�5      �5      
 p q "#���                  �5      �5       p ?&��5      �5       Q                      04      �4       U�4      �4       S�4      �4       �U�                    �4      �4      	 p  $ &��4      �4      	 x  $ &�                    �4      �4      	 p  $ &��4      �4       T                    0      :       T:      N       �T�                        :      A       TA      I      	 p t "#�@�I      M       PM      N       t ?&t "#�@�                     :      A       t ?&�A      I       PI      N       t ?&�                    ��       �       U �      ��       �U�                    ��      ��       V��      ��       V                         ��      �       0��      =�       P=�      ��       S��      ��       P��      ��       S                 �      ��       V��      ��       V                   �      =�       P=�      ��       S��      ��       S                          �#      X%       UX%      �'       S�'      �'       �U��'      )       S)      )       �U�                          �#      �$       T�$      �'       V�'      �'       �T��'      )       V)      )       �T�                      �#      >'       Q>'      �'       s�'      )       �Q�                       Q%      m%       0�m%      �%       1��%      �%       2��%      �'       3�                         �#      �$       t���$      �'       v���'      �'       �T#���'      )       v��)      )       �T#��                    �'      �'       P%(      )       P                    �#      �#       U�#      �#       �U�                      �#      �#       T�#      �#       S�#      �#       �T�                    �#      �#       Q�#      �#       �Q�                      �#      �#       R�#      �#       \�#      �#       �R�                      �#      �#       X�#      �#       V�#      �#       �X�                     �#      �#       R�#      �#       \�#      �#       �R�                        P      n       Un      �       S�      �       T�      �       �U�                    ]      �       V�      �       U                        p!      �!       U�!      b#       ^b#      g#       �U�g#      y#       U                 p!      r!       u�                        !      [#       S[#      f#       Tg#      q#       Sq#      y#       u�	                  �!      "       0�                  �!      �!       V                    �       �        U�       n!       �U�                      �       �        T�       h!       Sh!      n!       �T�                  �       m!       ]                            �       �        0��       �        \�       �        |��       	!       \"!      +!       0�+!      9!       V9!      B!       v�B!      S!       V                          �Y      �Z       U�Z       [       ��~ [      [       �U�[      [       U[      �g       ��~                            �Y      oZ       ToZ      �Z       S�Z      [       �T�[      [       T[      �[       S�[      �g       �T�                          �Y      �Z       Q�Z       [       ��} [      [       �Q�[      [       Q[      �g       ��}                          �Y      �Z       R�Z       [       ��~ [      [       �R�[      [       R[      �g       ��~                          �Y      �Z       X�Z       [       ��~ [      [       �X�[      [       X[      �g       ��~                            �Y      �Z       ][      �]       ]Ua      sa       ]�a      �a       ]�c      td       ]�d      e       ]                                      Z      �Z       \[      �]       \�]      Ua       ��~Ua      sa       \�a      �a       \�a      {b       ��~+c      �c       ��~�c      td       \td      �d       ��~�d      e       \e      �g       ��~                         Z      �Z       0��Z      �Z       P�Z      �Z       ��}�Z      [       0�[      <[       P<[      �g       ��}                       Z      �Z       0��Z      �Z       ��}�Z      Q[       0�Q[      u[       Pu[      �g       ��}                       Z      �Z       0��Z      �Z       w �Z      �[       0��[      �[       P�[      �g       w                         �[      �[       s p ��[      �\       s ��~�Ua      sa       s ��~��a      �a       s ��~�                          �\      ?]      
 ��~�
����a      �a      
 ��~�
����c      �c      
 ��~�
����d      �d      
 ��~�
����d      e      
 ��~�
���                                          �\      �\       P�\      ?]       S�]      0`       ��~�a      �a       PEb      {b       ��+c      �c       ��~�c      �c       S�c      �c       ��~�c      �c       ��~s �td      �d       ��~�d      e       S�e      �f       ��~�f      �f       ��~g      Bg       ��~                            �[      �[       v s ��[      ?]       VUa      sa       V�a      �a       V�c      �c       V�d      e       V                          �^      �^       P�^      Ua       ���a      Eb       ���c      td       Ve      �g       ��                                Z      +Z       0��]      �]       0��]      Ua       ��~�a      Ub       ��~\b      {b       P+c      �c       ��~td      �d       ��~e      �g       ��~                                                      ?]      k]       0�Q_      f_       0�f_      q_       t w ���_      �_       0��_      `       R�`      �`       0��`      Ua       T+c      8c       0�8c      `c       \`c      kc       0�kc      �c       \�d      �d       0��d      �d       \�e      �e       P�e      f       p�f      �f       P�f      �f       T�f      �f       P�f      g       T                
           Z      \       0�\      )\       P)\      Ua       ��~Ua      sa       Psa      �a       ��~�a      �a       0��a      �g       ��~                            Z      6\       0�6\      Z\       PZ\      Ua       ��~Ua      sa       0��a      �a       0��a      �a       P�a      �g       ��~                          Z      i\       0�i\      p\       Pp\      Ua       ��~Ua      sa       0��a      �a       0��a      �g       ��~                   Z      [       _[      �g       _                                Z      �Z       0�[      ?]       0�Ua      sa       0��a      �a       0�c      +c       ��~�c      �c       0��c      �c       P�c      td       ��~�d      e       0�                                           Z      �Z       0�[      �]       0��]      Ua       ��~Ua      sa       0��a      �a       0��a      �a       ��~�a      �a       0��a      {b       ��~+c      �c       ��~�c      td       0�td      �d       ��~�d      e       0�e      :g       ��~:g      Bg       PBg      �g       ��~                      �^      �^       ��~�^      ;`       S�e      �e       S:g      Bg       P                        Z      �^       0��^      _       ��~Ua      �a       0�b      e       0�g      Bg       0�                                     Z      3_       0�3_      6_       P6_      d_       Ud_      Ua       ��~Ua      �a       0��a       b       ��~ b      e       0�e      �e       ��~�e      �e       U�e      g       ��~g      Bg       0�Bg      �g       ��~                                       Z       ]       0� ]      "]       P"]      Ua       ��~Ua      �a       0��a      c       ��~c      +c       0�+c      �c       ��~�c      ,d       0�,d      7d       P7d      �d       ��~�d      �d       0��d      �d       P�d      �d       ��~�d      e       0�e      �g       ��~                                   Z      0]       0�0]      N]       PN]      Ua       ��~Ua      �a       0��a      c       ��~c      +c       0�+c      �c       ��~�c      id       0�id      td       Ptd      �d       ��~�d      e       0�e      �g       ��~                        ^      ^       p 
���^      v^       ~ 
���+c      �c       ~ 
���td      �d       ~ 
���                            ^       ^       p 
��� ^      �^       s 
���+c      �c       s 
���td      �d       s 
����d      �d       p 
����d      �d       s 
���                        y^      �^       P�^      �_       \�e      �e       \g      Bg       \                      �e      f       Zf      �f       Z�f      �f       Z                      �e      f       T f      �f       T�f      �f       T                            �e      �e       R�e      �e      9 p 3$��~"� $ &| p 3$��~"� $ &| ?&"#��@& $ &�Nf      �f       R�f      �f       R�f      �f      9 p 3$��~"� $ &| p 3$��~"� $ &| ?&"#��@& $ &��f      �f       R                          �e      �e       Q�e      �e      $ p 3$��~"� $ &| s "#��@& $ &�df      �f       Q�f      �f      $ p 3$��~"� $ &| s "#��@& $ &��f      �f       Q                   f      ,f       p 3$s ",f      7f      	 p 3$��~"                   0f      7f       Q7f      7f      
 q r "#���                  0f      7f       q ?&�7f      7f       R                  Nf      Qf       p 3$s "Qf      Uf      	 p 3$��~"                  Nf      Uf       QUf      Uf      
 q s "#���                  Nf      Uf       q ?&�Uf      Uf       S                    �_      �_       Q�_      �_       P                �_      �_      	 t 3$��~"                   �_      �_       Q�_      �_      
 q u "#���                  �_      �_       q ?&��_      �_       U                  �_      �_      	 t 3$��~"�_      �_       r ����3$��~"                   �_      �_       Q�_      �_      
 q t "#���                  �_      �_       q ?&��_      �_       T                              �`      �`       R�`      �`       x p "a      Ua       R�f      �f       R�f      g       Rg      	g       x p "g      g       R                        �`      �`       [a      Ua       [�f      �f       [�f      g       [                        �`      �`       Sa      Ua       S�f      �f       S�f      g       S                            �`      �`       Q�`      �`       p 1$v "#p 1$z "#�a      Oa       QOa      Sa       p 1$v "#p 1$z "#��f      �f       Q�f      g       Q                         `      Ua       ��}e      �e       ��}�f      �f       ��}�f      g       ��}Bg      �g       ��}                         `      Ua       w e      �e       w �f      �f       w �f      g       w Bg      �g       w                          `      Ua       ��}e      �e       ��}�f      �f       ��}�f      g       ��}Bg      �g       ��}                         `      Ua       Ve      �e       V�f      �f       V�f      g       VBg      �g       V                           O`      �`       \e      -e       \-e      je       ��je      pe       \pe      �e       [Bg      �g       ��                                  O`      �`       Ze      /e       Z/e      je       \je      �e       ZBg      Pg       \Pg      ug       Zug      �g       ~��g      �g       Z�g      �g       ~�                   e      �e       ]Bg      �g       ]                                   e      /e       ]/e      >e       QBe      he       Qhe      je       u�je      pe       ]pe      �e       SBg      ug       Qug      �g       S�g      �g       Q�g      �g       S                                    ;`      p`       \p`      x`       Qx`      �`       ]�`      �`       q��`      �`       Q�`      �`       \e      e       \e      e       ]e      Be       ^Be      Fe       ~�Oe      pe       ^                        ;`      �`       ��~�`      �`       Pe      �e       ��~Bg      �g       ��~                    /e      Be       Vae      je       V                    /e      Be       ��}ae      je       ��}                    /e      Be       ^ae      je       ^                      /e      >e       Qae      he       Qhe      je       u�                      /e      >e       T>e      Be       ~�ae      je       T                    /e      >e       Uae      je       U                 pe      �e       V                 pe      �e       ��}                 pe      �e       S                 pe      �e       Z                 pe      �e       \                        �e      �e       [�e      �e       [�e      �e       S�e      �e       S                  ^g      vg       V                  ^g      vg       ��}                  ^g      vg       ]                    ^g      ug       Qug      vg       S                    ^g      ug       Zug      vg       ~�                    ^g      ug       Uug      vg       s�                  g      �g       V                  g      �g       ��}                  g      �g       ]                  g      �g       S                    g      �g       T�g      �g       }�                      g      �g       \�g      �g       U�g      �g       ��                                        �=      >       U>      A>       SA>      �>       �U��>      �@       S�@      �B       ���B      �B       �U��B      �B       ���B      C       SC      `D       ��`D      E       SE      #E       ��#E      9E       S                                  �=      >       T>      >       Q>      >       _>      �>       �T��>      �?       _�?      �?       U�?      C       _C      	C       U	C      9E       _                                  �=      A>       V�>      �@       V�@      �B       ���B      �B       ���B      C       VC      `D       ��`D      E       VE      #E       ��#E      9E       V                                       �=      >       U>      A>       SA>      �>       �U��>      �@       S�@      �B       ���B      �B       �U��B      �B       ���B      C       SC      `D       ��`D      E       SE      #E       ��#E      9E       S                  �>      �>       ��~} �                      �?      O@      
 ��~�
����B      C      
 ��~�
���`D      �D      
 ��~�
���                                    �?      #@       R(@      8@       R8@      }A       ��~bB      �B       ��~�B      C       RC      �C       ��~�C      �C       ��~`D      �D       R�D      �D       ��~�D      �D       ��~z �E      9E       ��~                            JA      NA       QNA      bB       ���B      �B       ���C      �C       ���C      `D       ��yD      �D       ]                                  q@      �@       0��@      lB       ��~pB      �B       P�B      �B       0��B      �B       R�B      �B       Q�B      �B       ��~C      `D       ��~E      #E       ��~                                            �A      �A       0��A      �A       q��A      B       QB      B       q�C      5C       0�5C      _C       S_C      pC       0�pC      �C       S�C      �C       r��C      �C       0��C      �C       VD      #D       0�#D      RD       URD      `D       T                          �=      A>       0�Y>      #?       0�#?      2?       P2?      S?       ^S?      r?       Pr?      9E       ^                	          �=      A>       0�f>      }?       0�}?      �?       P�?      �?       ��~�?      �?       P�?      9E       ��~                
      �=      A>       0�s>      �?       0��?      �?       P�?      9E       ��~                   �=      �>       \�>      9E       \                               �=      A>       0��>      q@       0��B      �B       ��~�B      C       0�`D      �D       0��D      �D       P�D      E       ��~#E      9E       0�                                       �=      A>       0��>      �@       0��@      ,B       ��~,B      5B       0�5B      �B       ��~�B      �B       ��~�B      C       0�C      �C       ��~�C      �C       P�C      `D       ��~`D      E       0�E      #E       ��~#E      9E       0�                        pA      }A       ��~}A      NB       S�B      �B       S�C      �C       P�C      `D       S                                 �=      �A       0��A      �A       P�A      BB       VBB      �B       0��B      �B       P�B      �B       V�B      �C       0��C      D       PD      `D       V`D      9E       0�                                �=      A>       0�~>      W@       0�W@      [@       P[@      �B       ]�B      C       0�C      `D       ]`D      �D       0��D      �D       P�D      9E       ]                          �@      �@       p 
����@      -A      
 ��~�
���C      �C      
 ��~�
����C      �C      
 ��~�
���E      #E      
 ��~�
���                              �@      �@       p 
����@      A       s 
���C      0C       s 
���0C      �C      
 ���
����C      �C       p 
����C      �C       s 
���E      E       s 
���                        A      #A       P#A      }A       R�C      �C       R�C      �C       ��~                 #D      LD       t 3$} "                #D      8D       t 3$v "                   1D      8D       Q8D      8D      
 q r "#���                  1D      8D       q ?&�8D      8D       R                 �A      B       q 1$s "�
���                 �A      B       t 3$} "                �A       B       q 3$v "                   �A       B       R B       B      
 r y "#���                  �A       B       r ?&� B       B       Y                       !       u                            ��      �       U�      b�       Sb�      j�       �U�j�      ��       S��      ��       �U���      ��       S                              ��      �       T�      c�       Vc�      j�       �T�j�      ��       V��      ��       �T���      ��       T��      ��       V                               ��      �       6��      ��       P&�      5�       PN�      ]�       Pj�      {�       P|�      ��       P��      ��       6���      ��       P                   �      %�       s�	j�      {�       s�	                     �      
�       q
�      ]�       ]j�      r�       q                   �      %�       s�@%�j�      {�       s�@%�                  ��      ]�       \                 ��      %�       s�                  �      ]�       ^                            ��      �       U�      \�       ]\�      ]�       �U�]�      ��       ]��      ��       U��      à       ]                          ��      �       T�      +�       S+�      /�       s�/�      ]�       �T�]�      à       S                            ��      �       Q�      Z�       \Z�      ]�       �Q�]�      ��       \��      ��       Q��      à       \                       ��      �       0���      ��       0���      ��       P��      à       P                    �      R�       V]�      ��       V��      à       V                             �      �       0��      �       p��      �       P�      $�       p�$�      ;�       R]�      o�       0�                     �      ��       S��      R�       R]�      ��       R                            P�      ��       U��      ՝       ]՝      ڝ       �U�ڝ      D�       ]D�      N�       UN�      ��       ]                      P�      ��       T��      Н       Sڝ      ��       S                                  P�      ��       Q��      f�       _f�      ڝ       �Q�ڝ      +�       _+�      D�       �Q�D�      N�       QN�      ��       _��      ��       �Q���      ��       _                   ��      ��       }�	c�      ~�       }�	                        ��      ��       Vڝ      D�       Vc�      ��       V��      ��       V                           ��      ��       0���      ��       q���      Μ       QΜ      ݜ       q��      �       T�      �       T��      ��       0�                   |�      ӝ       \ڝ      ��       \                                  ��      ��      
 q 3$p "#���      Μ       q 3$p "�Μ      ۜ      
 q 3$p "#��      �       P�      3�       p q "�3�      7�       p q "#�7�      <�       p q "��      �       P�      !�       px�!�      +�       P                                 ��      ��       _��      ��      
 q 3$ "#���      Μ       q 3$ "�Μ      ݜ      
 q 3$ "#��      �       X�      3�       x q "�3�      7�       x q "#�7�      <�       x q "���      ��       _                         |�      f�       0�f�      j�       Pj�      ǝ       _ǝ      +�       0�+�      D�       _D�      ��       0�                      |�      ��       0�ɜ      Μ       1�.�      3�       1��      �       1�D�      ��       0�                   �      �       q @%��      �       }�@%�                   �      �       q @%����4$v"@��      �       }�@%����4$v"@�                  �      +�       Q                            Р      ��       U��      l�       ]l�      m�       �U�m�      ��       ]��      ��       U��      ӡ       ]                          Р      ��       T��      ;�       S;�      ?�       s�?�      m�       �T�m�      ӡ       S                            Р      ��       Q��      j�       \j�      m�       �Q�m�      ��       \��      ��       Q��      ӡ       \                       Р      ��       0���      ��       0���      ��       Pɡ      ӡ       P                    �      b�       Vm�      ��       V��      ӡ       V                            �      �       0��      #�       p�#�      +�       P+�      4�       p�4�      K�       Rm�      �       0�                     ��      �       S�      b�       Rm�      ��       R                                P�      ��       U��      Ȗ       \Ȗ      ϖ       �U�ϖ      �       \�      ��       U��      ̛       \̛      ,�       ^,�      I�       \                                           P�      ��       T��      L�       S��      ��       S��      #�       SA�      +�       S+�      k�       Vk�      ��       S��      ��       S��      ��       V��      �       S�      K�       VK�      қ       Sқ      '�       \'�      I�       S                                      P�      ��       Q��      	�       ^	�      ��       �Q���      ��       ^��      �       �Q��      ��       Q��      �       ^�      ��       �Q���      m�       ^m�      ��       �Q���      ɛ       ^ɛ      I�       ��~                        P�      ��       R��      �       �R��      ��       R��      I�       �R�                    ��      	�       |�	��      ��       |�	��      �       |�	                       ��      M�       _��      ��       _A�      m�       _��      I�       _                               ��      ȓ       0�&�      M�       0�M�      h�       Ph�      j�       p�j�      r�       P�      �       Q�      #�       P��      ��       0�                                      ��      �       0��      `�       ��~��      ��       0���      �       ��~�      �       0��      #�       ��~A�      y�       0�y�      ��       ��~��      m�       0�m�      ��       ��~��      ��       ��~��      I�       0�                        ��      ��       P��      �       ��~�      ��       P��      I�       ��~                        }�      ��       ��~ϖ      �       ��~#�      A�       ��~m�      ��       ��~                          }�      �       Y�      �       1���      ޗ       Yޗ      �       1�m�      ��       Y                        Ɣ      ܔ       r x "�ܔ      ��       r x "#���      �       r x "�ȗ      ޗ       P                        ��      Ɣ       PƔ      ܔ       p x "�ܔ      ��       p x "#���      �       p x "�                       ��      ��       x @%���      ��       X��      ��       x���      �       |�@%�                       `�      ��       \ϖ      �       \��      ��       \��      ��       \                        `�      ��       ^ϖ      �       ^��      ��       ^��      ��       ^                        `�      ��       R��      ��       }��      ��       R��      ��       }                      `�      ��       S��      ��       s���      ��       S                         `�      m�       Pm�      ��       ��~ϖ      �       ��~��      ��       ��~��      ��       P                    T�      X�       pX�      ^�       P �      �       ��~#                      \�      ��       R�      �       R��      ��       R                	                       `�      o�       0�o�      s�       p�s�      {�       P{�      ��       p���      ��       R      �       0�\�      `�       0�`�      ��       P��      ��       p���      ��       P�      �       0���      ��       P��      ��       0�                          �      �       1��      6�       R6�      9�       T9�      >�       Rϖ      ږ       R                        `�      `�       S`�      ו       Vו      \�       ��~ϖ       �       ��~ �      �       V��      ��       V                           �       ]�      \�       _ϖ       �       _                 f�      k�       r�u �                 f�      k�       Q                   u�      |�       Q|�      |�      
 q t "#���                  u�      |�       q ?&�|�      |�       T                   ��      ��       u r����      ��       T                 ��      ��       Q                        ��      m�       \��      ݚ       \�      ̛       \̛      ,�       ^,�      5�       \                       ��      �       P�      m�       ��~��      ݚ       ��~�      5�       ��~                 ��      ژ       ��~                 ��      �       |�	                        -�      _�       S��      ��       S�      K�       Sқ      $�       V                      ؛      �       0��      �       S�      �       s��      �       S                  ��      �       ��~                 ��      ��      
 ��~��~"�                 �      �      
 ��~��"�                 �      ��      
 ��~��"�                                        �      b�       Ub�      ��       ]��      �       �U��      �       U�      �       ]�      ,�       �U�,�      č       ]č      �       �U��      a�       ]a�      A�       ��~A�             ]      O�       �U�                        �      b�       Tb�      �       ��}�      �       T�      O�       ��}                          >�      ��       V�      �       V,�      Ս       V�             VӒ      �       V                        C�      b�       Pb�      �       ��~�      �       P�      O�       ��~                             N�      b�       0�b�      ��       ^�      ��       0���      ��       P��      �       ^,�      ��       ^A�      g�       ^                             ҋ      �       0��      5�       0���      ��       0��      a�       0�a�      �       _�      �       ��      A�       _A�      g�       0���             0�                  l�      {�       0���      ��       0�                               N�      ��       0�߈      �       P�      �       R�      �       0�,�      w�       0�w�      ~�       P~�      ΋       U΋      O�       ��~                    .�      {�       Uҋ      �       T                          �      $�       P$�      a�       Ua�      �       \)�      A�       \��             P                              l�      щ       Qщ      ؉       p ؉      ؉       q{�؉      �       Q�      ,�       Q�      Y�       [A�      M�       [M�      g�        ��~"��~"��~"��~"�                            _�      �       P�      ,�       P��      ��       ^��      }�       Si�      ��       Q��      ��       qP���      ��       Q                              l�      ��       P��      ��       px���      ��       P��      ��       ]��      ��       }x���      �       ])�      A�       ]                                Z�      l�       Pl�      ��       ���
��4$u"��      a�       Ra�      �       ^�      �       ~p��      A�       ^��      ��       P��             R                           N�      b�       0�b�      ��       ��~�      Ɋ       0�Ɋ      ��       s 
�� $| 
��2$# $)�,�      �       ��~�      �       ��~                          w�      ��       R��      ��       ��~,�      �       ��~�             ��~Ӓ      ��       ��~                          _�      ��       \��      �       \,�      ��       \��      }�       ��~A�      g�       \                          �      �       p ��      �       r ��      ,�       r ���      ��       _��      a�       \a�      e�       |~�e�      s�       \A�      g�       _                   w�      ��        ��      O�        �                      |�      ��       P��      ��       ��~�      O�       ��~                      ��      ��       P��      ��       ��~�      O�       ��~                      ��      ��       P��      ��       ��~�      O�       ��~                          ��      ��       P��      ��       ��~�      ,�       ��~,�      9�       P9�      O�       ��~                       ��      ��       | 5�����,�      ��       | 5�������      }�       ��~�5�����A�      g�       | 5�����                     N�      ��        0)��      �        0)�,�      ��        0)�                    u�      y�       Py�             ^                    Ս      ��       V      Ӓ       V                        ��      �       p ���      &�       p ��A�      M�       p ��      Ӓ       p ��                     Ս      &�       	��&�      ��       ^      Ӓ       	��                  .�      G�       0�l�      ��       0�                   ��      �       ]�      O�       ]                    ��      �       V�      O�       V                  ��      }�       ^                   ��      �       _�      O�       _                     ��      ��       r���      �       s��      ��       s�                      }�      �       ^�      �       ^�      O�       Q                        ��      ��       P��      �       ��~�      �       ��~�      O�       R                  �      {�       ��~                    ��      �       P�      �       ��~                  ��      ��       ��~                  ��      ׏       ��~                  *�      2�       P                            �      �       U�      I       ^I      L       �U�L      v       ^v      y       �U�y             U                      �      �       T�      y       �T�y             T                            �      �       Q�      K       _K      L       �Q�L      x       _x      y       �Q�y             Q                            �      �       R�      E       \E      L       �R�L      r       \r      y       �R�y             R                            �      �       X�      G       ]G      L       �X�L      t       ]t      y       �X�y             X                           �      �       0��      3       S3      8       s�8      B       SL      o       Sy             0�                           �      �       @<$��      �       P�      7       P8      n       Pn      y       0�y             @<$�                          ��      ��       U��      �       \�      )�       �U�)�      :�       \:�      V�       U                   ��      ��       u�	:�      A�       u�	                            ѣ      q�       ^q�      v�       ~p�v�      ��       ^)�      :�       ^A�      Q�       ^Q�      V�       y(                      أ      ��       S)�      :�       SA�      V�       S                           ��      ��       0���      v�       ��v�      {�       P{�      ��       ��)�      :�       ��:�      V�       0�                         ��      ��       0���      ��       ��)�      5�       ��5�      :�       P:�      V�       0�                       ��      ��       0���      ��       ��)�      :�       ��:�      V�       0�                        ��      ,�       ]G�      O�       PO�      ��       ])�      :�       ]                      ��      �       PP�      {�       P)�      :�       P                     ��      �       \�      (�       u�~�(�      )�       �U�                    `      h       Uh      y       �U�                    `      m       Tm      y       �T�                   `      h       uh      q       �U#                                                                          `      �       U�      �       u�{��      4       U4      E       u�z�E      O       UO      `       u�{�`      �       U�      �       u�z��      �       U�      	       u�{�	      A       UA      R       u�z�R      �       U�      �       u�z��      �       U�      �       p�|��             u�|�             U             p�{�      (       u�{�(      7       U7      <       p�y�<      H       u�z�H      �       U�      �       u�z��      �       U�      �       p�{��      �       u�{��             U                                             �      �       P�      �       P�      �       P�      �       P             P1      2       PQ      R       Pq      r       P�      �       P�      �       P�      �       P�      �       P�      �       P�      �       P             P                    ��      ��       U��      ��       �U�                    ��      ��       T��      ��       �T�                    ��      ��       Q��      ��       �Q�                    ��      ƴ       Uƴ      Ǵ       �U�                    ��      ƴ       Tƴ      Ǵ       �T�                    ��      ƴ       Qƴ      Ǵ       �Q�                          ��      ѳ       Uѳ      `�       S`�      f�       �U�f�      q�       Uq�      ��       S                                  ��      ѳ       Tѳ      ��       V��      
�       T
�      A�       VA�      f�       �T�f�      q�       Tq�      ��       V��      ��       T��      ��       V                                  ��      ѳ       Qѳ      ��       ]��      �       Q�      [�       ][�      f�       �Q�f�      q�       Qq�      ��       ]��      ��       Q��      ��       ]                                ��      ѳ       Rѳ      ��       �R���      �       R�      f�       �R�f�      q�       Rq�      ��       �R���      ��       R��      ��       �R�                           ��      [�       0�f�      }�       0�}�      �       P�      ��       0���      ��       P��      ��       0�                   �      ��       VG�      [�       V                   �      ��       0�D�      T�       Q                  U�      [�       P                    �      ��       T(�      T�       T                 1�      G�       V                     �      ��       t��      ��       Q��      ��       t                           �      d�       Ud�      ��       ^��      ��       �U���      ��       U��      ��       ^                         �      c�       Tc�      ��       �T���      ��       T��      ��       �T�                    ;�      q�       S��      )�       S                            M�      q�       ]��      D�       ]D�      H�       UH�      Q�       ]��      ��       U��      ȱ       ]                   M�      z�       V��      ��       V                    ^�      ��       ]ֱ      ��       ]                 �      �       T                    Ȱ      ٰ       Pٰ      �       _                          ��      ��       P��      ��       w ��      �       w �      K�       w R�      ϲ       w                       �       �       P �      ��       _��      ݱ       _                          )�      H�       PH�      ��       S��      ��       P��      �       S�      �       S                 �      ��       ]                  �      �       } ��      |�       } �                       �      �       t s "��      ��       T��      �       w s "��      �       w s "�                  �      �       ^�      |�       ^                  �      �       _�      |�       _                        ��      ��       P��      �       ���      K�       ��R�      ϲ       ��                 K�      R�       8�                      �      K�       SR�      ��       S��      ��       R                   n�      ��       s 
��4&3#���      ��       r 
��4&3#�                   n�      ��       s ?
��#���      ��       r ?
��#�                   n�      ��       1s ?
��#$1���      ��       1r ?
��#$1�                    ϲ      ޲       Xi�      |�       X                      ��      �       Y�      1�       ��1�      q�       Y                      ��      �       Q�      1�       ��1�      N�       Q                    :�      U�       PU�      l�       t 2$u "                 Q�      q�       Q                  �      8�       P                    PF      uF       UuF      ZK       �U�                        PF      }F       T}F      �F       \�F      �F       �T��F      ZK       \                        PF      }F       Q}F      �F       ]�F      �F       �Q��F      ZK       ]                    kF      �F       S�F      ZK       S                    yF      �F       V�F      ZK       V                    �F      �F       P�F      �F       P                      �F      �F       P�F      �G       ��H      4H       ��                                  CG      NG       0�NG      jG       QjG      �G       ���G      �G       Q4H      6I       ��;I      UI       PUI      lI       ��lI      K       w K      ZK       w                                           �H      �H       0��H      �H       w )I      1I       R<J      LJ       QLJ      vJ       ��vJ      �J       Q�J      �J       R�J      �J       Q�J      �J       ���J      K       QK      K       RK      %K       Q%K      IK       ��IK      ZK       Q                  �J      �J       x�                  �I      �I       ��                     yF      �F       ^�F      �G       ^H      4H       ^                  �I      ZK       ^                       yF      �F       0��F      �F       _�F      :G       0�:G      NG       PNG      ZK       _                  �H      �H       ^                  �H      �H       ��                  �H      �H       ��                  �H      I       P                  �J      �J       P                  &K      IK       P                    �;      �;       U�;      �=       �U�                      �;      �;       S�;      F<       SP<      �=       S                      �;      �;       ]�;      K<       ]P<      �=       ]                     �;      �;       \�;      I<       \P<      �=       \                    �<      �<       P�<      i=       _                      #<      '<       P'<      9<       VP<      �<       V                              0<      9<       P9<      P<       ��P<      U<       PU<      q<       Qq<      �<       ���<      �<       ^�<      �=       ��                      �<      �<       0��<      <=       w <=      A=       w �#�Y=      �=       w                           �<      �<       0��<      =       V\=      m=       Pm=      q=       _q=      w=       v�                          �2      �2       U�2      v3       ^v3      �3       �U��3      4       ^4      (4       �U�                    �2      �2       T�2      (4       �T�                          �2      �2       Q�2      v3       Vv3      �3       �Q��3      4       V4      (4       �Q�                          �2      �2       0��2      �2       P�2      v3       ]�3      4       ]4      4       T4      4       0�                      3      63       p ���3      �3       p ���3      �3       p ��                    3      v3       \�3      4       \                                3      3       0�3      O3       SO3      i3       Ri3      v3       S�3      �3       S�3      �3       R�3      �3       S�3      4       P                                    +3      63       0�63      G3       _G3      O3       �O3      v3       _�3      �3       0��3      �3       _�3      �3       ��3      �3       _�3      �3       0��3      4       _                    �2      �2       P�2      (4       ��                        �0      1       U1      �1       \�1      �1       �U��1      �2       \                            �0      1       T1      d1       Vd1      �1       �T��1      
2       V
2      �2       �T��2      �2       V                            �0      1       Q1      f1       Sf1      �1       �Q��1      
2       S
2      �2       �Q��2      �2       S                         �0      S1       0�S1      W1       PW1      �1       w 
2      �2       w �2      �2       0�                          1      "1       p ��"1      �1       ^�1      �2       ^�2      �2       p ���2      �2       ^                          1      �1       p ���1      �1        ���1      �1       P�1      �1       ��#2      #2        ��#2      72       ��                                   b1      k1       0�k1      �1       S�1      �1       s��1      �1       s��1      �1       S�1      �1       s��1      �1       S
2      2       ]2      #2       S#2      >2       s�>2      \2       s�\2      o2       So2      v2       s�v2      �2       S                        �1      �1       0��1      �1       	��2      #2       0�C2      \2       0�\2      �2       	��                     b1      k1       0�k1      �1       V
2      �2       V                      �0      k1       ]�1      
2       ]�2      �2       ]                         �      ?�       U?�      �       ]�      $�       �U�$�      ,�       ]                         �      %�       T%�      �       V�      $�       �T�$�      ,�       V                             �      ��       Q��      �       ��{�      $�       �Q�$�      ��       ��{��      ��       �Q���      ,�       ��{                                           �      ��       R��      �       S�      $�       �R�$�      '�       S'�      �       �R��      )�       S)�      ��       �R���      ��       S��      [�       �R�[�      ��       S��      �       �R��      �       S�      ,�       �R�                                    M�      �       0�$�      0�       P0�      B�       ^}�      ��       P��      ��       ^��      ��       P��      �       ^)�      ��       ^��      �       ^��      �       ^�      ,�       ^                       v�      ��       _$�      B�       _v�      #�       _�      �       _                 �      ��       v                    ��      ��       ��|���      ��       X��      ��       ��|�                    ��      ��       ��|���      ��       R��      ��       ��|�                  ��      ��       ��{��      ��       S                 ��      ��       v                
�      R�       ��{                
�      R�       ��|�0$0&�                   �      R�       PR�      R�      
 p r "#���                  �      R�       p ?&�R�      R�       R                l�      s�       ��{                l�      s�      
 ��|�
���                  l�      s�       ^s�      s�      
 p ~ "#���                  l�      s�       ~ ?&�s�      s�       P                ��      ��       ��|�0$0&�                   ��      ��       P��      ��      
 p r "#���                  ��      ��       p ?&���      ��       R                ��      ��      	 | �
���                  ��      ��       _��      ��      
 p  "#���                  ��      ��        ?&���      ��       P                       v�      �       ]$�      B�       ]v�      ��       ]�      �       ]                     v�      ��       R��      M�       S$�      $�       S�      �       S                   v�      M�       V$�      $�       V�      �       V                	 v�      ��       U                
   v�      ��       u���      ��       P                 v�      ��       X                      ��      ��       P��      M�       ^$�      $�       P�      �       ^                 ��      ��       \                ��      ��       ��{                ��      ��       ��}                   ��      ��       Q��      ��      
 q r "#���                  ��      ��       q ?&���      ��       R                ��      ��       _                ��      ��       ��~                   ��      ��       P��      ��      
 p q "#���                  ��      ��       p ?&���      ��       Q                          p�      ��       ��{)�      i�       ��{|�      ��       ��{��      ��       ��{�      [�       ��{��      �       ��{                          p�      ��       \)�      i�       \|�      ��       \��      ��       \�      [�       \��      �       \                            u�      i�       S)�      i�       S|�      ��       S��      ��       S�      [�       S��      �       S                      ��      ��       P��      ��       ��{)�      i�       P                            ��      ��       @<$���      ��       ��{)�      i�       ��{|�      ��       ��{��      ��       ��{�      [�       ��{��      �       ��{                          ��      ��       _)�      i�       _|�      ��       _��      ��       _�      [�       _��      �       _                     ��      ��       R��      ��       ��{)�      i�       R                   ��      ��       s�
p "���      ��       P                   <�      ��       ��{��      ��       ��{��      ��       q�                   <�      ��       y 
�����      ��       y 
���                   <�      ��       S��      ��       S                     <�      i�       0�i�      ��       P��      ��       0�                    <�      ��       0���      ��       0���      ��       s�
p "�                  <�      ��       s�
��      ��       s�
                   <�      ��       s�
#���      �       s�
#�                         �      C�       XQ�      l�       X��      ��       X+�      M�       XM�      [�       ��{                             ��      0�       R0�      C�       ��|V�      o�       Ro�      ��       � ��      ��       R��      ��       RV�      [�       R                    ��      �       P��      ��       P                    �      +�       Q+�      C�       s�#h                    D�      V�       P|�      ��       P                d�      ~�       ��{                 d�      s�       X                   s�      ~�       X~�      ~�      
 p x "#���                  s�      ~�       x ?&�~�      ~�       P                ��      ��       ��{                ��      ��       S��      ��       R                ��      ��       P                 ��      ��       \                        ��      ��       U��      :�       S:�      D�       �U�D�      ��       S                                  ��      
�       T
�      ;�       V;�      D�       �T�D�      M�       TM�      m�       Vm�      ��       T��      ?�       V?�      Z�       TZ�      ��       V                                  ��      
�       Q
�      A�       ^A�      D�       �Q�D�      M�       QM�      m�       ^m�      ��       Q��      M�       ^M�      |�       Q|�      ��       ^                              ��      ��       R��      
�       [D�      X�       [X�      m�       w m�      s�       �R�s�      ?�       [?�      ��       �R�                                  ��      
�       X
�      D�       �X�D�      M�       XM�      m�       �X�m�      ��       X��      ?�       �X�?�      |�       X|�      ��       ����      ��       �X�                   ��      =�       \D�      ��       \                   ��      C�       _D�      ��       _                    ��      "�       PO�      `�       P                                  ��      
�       { � $0.�
�      D�       �R� $0.�D�      M�       { � $0.�M�      m�       �R� $0.�m�      ��       { � $0.���      ?�       �R� $0.�?�      |�       { � $0.�|�      ��       ���� $0.���      ��       �R� $0.�                          ��      ��       P��      
�       w D�      M�       w m�      ��       w ?�      	�       w                             ��      ��       R��      ?�       ���      B�       RB�      ��       ����      ��       R��      ��       ��                               }�      ��       1���      F�       ��?�      5�       1�5�      B�       0�B�      ��       ����      ��       1���      ��       ����      ��       1�                     ��      ��       0��      5�       1���      ��       0�                     ��      ��       0�0�      5�       ����      ��       0�                           }�      .�       0�9�      `�       1�?�      _�       0�_�      e�       1�q�      ��       1���      ��       0���      ��       1���      ��       0�                          ?�      M�       { � $0.�_�      |�       { � $0.�|�      ��       ���� $0.���      ~�       �R� $0.���      �       �R� $0.���      ��       �R� $0.�                 ?�      M�       T                          ?�      ?�       0�?�      M�       P_�      l�       0���      ��       P��      ��       0���      �       P��      ��       0�                         _�      |�       { � $0.�|�      ��       ���� $0.���      e�       �R� $0.���      ��       �R� $0.���      ��       �R� $0.�                    i�      p�       Pp�      	�       ��                    p�      |�       P|�      	�       ��                        ��      	�       �� �      3�       Q3�      e�       ����      ��       ��                 p�      	�       ��#��                     ��      ~�       v����      �       v����      ��       v��                   �      ��       0��      ��       0�                   �      ��       ���      ��       ��                     �      3�       Q3�      ��       ���      ��       ��                   �      ��       ���      ��       ��                 Q�      ��       t�#                   ��      l�       �R� $0.���      �       �R� $0.�                     ��      ��       Q��      l�       V��      �       V                    ��      ��       X��      ��       ����      ��       ��                    ��      ��       R��      ��       ����      ��       ��                     ��      ��       P��      ��       0���      �       P                     _�      ��       r����      l�       ��#����      ��       r����      �       ��#��                     _�      ��       r����      l�       ��#����      ��       r����      �       ��#��                 ��      ��       P                 ��      ��       Q                 ��      ��       1�                 ��      ��       R                 ��      ��       2�                 ��      ��       R                 ��      ��       3�                 ��      ��       R                 ��      l�       V                 ��      l�       R                       �      -�       0�-�      I�       1�I�      e�       2�e�      l�       3�                 ��      ��       0�                 ��      ��       1�                 ��      ��       U                   ��      ��       u����      �       ��#��                    ��      ��       0���      ��       0�                  [�      m�       ]                                                �g      =h       U=h      \h       S\h      nh       �U�nh      �l       S�l      m       �U�m      z       Sz      ||       ^||      K}       SK}      y}       ^y}      �}       S�}      �}       ^�}      A~       SA~      �~       ^�~      �       S�      �       ^�      h�       S                                                    �g      h       Th      \h       \\h      nh       �T�nh      �h       T�h      �l       \�l      m       �T�m      �m       \�m      �o       �T��o      p       \p      �q       �T��q      ~r       \~r      	t       �T�	t      �y       \�y      y}       �T�y}      �}       \�}      �}       �T��}      A~       \A~      h�       �T�                                                                �g      Hh       QHh      \h       ]\h      nh       �Q�nh      �h       Q�h      �l       ]�l      m       �Q�m      �m       ]�m      �o       ��}�1��o      �o       �Q��o      :p       ]:p      �q       �Q��q      ~r       ]~r      	t       �Q�	t      �y       ]�y      ||       ��}�1�||      K}       �Q�K}      y}       ��}�1�y}      �}       ]�}      �}       ��}�1��}      �}       �Q��}      A~       ]A~      1�       ��}�1�1�      R�       ]R�      h�       ��}�1�                        �g      Lh       RLh      nh       �R�nh      �h       R�h      h�       �R�                                    0h      9h       T9h      \h       w h      �l       w m      �m       w �o      �p       w �q      �r       w 	t      �y       w y}      �}       w �}      A~       w 1�      R�       w                    0h      9h       u#X#h      �h       ��|                               �h      �h       P�h      �l       ��|m      Um       0�Um      �m       ��|�o      Or       ��|~r      0t       ��|||      K}       ��|�}      �}       ��|                                           �g      \h       Vnh      �l       Vm      �m       V�m      �o       ��|�o      z       Vz      ||       ��|||      K}       VK}      y}       ��|y}      �}       V�}      �}       ��|�}      A~       VA~      1�       ��|1�      R�       VR�      h�       ��|                                        �g      �g       P�g      =h       u=h      Lh       sLh      \h       ��|nh      �h       s�h      �l       ��|m      �m       ��|�o      z       ��|||      K}       ��|y}      �}       ��|�}      A~       ��|1�      R�       ��|                               �g      \h       0�nh      �l       0�m      �o       0��o      p       1�p      �q       0��q      ~r       1�~r      	t       0�	t      �t       1��t      �}       0��}      $~       1�$~      h�       0�                         �g      \h       0�nh      �h       0��h      m       ��|m      m       0�m      Um       1�Um      h�       ��|                        r      mr       ^	t      �y       ^y}      �}       ^�}      A~       ^                          �m      �o       ��|�0$0&�\t      ft      	 t 0$0&�ft      ||       ��|�0$0&�K}      �}       ��|�0$0&�$~      h�       ��|�0$0&�                          �m      �o       ��}�0$0&�at      ft      	 p 0$0&�ft      ||       ��}�0$0&�K}      �}       ��}�0$0&�$~      h�       ��}�0$0&�                          �m      �o       ��|�t      �t       P�t      ||       ��|K}      �}       ��|$~      h�       ��|                  �}      ~       P                    	t      t       Qt      0t       P                                  �u      �u       0��u      �u       P�u      v       p�v      v       Pv      Pv       RPv      Sv       p�Sv      |v       ��|�#�|v      �v       T�v      w       P<w      >w       0�>w      \w       Q\w      dw       q�dw      yw       Q                      �t      �t       P�t      1v       ��|y}      �}       ��|                        �u      �u       U�u      �u       uP��u      v       U<w      qw       P                     �t      u       0�u      8u       P8u      #v       ��|                     �t      Du       0�Du      lu       Plu      -x       _                     �t      zu       0�zu      �u       P�u      w       ��|                             �t      �u       0��u      �u       P�u      w       Yw      -x       ��|=x      Ax       YAx      �x       ��|�x      �x       0�y}      �}       0�                   �y      z       0�1�      R�       0�                      �z      �z       Z�z      �{       ��|�      �       ��|                               �y      z       0�gz      vz       Rvz      vz       0�vz      �z       |� } "�{      �{       RK}      e}       Re}      y}       ��|V~      �~       R�      �       R1�      R�       0�                                         �m      �o       ��|�y      z       ��|�0$0&�z      vz       ��|vz      �{       ��|�0$0&��{      �{       T�{      ||       ��|K}      y}       ��|�}      �}       ��|A~      �       ��|�      �       ��|�0$0&��      1�       ��|1�      R�       ��|�0$0&�R�      h�       ��|                    �y      �y       ^1�      R�       ^                    �y      z       \1�      R�       \                            �m      �o       ��|�y      �y       P�y      ||       ��|K}      y}       ��|�}      �}       ��|A~      h�       ��|                            �m      �o       ��|�y      �y       P�y      ||       ��|K}      y}       ��|�}      �}       ��|A~      h�       ��|                                      �z      �z       V��8�z      �z       V�S��0�z      �z       V�S�_�u��� �z      �{       V�S�_���|�� �{      �{       �S�_���|�� �{      �{      
 �S�_��(�{      �{       �S��0K}      \}       �S�_���|�� \}      y}      
 �S�_��(�      �       V�S�_���|�� �      �       �S�_���|��                  �z      �z       ��|                     �z      �{       ��|K}      a}       ��|�      �       ��|                     �{      �{       ZK}      e}       Ze}      y}       ��|                           z      \z       ��|�0$0&��{      ||       ��|�0$0&�K}      y}       ��|�0$0&��}      �}       ��|�0$0&�A~      Q~       ��|�0$0&��      �       ��|�0$0&�                     �{      �{       RK}      e}       Re}      y}       ��|                           z      \z       ^�{      ||       ^K}      y}       ^�}      �}       ^A~      Q~       ^�      �       ^                          z      Pz       V�{      �{       VK}      y}       VA~      Q~       V�      �       V                   �{      �{       p �0$0.�K}      e}       p �0$0.�                                 Lz      \z       _�{      �{      	   $ &��{      |       _.|      k|       _k|      o|       `�o|      ||       _�}      �}       _�      �      	   $ &��      �       _                                 Pz      \z       S�{      �{      	 s  $ &��{      +|       SD|      s|       Ss|      w|       s`�w|      ||       S�}      �}       S�      �      	 s  $ &��      �       S                       z      z       v�0$0&�z      1z       P1z      Pz       v�0$0&�A~      Q~       P                   z      Ez       _A~      Q~       _                    z      z       Sz      Iz       SA~      Q~       S                  ?z      Pz       P                  Bz      Pz       Q                  |      ||       t                 |      ||       t                |      |       t                 |      |       _                   |      |       _|      |      
 p  "#���                  |      |        ?&�|      |       P                .|      5|       t                  .|      5|       S5|      5|      
 p s "#���                  .|      5|       s ?&�5|      5|       P                 N|      ||       ~                  N|      ||       ~ #�                  �      �       P                  �      �       P                  �      �       _�      �      
 q  "#���                  �      �        ?&��      �       Q                �      �       S�      �      
 p s "#���                �      �       P                       �m      �o       ��}�0$0&��~      �       ��}�0$0&��      1�       ��}�0$0&�R�      h�       ��}�0$0&�                       �m      �o       ��|�0$0&��~      �       ��|�0$0&��      1�       ��|�0$0&�R�      h�       ��|�0$0&�                       �m      �o       S�~      �       S�      1�       SR�      h�       S                    �~      u       |��      1�       |�                     Qo      So       0�So      ao       Qdo      �o       Q                      �m      �o       \u      �       \R�      h�       \                    n      �o       ]R�      h�       ]                     n      jn       s #�R�      c�       q�c�      h�       s #�                 �n      Qo       ��}�0$0&�                 �n      Qo       ��|�0$0&�                 �n      Qo       r�                 �n      Qo       s��                   r      +r       ]+r      Dr       P                                               �m      �o       s��r      Sr       RSr      br       ��|br      mr       s��	t      4t       R4t      z       s��z      ||       ~��K}      y}       ~��y}      �}       s���}      �}       ~���}      �}       ��|�}      A~       s��A~      �~       ~���~      �       s���      �       ~���      h�       s��                       r      <r       Q?r      Sr       Q	t      4t       Q4t      Gt       ��|                �x      �x       w                 �x      �x       s�                    �x      �x       P�x      �x      
 p r "#���                  �x      �x       p ?&��x      �x       R                �x      �x       w                 �x      �x       s�                   �x      �x       P�x      �x      
 p r "#���                  �x      �x       p ?&��x      �x       R                �x      y       w                 �x      y       s�                   y      y       Py      y      
 p r "#���                  y      y       p ?&�y      y       R                )y      ;y       ��|                )y      ;y       s�                   4y      ;y       P;y      ;y      
 p u "#���                  4y      ;y       p ?&�;y      ;y       U                Py      by       w                 Py      by       s�                   [y      by       Tby      by      
 p t "#���                  [y      by       t ?&�by      by       P                wy      �y       ��|                wy      �y       s�                   �y      �y       R�y      �y      
 p r "#���                  �y      �y       r ?&��y      �y       P                 �h      �i       \                 �h      �i       S                  �h      �i       _                  ~i      �i       P                   �h      i       Zi      �i       ��|                    3i      Ii       PIi      �i       ��|                    3i      ;i       ��}�;i      Ii       XIi      Ji       ��}�                    3i      Ci       ��}�Ci      Ii       RIi      Ji       ��}�                3i      Ji       \                3i      Ji       _                �k      �k       w                 �k      �k       s�                    �k      �k       P�k      �k      
 p r "#���                  �k      �k       p ?&��k      �k       R                il      pl       ��|                il      pl       s�                  il      pl       Rpl      pl      
 p r "#���                  il      pl       r ?&�pl      pl       P                l      "l       w                 l      "l       s�                   l      "l       P"l      "l      
 p r "#���                  l      "l       p ?&�"l      "l       R                7l      Il       w                 7l      Il       s�                   Bl      Il       PIl      Il      
 p r "#���                  Bl      Il       p ?&�Il      Il       R                �l      �l       w                 �l      �l       s�                  �l      �l       Q�l      �l      
 p q "#���                  �l      �l       q ?&��l      �l       P                �l      �l       ��|                �l      �l       s�                   �l      �l       P�l      �l      
 p q "#���                  �l      �l       p ?&��l      �l       Q                       p      �q       S~r      	t       S||      K}       S�}      �}       S                        p      �q       \~r      s       \�s      �s       \�|      K}       \                       7p      �q       |� �~r      s       |� ��s      �s       |� ��|      K}       |� �                   7p      �p       ^~r      s       ^                        7p      �q       _~r      	t       _||      K}       _�}      �}       _                                7p      �p       0��p      �p       Y�q      �q       Y�q      �q       0�~r      �r       0��r      �r       P�r      s       w �|      .}       Y.}      K}       w                                �p      7q       |� 7q      >q       P>q      ~q       pp�~q      �q       P�s      �s       |� �s      �s       P�s      �s       pp��s      	t       P                              �p      q       t x "�q      �q       X�q      �q       t } "#@�s      �s       t } "#@��s      	t       X||      �|       t } "#@��}      �}       t } "#@�                       �p      q       0�q      1q       R1q      7q       p�s      �s       R                       �p      q       0�q      4q       Q4q      7q       p�s      �s       Q                   �p      q       0�q      �q       1��s      	t       1�                  7q      >q       p >q      Iq       pp                   Bq      Iq       ZIq      Iq      
 z { "#���                  Bq      Iq       z ?&�Iq      Iq       [                   dq      kq       Zkq      kq      
 z { "#���                  dq      kq       z ?&�kq      kq       [                        �s      �s       Y�s      �s       R�s      �s       rp��s      	t       R                  �s      �s       r �s      �s       rp                   �s      �s       Q�s      �s      
 q { "#���                  �s      �s       q ?&��s      �s       [                   �s      �s       Q�s      �s      
 q { "#���                  �s      �s       q ?&��s      �s       [                 �|      "}       0�                 �|      "}       |� �                 �|      "}       s��                    �      �       0��             0�      "       q�                  �      �       0��             0�      "       q�                      �      �       0��      %       0�%      F       x q �U      W       x q �                     �      �       u #��             Q      \       u #�                             ,      C,       UC,      .       S.      .       �U�.      $0       S$0      .0       �U�.0      i0       S                     ,      ,       T,      i0       �T�                  ,      ,       u                       %,      .       V.      %0       V.0      i0       V                           %,      C,       u��C,      .       s��.      .       �U#��.      $0       s��$0      .0       �U#��.0      i0       s��                      0,      .       \.      '0       \.0      i0       \                  �/      �/       P                   .      6.       s6.      �.       P                  /.      �/       �^��                 D.      `.       \                 D.      `.       _                 D.      `.       3�                 D.      `.       U                 �.      �/       U                 �.      �.       0�                 �.      �.       3�                 �.      �.       U                 �.      �/       u��                        `K      �K       U�K      �L       w �L      �L       ���L      �N       w                           �K      1L       XCL      _L       P_L      �L       X�L      xN       XxN      �N       ���N      �N       X                                        {K      �K       ^�K      �K       U�K      �K       u��K      �K       T�K      rL       ^rL      �L       ~��L      �L       U�L      	M       T	M      &M       t�&M      1M       ~~�1M      BM       ^BM      TM       UTM      hM       u�hM      �M       T�M      �M       U�M      �M       u��M      �M       T�M      �M       t��M      N       t�N      N       t�N      N       ~~�N      -N       ^-N      -N       U-N      <N       u�<N      RN       TRN      �N       ^                    �K      �L       V�L      �N       V                    �K      �L       S�L      kN       S                    �K      �L       \�L      �N       \                      �K      1L       PjL      �L       P�L      xN       P                       �K      �K       0��K      L       ]L      +L       �+L      �L       ]�L      �N       ]                               �K      L       @<$�L      1L       R�L      1M       @<$�1M      BM       R�M      �M       @<$��M      -N       RDN      _N       @<$�_N      xN       R                             �K      L       0�L      1L       Y�L      BM       0��M      N       0�N      -N       YDN      _N       0�_N      xN       Y                               �K      L       @<$�L      L       RL      1L       T�L      =M       @<$�=M      BM       T�M      (N       @<$�(N      -N       TDN      _N       @<$�_N      xN       T                               �K      L       0�L      1L       U�L      BM       0��M      N       0�N      -N       UDN      _N       0�_N      tN       UtN      xN       p                            �K      �K       R�L      �L       2��L      �L       R�L      �L       	�0t 0$0)( 	�#��M      �M       R�M      �M       	�0t 0$0)( 	�#�                 pN      xN       s0                                  �5      �5       U�5      �8       V�8      �8       U�8      �8       V�8      �8       �U��8      9       U9      9       V9      (9       U(9      p:       V                             Z7      x7       P�7      �8       0�19      ?9       P^9      h9       Ph9      �9       0��9      �9       F��9      p:       0�                                                        �5      �5       R6      46       r�R6      �6       S�6      Y7       ZY7      �7       ���7      �7       Y�7      8       T8      48       U48      98       TN8      y8       Ry8      �8       [�8      �8       R�8      �8       T�8      �8       R�8      �8       R�8      9       r�9      09       R09      ?9       w h9      n9       Tn9      }9       U}9      �9       Y�9      �9       [�9      �9       Z�9      �9       R�9      �9       T�9      +:       R+:      F:       TF:      `:       R`:      p:       Y                    �5      �8       ]�8      p:       ]                    �5      �8       \�8      p:       \                    �5      �8       ^�8      p:       ^                     �7      �8       |� �h9      �9       |� ��9      p:       |� �                    7      �8       Sh9      p:       S                       �6      �6       0��6      �6       ��6      �6       _?9      J9       0�                                      �7      �7       X�7      98       PE8      g8       |� g8      �8       Qh9      �9       P�9      �9       Q�9      �9       Q�9      	:       Y	:      :       y�:      F:       Y`:      h:       Xh:      p:       P                      �7      g8       [h9      �9       [`:      p:       [                             �7      �7       Q�7      8       x 8      8       p8      (8       t (8      48       Qh9      �9       Qh:      p:       Q                    �9      �9       u h:      p:       u                           >8      g8       Ug8      �8       P�9      �9       P�9      �9       P�9      `:       U                      E8      �8       Z�9      �9       Z�9      `:       Z                       E8      g8       0�g8      �8       X�8      �8       X�9      �9       X                    �9      �9       Q:      A:       Q                           �5      46       |� 46      A6       XA6      �6       Q�8      �8       X�8      9       X?9      B9       Q                          �5      6       ~ 0$0&1$|� "�6      
6      
 p 1$|� "�
6      �6       U�8      �8       X�8      9       X?9      Y9       U                       +6      n6       Pn6      �6       T�6      �6       T9      9       P                               g8      8       0�8      �8       R�8      �8       0��8      �8       r ��8$r��!0$0&��8      �8       { 8$r��!0$0&��8      �8       { 8$t��!0$0&��8      �8       t~��8$t��!0$0&��9      �9       R�9      �9       r ��9      �9      	 {���                          g8      |8       T|8      �8       q �8      �8       T�8      �8       q �9      �9       q                            �9      �9       0��9      �9       R�9      �9       r �:      +:       0�+:      /:       r ��8$r��!0$0&�/:      3:       x 8$r��!0$0&�3:      7:       x 8$t��!0$0&�7:      >:       t~��8$t��!0$0&�                    �9      :       P:      F:       P                    �       �        Q�              q�      "       q�"      9       q�9      P       q�P      p       Rp      q       u�                 �       q       u�                    �0      �0       U�0      �0       �U�                   �0      �0       u0�0      �0       U                          p0      �0       U�0      �0       V�0      �0       �U��0      �0       V�0      �0       �U�                    p0      u0       Tu0      �0       �T�                    p0      �0       Q�0      �0       �Q�                          p0      �0       R�0      �0       \�0      �0       �R��0      �0       \�0      �0       �R�                    �0      �0       P�0      �0       P                    �0      �0       S�0      �0       S                        @       �        U�       �        S�       �        �U��       �        U                      @       �        T�       �        �T��       �        T                   @       `        u �       �        u                    @       �        0��       �        w �       �        0�                   @       �        0��       �        �`�       �        0�                  �       �        P                              0�      ��       U��      ��       T��      ��       �U���      ��       U��      ��       T��      ��       �U���      &       U                                      0�      7�       T7�      ��       P��      ��       �T���      ��       P��      ��       �T���             P             �T�             P             �T�      %       P%      &       �T�                          0�      ��       Q��      ��       �Q���      ��       Q��      ��       �Q���      &       Q                              0�      z�       Rz�      ��       R��      ��       r 9!���      ��       x 9!���      ��       X��      ��       R��      ��       R��      &       R                             0�      ��       U��      ��       T��      ��       �U���      ��       U��      ��       T��      ��       �U���      &       U                                      3�      7�       T7�      ��       P��      ��       �T���      ��       P��      ��       �T���             P             �T�             P             �T�      %       P%      &       �T�                                    7�      i�       Ti�      ��       u��      ��       t��      ��       T��      ��       u��      ��       t��      ��       u��      ��       T��      ��       u��      &       T                                        U      6       S6      7       �U�7      R       SR      S       �U�                               $       T$      7       �T�7      D       TD      S       �T�                          $       U7      D       U                             6       S6      7       �U�7      R       SR      S       �U�                           %       0�%      7       P7      S       0�                       $       u�                                    s�      $       Q$      6       s�6      7       �U#�                              $        U$       .        �U�.       3        U                              $        T$       .        �T�.       3        T                              $        Q$       .        �Q�.       3        Q                                $        R$       -        S-       .        �R�.       3        R                             $        U$       .        �U�.       3        U                             $        P.       2        P2       3        u�                    �N      �N       U�N      �N       X                  �N      �N       T                    �N      �N       U�N      �N       X                   �N      �N       u� �N      �N       x�                  �N      �N       Q                      P      e       Te      k       Pk      x       T                        P      `       Q`      e       �Q�e      p       Qp      x       �Q�                  w      x       P                          �N      �N       U�N      �N       �U��N      O       UO      'O       �U�'O      LO       U                              �N      �N       T�N      �N       Q�N      �N       �T��N      O       TO      'O       �T�'O      JO       TJO      LO       �T�                      �N      �N       Q�N      �N       �Q��N      LO       Q                          �N      �N       R�N      �N       �R��N      O       RO      'O       �R�'O      LO       R                      �N      �N       X�N      �N       �X��N      LO       X                    'O      JO       TJO      LO       �T�                  'O      LO       X                  'O      LO       R                  'O      LO       Q                  'O      LO       U                            PO      �O       U�O      �O       \�O      �O       �U��O      
P       U
P      BP       \BP      lP       U                          PO      �O       T�O      �O       �T��O      
P       S
P      BP       �T�BP      lP       S                          PO      �O       Q�O      �O       �Q��O      
P       Q
P      BP       �Q�BP      lP       Q                    PO      oO       RoO      lP       �R�                          PO      �O       X�O      �O       �X��O      
P       X
P      BP       �X�BP      lP       X                    �O      �O       0��O      �O       1�                           _O      �O       U�O      �O       \�O      �O       �U��O      
P       U
P      BP       \BP      lP       U                    �O      BP       �R�WP      lP       �R�                      �O      
P       X
P      BP       �X�WP      lP       X                      �O      
P       Q
P      BP       �Q�WP      lP       Q                      �O      
P       S
P      BP       �T�WP      lP       S                      �O      
P       U
P      BP       \WP      lP       U                    �O      ;P       0�;P      BP       1�                
P      2P       ^                
P      2P       ]                    
P      (P       S(P      1P       Q1P      2P       s�                
P      2P       \                      pP      �P       U�P      �P       �U��P      �P       U                      pP      �P       T�P      �P       �T��P      �P       T                      pP      �P       Q�P      �P       �Q��P      �P       Q                  �P      �P       U                  �P      �P       R                  �P      �P       X                  �P      �P       Q                  �P      �P       T                 �P      =Q       t $ &#04$u "#�                        R      !R       Q!R      *R       �Q�*R      8R       Q8R      GR       �Q�                           R      R      	 p t "	��R      !R       q t "# 	��!R      %R       �Qt "# 	��%R      )R       P)R      *R       �Qt "# 	��FR      GR       P                  *R      GR       U                    *R      8R       Q8R      GR       �Q�                  *R      GR       T                         *R      3R      
 p t 	��3R      8R       q t # 	��8R      ?R       �Qt # 	��?R      FR       PFR      GR       �Qt # 	��                        PR      ^R       Q^R      kR       �Q�kR      sR       QsR      �R       �Q�                      bR      fR       p �fR      jR       PjR      kR       �Qt "	�# �                  kR      �R       U                    kR      sR       QsR      �R       �Q�                  kR      �R       T                    �R      �R       P�R      �R       r q �                          �R      �R       Q�R      �R       �Q��R      �R       Q�R      �R       P�R      �R       �Q�                         �R      �R      	 t q "	���R      �R      
 t �Q"	���R      �R       P�R      �R      
 t �Q"	���R      �R       P                  �R      �R       U                      �R      �R       Q�R      �R       P�R      �R       �Q�                  �R      �R       T                         �R      �R      
 q t 	���R      �R      
 p t 	���R      �R       �Qt 	���R      �R       P�R      �R       �Qt 	��                        �R      �R       Q�R      �R       �Q��R      �R       Q�R      S       �Q�                           �R      �R      	 p t "	���R      �R       q t "#?	���R      �R       �Qt "#?	���R      �R       P�R      �R       �Qt "#?	��S      S       P                  �R      S       U                    �R      �R       Q�R      S       �Q�                  �R      S       T                         �R      �R      
 p t 	���R      �R       q t #?	���R      �R       �Qt #?	���R      S       PS      S       �Qt #?	��                        S      !S       Q!S      *S       �Q�*S      8S       Q8S      GS       �Q�                           S      S      	 p t "	��S      !S       q t "#	��!S      %S       �Qt "#	��%S      )S       P)S      *S       �Qt "#	��FS      GS       P                  *S      GS       U                    *S      8S       Q8S      GS       �Q�                  *S      GS       T                         *S      3S      
 p t 	��3S      8S       q t #	��8S      ?S       �Qt #	��?S      FS       PFS      GS       �Qt #	��                         sS      vS      	 r t "p �vS      yS       u�q "t "x p �yS      S       r x "�S      �S       P�S      �S       r x "�                  �S      �S       Q                  �S      �S       T                  �S      �S       U                           �S      �S      
 r t p ��S      �S       u�q "t x p ��S      �S       u�q "t x u���S      �S       u�t u�q "u���S      �S       P�S      �S      	 r u��                        �S      �S       Q�S      �S       �Q��S      �S       Q�S      �S       �Q�                           �S      �S       p t "r r ��S      �S       u�q "t "x r r ��S      �S       u�t "x �Q"r r ��S      �S       p x "��S      �S       P�S      �S       u�t "x �Q"r r x "�                    �S      �S       Q�S      �S       �Q�                  �S      �S       T                  �S      �S       U                           �S      �S       p t r r ��S      �S       u�q "t x r r ��S      �S       u�t x �Q"r r ��S      �S       u�t u��Q"r r ��S      �S       P�S      �S       u�t u��Q"r r u��                  `T      �T       T                  `T      �T       U                      �T      U       TU      U       �T�U      =U       T                    �T      U       QU      =U       Q                    �T      U       XU      =U       X                    �T      U       RU      =U       R                    �T      U       TU      =U       T                    �T      U       UU      =U       U                        @U      �U       U�U      �V       S�V      �V       �U��V      �W       S                     @U      @U       0�@U      �U       T�V      �V       TW      FW       T                              �U      >V       _vV      �V       P�V      W       _�W      �W       P�W      �W       _�W      �W       P�W      �W       _                        ,V      >V       P>V      �V       ^W      W       ^�W      �W       ^                 @U      BU       u�                    �U      �U       T�U      �U       u�v "�                 �U      �U       P                     �V      �V       p 3�#<3$s "#�V      W       s��3�#<3$s "#�W      �W       s��3�#<3$s "#                   �V      W       _�W      �W       _                   �V      W       S�W      �W       S                      �V      �V        q "��V      W       ^�W      �W        q ��W      �W       _                      <W      JW       QJW      �W       s�v "��W      �W       s�v "�                     <W      pW       PpW      �W       s��
��4$s� "��W      �W       P                       wW      {W       p t "#��@& $ &���{W      �W      ( p t "#��@& $ &��q u "#��@& $ &���W      �W      ; s�v "�z  $ &x p "#��@& $ &��q u "#��@& $ &���W      �W      Y s�v "�z  $ &x p "#��@& $ &��s�v "#�y  $ &s�� $ &u "#��@& $ &���W      �W      z s�v "�z  $ &x p "#��@& $ &��s�v "#�y  $ &s�� $ &s�v "#�y  $ &s�� $ &?&"#��@& $ &��                SW      wW       X                    SW      VW       t z �VW      iW       TiW      wW       s�v "�z �                   iW      wW       TwW      wW      
 p t "#���                  iW      wW       t ?&�wW      wW       P                  wW      {W       Q{W      {W      
 q u "#���                  wW      {W       q ?&�{W      {W       U                �W      �W       s�                 �W      �W       P                   �W      �W       P�W      �W      
 p q "#���                  �W      �W       p ?&��W      �W       Q                         X      X       UX      +X       P+X      EX       [EX      �Y       �U�                     X      EX       TEX      �Y       ��                                 X      X       QX      EX       ]EX      ~X       X�X      �X       Z�X      �X       ��4Y      vY       X�Y      �Y       X�Y      �Y       Z                               X      EX       REX      ~X       Z�X      �X       X�X      �X       ��4Y      vY       Z�Y      �Y       Z�Y      �Y       P                       X      %X       X%X      RY       ^UY      �Y       ^                           X      QX       YQX      �X       Y�X      �X       ��4Y      vY       Y�Y      �Y       Y                    �X      �X       T�X      �X       ��fY      vY       ��                  X      EX       0�                          �X      Y       PY      4Y       PvY      �Y       P�Y      �Y       q �Y      �Y       P                         �X      �X       \�X      KY       SUY      �Y       S�Y      �Y       x  $ &4$~ "�Y      �Y       z  $ &4$~ "                           �X      �X       S�X      �X       Q�X      NY       \UY      �Y       \�Y      �Y       z  $ &4$~ "�Y      �Y       p  $ &4$~ "                         �X      �X       Q�X      �X       w UY      vY       x  $ &4$y "�Y      �Y       x  $ &4$y "�Y      �Y       z  $ &4$y "                     UY      vY       z  $ &4$y "�Y      �Y       z  $ &4$y "�Y      �Y       p  $ &4$y "                         �X      �X       _�X      �X       ]UY      vY       x  $ &4$y "x  $ &4$~ "��Y      �Y       x  $ &4$y "x  $ &4$~ "��Y      �Y       z  $ &4$y "z  $ &4$~ "�                         �X      �X       ]�X      �X       RUY      vY       z  $ &4$y "z  $ &4$~ "��Y      �Y       z  $ &4$y "z  $ &4$~ "��Y      �Y       p  $ &4$y "p  $ &4$~ "�                    �X      �X       PfY      vY       0�                   vY      �Y       p s ��Y      �Y       P                   �Y      �Y       P�Y      �Y      
 p { "#���                  �Y      �Y       p ?&��Y      �Y       [                        p�      ��       U��      Q�       ^Q�      T�       �U�T�      ,�       ^                          p�      ��       T��      �       S�      T�       �T�T�      l�       Sl�      ,�       �T�                        p�      ̀       Q̀      M�       \M�      T�       �Q�T�      ,�       \                    p�      }�       R}�      ��       �R�                    p�      ��       X��      ��       �X�                    �      J�       ST�      ,�       S                        ��      ��       Y��      ��       P��      �       YT�      g�       Y                        ��      �       Z�      E�       ��T�      l�       Z��      ,�       ��                    ɀ      O�       ]T�      ,�       ]                        ̀      	�       Q	�      E�       _T�      ��       Q��      ,�       _                     ̀      �       _�      �       VT�      ��       _                            ׀      ݀       X݀      �       [�      I�       w I�      T�       ��T�      ��       [��      ,�       w                     ڀ      �       RT�      ��       R                        ݀      �       X�      E�       w  �T�      ��       X��      ,�       w  �                        �      �       0��      E�       Z��      �       Z�      ,�       P                          �      �       0��      E�       [��      ��       [��      ׁ       1�ׁ      �       [�      ,�       1�                        �      "�       P,�      E�       P��      ��       Pҁ      �       P                ��      ��       Z                ��      ��       ~v "y �                   ��      ��       P��      ��      
 p { "#���                  ��      ��       p ?&���      ��       [                  g�      ��       Y                              P�      a�       Ua�      ��       S��      ��       �U���      �       S�      �       �U��      ,�       S,�      2�       �U�                                P�      x�       Tx�      ��       \��      ��       �T���      ��       T��      �       \�      �       �T��      1�       \1�      2�       �T�                             P�      a�       Ua�      ��       S��      ��       �U���      �       S�      �       �U��      ,�       S,�      2�       �U�                             P�      {�       0�{�      ��       P��      ��       V��      ��       0���      ą       V�      $�       P$�      +�       V                 g�      x�       U                 g�      x�       u�                    ��      �       \�      �       �T�                    ��      �       S�      �       �U�                      ą      ̅       P̅      �       V�      �       P                  ޅ      �       Q                        @�      f�       Tf�      j�       �T�j�      z�       Tz�      �       ��                          @�      z�       Qz�      �       ]�      ��       �Q���      ��       ]��      �       �Q�                        @�      ]�       R]�      ��       ^��      ��       �R���      �       ^                   @�      z�       Uz�      �       ��                    U�      ��       V��      �       V                                       j�      z�       0�z�      ��       _��      ��       ���      ކ       _ކ      �       ��      �       ��0�      ��       ]��      ��       _��      Շ       ]Շ      ��       }���      �       ]�      �       S�      �       0�                          0�      e�       1�e�      {�       T{�      �       X�      ��       T��      ʇ       T                       j�      φ       Sφ      ކ       sP�ކ      �       S��      ��       S                        0�      ��       \��      ه       \ه      ��       |p���      �       \�      �       ��#8                          z�      ��       U��      ��       P��      ��        3$} "��      ˆ       U��      ��       U                          �      1�       T1�      y�       _y�      z�       �T�z�      ��       _��      ��       T                      �      �       Q�      ��       P��      ��       �Q�                      �      1�       R1�      ��       �R���      ��       R                    �      �       P�      ��       ��                        �      1�       s 1$��#"�1�      ��       ��1$��"���      ��       s 1$��#"���      ��       ��1$��#"�                           �      1�       0�1�      (�       \(�      <�       |�<�      p�       \p�      z�       ���#�z�      ��       \��      ��       0�                       Z�      l�       0�l�      �       ^z�      ��       ^��      ��       0�                       �      1�       0�1�      O�       ��z�      ��       ����      ��       0�                 <�      D�       p q "#��@& $ &�                 �      z�       ����"1$��"�0$0&@$�                           1�      l�       @<$�l�      ��       P��      �       P�      �       Pz�      ��       P��      ��       @<$�                        K�      O�       t 2$p"O�      V�       t 2$p "V�      l�       t 2$��#"��      ��       t 2$��#"                    Z�      h�       Sz�      ��       S                �      <�       ����"1$��"�0$0&@$�                   :�      <�       P<�      <�      
 p q "#���                  :�      <�       p ?&�<�      <�       Q                      �      ��       U��      �       S�      �       �U�                      �      ��       T��      �       V�      �       �T�                    �      ��       Q��      �       �Q�                  ��      �       P                  ��      �       �Q�                  ��      �       V                  ��      �       S                            д      ڴ       Uڴ      �       \�      ��       �U���      0�       \0�      1�       U1�      2�       �U�                            д      �       T�      �       V�      ��       �T���      *�       V*�      1�       T1�      2�       �T�                        �      �       P�      �       S�      �       P�      #�       S                      ��      *�       V*�      1�       T1�      2�       �T�                      ��      0�       \0�      1�       U1�      2�       �U�                  �      �       U                  �      �       P                  �      .�       P                                @�      Q�       UQ�      q�       Vq�      r�       �U�r�      ��       V��      ��       �U���      ��       V��      ��       �U���      ��       V                  @�      W�       T                          @�      ��       Q��      ��       �Q���      ��       Q��      ��       U��      ��       �Q�                    @�      K�       RK�      ��       �R�                               F�      Q�       UQ�      q�       Vq�      r�       �U�r�      ��       V��      ��       �U���      ��       V��      ��       �U���      ��       V                  {�      ��       �T�                    {�      ��       P��      ��       P                            {�      �       U�      ��       Q��      ��       �Q���      ��       Q��      ��       U��      ��       �Q�                          {�      ��       V��      ��       �U���      ��       V��      ��       �U���      ��       V                          ��      ��       P��      ��       P��      ��       v� ��      ��       �U#x��      ��       P                 �      ��       Q                     ��      ��       Q��      ��       U��      ��       �Q�                      ��      ӵ       Uӵ      ܵ       u ܵ      �       �U�                    ��      ܵ       Tܵ      �       �T�                             �      z�       Uz�      ��       �U���      ��       U��      ��       �U���      ö       Uö      ʶ       �U�                             �      c�       Tc�      ��       �T���      ��       T��      ��       �T���      ��       T��      ʶ       �T�                             �      `�       Q`�      ��       �Q���      ��       Q��      ��       �Q���      ��       Q��      ʶ       �Q�                         �      ��       R��      ��       Q��      ��       �R���      ʶ       R                              Y�      z�       Yz�      }�       P}�      ��       U��      ��       Y��      ��       U��      Ŷ       YŶ      ʶ       U                          f�      t�       Qt�      ��       Y��      ��       Q��      ��       T��      Ŷ       QŶ      ʶ       Y                   t�      ��       QŶ      ʶ       Q                                D�      V�       XV�      `�       q 
��4$u�"�`�      z�       �Q
��4$u�"�z�      ��       �Q
��4$�U#�"���      ��       �Q
��4$u�"���      ��       �Q
��4$�U#�"���      ö       �Q
��4$u�"�ö      ʶ       �Q
��4$�U#�"�                                O�      ]�       P]�      c�       t 
��4$u�"�c�      z�       �T
��4$u�"�z�      ��       �T
��4$�U#�"���      ��       �T
��4$u�"���      ��       �T
��4$�U#�"���      ö       �T
��4$u�"�ö      ʶ       �T
��4$�U#�"�                            �      z�       u�z�      ��       �U#���      ��       u���      ��       �U#���      ö       u�ö      ʶ       �U#�                        z�      ��       R��      ��       R��      ��       Q��      ��       �R�ö      ʶ       R                        z�      ��       R��      ��       R��      ��       Q��      ��       �R�ö      ʶ       R                      z�      ��       Y��      ��       Tö      Ŷ       QŶ      ʶ       Y                        z�      }�       P}�      ��       U��      ��       Uö      Ŷ       YŶ      ʶ       U                    ��      ��       T��      ��       T                    ��      ��       Q��      ��       Q                    ��      ��       R��      ��       R                    ��      ��       U��      ��       U                        �&      �&       U�&      �&       V�&      �&       �U��&      �&       V                        �&      �&       T�&      �&       S�&      �&       �T��&      �&       S                        �&      �&       Q�&      �&       \�&      �&       �Q��&      �&       \                      �&      �&       P�&      �&       ]�&      �&       ]                    �&      �&       P�&      �&       Q                 �      8       U                     \      $\       U$\      �`       �U�                                 \      )\       T)\      J_       SJ_      R_       �T�R_      �_       S�_      �_       �T��_      C`       SC`      N`       �T�N`      �`       S                           \      \       Q\      �\       V�\      �_       �Q��_      �_       V�_      �`       �Q�                     \      -\       R-\      �`       �R�                     \      -\       X-\      �`       �X�                                \      )\       T)\      J_       SJ_      R_       �T�R_      �_       S�_      �_       �T��_      C`       SC`      N`       �T�N`      �`       S                                            �\      �\       P�\      ^       ]^      �^       P�^      �^       0��^      �^       P�^      �^       ]�^      ?_       0�?_      B_       VR_      �_       ]�_      `       ]`      5`       0�5`      N`       6�N`      X`       Pi`      �`       ]�`      �`       0�                           =\      D\       PD\      �^       \R_      �_       \�_      `       \5`      I`       \N`      �`       \                             T\      g\       Pg\      Q_       ^R_      �_       ^�_      �_       P�_      �_       �T#��_      M`       ^N`      �`       ^                                \      )\       t��)\      J_       s��J_      R_       �T#��R_      �_       s���_      �_       �T#���_      C`       s��C`      N`       �T#��N`      �`       s��                                \      )\       t��)\      J_       s��J_      R_       �T#��R_      �_       s���_      �_       �T#���_      C`       s��C`      N`       �T#��N`      �`       s��                   \      )\       t�)\      -\       U                            =\      D\       PD\      �^       \R_      �_       \�_      `       \5`      I`       \N`      �`       \                       �\      B_       SR_      �_       S�_      5`       SN`      �`       S                          ]      y]       Q�_      �_       Q�_      �_       q��_      �_       Q�_      �_       q��_      �_       Qi`      �`       Q                     ]      y]       R�_      �_       Ri`      �`       R                   X]      `]       1�i`      �`       0�                     �^      B_       S`      5`       S�`      �`       S                      �^      B_       \`      5`       \�`      �`       \                       �^      ,_       0�,_      <_       U`      0`       0�0`      5`       U�`      �`       0��`      �`       U�`      �`       0��`      �`       U                        �      �       U�      �        S�       �        �U��       !       U                       �      �       U�      �        S�       �        �U��       !       U                  �      �        V                     �      �       u���      �        s���       �        �U#��                         �        s���       �        �U#��                      P      y       Uy      �       S�      �       �U�                      Z      m       Pm      y       uy      }       s                  a      �       V                  ~      �       P                  �      �       P                      �G      �G       U�G      H       SH      H       �U�                      �G      �G       T�G      H       \H      H       �T�                     �G      �G       U�G      H       SH      H       �U�                    �G      �G       P�G      H       V                       H      +H       U+H      gH       SgH      hH       �U�                      H      +H       U+H      gH       SgH      hH       �U�                    H      RH       0�RH      bH       P                    3H      5H       P5H      QH       R                  =H      QH       P                                    �N      �N       U�N      �O       ^�O      �P       �U��P      Q       ^Q      9Q       �U�9Q      VW       ^VW      �W       �U��W      1Y       ^1Y      -Z       ��y-Z      VZ       �U�VZ      �[       ^                     O      �P       S�P      �P       ��y��P      �[       S                                   �N      �N       u���N      �O       ~���O      �P       �U#���P      Q       ~��Q      9Q       �U#��9Q      VW       ~��VW      �W       �U#���W      1Y       ~��1Y      -Z       ��y#��-Z      VZ       �U#��VZ      �[       ~��                                   �N      �N       u���N      �O       ~���O      �P       �U#���P      Q       ~��Q      9Q       �U#��9Q      VW       ~��VW      �W       �U#���W      1Y       ~��1Y      -Z       ��y#��-Z      VZ       �U#��VZ      �[       ~��                                  �N      �O       V�P      Q       V9Q      �T       V�W      �W       V�W      �W       V�W      bX       ��ybX      �X       V�Z      }[       ��y�[      �[       V                  �U      V       0�                 �Z      �Z       ~�                            �X      =Y       0�=Y      SY       ��ySY      �Y       \�Y      "Z       ��y�1�"Z      -Z       ��y}[      �[       0�                        �Y      �Y       0��Y      �Y       |��Y      �Y       \Z      Z       |�                    �X      VZ       0�}[      �[       0�                        �X      =Y       0�=Y      Z       ��yZ      -Z       ��y}[      �[       0�                    =Y      SY       ]^Y      -Z       ]                      �Y      �Y       V�Y      �Y       VZ      "Z       V                                   �N      �N       U�N      �O       ^�O      �P       �U��P      Q       ^Q      9Q       �U�9Q      VW       ^VW      �W       �U��W      1Y       ^1Y      -Z       ��y-Z      VZ       �U�VZ      �[       ^                   �N      �N       ��y��N      �N       S                                 O      �O       V�P      Q       V9Q      �T       V�W      �W       V�W      �W       V�W      bX       ��ybX      �X       V�Z      }[       ��y�[      �[       V                         O      O       RO      �O       _�P      Q       _9Q      `Q       _{Q      R       _bX      �X       _                       O      �O       \�P      Q       \9Q      `Q       \{Q      R       \bX      �X       \                       O      �O       S�P      Q       S9Q      `Q       S{Q      R       SbX      �X       S                   �O      yP       SQ      9Q       S                   �O      yP       SQ      9Q       S                  �O      9P       V                   MP      yP       SQ      9Q       S                   MP      yP       VQ      9Q       V                           "R      �T       V�W      �W       V�W      �W       V�W      bX       ��y�Z      }[       ��y�[      �[       V                     "R      VU       S�W      UX       S�Z      }[       S�[      �[       S                       2R      [R       \[R      aR       ��{�W      UX       \�Z      }[       \                         BR      �T       _�W      �W       _�W      UX       _�Z      [       _�[      �[       _                               [R      aR       RaR      �R       \�R      �R       |v��R      �R       P�R      'S       P'S      =S       s HS      �T       ]�W      �W       \�[      �[       ]                          _R      �R       P�R      CS       \HS      �T       \�W      �W       \�W      �W       P�[      �[       \                      cS      �S       P�S      �S       ��y�[      �[       P                  �S      �S       p  $0.�                     �W      �W       P�W      UX       ��y�Z      }[       ��y                    �!      �!       U�!      w&       ��                                �!      �!       T�!      �"       _�"      �"       �T��"      �%       _�%      �%       U�%      �%       _�%      �%       U�%      w&       _                    �!      �!       Q�!      w&       �Q�                    �!      �!       R�!      w&       �R�                               �!      �!       T�!      �"       _�"      �"       �T��"      �%       _�%      �%       U�%      �%       _�%      �%       U�%      w&       _                     �!      �"       S�"      �"       �Q�R"��"      w&       S                       �!      �!       0��!      �"       V�"       #       V #      A#       ^A#      w&       V                           �!      �!       0��!      1"       \4"      �"       \�"      <#       \A#      �#       \ %      C%       \                                 �!      1"       ^C"      �"       ^�"      #       ^#      #       ~s�#      �#       ^�#       %       \ %      C%       ^C%      w%       \|%      w&       \                      $      ?$       Q?$       %       ��C%      w&       ��                            ?$       %       ^C%      �%       ^�%      �%       T�%      �%       ^�%      �%       T�%      w&       ^                    ?$      f$       Xf$      �$       ��                              �$      �$       P�$       %      
 ��1#�C%      S%      
 ��1#�|%      �%      
 ��1#��%      �%      
 u��1#��%      �%      
 u��1#��%      w&      
 ��1#�                            �$       %       ^C%      X%       ^|%      �%       ^�%      �%       T�%      �%       ^�%      �%       T�%      w&       ^                            �$       %       _C%      X%       _|%      �%       _�%      �%       U�%      �%       _�%      �%       U�%      w&       _                    �$       %       ��C%      X%       ��|%      w&       ��                     X%      X%       P�%      �%       P�%      �%       P                                      �%      �%       ����%      �%       Q�%      �%       Q�%      �%       ����%      �%       Q�%      �%       ����%      �%       Q&      &       Q&      &       Q&      &&       ���&&      +&       Q<&      H&       ���H&      O&       Q`&      p&       ���p&      w&       Q                                  �%      �%       0��%      �%       R�%      �%       R�%      �%       0��%      �%       0��%      �%       R&      &       0�&      &       0�&      +&       0�<&      J&       0�J&      O&       R`&      r&       0�r&      w&       R                                �$      �$       Q�$       %       PC%      S%       P|%      �%       P�%      �%       P�%      �%       P&      	&       P&      w&       P                             (      N(       UN(      *,       \*,      1,       �U�1,      �,       \�,      �,       �U��,      �.       \                             (      U(       TU(      .,       ^.,      1,       �T�1,      �,       ^�,      �,       �T��,      �.       ^                            (      U(       TU(      .,       ^.,      1,       �T�1,      �,       ^�,      �,       �T��,      �.       ^                                    (      U(       t��U(      �(       ~���(      �(       P�(      ",       ��",      .,       ~��.,      1,       �T#��1,      �,       ���,      �,       ~���,      �,       �T#���,      �.       ��                                    (      U(       t��U(      �(       ~���(      �(       P�(      ",       ��",      .,       ~��.,      1,       �T#��1,      �,       ���,      �,       ~���,      �,       �T#���,      �.       ��                                      (      U(       t��U(      �(       ~���(      �(       P�(      ",       ��",      .,       ~��.,      1,       �T#��1,      �,       ���,      �,       ~���,      �,       �T#���,      �,       P�,      �.       ��                      D(      K(       PK(      U(       t U(      �.       ��~                   �,      �,       3��.      �.       P                    S(      U(       PU(      �.       ��~                                   S(      �(       ]�(      _)       __)      �)       ��)      �)       Q�)      j*       ��*      �+       _1,      P,       �],      �,       _�,      �,       ]%-      M-       _M-      Z-       ~                      S(      !+       S1,      �,       S�,      �-       S                      �(      ",       ]1,      �,       ]%-      �.       ]                        V(      e(       Pe(      (,       V1,      �,       V�,      �.       V                           S(      �(       0��(      &*       ��+*      ",       ��1,      �,       ���,      %-       0�%-      �.       ��                         S(      �(       0��(      ",       ��1,      �,       ���,      %-       0�%-      �.       ��                     _)      �)         x "��)      �)      
   ��~�"��)      �)      	 ��~�q �                     L*      j*       0�j*      n*       Pn*      �*       _�*      �*       0�                                �.      �.       U�.      l1       Vl1      u1       �U�u1      �1       V�1      �1       �U��1      �1       V�1      �1       �U��1      �1       V                                  �.      �.       T�.      t1       _t1      u1       �T�u1      {1       U{1      �1       _�1      �1       �T��1      �1       _�1      �1       �T��1      �1       _                                 �.      �.       T�.      t1       _t1      u1       �T�u1      {1       U{1      �1       _�1      �1       �T��1      �1       _�1      �1       �T��1      �1       _                                 �.      �.       t���.      t1       ��t1      u1       �T#��u1      {1       u��{1      �1       ���1      �1       �T#���1      �1       ���1      �1       �T#���1      �1       ��                        �.      r1       ^u1      �1       ^�1      �1       ^�1      �1       ^                              /       /       P /      5/       ��5/      ;/       Q;/      f1       ���1      �1       ���1      �1       Q�1      �1      	 r 3&�                      �/      �/       0��/      P1       \�1      �1       \                    �.      �.       P�.      �1       ��                         �/      Q0       S�0      �0       P�0      
1       S1      P1       S�1      �1       S                       �/      �/       0��/      �/       P�/      00       ]00      40       0��1      �1       0�                                            �      �       U�      D       VD      S       �U�S      =       V=      F       �U�F      �       V�      �       �U��      �       V�      6       ��6      N       VN      W       �U�W             V      h       ��h      z       �U�z      �       ��                                    �      �       T�      R       _R      S       �T�S      E       _E      F       ����F      �       _�      �       �T��      V       _V      W       �T�W      �       _                                   �      �       T�      R       _R      S       �T�S      E       _E      F       ����F      �       _�      �       �T��      V       _V      W       �T�W      �       _                                                       �      -       ^S      C       ^�      �       ^�      �        �      �       �T�      �       ^�      �       V�      �       ]�      6       VW             ^      �       V�      �       ]�      �       V�      &       ]&      V       Vh      z       ^z      �       V�      �       ]�      �       ^�      �       V�      �       ]                             �      D       SS      <       SF      �       S�      B       SB      r       w 6      M       SW             S                          �      D       ]S      A       ]F      �       ]�      6       ]6      R       ]W             ]                               S      =       v��=      F       �U#���      �       v���      6       ��#��W             v��      h       ��#��h      z       �U#��z      �       ��#��                   �      �       PW             
 �                              �      �       P�      ?       \?      F       ���      �       \�      6       ��r             
 �      h       ��z      �       ��                                   3      I       0�I      U       SU      h       Th      i       s�i      r       Sr      �       0��      6       w       !       w &      h       w z      �       w                        S      E       ��E      F       ���      6       ��W      �       ��                          `      t       Rt      ;       w ;      F       ���      ?       w W             R                   `      �       0�W      W       0�W             1�                        �      �       \      �       w �      �       R�      �       \                     �      �       p } ��      �       P�             V                          �2      �2       U�2      �3       S�3      �3       �U��3      4       S4      4       �U�                          �2      �2       T�2      �3       V�3      �3       �T��3      4       V4      4       �T�                          �2      �2       T�2      �3       V�3      �3       �T��3      4       V4      4       �T�                          �2      �2       u���2      �3       s���3      �3       �U#���3      4       s��4      4       �U#��                         �2      �2       u���2      �3       s���3      �3       �U#���3      4       s��4      4       �U#��                         �2      �2       U�2      �3       S�3      �3       �U��3      4       S4      4       �U�                  �2      3       p �                  �2      �2       P                                0       U0      �       S�      �       �U��      �       S�      �       �U�                                0       T0      �       ]�      �       �T��      �       ]�      �       �T�                                0       Q0      �       ^�      �       �Q��      �       ^�      �       �Q�                          0       R0      �       �R�                    4      <       P<      I       s                   .      e       V                    P      R       PR             _                      �      �       U�      �       S�      �       �U�                      �      �       T�      �       P�      �       �T�                            �      �       U�      �       V�      �       �U��      0       V0      �       �U��      �       V                        �      �       T�      �       S�      �       �T��      �       S                         �      �       0��      �       P�      
       0�
             P      �       0�                        �      �       T�      �       S�      �       �T��      �       S                    �      �       _�      �       _                   0      =       \=      p       |h�                    !      0       0�0      f       Vf      j       v��      �       0�                          �       ^�      �       ^                        !      %       P%      )       s)      �       ��|�      �       P                      P      v       Uv             S      W       �U�                          P      �       T�      �       U�      J       _J      K       �T�K      W       _                         �      �       T�      �       U�      J       _J      K       �T�K      W       _                    �             V             s�                     �             0�             ��z      $       P                      �      �       P�      �        �      5       ��z                    �      �       P�      5       ��z                    �      �       P�      W       ��z                              ��z                   �      �       0��      �       ^                     �      �       }h��      �       ]�             }h�                      �      �       U�             S      E       ��{                          �      �       T�      �       U�      -       _-      .       �T�.      E       _                          *       0�e      �       ��{�      �       ��{                          �      �       T�      �       U�      -       _-      .       �T�.      E       _                         �      �       0��      �       P�             0�      .       P.      E       0�                   �      �       s��      �       S                                     P      *        *             ��{.      >       ��{                              %       P%      *       *             ��{.      >       ��{                                 *       0�*      e       ��{e      �       0��      
       P
             ��{.      >       ��{                   *      �       ��{.      >       ��{                   �      �       0��      �       ]                   �      �       V�      �       vh�                      �&      '       U'      {'       S{'      (       �U�                          �&      '       T'      !'       U!'      (       ](      (       �T�(      (       ]                     j'      {'       0�{'      �'       V�'      �'       V                 �'      �'       3�                    c'      �'       \(      (       \                    j'      �'       ^(      (       ^                       {'      �'       _�'      �'       h��'      �'       _(      (       h�                   �'      �'       T�'      �'       R                      {'      �'       S�'      �'       S(      (       S                        �      �       U�      =       ]=      L       �U�L      �       ]                 �      �       u�                    �             SL      �       S                    �      �       ^L      �       ^                    �      �       VL      �       V                         �      	       1�p      �       P�      �       p��      �       0�L      �       1��      �       0��      �       1�                                vx�      #       v`�                      @A      fA       UfA      �A       �U��A      B       U                          @A      oA       ToA      �A       \�A      �A       |��A      �A       �T��A      B       T                        @A      iA       QiA      �A       ]�A      �A       �Q��A      B       Q                        SA      �A       V�A      �A       v�~��A      �A       V�A      B       u�                       �A      �A       0��A      �A       S�A      �A       s��A      �A       ^                   wA      �A       \�A      �A       ^                      �F      �F       U�F      0G       ]0G      3G       �U�                      �F      �F       T�F      ,G       V,G      3G       �T4�T����4,( �                      �F      �F       Q�F      G       ^G      3G       �Q�                     �F      �F       0��F      G       SG      G       s�                    �G      �G       U�G      �G       �U�                    �G      �G       T�G      �G       �T�                               E      hE       UhE      F       ��~F      0F       �U�0F      �F       ��~�F      �F       U�F      �F       ��~�F      �F       U                         E      HE       THE      F       \0F      �F       \�F      �F       T                               E      hE       QhE      F       ]F      0F       �Q�0F      �F       ]�F      �F       Q�F      �F       ]�F      �F       Q                    F      F       P�F      �F       P                    8E      -F       ^0F      �F       ^                         WE      hE       0�hE      �E       S�E      �E       s�0F      �F       S�F      �F       0�                          �E      �E       0��E      �E       P�E      �E       X�E      �E       P0F      3F       P^F      zF       P                      �E      �E       U0F      8F       UYF      vF       U                      �E      F       P6F      8F       P{F      �F       P                     hE      �E       V�E      F       vh�0F      �F       V                    tE      �E       Y0F      zF       Y                        xE      �E       [0F      3F       [3F      8F       v8F      zF       [                          xE      �E       	���E      �E       X�E      �E       	���E      �E       X0F      3F       X8F      ^F       	��^F      zF       X                    xE      �E       	��0F      3F       	��8F      ^F       	��^F      zF       P                          �E      �E       y �E      �E       R�E      �E       y 0F      3F       R^F      dF       RdF      hF       y q "8                      @      R       UR      �       �U��      �       U                      @      �       Q�      �       �Q��      �       Q                            G      n       Pn      �       �U#��      �       P�      �       �U#��      �       P�      �       u�                          Z      p       0�p      s       p�s      {       P{      �       p��      �       R                      @      j       Uj      �       �U��      6       U                      @      q       Tq      �       �T��      6       T                          @      u       Qu      �       �Q��      �       Q�      +       �Q�+      6       Q                  G      6       X                                 Y      u       0�u      {       p�{      �       P�      �       p��      �       0��      �       p��      �       P�      �       p��      �       S                        �             S             x �t x �t ����,( �      *       S*      +       x �t x �t ����,( �                      �@      �@       U�@      )A       �U�)A      <A       U                          �@      �@       T�@      �@       [�@      �@       {��@      )A       �T�)A      <A       T                        �@      �@       Q�@      'A       S'A      )A       �Q�)A      <A       Q                      �@      (A       V)A      ;A       V;A      <A       u�                       �@      �@       0��@      �@       P�@      �@       p��@      
A       Q                     �@      �@       [�@      
A       Q
A      (A       v��Tv��T����,( �                    B      9B       U9B      �C       �U�                            B      5B       T5B      KB       VKB      RB       �T�RB      �C       V�C      �C       �T��C      �C       V                    )B      BB       ZRB      tB       Z                           )B      BB       0�RB      xB       0�xB      |B       P|B      �C       ^�C      �C       �T�C      �C       ^                    �B      �B       0�VC      ^C       0�^C      nC       \                        0B      JB       SRB      QC       SQC      ^C       s�~��C      �C       S                           2      62       U62      `2       �U�`2      h2       Uh2      �2       �U��2      �2       U                         2      �2       T�2      �2       U�2      �2       �T��2      �2       T                    2      =2       1��2      �2       1�                      �       �        U�       5       �U�5      >       U                  �       >       R                   �       �        0��              Q                   �       -       p t "#�-      2       p t "@�                   �       -      	 r p "#��-      2      	 r p "#��                                  �	      
       U
      
       V
      2
       �U�2
             V      �       v�z��      �       �U��      �       U�             V      ~       �U�                            �	      
       T
      +
       \+
      2
       �T�2
      �       \�      �       T�      ~       \                              �	      
       Q
      -
       ]-
      2
       �Q�2
      �       ]�      �       s�      �       Q�             ]      4       s                         �	      (
       S2
      �       S�      �       S�      �       P�      ~       S                      �	      1
       _2
      �       _�      ~       _                 
      2
       3�                 (      B       2�                  D      `       1�                        �      C       UC      �       S�      �       �U��      �       S                                    �      k       Tk      �       ^�      �       �T��      �       T�      G       ^G      �       �T��      �       ^�      �       T�      Q       �T�Q      �       ^                                  �      !       Q!      j       _j      �       �Q��      �       Q�      �       _�      �       �Q��      �       _�      �       Q�      �       �Q�                            �      $       R$      �       ]�      �       R�      �       ]�      �       ]�      �       R                       �      C       UC      �       S�      �       �U��      �       S                                  �      �       P�      F       \F      V       PV      �       \�      _       \_      �       0��      �       P�      �       \�      �       \                    �      �       V�      �       V                               ]      _      
 p 3 $0)�_      |      
 } 3 $0)�|      �       T�      �       s��      �       ��g�      �       ��g�      �      
 } 3 $0)��      �       ��g                   �      �       v���      �       v��                     �      P       v��      �       v��      �       v�                              �             P      P       v�#P             ��g�      �       v�#�      G       ��g�      �       ��g�      �       v�#                       �      �       _�T��      �       _���g��      �       _���g��      �       _���g�                     �      �       0��      �       1��      �       0��      �       1��      �       0�                         �      N       0�N      �       1��      �       0��      �       1��      �       0��      �       1�                  �      G       ]                   �      �       s0��      �       s0�                  �      �      	 q 0$0&�                   �      X       ��h�      Q       ��h                         �             ��h#�      �       ��h#�             P      G       pp�G      Q       P                   �             s��      �       s�                   �             s��      �       s�                      %       s�                          %       T%      %      
 p t "#���                        %       t ?&�%      %       P                7      F       s�                    ?      F       RF      F      
 p r "#���                  ?      F       r ?&�F      F       P                  �             p              pp                                Q            
 q x "#���                               q ?&�             X                   -      4       Q4      4      
 q x "#���                  -      4       q ?&�4      4       X                {      �       ��g                {      �       s�                    �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       ��g                �      �       s�                    �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                          p      �       U�      �       T�      �	       ]�	      �	       �U��	      �	       U                        p      �       T�      C	       VC	      �	       �T��	      �	       T                        p      �       Q�      A	       \A	      �	       �Q��	      �	       Q                    p      �       R�      �	       �R�                          p      �       X�      C	       SC	      �	       �X��	      �	       S�	      �	       X                         p      �       U�      �       T�      �	       ]�	      �	       �U��	      �	       U                         p      �       u���      �       t���      �	       }���	      �	       �U#���	      �	       u��                 p      r       u�                     9	      R	       0�R	      [	       1�[	      �	       0��	      �	       1��	      �	       0�                      �      �       PC	      [	       Pg	      {	       P                        @      �       U�      �       T�      Z       VZ      a       �U�                      @      j       Tj      \       \\      a       �T�                      �      �       P�      ^       ]^      a       P                                0�      B       S                       @      �       u���      �       t���      Z       v��Z      a       �U#��                  `      `       ^                      �      �       U�      0       S0      1       �U�                    �      �       T�      1       �T�                   �      &       P&      +       �L                        &       s                        �      C       UC      �       S�      �       �U��      �       S                          �      G       TG      �       ]�      �       �T��      �       ]�      �       T                        �      �       Q�      �       _�      �       �Q��      �       _                      �      G       RG      �       ��k�      �       R                    �      �       V�      �       V                   �      �       v���      �       v��                             �      H       0�H      ]       P�      �       P�             PQ      �       P�      �       P�      �       0�                    �      �       ^�      �       ^                        �      �       P�             w       �       ��k�      �       w                     �      �       \�      �       \                    �>      ?       U?      r?       �U�                    �>      �>       T�>      r?       �T�                    �>      ?       Q?      r?       �Q�                   �>      ?       U?      r?       �U�                       �>      �>       P�>      ?       u�?      W?       �U#�Z?      r?       �U#�                       �>      �>       P�>      ?       u�?      W?       �U#�Z?      r?       �U#�                   �>      W?       RZ?      r?       R                      �>      ?       Q?      W?       �Q�Z?      r?       �Q�                      �>      �>       T�>      W?       �T�Z?      r?       �T�                   ?      W?       XZ?      r?       X                      ?      ?       P7?      W?       PZ?      h?       P                      ?      ?       x p "�?      ?       TI?      W?       T                      ?      W?       QZ?      d?       Qd?      r?       �T����@$�Q����!�                      ?      ?       UD?      W?       UZ?      r?       U                    4      4       U4      4       �U�                    4      4       T4      4       �T�                                      �4      #5       U#5      =5       �U�=5      6       U6      66       �U�66      B8       UB8      �8       \�8      �8       �U��8      9       U9      9       \9      I9       �U�I9      �>       U                    �4      5       T5      �>       �T�                                      �4      #5       Q=5      6       Q6      66       �Q�66      K8       QK8      W8       �Q�W8      \8       p �8      9       Q9      I9       �Q�I9      �9       Q�9      �9       P�9      �>       Q                                        �4      #5       R#5      =5       �R�=5      6       R6      66       �H66      K8       RK8      \8       �H\8      �8       �R��8      9       R9      (9       �H(9      >9       R>9      I9       �HI9      �>       R                                  �4      #5       X#5      =5       �X�=5      6       X6      66       �X�66      K8       XK8      �8       �X��8      9       X9      I9       �X�I9      �>       X                                                                                                                       �4      #5       0�=5      =5       0�=5      d5       2�d5      d5       0�d5      �5       2��5      �5       0��5      �5       2��5      �5       0��5      �5       1��5      6       0�6      6       p�6      66       V66      �6       0��6      �6       8��6      �6       0��6      7       8�7      )7       0�)7      S7       2�S7      S7       0�S7      }7       1�}7      }7       0�}7      �7       4��7      �7       0��7      �7       1��7      �7       0��7      �7       2��7      �7       0��7      '8       2�'8      }8       0�}8      �8       V�8      �8       P�8      �8       0��8      �8       4��8      9       0�9      9       p�9      I9       VI9      I9       0�I9      u9       4�u9      �9       0��9      �9       V�9      �9       0��9      :       4�:      :       0�:      -:       4�-:      P:       0�P:      u:       1�u:      �:       0��:      �:       8��:      �:       0��:      �:       1��:      �:       0��:      ;       8�;      ;       0�;      K;       8�K;      K;       0�K;      u;       1�u;      u;       0�u;      �;       1��;      �;       0��;      �;       2��;      �;       0��;      <       1�<      <       0�<      -<       4�-<      -<       0�-<      O<       8�O<      _<       0�_<      �<       2��<      �<       0��<      �<       1��<      �<       0��<      �<       2��<      =       0�=      1=       2�1=      1=       0�1=      ]=       1�]=      ]=       0�]=      �=       4��=      �=       0��=      �=       2��=      �=       0��=      �=       1��=      �=       0��=      >       2�>      3>       1�3>      B>       2�B>      R>       4�R>      �>       8�                              5      75       S75      =5       �X0�X0*( �=5      �8       S�8      �8       �X0�X0*( ��8      *>       S*>      3>       x 0x 0*( �3>      �>       S                                     5      #5       U#5      =5       �U�=5      6       U6      66       �U�66      B8       UB8      �8       \�8      �8       �U��8      9       U9      9       \9      I9       �U�I9      �>       U                                     5      #5       u��#5      =5       �U#��=5      6       u��6      66       �U#��66      B8       u��B8      �8       |���8      �8       �U#���8      9       u��9      9       |��9      I9       �U#��I9      �>       u��                               ;      F;       0�F;      K;       PR>      Y>       0�Y>      ^>       P^>      e>       0�e>      j>       Pj>      q>       0�q>      v>       P                               �:      �:       0��:      �:       Pv>      }>       0�}>      �>       P�>      �>       0��>      �>       P�>      �>       0��>      �>       P                   5      #5       0�'8      W8       0�W8      \8       1�                  L8      \8       P                      �       �        U�       �        t�}��       �        �U�                        �       �        T�       �        P�       �        U�       �        �T�                      !      6!       U6!      }!       �U�}!      �!       U                            !      6!       T6!      d!       Vd!      i!       �T�i!      x!       Vx!      }!       �T�}!      �!       T                           !      6!       0�6!      L!       s�L!      c!       Sc!      i!       Pi!      w!       s�}!      �!       0�                 L!      W!       s 3$| "                    �>      �>       U�>      �>       �U�                    �>      �>       T�>      �>       �T�                      �>      �>       Q�>      �>       P�>      �>       �Q�                      �>      �>       R�>      �>       Q�>      �>       �R�                       4      T4       UT4      �4       �U��4      �4       U                           4      T4       TT4      �4       ^�4      �4       �T��4      �4       ^�4      �4       T                           4      T4       QT4      �4       ]�4      �4       �Q��4      �4       ]�4      �4       Q                           4      T4       RT4      �4       _�4      �4       �R��4      �4       _�4      �4       R                      54      �4       \�4      �4       \�4      �4       u�                      L4      T4       0�T4      �4       S�4      �4       S                      T4      i4       Vx4      �4       V�4      �4       V                        `I      �I       U�I      �I       S�I      �I       �U��I      �M       S                        `I      I       TI      �I       _�I      �I       �T��I      �M       _                       =J      �J       ]�J      �J       ]�K      �L       ]�M      �M       ]                    xI      �I       \�I      �M       \                           xI      �I       0��I      �I       P�I      �I       V�I      �I       P�I      �K       V�K      �K       0��K      �M       V                       �I      �I       U�I      �I       S�I      �I       �U��I      �M       S                       �I      �I       u���I      �I       s���I      �I       �U#���I      �M       s��                       iJ      �J       � �K      *L       Q*L      mL       � �M      �M       �                  �K      �M       V                   �K      sM       _�M      �M       _�M      �M       _                   �K      sM       S�M      �M       S�M      �M       S                          �K      �K       P�K      mL       8mL      sM       ��~�M      �M       8�M      �M       ��~�M      �M       ��~                	     �K      *L       Q*L      mL       � �M      �M       �                 
         �K      ZL       RZL      mL       � �L      sM       ]�M      �M       R�M      �M       ]                           �K      �K       q� ��K      
L       P
L      L       p�L      7L       P7L      :L       ~~�:L      �L       ^�L      0M       ~|�0M      sM       ^�M      �M       ^                         �L      �L       P�L      �L       Q�L      0M       ��0M      IM       Q�M      �M       Q�M      �M       ��                       �K      �K       q� ��8$q� ��!
����K      �K       p 8$q� ��!
����K      *L       q� ��8$q� ��!
���*L      :L       � #d��8$� #c��!
���                          �L      �L       P�L      �L       s��L      sM       ���M      �M       s��M      �M       ��                       �L      �L       0��L      �L       T�L      �L       p �L      �L       T�M      �M       T                 �L      �L       0�                         )        U                         )        T                         )        R                           %        Q%       )        t �����@$t�����!�                        `      t       Ut      �       V�      �       U�      �       �U�                        `      p       Tp      �       S�      �       T�      �       �T�                    �?      7@       Q\@      �@       Q                    �?      7@       T\@      �@       T                    �?      7@       U\@      �@       U                           D      %D       T%D      (D       �T�(D      QD       TQD      E       XE      E       T                    D      QD       UE      E       U                           (D      QD       0�[D      �D       V�D      �D       v��D      �D       z��D      �D       V�D      E       v�                          [D      iD       0�iD      �D       R�D      �D       r��D      �D       R�D      �D       r��D      �D       R                        D      QD       0�[D      �D       �G�D      �D       1��D      E       �GE      E       0�                        [D      iD       @<$�iD      �D       P�D      �D       P�D      �D       P                      tD      �D       T�D      �D       u r 3$q " v  $0)( ��D      �D       T                   �D      �D       T�D      �D       u r 3$q " v  $0)( �                 �D      �D       P                      �D      �D       P�D      �D      
 p t "#����D      �D       P                   �D      �D       p ?&��D      �D       T                      @G      NG       UNG      oG       SoG      qG       �U�                      @G      RG       TRG      pG       VpG      qG       �T�                    @G      [G       Q[G      qG       �Q�                  SG      qG       P                    WG      [G       Q[G      nG       �Q�                  WG      nG       V                  WG      nG       S                 �G      �G       U                    �G      �G       S�G      �G       S                    �G      �G       P�G      �G       P                        pH      �H       U�H      �H       S�H      �H       �U��H      �H       U                       pH      �H       U�H      �H       S�H      �H       �U��H      �H       U                      ~H      �H       U�H      �H       S�H      �H       �U�                  �H      �H       P                        �H      �H       U�H      5I       ^5I      GI       �U�GI      UI       ^                        �H      �H       T�H      5I       ��5I      GI       �T�GI      UI       ��                    �H      �H       Q�H      UI       �Q�                   �H      �H       Q�H      UI       �Q�                        �H      �H       0��H      �H       s�I      5I       SGI      UI       s�                     �H      �H       VI      5I       VGI      UI       V                          �M      �M       U�M      N       SN      N       �U�N      rN       SrN      vN       �U�                          �M      �M       T�M      N       \N      N       �T�N      uN       \uN      vN       �T�                          �M      �M       Q�M      N       VN      N       �Q�N      sN       VsN      vN       �Q�                         �M      N       PN      0N       P1N      ?N       P@N      RN       PmN      vN       P                 DN      mN       V                 DN      mN       \                 DN      mN       S                      DN      dN       0�dN      hN       PhN      mN       �LmN      mN       P                 �             U                        @1      i1       Ui1      �3       V�3      �3       �U��3      �3       U                       @1      i1       Ui1      �3       V�3      �3       �U��3      �3       U                  b1      �3       ^                 b1      i1       P                  q1      �3       S                 z1      �3       S                  �1      �3       \                    �1      �1       ]�1      �1       }�                  �1      �1       T                  �1      �1       \                 �1      &2       s��                 *2      12       P                  *2      �2       s�
�                 *2      �2       ]                 *2      �3       s�
�                 *2      Q2       ]                     �2      �2       s���2      �2       T�2      �2       s��                 �2      �2       \                 �2      �2       s                 �2      �2       s�&�                 �3      �3       V                  �3      �3       P                                                                        �H      I       UI      fJ       SfJ      {J       �U�{J      O       SO      pO       \pO      QS       SQS      �U       �U��U      PV       SPV      CZ       �U�CZ      xZ       SxZ      �[       �U��[      �[       S�[      G^       �U�G^      �i       S�i      �i       ]�i      <j       S<j      Mj       \Mj      �j       S�j      >k       ]>k      "m       S"m      0m       ]0m      �n       S�n      �n       \�n      �n       S�n      �n       \�n      �n       S�n      �n       \�n      o       S                                                              �H      �H       T�H      WJ       ]WJ      {J       �T�{J      �M       ]�M      �P       �T��P      �R       ]�R      �U       �T��U      PV       ]PV      CZ       �T�CZ      xZ       ]xZ      �[       �T��[      �[       ]�[      G^       �T�G^      �^       ]�^      _       �T�_      �_       ]�_      Rj       �T�Rj      �j       ]�j      uk       ��}uk      m       �T�m      "m       ]"m      :m       ��}:m      o       �T�                                                              �H      
I       Q
I      WJ       ^WJ      {J       �Q�{J      �M       ^�M      �P       �Q��P      �R       ^�R      �U       �Q��U      PV       ^PV      CZ       �Q�CZ      xZ       ^xZ      �[       �Q��[      �[       ^�[      G^       �Q�G^      �^       ^�^      _       �Q�_      �_       ^�_      Rj       �Q�Rj      �j       ^�j      l       ��}l      m       �Q�m      "m       ^"m      :m       ��}:m      o       �Q�                              �H      
I       R
I      J       ��}J      {J       �R�{J      �J       ��}�J      �P       �R��P      �P       ��}�P      o       �R�                                  �H      
I       X
I      WJ       ��}WJ      {J       �X�{J      �J       ��}�J      �P       �X��P      Q       ��}Q      �U       �X��U      +V       ��}+V      o       �X�                                                             �H      �H       T�H      WJ       ]WJ      {J       �T�{J      �M       ]�M      �P       �T��P      �R       ]�R      �U       �T��U      PV       ]PV      CZ       �T�CZ      xZ       ]xZ      �[       �T��[      �[       ]�[      G^       �T�G^      �^       ]�^      _       �T�_      �_       ]�_      Rj       �T�Rj      �j       ]�j      uk       ��}uk      m       �T�m      "m       ]"m      :m       ��}:m      o       �T�                   WJ      fJ       ;�>Z      CZ       P                          I      ,I       P,I      PJ       \{J      �J       \�P      Q       \�U      &V       \                         :I      >I       P>I      WJ       ��}{J      K       ��}�P      Q       ��}�U      +V       ��}                          LI      PI       PPI      WJ       ��}{J      K       ��}�P      Q       ��}�U      +V       ��}                  QI      vI       P                         �I      �I       P�I      WJ       ��}{J      K       ��}�P      Q       ��}�U      +V       ��}                	           �H      J       1�J      WJ       ��}{J      �J       1��J      K       ��}�P      �P       1��P      Q       0��U      +V       ��}                
                                                               �H      BJ       0�BJ      WJ       1�{J      �J       0��J      �M       \�M      �P       ��~�P      Q       0�Q      �R       \�U      +V       0�+V      PV       \CZ      xZ       \�[      �[       \G^      �^       \�^      _       ��~_      �_       \�_      �`       ��~�b      �b       ��~.f      �f       ��~�f      ,h       ��~�h      �h       ��~�h      �i       ��~j      j       ��~<j      Rj       ��~Rj      �j       \�j      �j       ��~�j      Ck       ^Ck      jk       ��~jk      l       \l      m       ��}m      "m       \"m      5m       ^5m      Vm       ��~Vm      �m       ��}�m      o       ��~                         �H      �I       0��I      WJ       1�{J      �J       0��J      K       ��~�P      Q       1��U      +V       1�                        �H      WJ       V{J      L       V�P      ,Q       V�U      +V       V                 (I      ,I       U                          :I      >I       P>I      WJ       ��}{J      K       ��}�P      Q       ��}�U      +V       ��}                 aI      vI       }�                          �I      �I       P�I      WJ       ��}{J      K       ��}�P      Q       ��}�U      +V       ��}                           �J      �J       0��J      �J       P�J      K       RK      DK       [DK      �K       ��}Q      Q       ��}                   S      YS       {��YS      �S       ��}#��                    �J      �J       P�J      K       ��}                           �W      X       
�X      X       PX      5X       0�5X      uX       s ��uX      �X       S�X      �X       S�X      �X       }                      �S      
T       P
T      T       {�T      )T       s                  )S      YS       }�                   )S      YS       }�YS      �S       S                   )S      ;S       ~ @%�;S      �S       ^                        �S      �U       VPV      CZ       VxZ      �[       V�[      G^       V                         �S      �S       {���S      �U       v0�PV      CZ       v0�xZ      �[       v0��[      G^       v0�                         �S      �S       {���S      �U       v(�PV      CZ       v(�xZ      �[       v(��[      G^       v(�                    �S      T       S�Z      �[       S                      )T      �T       \�T      �U       \PV      XV       \                     )T      �T       ���T      �U       ��PV      XV       ��                     �T      �T       |� �MU      �U       |� �PV      XV       |� �                     �T      �T       |� �MU      �U       |� �PV      XV       |� �                     �T      �T       |� �MU      �U       |� �PV      XV       |� �                      �T      �T       ^iU      �U       ^PV      XV       ^                  bT      �T       ^                       jV      �W       0��[      :]       0�W]      |]       0�|]      �]       P�]      G^       \                  �[      	\       P                 \      	\       P                  \      	\       U	\      
\       ��}                 
\      
\       P                  �W      �W       P                         �W      �W       P\      \       P\       \       p� \      -\       P-\      1\       p�1\      6\       PW]      t]       P                      �W      �W       T\      6\       TW]      h]       T                 p]      t]       T                  p]      t]       Ut]      |]       ��}                 |]      |]       P                   |]      �]       P�]      G^       \                 |]      G^       S                  �]      G^       ^                  �]      �]       P                                  �]      �]       1��]      �]       2q ��]      �]       2q ��]      �]       r��]      ^       R^      ^       p�^      -^       P;^      ?^       P?^      G^       R                  ]      +]       P                 ]      +]       P                ]      ,]       ��}                 ,]      ,]       P                  :X      SX       P                �W      �W      
 �F     �                  �W      �W       U�W      �W       ��}                 �W      �W       P                         \\      e\       Pe\      g\       Ug\      �\       X�\      �\       R�\      �\       X                         \\      �\       0��\      �\       q x #��\      �\       q x ��\      �\       q x #��\      �\       7��\      �\       r x #�                  k\      �\       U                         k\      �\       1��\      �\       Z�\      �\       Z�\      �\       0��\      �\       Z�\      �\       1�                        �X      Y       QY      Y       }� Y      /Y       R/Y      EY       }�                        �X      Y       0�Y      EY       QuY      �Y       S�Y      �Y       S�Z      �Z       0�                  �X      �X       {���Z      �Z       {��                   %Z      CZ      
 ��F     ��[      �[      
 ��F     �R]      W]      
 ��F     �                                                                       �J      �M       \�M      �P       ��~Q      �R       \+V      PV       \CZ      \Z       \G^      �^       \�^      �^       \�^      _       ��~_      �_       \�_      �`       ��~�b      �b       ��~.f      �f       ��~�f      ,h       ��~�h      �h       ��~�h      �i       ��~j      j       ��~<j      Rj       ��~Rj      �j       \�j      �j       ��~�j      Ck       ^Ck      jk       ��~jk      l       \l      m       ��}m      "m       \"m      5m       ^5m      Vm       ��~Vm      �m       ��}�m      o       ��~                 �J      K       ��}                                               �J      �M       ]�M      �P       �T�Q      �R       ]+V      PV       ]CZ      \Z       ]G^      �^       ]�^      �^       ]�^      _       �T�_      �_       ]�_      Rj       �T�Rj      �j       ]�j      uk       ��}uk      m       �T�m      "m       ]"m      :m       ��}:m      o       �T�                         �J      �J       P�J      K       RK      DK       [DK      �K       ��}Q      Q       ��}                                               �J      �M       ^�M      �P       �Q�Q      �R       ^+V      PV       ^CZ      \Z       ^G^      �^       ^�^      �^       ^�^      _       �Q�_      �_       ^�_      Rj       �Q�Rj      �j       ^�j      l       ��}l      m       �Q�m      "m       ^"m      :m       ��}:m      o       �Q�                                                           �J      O       SO      pO       \pO      �P       SQ      �R       S+V      PV       SCZ      \Z       SG^      �^       S�^      �i       S�i      �i       ]�i      <j       S<j      Mj       \Mj      �j       S�j      >k       ]>k      "m       S"m      0m       ]0m      �n       S�n      �n       \�n      �n       S�n      �n       \�n      �n       S�n      �n       \�n      o       S                   �J      L       VQ      ,Q       V                 �J      K       ��}                          \K      vK       PvK      )L       ��}Q      �R       ��}+V      PV       ��}]^      v^       ��}                   =K      �K       ��}#��Q      Q       ��}#��                                           �L      �L       R�L      �P       ��~CZ      \Z       ��~G^      ]^       0�v^      �^       R�^      �^       ��}�^      �`       ��~�b      �b       ��~.f      �f       ��~�f      ,h       ��~�h      �h       ��~�h      �i       ��~j      j       ��~<j      o       ��~                          �M      �N       0��N      �N       P"O      ,O       v�3$s "�^      �_       0�Rj      :m       0�Vm      o       0�                            �N      �N       R�N      �N       r��N      "O       R"O      AO       VAO      EO       Q`O      �O       V                    �M      �M       P_      %_       P                         �M      &N       ��}�^      �^       ��}_      �_       ��}Rj      :m       ��}Vm      o       ��}                                             �M      &N       S�^      �^       S_      �_       SRj      �j       S�j      >k       ]>k      "m       S"m      0m       ]0m      :m       SVm      �n       S�n      �n       \�n      �n       S�n      �n       \�n      �n       S�n      �n       \�n      o       S                      �M      �M       {�'�_      %_       {�'�%_      G_       ��}#�'�                             �M      �M       R�M      &N       ��}�^      �^       ��}_      _       R_      �_       ��}Rj      :m       ��}Vm      o       ��}                                      �M      �M       0��M      �M       ��}N      N       TN      N       ��}N      &N       0��^      �^       0�_      �_       0�Rj      �j       0��j      �j       P�j      m       ��}m      "m       0�"m      :m       ��}Vm      o       ��}                                    �j      l       Vl      m       ��~"m      :m       VVm      nm       ��~nm      �m       P�m      �m       ��~�m      �n       ��}�n      �n       P�n      �n       ��}o      o       ��}                           dl      �l       \�l      m       \�n      �n       S�n      �n       S�n      �n       T�n      �n       S                      {_      �_       ��}Rj      l       ��}"m      :m       ��}                  �_      �_       p 
���                      tj      �j       P�j      �k       ��~"m      :m       ��~                    Cl      m       ]Vm      dm       ]                 rl      �l       V                  wl      �l       ��~                  �l      �l       ��~                  �l      �l       P                  �m      �m      
 v 4$��}"�                  �O      �O       T                      �O      �O       U�O      fP       S:m      Vm       S                    �O      fP       V:m      Vm       V                    �O      P       ��}#�&�Jm      Vm       ��}#�&�                    �O      P       PJm      Vm       P                    P      #P       p 
���#P      .P       P                  %Q      _Q       P                                `      !`       p ����
��.��}�0.�!`      �`       ��}�
��.��}�0.��b      �b       ��}�
��.��}�0.�.f      �f       ��}�
��.��}�0.��f      ,h       ��}�
��.��}�0.��h      �h       ��}�
��.��}�0.��h      �i       ��}�
��.��}�0.�j      j       ��}�
��.��}�0.�                              !`      �`       ��}�
��.��}�0.��b      �b       ��}�
��.��}�0.�.f      �f       ��}�
��.��}�0.��f      ,h       ��}�
��.��}�0.��h      �h       ��}�
��.��}�0.��h      �i       ��}�
��.��}�0.�j      j       ��}�
��.��}�0.�                        !`      �`       P.f      af       P�f      �f       P�h      'i       P                              !`      �`       ��}�b      �b       ��}.f      �f       ��}�f      ,h       ��}�h      �h       ��}�h      �i       ��}j      j       ��}                          !`      a       S�b      �b       S.f      �h       S�h      �i       S�i      �i       ]�i      <j       S                      !`      a       \�b      �b       \.f      �h       \�h      <j       \                              !`      �`       ��}�b      �b       ��}.f      �f       ��}�f      ,h       ��}�h      �h       ��}�h      �i       ��}j      j       ��}                                          &`      y`       Ry`      �`       U�`      �`       ��}�b      �b       ��}.f      Sf       RSf      �f       ��}�f      �f       R�f      ,h       ��}�h      �h       ��}�h      �h       ��}�h      i       Ri      �i       ��}j      j       ��}                          �g      �g       P�g      �g       ^�g      h       ~ r "�h      h       Ph      )h       ^                          �g      �g       ]�g      �g       }��g      $h       ]Vi      ^i       ]�i      �i       v�                        �g      �g       P�g      �g       T�g      h       Ph      h       P                   �g      �g       0��g      h       R                          ea      �a       Q�a      b       {��b      �b       Q�b      7c       {�7c      Rc       Q                         ea      �a       ��}�b      �b       ��}�b      c       ��}7c      �c       ��}�e      f       ��}                        ea      �b       S�b      �b       S�b      �b       S�b      .f       S                        ea      �b       \�b      �b       \�b      �b       \�b      .f       \                          ea      b       {��b      �b       ��}#���b      Rc       {��Rc      �c       ��}#���e      �e       ��}#��                                  �b      �b       ��}�c      �c       p ���c      �d       v ���d      e       v ��e      e       Pe      �e       ��}�e      �e       p ���e      f       v ��f      .f       ��}                                    *b      Sb       p�Sb      Wb       P_b      �b       p��b      �b       R�c      �c       0��c      �d       ��}�d      �d       ��}e      �e       ��}�e      �e       1��e      f       Qf      )f       ��}                    Re      �e       Pf      .f       P                           d      (d       Q(d      \d       ��}\d      �d       QAe      ce       v ���e      �e       t p "����e      �e       t r "1���                          *b      :b       R:b      >b       Q>b      Lb       p 1${ "#��
���kb      ob       Rob      zb       p 1${ "#��
���                   *b      >b       0�>b      Sb       q 
���kb      ob       0�                    *b      :b       R:b      >b       Q>b      >b       p 1${ "#��
���                  *b      >b       0�>b      >b       q 
���                  4d      \d       P                       �c      �c       1��c      �d       ��}�d      �d       U�d      �d       ��}                  \d      �d       R                     qe      se       0�se      �e       Rf      .f       R                        �e      �e       T�e      �e       t p "��e      �e       t p "#��e      f       t r "�f      f       t p "�                            @       U@      [       S[      d       �U�                            4       P4      @       u@      D       s                         4       p�	4      D       Q                  (      c       V                  E      O       P                  P      [       P                          �      �       U�      �       V�      �       �U��             V             �U�                          �      �       T�      l       Sl      �       �T��      
       S
             �T�                         �      �       U�      �       V�      �       �U��             V             �U�                    (      5       P5      �       ]                 �      �       U                 �      �       u�                 1      ]       v                   I      �       ^                  P      �       _                  W      �       \                  e      r       P                   r      �       P�      �       ~ s "#�                      r      �       R�      �       ���      �       R                       �      �       P�      �       w �      �       Y�      �       Y                    �      �       Q�      �       Q                      @      X       UX      (       V(      1       �U�                    @      \       T\      1       �T�                     @      X       UX      (       V(      1       �U�                    f      v       Pv              ]                 r      �       v                   �              ^                  �              _                  �              \                  �      �       P                   �      �       P              ~ s "#�                      �      �       R�      �       ��              R                       �      �       P�      �       w �      �       Y              Y                    �      �       Q              Q                               7       U7      �       V�      �       �U��      ^       V                              7       U7      �       V�      �       �U��      ^       V                          D      T       PT      �       \�      4       \4      =       PK      ^       \                  T      p       P                      l      �       ]�      4       ]K      ^       ]                           l      ~       0�~      �       P�      �       P�      �       _�      4       ��}K      ^       ��}                 l      p       U                  �      �       P                 �             } s "#�                    p      }       U}      �       Q                    s      }       u��}      �       q��                                              �      �       0��      �       P�      �       p��      �       0��      �       P�      �       p��      �       0��      �       P�             p�             0�      -       P-      1       p�~      �       0��      �       P�      �       p��      �       0��      �       P�      �       p�                            �      �       U�      �       U�             U      w       U~      �       U�      �       U                      @      Y       UY      �       �U��      �       U                 @      B       u #�                     @      Y       UY      �       �U��      �       U                 @      B       u                  @      B       u #�	                        Q      �       V�      �       T�      �       V�      �       p                     o      z       Pz      �       \                    �      �       P�      �       s�                        �D      ,E       U,E      �F       ^�F      �F       �U��F      �H       ^                                        �D      VE       TVE      �F       V�F      �F       �T��F      �F       V�F      �F       �T��F      �G       V�G      XH       �T�XH      qH       VqH      �H       �T��H      �H       V�H      �H       �T��H      �H       V                          �D      E       QE      �E       ��~�E      �F       �Q��F      �F       ��~�F      �H       �Q�                        �D      �D       R�D      �F       \�F      �F       �R��F      �H       \                          �D      E       XE      �E       ��~�E      �F       �X��F      �F       ��~�F      �H       �X�                      �D      wE       YwE      �E       ���E      �H       �Y�                    �D      �E       � �F      �F       �                     �D      �E       ��F      �F       �                                                     �E      �E       R�E      fF       0�fF      qF       PqF      �F       _�F      �F       _�F      �F       P�F      �F       0��F      G       PG      G       _G      +G       P+G      +G       0�@G      CG       PCG      wG       _wG      �G       P�G      H       _H      1H       P1H      5H       _5H      OH       POH      SH       _XH      �H       _�H      �H       P                     5E      �F       ^�F      �F       �U��F      �H       ^                     5E      �F       ~���F      �F       �U#���F      �H       ~��                        @E      HE       PHE      �E       �#��E      �E       ��~�F      �F       ��~                   @E      �F       s  $0)��F      �H       s  $0)�                        SE      �E       _�E      �F       	�0s  $0)( 
�#`��F      �F       _�F      �F       	�0s  $0)( 
�#`��F      �H       	�0s  $0)( 
�#`�                  �H      �H       V                  VE      �E       0��F      �F       0�                    VE      �E       _�F      �F       _�F      �F       	�0s  $0)( 
�#`�                    VE      eE       TeE      �E       �                   VE      �E       ^�F      �F       ^                      VE      wE       YwE      �E       ���E      �E       �Y��F      �F       �Y�                  VE      �E       ��~��F      �F       ��~�                  [E      �E       ]�F      �F       ]                   yF      �F       VXH      qH       V                   yF      �F       ]XH      qH       ]                 XH      kH       v                  �F      �F       ��~�                 �F      �F       ��~                          �8      9       U9      9       �U�9      69       U69      �9       t��9      };       ]                              �8      9       T9      9       �T�9      �9       T�9      :       z�:      �:       \�:      �:       T�:      };       \                                  �8      9       Q9      9       �Q�9      �9       Q�9      �9       t��9      :       z�:      �:       �Q��:      �:       Q�:      �:       t��:      };       �Q�                                    �8      9       R9      9       �R�9      99       R99      �9       Y�9      �9       t��9      :       z�:      �:       �R��:      �:       Y�:      �:       t��:      };       �R�                                     �8      9       0�9      >:       0�>:      Q:       PQ:      T:       VT:      \:       P\:      �:       V�:      �:       0��:      �:       P�:      �:       V�:      �:       P�:      };       V                             �8      9       T9      9       �T�9      �9       T�9      :       z�:      �:       \�:      �:       T�:      };       \                             �8      9       t��9      9       �T#��9      �9       t���9      :       z�#��:      �:       |���:      �:       t���:      };       |��                    �8      9       S9      };       S                    �9      �9       a��:      �:       [                    �9      �9       t��9      :       zn                    �9      �9       t��9      :       zl                  �9      (:       V�:      �:       V                    �9      �9       Q�9      :       ��~                      �9      �9       t���9      :       z�#��:      (:       |���:      �:       |��                    �9      �9       Y�9      :       ��                  �9      (:       ��~��:      �:       ��~�                  �9      (:       ^�:      �:       ^                a:      }:       \                 }:      �:       ��~�                 }:      �:       ��~                    P      Y       UY      Z       �U�                    P      Y       TY      Z       �T�                    P      Y       QY      Z       �Q�                    P      Y       RY      Z       �R�                    P      Y       XY      Z       �X�                 P      Y       u�                    @      h       Uh      {       �U�                    @      e       Te      {       �T�                    @      l       Ql      {       �Q�                    @      p       Rp      {       �R�                                �      �       U�      �       �U��             U      i       ]i      k       Xk      �       �U��      �       U�      Y       �U�                            �      �       T�      �       �T��             T      �       ���      �       T�      Y       ��                            �      �       Q�      �       �Q��      �       Q�      �       ���      �       Q�      Y       ��                            �      �       R�      �       �R��             R      �       ���      �       R�      Y       ��                 �      �       3�                   �      �       u#�      �       u#                                !       R!      k       Sk      �       ��~�#��      �       ��~�#�             ��~�#�                     �             u#�'�      %       }#�'��      �       u#�'�                    �      %       P%      V       ��~                           <      k       0�k      �       V�      �       v��      �       V�      �       V�      �       v�             V                 �             0�                   z      �       P�             P                              #       U#      Z        s "��      �        s "�              s "�                  �      �       P                 d      z       t                    s      z       Qz      z      
 p q "#���                  s      z       q ?&�z      z       P                      P      r       Ur      �       S�             �U�                      P      d       Td             ]             �T�                            i      r       0�r      �       V�      �       v��      �       V�      �       0��      �       \�      �       |��      �       \                          P      �       U�      �       V�             �U�             U      4       V                          P      �       T�      �       \�             �T�             T      4       \                            P      �       Q�      �       Z�             �Q�             Q      %       Z%      4       �Q�                    v      �       0�      4       0�                  �      �       Q                     e      �       0��      �       S      4       0�                         p      &       0�&      '       P'      4       0�4      5       P5      ;       0�;      I       P                       �      �       Q�      �       q��      �       q��      �       R�      �       r��             R5      I       R                    �             Z5      I       Z                      �      �       P�      �       r �             P5      I       P                        �      �       X�             Y             Q5      ;       X;      I       Y                          �             Y             Q             Y5      ;       Y;      >       Q                                �       �        U�       0!       S0!      2!       �U�2!      B!       SB!      D!       �U�D!      ^!       S^!      `!       �U�`!      t!       S                    �       �        T�       t!       �T�                                 �       �        u8��       �        U�       0!       s8�0!      2!       �U#8�2!      B!       s8�B!      D!       �U#8�D!      ^!       s8�^!      `!       �U#8�`!      t!       s8�                 �       
!       V                               �       
!       0�
!      !       P!      1!       V1!      2!       P2!      D!       0�D!      _!       V_!      `!       P`!      t!       V                       !!      0!       s8�0!      2!       �U#8�D!      ^!       s8�^!      `!       �U#8�                       !!      0!       s8�0!      2!       �U#8�D!      ^!       s8�^!      `!       �U#8�                       !!      2!       �P�D!      Q!       �P�Q!      U!       TU!      `!       �P�                 D!      U!       s8                            �             U      �       S�      �       �U��      �       S�      �       �U��      �        S                          �      �       T�             V      +       v  ��      �       V�      h        V                              �      	       Q	      �       ^�      �       �Q��      �       ^�      �       �Q��      �       Q�      �        ^                          �      A       RA      �       �R��      �       R�      4        ��4       �        �R�                  �       �        P                      �      �       _�      �       _�      �        _                              �       \�      �       \               P       �        \                                 �      +       0�+      9       P<      V       P\      i       P�      �       0��      4        0�4       A        PY       h        P�       �        P                 �      �       s��v �����                        `      �       U�      �       S�      �       �U��      p       S                            `      �       T�      �       ^�      �       �T��      >       ^>      h       Th      p       ^                                `      �       Q�      >       �Q�>      c       Qc      {       Z{      �       ���      �       �Q��      �       ���      p       �Q�                            `      �       R�      �       w �      �       ���      >       w >      p       Rp      p       w                        �      �       \�      X       \>      �       \�      p       \                                 �      �       0��      �       0��      �       P�      >       ��>      �       0��      �       ���      �       0��      �       ���      p       0�                               �      �       0��      $       0�$      (       P(      E       _>      �       0��      �       0��      �       _�      p       0�                   �      �       } ����s("��      �       } ����s("�                            =      Z       1�Z      �       ]�             }�             ]�      �       ]�      �       1��      �       1�                         :      :       s01�:      Z       0�Z      �       T�             T�      �       T�      �       s01��      �       0��      �       0�                          .      Z       0�Z      �       R�      �       ���             R�      �       R�      �       0��      �       0�                      :      Z       Y�      �       Y�      �       Y                         Z      �       V�      �       V�             T�      �       V�      �       T                     E      �       S�      �       S�      �       S�      p       S                     M      �       _�      �       _�      �       _�      p       _                     M      �       \�      �       \�      �       \�      p       \                        w      {       P{      �       ���      �       ���      �       ���      p       ��                            w      {      	 p �r �{      �       ����v ��      �       }����������             ����v �      �       }����������      �       }����������      p       }���������                                   #      a       P�      �       P�             p~�      $       P$      ,       p r "�,      0       p r "#�0      :       p r "�:      N       PN      ^       p}�^      p       P                          '      a       Ta      m       � v "��      $       T$      :       p v "�:      p       T                                        #      T       QT      \       qx�\      a       Q�      �       Q�             qx�      $       Q$      ,       r 3$q "�,      0      
 r 3$q "#�0      :      
 r3$q "#�:      R       QR      f       qx�f      p       Q                               #       U#      P       SP      `       �U�`      a       U                       '       P                        _       V                                �!      �!       U�!      	"       S	"      "       �U�"      ="       S="      G"       �U�G"      #       S#      #       �U�#      %#       S                                  �!      �!       T�!      "       ]"      "       �T�"      B"       ]B"      G"       �T�G"      T"       UT"      #       ]#      #       �T�#      %#       ]                    �!      �!       Q�!      %#       �Q�                    �!      �!       R�!      %#       �R�                        �!      
"       V"      >"       VG"      #       V#      %#       V                           �!       "       P "      "       ^"       "       ^U"      a"       p 
���a"      #       ^#      %#       ^                    x"      �"       P�"      �"       s                         �"      �"       T�"      �"       s�#����p ��"      �"       P�"      �"       T#      #       T                    P      d       Ud      e       �U�                            p5      �5       U�5      �6       ]�6      �6       �U��6      �8       ]�8      �8       �U��8      �8       ]                    p5      �5       T�5      �8       �T�                              p5      �5       Q�5      �5       P�5      �6       w �6      �6       ���6      �8       w �8      �8       ���8      �8       w                                                          |5      �5       T�5      �5       \�5      �5       rx
6      t6       \�6      �6       \�6      7       |�7      e7       \e7      �7       Q�7      �7       \�7      �7       |��7      �7       q #��7      8       \8      8       |�8      8       q #�8      8       \8      (8       |�(8      78       P78      X8       |�X8      |8       p�|8      �8       |��8      �8       p~��8      �8       p��8      �8       \�8      �8       |��8      �8      	 }(8#�                      |5      �6       0��6      67       0�67      ?7       P?7      �8       0�                                        �5      �5       P6      E6       P\7      u7       P�7      �7       P8      (8       P78      F8       p 4%��F8      I8       p ?��I8      X8      
 |�?��X8      d8       }(8#�?��d8      u8       q 4%��u8      x8       q ?��x8      |8      
 p�?��|8      �8      
 |�?���8      �8       }(8#�?��                           <6      E6       PE6      I6       }4�p !�I6      t6       P�6      �6       P?7      L7       P\7      u7       P{7      �7       P                               96      t6      
 }(} 8��6      �6      
 }(} 8�7      7      
 }(} 8�,7      57      
 }(} 8�?7      V7      
 }(} 8�\7      �7      
 }(} 8��7      �7      
 }(} 8��7      �7       R                             E6      _6      
  �F     �_6      t6       S�6      �6       S7      &7       S,7      ?7       S?7      L7      
  �F     ��7      8       S                           �6      �6       P7      ,7       PW7      \7       P�7      �7       0��7      8       _�8      �8       P                        �6      ?7       VD7      \7       V�7      8       V�8      �8       V                   �7      �7       s�����p "��7      �7       q ����p "�                   �7      �7       } �7      8       ^                 �6      �6       }                  �6      �6       3�                 �6      �6       ]                 7      7       }                  7      7       ]                      �;      �;       U�;      �;       �U��;      �;       U                      �;      �;       S�;      �;       S�;      �;       u8                   �;      �;       u �;      �;       u #��;      �;       u                    �;      �;       0��;      �;       3�                          @=      �=       U�=      s?       ]s?      �?       �U��?      Q@       ]Q@      ^@       U                      D=      �=       PQ@      ]@       P]@      ^@       u8                   {=      w?       _�?      Q@       _                      �=      �=       S�=      w?       ���?      Q@       ��                  �=      �=       P                   �=      �=       Pa?      a?       ��a?      x?       P                   �=      K>       V�?      Q@       V                  �=      a?       ]�?      Q@       ]                  �=      a?       _�?      Q@       _                          @>      K>       PK>      �>       ���>      �>       P�>      �>       ^C?      Q?       ^                 9>      K>       S                   @>      C?       0�C?      Q?       1�                       o>      �>       1��>      �>       p ���#��>      �>      	 ~ �����>      �>       ~ ���#�                        >      />       [/>      K>       v 2$v "��?      �?       [�?      Q@       ��                	   �=      w?       ���?      Q@       ��                    �=      />       U�?      �?       U                    �=      K>       \�?      Q@       \                    >      2>       S�?      Q@       S                      e>      �>       V�>      �>       v|��>      Q?       V                      o>      �>       Q�>      �>       w �>      Q?       Q                  �?      Q@       ^                    �?      �?       Z�?      Q@       w                   @      Q@       P                   @      *@       } *@      Q@       Q                      �;      �;       U�;      �;       �U��;      �;       U                      �;      �;       S�;      �;       S�;      �;       u8                   �;      �;       u �;      �;       u #��;      �;       u                  �;      �;       q��                 �;      �;       0�                       <      &<       U&<      Y<       SY<      ^<       �U�                  <      <       u8                  <      <       V<      6<       v�6<      Y<       v�                 <      W<       ��W<      Y<       0�                      `<      �<       U�<      �<       S�<      �<       �U�                 `<      y<       u8                `<      �<       ��                    �<      �<       P�<      �<       R                          �<      �<       U�<      )=       S)=      -=       �U�-=      1=       S1=      :=       �U�                 �<      �<       u8                        �<      �<       V�<      �<       u �<      �<       V�<      *=       v�-=      7=       v�                   �<      &=       ��&=      -=       0�-=      :=       ��                         =      =       P=      (=       P(=      ,=       |�-=      6=       P                      �4      �4       U�4      5       V5      5       �U�                 �4      �4       u8                 �4      �4       u8#��                  �4      �4       S�4      �4       s��4      �4       s��4      5       s�                 �4      5       ��5      5       0�                 �4      �4       S�4      �4       s��4      �4       s��4      5       s�                    �4      �4       U�4      �4       V                 �4      �4       s��4      �4       s��4      5       s�                 �4      �4       V                 �4      �4       s��4      5       s�                 �4      �4       V                 �4      5       s�                 �4      5       V                        `@      �@       U�@      �A       V�A      �A       �U��A      �C       V                 `@      b@       u8                 `@      b@       u8#@�                 `@      b@       u8#p�                 `@      b@       u8#h�                              w@      �@       ^�@      BA       ~  "#�BA      HA       ~  "�HA      �A       ~  "#��A      �A       ~  "��A      B       ~  "#�B      AC       ~  "�AC      �C       ~  "#�                     �@      �@      
 ���������@      �A       \�A      �C       \                         �@      �@      
 �       ��@      �A       S�A      �B       S�B      C       s �C      �C       S                 �@      �@       0�                                BB      ZB       PZB      cB       � r "�qB      �B       P�B      �B       � r "�C      C       PC      $C       � r "�)C      3C       P3C      <C       � r "�                      BB      cB       T�B      �B       TC      AC       T                                BB      \B       Q\B      cB       t 1&��B      �B       Q�B      �B       t 1&�C      C       QC      )C       t 1&�)C      5C       Q5C      AC       t 1&�                             �@      BA       ~  "�BA      HA       ~  "8�LA      �A       ~  "��A      �A       ~  "8��A      B       ~  "�B      AC       ~  "8�AC      �C       ~  "�                        �@      "A       VLA      �A       V�A      B       VAC      �C       V                          �@      �@       P�@      !A       U`A      yA       PyA      �A       UAC      �C       P                                  �@      �@       5��@      �@       6��@      �@       7��@      �@       8��@      A       9�AC      WC       5�WC      uC       6�uC      �C       7��C      �C       8�                                      `	      �	       U�	       
       �U� 
      &       U&      ;       �U�;      �       U�      �       �U��      �       U�      �       �U��             U              �U�       ;       U                    `	      �	       T�	      ;       �T�                                        `	      �	       Q�	       
       �Q� 
      �
       Q�
      �
       �Q��
             Q      ;       �Q�;      t       Qt      �       �Q��      �       Q�              �Q�       +       Q+      ;       �Q�                        `	      �	       R�	      �	       V�	       
       �R� 
      ;       V                           `	      �	       T 
      
       T;      �       T�      �       T�      �       T       ;       T                                �	      �	       Z 
             Z1      f       Z�      .       Z;      �       Z�      �       Z�             Z       ;       Z                             �	      �	       R�	      �	       R 
      m
       R�
      -       R1      �       R�      �       R�      �       _;      M       _                                �	      �	       X�	      �	       p ��
      �
       X6      ;       P�      �       P�      �       P�      �       X              P                                              �	      �	       X 
      
       X"
      ,
       X7
      �
       X�
      �
       X�
      �
       P�
      �
       X�
      �       X�      .       X;      S       XX      �       X�      �       X�      �       X�      �       X�      �       P       6       X6      ;       P                                     a
      m
       0�t
      �
       ]�
      �
       [�
      �
       ^�
      �
       [      H       [O      `       [�      �       [�      �       { ��      �       [;      M       [X      �       ]�      ;       ]                       `	      �	       0��	      �	       S 
      
       S
      ;       S                             `	      �	       0� 
      m
       0��
             0�      ^       ^`      �       0��      �       ^;      M       ^                        �	      �	       P 
      p
       P�
      �       P;      M       P                   "
      3
       y�3
      <
       Y                                           M
      �
       \�
      �
       Y�
      `       \f      �       \�      .       Y;      M       \X      X       \X      t       | } �t      �       \�      �       | ��      �       Y�      �       Y�      �       \�      �       9�       )       | } �6      ;       \                  �
      �
       P                  �
      �
       Q                  �	      �	       U�	      �	       U                  �	      �	       T�	      �	       T                  �	      �	       T�	      �	       T                              U                              T                              T                 n      x       U                 n      x       T                 n      x       T                 �      �       T�      I       t�                                  �      �       Q�      �       t ����      �       Q�             t ���             Q      (       t ���(      ;       Q;      B       q��B      I       t ���                                 �      �       0��      �       P�      �       0��      �       P�             0�      '       0�'      (       P(      H       0�H      I       P                 �      �       U                 �      �       t�                   �      �       t��      �       Q                 �             U                 �             t�                 �      �       t�                       (       U                       (       t�                                t�             Q                 (      I       U                 (      I       t�                 (      5       t�                        �#      B$       UB$      S$       SS$      ]$       �U�]$      �.       S                                          �#      B$       TB$      H$       \H$      ]$       �T�]$      �$       T�$      �)       \�)      *       T*      B+       \B+      !-       �T�!-      =-       \=-      [-       �T�[-      �-       \�-      �-       �T��-      �.       \                                �#      B$       QB$      ]$       ��i]$      j$       Qj$      �)       ��i�)      *       Q*      *       ��i*      *       �Q�*      *       P*      �.       ��i                                        �#      B$       RB$      H$       V]$      �$       R�$      c)       Vc)      �)       �R3!�R�R
  $0.( ��)      *       R*      C-       VC-      [-       �R3!�R�R
  $0.( �[-      -.       V-.      q.       �R3!�R�R
  $0.( �q.      �.       V�.      �.       �R3!�R�R
  $0.( �                                                   &      &       P&      /&       _/&      P&       PP&      m&       _m&      �&       P�&      �&       _�&      �&       0�%'      T'       P�(      �(       P�(      �)       _*      $*       P$*      H*       _H*      R*       P�-      .       _.      .       0�-.      q.       _q.      �.       P�.      �.       _                        $      H$       ^]$      �+       ^!-      =-       ^[-      �.       ^                          �%      �%       R�%      �'       ��i*      *       ��i*      R*       0�R*      -.       ��iq.      �.       ��i                                   $      H$       0�]$      Y%       0�Y%      �'       ��i�'      |(       0�|(      �(       1��(      *       0�*      *       ��i*      R*       1�R*      -.       ��i-.      q.       0�q.      �.       ��i�.      �.       0�                        $      H$       ]]$      �+       ]!-      =-       ][-      �.       ]                       $      B$       ~�]$      �$       ~��(      �(       ~��)      *       ~�                       $      B$       ~�#P]$      �$       ~�#P�(      �(       ~�#P�)      *       ~�#P                                   M%      T%       P��T%      Y%       }���Y%      �'      
 ��i���h�-(      2(       T��2(      H(       T�P�H(      Q(       ��i�P�Q(      �(      
 ��i���h�*      V-      
 ��i���h�[-      -.      
 ��i���h�q.      �.      
 ��i���h�                     �$      �$       | �(      �(       Q�(      �(       |                      �$      �$       | #��(      �(       q��(      �(       | #�                     �$      �$       | #��(      �(       q��(      �(       | #�                      �)      �)       1�-.      X.       0��.      �.       0�                  �'      �(       _                    (      Q(       XQ(      �(       ��h                  �'      �'       P�'      �'       q�                 �-      .       }�
�                  q'      �'       P                   R*      �-       s0�.      -.       s0�                      �*      �*       0�[-      �-       1�.      -.       0�                  �,      �,      	 q 0$0&�                   �+      B,       s���,      !-       s��                         �+       ,       s��,      �,       s��,      �,       P�,      -       pp�-      !-       P                   �+       ,       s��,      �,       s�                   �+       ,       s��,      �,       s�                 ,      ,       s�                    ,      ,       R,      ,      
 p r "#���                  ,      ,       r ?&�,      ,       P                !,      0,       s�                    ),      0,       T0,      0,      
 p t "#���                  ),      0,       t ?&�0,      0,       P                  �,      �,       p �,      �,       pp                   �,      �,       Q�,      �,      
 q x "#���                  �,      �,       q ?&��,      �,       X                   �,      -       Q-      -      
 q x "#���                  �,      -       q ?&�-      -       X                `+      o+       ��i                `+      o+       s�                    m+      o+       Po+      o+      
 p q "#���                  m+      o+       p ?&�o+      o+       Q                �+      �+       ��i                �+      �+       s�                    �+      �+       P�+      �+      
 p q "#���                  �+      �+       p ?&��+      �+       Q                   5$      B$       }�
��)      *       }�
�                      5$      B$       Q�)      *       Q*      *       ��i*      *       �Q�                    5$      B$       0��)      *       0�*      *       P                    �      �       U�      �       �U�                 �      �       u�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                 �      �       u�                    p      y       Uy      z       �U�                    p      y       Ty      z       �T�                 p      y       u�                    `      i       Ui      j       �U�                    `      i       Ti      j       �T�                    `      i       Qi      j       �Q�                 `      i       u�                    P      Y       UY      Z       �U�                    P      Y       TY      Z       �T�                    P      Y       QY      Z       �Q�                 P      Y       u�                    @      I       UI      J       �U�                    @      I       TI      J       �T�                 @      I       u�                    0      9       U9      :       �U�                    0      9       T9      :       �T�                    0      9       Q9      :       �Q�                 0      9       u�                           )       U)      *       �U�                           )       T)      *       �T�                           )       Q)      *       �Q�                        )       u�                                 U             �U�                                 T             �T�                                 Q             �Q�                              u�                           	       U	      
       �U�                           	       T	      
       �T�                           	       Q	      
       �Q�                        	       u�                      �      �       R�      �       u�	�      �       R                       �      �       t ����1$r�
"�
����      �       t ����1$r "�
����      �       t 1$r "�
����      �       t 1$u�	#�
"�
���                   �      �       r���      �       u�	#��                  �      �       P                 �      �       p��                    �      �       U�      �       �U�                          �             T      F       ]F      S       �T�S      b       Tb      �       ]                          �             Q      F       \F      S       �Q�S      i       Qi      �       \                          �             R      F       VF      S       �R�S      i       Ri      �       V                     �      H       0�S      _       6�_      �       0�                    �      M       SS      �       S                   �      F       s��S      �       s��                              p      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U��      �       U                              p      �       T�      �       V�      �       T�      �       �T��      �       V�      �       �T��      �       T                             p      �       U�      �       S�      �       U�      �       �U��      �       S�      �       �U��      �       U                   p      �       u �      �       u                    p      �      	 u #�#�      �      	 u #�#                  �      �       P                  �      �       P                            �      	       U	      	       �U�	      3	       U3	      \	       S\	      ^	       U^	      _	       �U�                    �      	       V	      ]	       V                     �      	       u�	      3	       u�3	      7	       s�                 *	      7	       p                  8	      F	       P                  G	      O	       P                        �              U              �U�             U      �       �U�                          �              T              V             �T�      )       T)      �       V                    �             \      �       \                       �       |��                           1       0�1      5       P5      �       S                                u�      -       U                  N      _       P                    `      u       Pu      �       }y�                    v      �       P�      �       P                    {      �       ]�      �       ]                        �      �       U�      �       �U��             U      �       �U�                        �      �       T�      �       S�      �       �T��      �       S                    �      �       \�      �       \                 �      �       |��                     �             0�             P      �       V                   �             u�             U                                @      ^       U^      {       V{      �       �U��             V      1       �U�1      D       VD      I       UI      J       �U�                            @      s       Ts      +       S+      1       �T�1      C       SC      I       TI      J       �T�                    W      0       ]1      H       ]                   W      0       }�
�1      H       }�
�                   {      �       P�      �       V                    �      �       T�      �       P                        �      �       U�      �       p 1$q "�      �       | ����1$q "�      �       U                    �      �       0��      �       \                   �      �       u�      �       U                  �             P                               P                 i      w       v�                    {      �       P�      �       V                 �      �       ]                  �      �       U                                 /      t/       Ut/      �/       \�/      �/       �U��/      �/       U�/      &0       \&0      -0       �U�-0      p0       Up0      �0       \                               /      */       T*/      t/       St/      �/       �T��/      �/       S�/      -0       �T�-0      p0       Sp0      �0       �T�                             /      t/       Qt/      �/       �Q��/      �/       Q�/      -0       �Q�-0      p0       Qp0      �0       �Q�                               /      t/       Rt/      �/       �R��/      �/       R�/      �/       R�/      (0       ]-0      p0       Rp0      �0       �R�                               /      t/       Xt/      �/       �X��/      �/       X�/      �/       V�/      -0       �X�-0      p0       Xp0      �0       �X�                             _/      �/       0��/      �/       1��/      �/       0��/      0       1�0      -0       0�W0      �0       0��0      �0       1�                          /      �/       0��/      �/       P�/      0       0�0      -0       P-0      �0       0�                          /      j/       _j/      t/       u��/      ,0       _-0      f0       _f0      p0       u�                       &/      t/       Ut/      �/       \-0      p0       Up0      �0       \                              �.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U                              �.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T                              �.      �.       Q�.      �.       �Q��.      �.       Q�.      �.       �Q��.      �.       Q�.      �.       �Q��.      �.       Q                              �.      �.       R�.      �.       �R��.      �.       R�.      �.       �R��.      �.       R�.      �.       �R3!��.      �.       R                             �.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U�.      �.       �U��.      �.       U                             �.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T�.      �.       �T��.      �.       T                      0      T       UT      ^       �U�^      c       U                      0      T       TT      ^       �T�^      c       T                      0      T       QT      ^       �Q�^      c       Q                        0      T       RT      ]       S]      ^       �R�^      c       R                     0      T       UT      ^       �U�^      c       U                      7      T       P^      b       Pb      c       u�                          #       U#      $       �U�                          #       T#      $       �T�                       #       u                        #       u #�	                       #      
 u #�	#�&                    �              U             �U�                    �              T             �T�                 �              u                  �              u #�	                 �             
 u #�	#�&                             2       U2      G       SG      H       �U�                        !       u                         !       u #�                        �       �        U�       �        T�       �        �U��       �        T                    �       �        T�       �        �T�                    �       �        Y�       �        Y                   �       �        y��       �        y�                          �       �        P�       �        P�       �        y�	�       �        P�       �        y�	                         �       �        p�
��       �        p�
��       �        y�	#�
��       �        p�
��       �        y�	#�
�                      �       �        Q�       �        p�&�       �        Q                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  �      �       U                 �      �       u�
�                     �      �       t ����1$u�
"�
����      �       t 1$u�
"�
����      �       �T����1$u�
"�
���                     P       t        0�t       x        Px       �        0��       �        P                  R       i        Q                     b       i        q�i       x        Qx       |        q��       �        Q                    0       D        TD       E        �T�                 0       D        0�                                 u                                  u #�	                                 u #�	#��                      `      n       Un      o       �U�o      q       U                    g      n       Po      q       P                      p      �       U�      �       �U��      �       U                            p      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T�                    �      �       T�      �       �T�                  �      �       U                 �      �       U                  �      �       T                 �             U                 �      �       u�	                          *       S,      3       S                          +       P,      2       P                      `      o       Qo      �       V�      �       �Q�                      y      �       P�      �       v �      �       �Q                 `      x       U                     `      �       0��      �       Q�      �       Q                          �       0��      �       R                        0#      P#       UP#      o#       �U�o#      w#       Uw#      �#       �U�                        0#      W#       TW#      o#       �T�o#      �#       T�#      �#       �T�                            0#      V#       QV#      m#       Sm#      o#       �Q�o#      �#       Q�#      �#       S�#      �#       �Q�                            0#      W#       RW#      n#       Vn#      o#       �R�o#      �#       R�#      �#       V�#      �#       �R�                  X#      o#       P                    o#      �#       R�#      �#       V                    o#      �#       Q�#      �#       S                    o#      �#       T�#      �#       �T�                    o#      w#       Uw#      �#       �U�                     o#      w#       u�	w#      ~#       U~#      �#       u�u�                        �#      �#       U�#      �#       �U��#      �#       U�#      �#       �U�                        �#      �#       T�#      �#       �T��#      �#       T�#      �#       �T�                        �#      �#       Q�#      �#       �Q��#      �#       Q�#      �#       �Q�                    �#      �#       Q�#      �#       �Q�                    �#      �#       T�#      �#       �T�                    �#      �#       U�#      �#       �U�                  �#      �#       P                 �#      �#       p�
�                   �#      �#       T�#      �#       �T�                 �#      �#       p�
                      �0      �0       U�0      61       V61      71       �U�                      �0      �0       T�0      51       S51      71       �T�                      �3      V4       UV4      W4       �U�W4      u4       U                          �3      �3       Q�3      M4       YM4      V4       QV4      W4       �Q�W4      u4       Y                          �3      �3       P�3      %4       R%4      24       P24      M4       RW4      u4       R                     5      d5       Ud5      n5       �U�                          �C      �C       U�C      �C       \�C      �C       �U��C      D       \D      	D       �U�                            �C      �C       T�C      �C       V�C      �C       �T��C      D       VD      D       TD      	D       �T�                        �C      �C       P�C      �C       S�C      �C       P�C      �C       S                      �C      D       VD      D       TD      	D       �T�                    �C      D       \D      	D       �U�                  �C      �C       U                  �C      D       P                                D      ,D       U,D      iD       ViD      nD       �U�nD      �D       V�D      �D       �U��D      �D       V�D      �D       U�D      �D       �U�                            D      GD       TGD      ID       SID      nD       �T�nD      |D       T|D      �D       S�D      �D       �T�                                  D      MD       QMD      mD       ]mD      nD       �Q�nD      �D       Q�D      �D       ]�D      �D       �Q��D      �D       ]�D      �D       Q�D      �D       �Q�                                  D      MD       RMD      kD       \kD      nD       �R�nD      �D       R�D      �D       \�D      �D       �R��D      �D       \�D      �D       R�D      �D       �R�                      ,D      MD       UnD      �D       U�D      �D       v�	                  ND      `D       P                   <D      ID       s ����1$u�
"ID      MD       �T����1$u�
"                          nD      �D       R�D      �D       \�D      �D       \�D      �D       R�D      �D       �R�                          nD      �D       Q�D      �D       ]�D      �D       ]�D      �D       Q�D      �D       �Q�                      nD      �D       S�D      �D       S�D      �D       T                        nD      �D       V�D      �D       V�D      �D       U�D      �D       �U�                 nD      �D       v�#                  �D      �D       P                    �D      �D       P�D      �D       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u��                                 P             u�                 p       �        U                        �      &       U&      �       S�      �       �U��      �       U                       �      &       U&      �       S�      �       �U��      �       U                        �       ]                           &       u��&      �       s���      �       �U#��                           &       u��&      �       s���      �       �U#��                            &       0�&      p       \p      t       |�                  :      }       V                      �      �       U�             S             �U�                    �      �       T�             �T�                  �      �       P                                   U      h       Sh      i       �U�                                  U      h       Sh      i       �U�                         S       0�S      c       P                    #      %       P%      R       X                    -      P       QP      R       s                    -      P       q
Pq�"�P      R       r 
Ps #�"�                   -      P       q
Pq�"�P      R       r 
Ps #�"�                      �      �       U�             S             �U�                      �      �       P�      �       u�      �       s                  �             V                  �             P                  	             P                              /        U/       B        �U�B       I        U                                        T       1        Q1       B        �T�B       I        T                  ,       A        S                        p      �       U�      �       \�      �       �U��      z       \                    p      �       T�      z       �T�                       p      �       u���      �       |���      �       �U#���      z       |��                    �      �       V�      z       V                    �      �       ]�      z       ]                      �      �       P�      �       S�      z       S                       1       0�                   1      F       q|�F      z       q�}�                      �      $       U$      K       \K      X       �U�X      i       \                      �      !       T!      K       VK      X       �T�X      i       V                        �       s  $ &
P} "�                     �      $       U$      K       \K      X       �U�X      i       \                  5      b       p �                       �       s  $ &
P} "#��                       �       s  $ &
P} "#��                  '      5       P                               �       U�      �       S�      �       �U��      �       S                                     �       T�      �
       ]�
      �       �T��             T      �       ]�      �       �T��      �       ]                                     ]       Q]      @	       ^@	      �       �Q��             ^      �       �Q��      �       ^�      �       �Q�                                   �       R�      �       V�      �       R�      '       V�      �       V�      �       V                              �       U�      �       S�      �       �U��      �       S                                  �      �       P�      	       _	      .	       P.	      �       _      u       _u      �       0��      �       P�      �       _�      �       0��      �       _                    ;      2
       \�      �       \                              �      �       Q�      �       u�D	      K	       PK	      �	       s��	      �       ��g      �       ��g�      �       ��g                          O	      W	       PW	      �	       s��	      �       ��g      �       ��g�      �       ��g                       ;      �       |��      �       ��g�             |�      �       ��g                       �	      �	       ��g�^��	      �       �^�      �       �^��      �       �^�                       ;      �       0��      �	       1��	      �       0��      �       0��      �       1��      �       0�                  '      �       V                   �	      �       s0��      �       s0�                  �
            	 q 0$0&�                   �
      �       ��h�      �       ��h                         �
             ��h#             P      O       pp�O      T       P�      �       ��h#                   �
             s��      �       s�                   �
             s��      �       s�                               p              pp                                Q            
 q y "#���                               q ?&�             Y                   5      <       Q<      <      
 q y "#���                  5      <       q ?&�<      <       Y                T      c       s�                    \      c       Uc      c      
 p u "#���                  \      c       u ?&�c      c       P                u      �       s�                    }      �       T�      �      
 p t "#���                  }      �       t ?&��      �       P                P
      _
       ��g                P
      _
       s�                    ]
      _
       P_
      _
      
 p q "#���                  ]
      _
       p ?&�_
      _
       Q                u
      �
       ��g                u
      �
       s�                    ~
      �
       P�
      �
      
 p q "#���                  ~
      �
       p ?&��
      �
       Q                                   }       U}             V      (       �U�(      ;       V;      N       UN              V                               �       T�      ;       ��k;      a       Ta              ��k                          8      .       _�      �       _(      ]       _]      k       U�              _                         8      .       ���      �       ��(      ]       ��]      k       u���              ��                            �      �       P�      �       P�      �       Q�      �       x� �             P      &       P�      �       P              Q                    �      F       S�      ;       S�             S                      J      �       X;      r       Xr      �       ��k                                   R      �       0��             ]      3       0�3      �       ]�             0�      5       P5      ;       ];      �       0��      �       P�      �       ]�              0�                        V      ]       P]             w       (       ��k(              w                                   V      �       0��      �       ��k(      5       0�5      �       ��k�             0�      
       P
      ;       ��k;      �       0��             0�              0�                          b      i       Pi      �       ��      ;       ��k;      r       �r              ��k                           b      .       0�.      �       \�      �       0��      !       \(      �       0��      �       1��              0�                    m      %       ^(              ^                   �      �       T�      �       T                  �      �       ��  �      �       ��                       �      �       0��      �       S�      �       0�                   �      �       P�      �       P                    Z      �       S             S                         U       RU      �       ��k                  L      �       \�             0�                   �      �       T              T                  �      �       ��                ��                       �      �       0��      �       S              0�                    �      �       Q�      �       q��      �       Q              Q                     �             Q             ��      �       Q                   �             ��  �             ��                      �             0�             R�             0�                    �             P             p�             P�      �       P                      L       �                      L       ��                          &       0�&      L       \                        4       P4      <       p�<      L       P                      W      .       S�      �       S5      v       S                          !       P!      F      
 s 4$�"�                      �      �       P�      �       ��k�      �       P                 �      �       U                    �      �       S�      �       S                    �      �       P�      �       P                        p      �       U�      �       S�      �       �U��      �       U                       p      �       U�      �       S�      �       �U��      �       U                      ~      �       U�      �       S�      �       �U�                  �      �       P                                    �      �       U�      �       S�             �U�      �       S�      �       �U��      �       S�      E       �U�E      �       S�      �       �U��              S       �%       �U�                                                          �      �       T�      �       ]�             �T�      �       ]�      �       �T��      �       ]�      &       ��{&      8       �T�8      �       ��{�      �       �T��             ��{      E       �T�E      T       TT      �       ]�      �       ��{�      �       �T��              ]       &        �T�&       5        ��{5       �        �T��       �        ��{�       �%       �T�                        �      �       Q�      E       ��{E      \       Q\      �%       ��{                        �      �       R�      E       �R�E      \       R\      �%       �R�                        �      �       X�      E       �X�E      \       X\      �%       �X�                                                         �      �       T�      �       ]�             �T�      �       ]�      �       �T��      �       ]�      &       ��{&      8       �T�8      �       ��{�      �       �T��             ��{      E       �T�E      T       TT      �       ]�      �       ��{�      �       �T��              ]       &        �T�&       5        ��{5       �        �T��       �        ��{�       �%       �T�                        �      �       P             P      _       X      +       6�                         �      �       t�E      T       t�T      \       }�]      {       P�              P                    �      �       t�u      {       }��      �       P                                �       S�      �       �U��      �       S�      E       �U��      �       �U�       �%       �U�                            E       �R��      �       �R�       �%       �R�                            E       �X��      �       �X�       �%       �X�                            E       ��{�      �       ��{       �%       ��{                                                    �       ]�      �       �T��      �       ]�      &       ��{&      8       �T�8      �       ��{�      �       �T��             ��{      E       �T��      �       ��{�      �       �T�       &        �T�&       5        ��{5       �        �T��       �        ��{�       �%       �T�                            �      �       X�      �       X      E       X�      &       X&      +       ��{�      �       X                                 �       ��{�      �       ��{�             ��{�      �       ��{+      �       ��{       �%       ��{                                                 �       ]�      �       �T��      �       ]�      &       ��{&      8       �T�8      �       ��{�             ��{             �T��      �       ��{+      �       �T�       &        �T�&       5        ��{5       �        �T��       �        ��{�       �%       �T�                               V      _       U_      E       ^�      �       ^�      �       U�      �       ^       �        ^�       !       U!      �%       ^                                   V      _       R_      �       ��{�      �       ��{�             ��{�      �       ��{+      �       ��{       �!       ��{$      M$       ��{W$      i$       ��{(%      ,%       ��{                 "      P       0�                                             V      �       }���      �       �T#���      �       }���      &       ��{#��&      8       �T#��8      �       ��{#���      �       �T#���             ��{#��      E       �T#���      �       ��{#���      �       �T#��       &        �T#��&       5        ��{#��5       �        �T#���       �        ��{#���       �%       �T#��                      "      �       U	!      !       U!      h!      	 }��                   "      �       x { " $ &�	!      E!       x { " $ &�                                             V      �       ]�      �       �T��      �       ]�      &       ��{&      8       �T�8      �       ��{�      �       �T��             ��{      E       �T��      �       ��{�      �       �T�       &        �T�&       5        ��{5       �        �T��       �        ��{�       �%       �T�                	V      V       U                   V      ^       Q^      _       }�                           V      _       R_      �       ��{�      �       ��{8      �       ��{�             ��{�      �       ��{&       5        ��{�       �        ��{                           V      �       V�      �       U�      �       V8      �       V�             V�      �       V&       5        V�       �        V                           V      _       U_      �       ^�      �       ^8      �       ^�             ^�      �       ^&       5        ^�       �        ^                                  �      �       P�      �       2��      �       0�"      7       P�      �       P�             P�      �       0��      �       P�      �       P�      �       3�0       5        3��       �        0�                            }      �       P�      �       ��{�      �       ��{8      �       ��{�             ��{�      �       ��{&       5        ��{�       �        ��{                                  �      �       ]�      �       P�      �       w 8      q       ]q      v       Pv      �       ]�      �       }�~��      �       ]�             w �      �       w &       +        ]�       �        w                           �      �       S�             ��}      �      	 w ��{��            	 w ��{��      �      	 w ��{��       �       	 w ��{�                        I      n       _�      �       Q�      �       _�      �       ~                                <      �       YD      l       \l      n       ��{n      �       |	�8      �       Y�             |	��      �       }�&       5        Y�       �        |	�                                       X      n       ��{n      �       X�      �       S�      �       X�             X                      .      �       S�      �       _�      �       S�             S�       �        S                        �      �       
	��             S      �       _8      �       _�      �       
 �                         �      �       0��      �       w 8      q       w v      �       w �      �       9�&       5        w                             �      �       ��}��      <       \<      P       Pc      �       Pv      �       P�      �       ��}��      �       \&       0        P                    
              p �             _                 �       �        P                 �      �       ^                 �      �       ^                 �      �       ^                 �      �       ��|                        &       ��}                        &       \                                        �       ^+      �       ^�      �       U�      �       ^�       �        ^�       !       U!      	!       ^$      D$       ^W$      i$       ^                        &       ]                                         8       ^+      �       ^�      �       U�      �       ^�      �       ^       &        ^5       �        ^�       �        ^�       !       U!      �%       ^                                       "      [       \d             \�      �       \�      �       V+      =       \=      {       V{             v�      �       P�      �       v��      �       V�       �        v��       	!       v�$      D$       v�W$      i$       v�                               "      &       S&      �       w #�+      �       w #�w      �       w #��       �        w #��       	!       w #�$      D$       w #�W$      i$       w #�                    T      �       P4      I       P                            �      �       Q�      �       ��{�       �        ��{�       	!       ��{$      D$       ��{W$      i$       ��{                                    �      A       ]A      �       _�      �       T�      �       _�      �       ]�       �        _�       !       T!      	!       _$      D$       _W$      i$       _                      �      <       S�      �       S�      �       }                                     1�      )       P/      4       P                             A      �       _�      �       T�      �       _�       �        _�       !       T!      	!       _$      D$       _W$      W$       _                             A      �       ^�      �       U�      �       ^�       �        ^�       !       U!      	!       ^$      D$       ^W$      W$       ^                       A      �       ]�       �        ]�       	!       ]$      D$       ]W$      W$       ]                      �      �       P!      	!       P'$      ,$       PW$      W$       ��                             A      �       ^�      �       U�      �       ^�       �        ^�       !       U!      	!       ^$      D$       ^W$      W$       ^                        z      �       P�       !       P3$      8$       P?$      D$       P                       A      �       }���       �        }���       	!       }��$      D$       }��W$      W$       }��                  �       �        P                             �      �       ]�      8       w �      w       w        &        w 5       R        w �       �        w D$      M$       w                   �      �       T                  �      �       \                    |      �       P�      �       V                         �      8       S�      w       S       &        S5       R        S�       �        SD$      H$       S                      �      �       PH      W       PR       R        0�D$      H$       P                                      �      �       ��}��      �       P�      �       Q�      �       q��      8       Q�             QP      `       ��}�`      n       Rn      w       Q               Q5       E        QE       I        q�I       R        Q�       �        Q                     �      �       ��}��      �       Pc      i      
 � p "
P�                                  �      �       V�      �       U�      8       V�             V             U      w       V       &        V5       N        V�       �        VD$      H$       V                          �      8       \�      w       \       &        \5       R        \�       �        \D$      H$       \                      �      �       R4      8       R�             R                                 �      �       1��      �       ]�      �       R�      8       ]�      w       ]               ]5       R        ]�       �        ]D$      H$       ]                                �      �       0��      �       T�      8       0��             T      w       0�       &        0�5       N        0��       �        0�D$      H$       0�                           4       P4      n       _D$      H$       _                           "       q p �"      C       QC      G       s �                     P      �       r���      �       r�|��      �       r��                       8!      $       ]M$      W$       ]i$      %       ](%      �%       ]                     8!      $       }��M$      W$       }��i$      �%       }��                          _!      h!       Uh!      $       w M$      W$       w i$      %       w (%      �%       w                        _!      $       _M$      W$       _i$      %       _(%      �%       _                                    �!      $       ��{$      $       ��{�#�M$      W$       ��{i$      �$       ��{�$      �$       0��$      �$       \,%      `%       ��{`%      i%       0�i%      n%       Pn%      �%       ��{                        �!      $       ��{M$      W$       ��{i$      %       ��{,%      �%       ��{                             _!      �!       0��!      $       ��{M$      W$       ��{i$      %       ��{(%      ,%       0�,%      v%       ��{v%      �%       R                                   _!      �!       0��!      "       \"      -"       P-"      $       \M$      W$       \i$      w$       \w$      %       S%      %       0�(%      ,%       0�,%      `%       \`%      i%       Si%      �%       \�%      �%       S                          d!      h!       Ph!      $       ��{M$      W$       ��{i$      %       ��{(%      �%       ��{                          �!      P#       SM$      W$       Si$      w$       Sv%      �%       S�%      �%       }�{ "�                                 �!      "       s"      $       ��{M$      W$       ��{i$      %       ��{,%      i%       ��{n%      v%       ��{v%      �%       s�%      �%      	 }�{ "#�%      �%       ��{                            �"      �"       0��"      �"       T�"      �"       1��#      �#       p��#      �#       p�M$      W$       T9%      T%       S                            �!      $       VM$      W$       Vi$      �$       V�$      %       ��{�1�,%      i%       Vn%      �%       V                 #      1#       ��{                     �"      �"       P�"      �"       XM$      W$       P                      �!      "       P"      -"       ��{v%      �%       P                    �"      �"       s�M$      W$       s�                   �"      �"       �^/  M$      W$       �^/                       �"      �"       0��"      �"       QM$      W$       0�                    �"      �"       P�"      �"       p��"      �"       PM$      W$       P                 �#      �#       p3$| "p 3$| "�                   9%      T%       s3$| "s 3$| "�T%      V%       s 3$| "s3$| "�                               �       }���      �       }��      E       }���             }���      �       }��                               �       }���      �       }��      E       }���             }���      �       }��                          g      �       T      (       T(      ,       t�,      8       T8      @       t�@      E       T�      �       T                     g      �       Q      E       Q�      �       Q                        �             U             �U�      �       U�      �       �U�                            �      �       T�             T      (       0�d      w       0��      �       T�      �       �T1�                              �             Q             Q      &       Q&      (       �Q�d      q       Qq      s       �Q�s      }       Q�      �       0�                              �      �       R�             \             �R�      (       R(      d       \d      n       Rn      �       \                       �             U             �U�      �       U�      �       �U�                           �             0�      �       0��      �       P�      �       P�      �       �L�      �       P                       �             u��             �U#��      �       u���      �       �U#��                        /      =       p t "=      @       V@      d       u�t "�      �       u�t "                       /      =       p q "=      d       u�q "�      �       u�q "�      �      
 �U#�q "                    B      d       V�      �       V                   B      d       S�      �       S                     B      d       u��      �       u��      �       �U#�                      �             Q      �       s����      �       s���                    �      �       X�      �       X                                   R      �      2 @K$Os��(  / 0@K$(	 1$#/��O'�%��      �      2 @K$Os��(  / 0@K$(	 1$#/��O'�%�                          �       T�      �       T                                      q r �             Q             s��r �      �      : s��@K$Os��(  / 0@K$(	 1$#/��O'�%��      �      : s��@K$Os��(  / 0@K$(	 1$#/��O'�%�                             8       U8      �       }� �      �       U�      �       }�                          �       y �0.��      �       y �0.�                         �       { �0.��      �       { �0.�                                             ,       Q,      F       ZF      V       QV      `       Zl      �       Q�      �       Z�      �       }� �      �       Z�      �       Q�      �       Z�      �       }� �      �       Z                            0      F       QX      `       R�      �       R�      �       Q�      �       Q�      �       Q                  �      �       R                              �      �       U�      A       SA      `       �U�`      �"       S�"      f#       �U�f#      K%       SK%      �&       �U�                              �      �       T�      A       _A      `       �T�`      �       T�      v%       _v%      �%       �T��%      &       _&      �&       �T�                                              �      �       Q�             V      A       �Q�Q $0.�A      N       VN      `       �Q�Q $0.�`      \       V\      p       �Q�Q $0.�p      #       V#      f#       �Q�Q $0.�f#      K%       VK%      �%       �Q�Q $0.��%      �%       V�%      &       �Q�Q $0.�&      *&       V*&      �&       �Q�Q $0.�                                        �      �       R�      �       ^�      `       �R�`      }       R}      \       ^\      p       �R�p      �"       ^�"      f#       �R�f#      K%       ^K%      �%       �R��%      &       ^&      �&       �R�                             �      �       U�      A       SA      `       �U�`      �"       S�"      f#       �U�f#      K%       SK%      �&       �U�                             �      �       T�      A       _A      `       �T�`      �       T�      v%       _v%      �%       �T��%      &       _&      �&       �T�                        x      �       P�      A       \\      p       \%      �%       0�                        �      �       ]`      �       ]�      �       ���      �       ��                    
      A       V\      p       V                             �      �       u���      A       s��A      `       �U#��`      �"       s���"      f#       �U#��f#      K%       s��K%      �&       �U#��                      @      M       QM      A       ��\      p       ��                   �      A       s0�\      p       s0�                                   P      Y       P\      p       P                              Q                              T                    �      A       ~  $0)�\      p       ~  $0)�                 Y      t       0�                 K      t                         K      t       (                      Y             P      �       pp��      �       P                  t             p       �       pp                   �      �       Q�      �      
 q y "#���                  �      �       q ?&��      �       Y                   �      �       Q�      �      
 q y "#���                  �      �       q ?&��      �       Y                �      �       X                   �      �       U�      �      
 p u "#���                  �      �       u ?&��      �       P                  �      �       T�      �      
 p t "#���                  �      �       t ?&��      �       P                    I      M       XM      x       ��~                  I      x       \                    I      M       QM      x       ��                    I      M       TM      x       w                       I      p       s��p      t       Ut      x       s��                               `      }       r @B$ $0.�}      \       ~ @B$ $0.�p      �"       ~ @B$ $0.��"      f#       �R@B$ $0.�f#      K%       ~ @B$ $0.�K%      %       �R@B$ $0.��%      &       ~ @B$ $0.�&      �&       �R@B$ $0.�                                 `      \       Vp      #       V#      f#       �Q�Q $0.�f#      K%       VK%      %       �Q�Q $0.��%      �%       V�%      &       �Q�Q $0.�&      *&       V*&      �&       �Q�Q $0.�                         `      �       T�      \       _p      v%       _v%      %       �T��%      &       _&      �&       �T�                           `      \       Sp      �"       S�"      f#       �U�f#      K%       SK%      %       �U��%      �&       �U�                                        �             P      (       Pp      �       0�u       �        P�       �        P�       Z!       \Z!      w"       0�w"      �"       P�"      f#       \f#      �#       0��#      *%       \K%      v%       \v%      %       0��%      �&       \                     `      �       ]�      �       ���      �       ��                 `      �       }�                     `      �       }���      �       ��#���      �       ��#��                    �      m        \8%      =%       \                        p      �       ���      Q"       ��f#      =%       ��F%      K%       ��                 `      �       v ����4$}�"�                      n      �       \�      �       ���      �       ��                 n      �       0�                         �      �       4��      �       Q�      �       |�1r  $0)#��      �       Q�      V       ��~                     L      \       �t  �      �       �t  *%      K%       �t                       L      \       �t  �      �       �t  *%      K%       �t                       L      \       Y�      �       Y*%      K%       Y                     L      �       |��      �       ��#��      �       ��#�                   L             T�      �       T                     L      \       [�      �       [*%      K%       [                            \       U�      �       U*%      K%       U                                       T      &       Q&      \       T�      �       T*%      K%       T                       L      a       4�a      \       X�      �       X*%      K%       X                     L      �       u 1��      	       ��~�1��      �       ��~�1�                                  &       \4      D       RD      \       \�      �       \�      �       |�*%      *%       \*%      -%       |�=%      K%       \                      �      �       [�      �       Q�      �       Q                    �             U�      �       U                      �      �       P�      �       P�      �       P                       �      �       	���      �       R�      �       P�      �       R�      �       P                                &       Q.      \       Q�      �       Q�      �       u t "1%�*%      K%       u t "1%�                            &       PP      \       P�      �       P                       p      �       [       V!       0�V!      f"       [f#      �#       [�#      *%       0�                       p      �       ��       V!       0�V!      Y"       ��f#      �#       ���#      *%       0�                                 p      �       ��~'       7        P8       Y        Pf       t        Pt       V!       ��~V!      b"       ��~f#      �$       ��~�$      �$       ��~�$      %%       ��~                         p      �       Q       V!       0�V!      �!       Q�!      f"       s�f#      �#       Q�#      *%       0�                         p      �       P       V!       0�V!      �!       P�!      f"       s�f#      �#       P�#      *%       0�                              p      �       z ��       Z!       0�Z!      f"       z ��f"      f#      	 ��~���f#      �#       z ���#      *%       0�K%      v%      	 ��~����%      �&      	 ��~���                                             p      �       Y�       �        P�       !       t� !      Z!       w #@Z!      f"       Yf"      f#       ��f#      �#       Y�#      $       w #@$      $       P$      $$       t� $$      Z$       PZ$      k$       w #@k$      �$       P�$      �$       t� �$      *%       w #@K%      v%       ���%      �&       ��                   �       Z!       �dv  �#      *%       �dv                     �       Z!       �=v  �#      *%       �=v                     �       Z!       �Wv  �#      *%       �Wv                     �       Z!       �Jv  �#      *%       �Jv                     �       Z!       �0v  �#      *%       �0v                     �       Z!       �#v  �#      *%       �#v                          �       V!       ��~�#      �$       ��~�$      �$       ��~�$      %%       ��~                               �       V!       RV!      Z!       w #H�#      �$       R�$      �$       w #H�$      �$       R�$      �$       w #H�$      %       R%      *%       w #H                   �       Z!       �qv  �#      *%       �qv                    �       Z!       0��#      *%       0�                                 �       !       Z!      	!       z 2%�	!      !       T!      .!       z 2%�.!      5!       z 4%�5!      8!       T8!      Z!       z 4%�Z!      Z!       w #@�4%��#      $       z 2%�$      �$       Z�$      *%       z 4%�                           �       �        P�       �        [�       !       t� #�#      �#       P�#      �#       Q�#      �#       t                                      �       �        P�       �        Q�       �        p��       Z!       Y�#      �#       Y�#      �#       T�#      �#       Y�#      �#       y��#      �#       u~��#      �#       U�#      �#       Y�#      �#       y��#      $       T$      $       p�$      $       p�$      $$       Y$$      1$       p�1$      R$       p�R$      k$       Yk$      x$       p�x$      �$       p��$      �$       t� #��$      �$       Y�$      �$       T�$      �$       Y�$      �$       T�$      %       Y%      *%       T                                �       �        0��       Z!       [�#      $       [$      $       0�$      $$       [$$      R$       0�R$      k$       [k$      �$       0��$      *%       [                                  �       !       0�!      !       P!      Z!       ���#      $       ��$      $       0�$      $$       P$$      f$       0�f$      k$       Pk$      �$       0��$      �$       P�$      *%       ��                              �       V!       0�V!      Z!       ��~�#      �$       0��$      �$       U�$      �$       0��$      �$       U�$      %%       0�%%      *%       U                                  �       .!       0�.!      Z!       Q�#      �#       0��#      �#       Q�#      �#       0��#      �#       Q�#      �#       0��#      $       Q$      �$       0��$      *%       Q                                �       .!       0�.!      Z!       P�#      �#       0��#      �#       P�#      �#       0��#      �#       P�#      �#       0��#      $       P$      �$       0��$      *%       P                      �"      �"       s���"      f#       �U#��K%      v%       �U#���%      �&       �U#��                     �"      �"       }��2 $0.��%      �%       }��2 $0.�&      &       }��2 $0.�                    �"      f#      	 ��~���K%      v%      	 ��~����%      �&      	 ��~���                            �"      #       Y#      f#       ��K%      v%       ���%      �%       Y�%      &       ��&      5&       Y5&      �&       ��                    �"      f#       0�K%      v%       0��%      �&       0�                                               �"      �"       P���"      �"       P�R���"      �"      
 P�s����"      �"      
 P�s����"      #       P�R��#      #       ]�R��#      "#       P�R��"#      f#       ]�R��K%      v%       ]�R���%      �%       P�R���%      �%       [�R���%      �%       P�R���%      &       [�R��&      5&       P�R��5&      =&       ]�R��=&      K&       P�R��K&      �&       ]�R��                 �"      �"       }��2 $0.�                   �"      �"       s���"      �"       �U#��                 �"      �"       �x                     #      f#       YK%      v%       Y                   #      f#       SK%      v%       S                   #      f#       XK%      v%       X                   #      f#       UK%      v%       U                       #      (#       V/#      2#       v ��2#      f#       VK%      v%       V                       #      #       [#      "#       T"#      I#       [I#      M#       {�M#      f#       [K%      v%       [                    #      #       P#      f#       PK%      v%       P                       #      #       z 1%�#      "#       ��"#      I#       ZI#      R#       z 1%�R#      W#       ZW#      f#       ��K%      v%       Z                     #      #       ^#      "#       0�"#      W#       ^W#      f#       0�K%      v%       ^                   �%      �%       Y�%      �%       y��%      &       Y                 �%      &       �x                      �%      �%       Q�%      &       U                  �%      &       S                       �%      �%       T�%      �%       Z�%      �%       T�%      �%       Z�%      �%       z��%      &       Z                  �%      �%       P�%      &       P                         �%      �%       ���%      �%       x 1%��%      �%       ���%      �%       X�%      �%       x 1%��%      �%       X�%      �%       ���%      &       X                   �%      �%       0��%      &       ]                       �%      �%       0��%      �%       Q�%      �%       0��%      �%       Q�%      �%       0��%      &       Q                      5&      [&       Yc&      �&       Y�&      �&       y��&      �&       Y                         [&      h&       [�&      �&       1��&      �&       [�&      �&       0��&      �&       [�&      �&       [                     5&      �&       X�&      �&       X�&      �&       X                        5&      [&       �^�c&      �&       �^��&      �&       �^��&      �&       �^�                  5&      �&       U                      5&      Q&       VX&      [&       v ��[&      �&       V                      5&      8&       S8&      K&       TK&      h&       Sh&      k&       s�k&      �&       S                   5&      =&       P=&      �&       P                        5&      8&       z 1%�8&      K&       ��K&      h&       Zh&      p&       z 1%�p&      u&       Zu&      �&       ���&      �&       Z                      5&      =&       _=&      K&       0�K&      u&       _u&      �&       0��&      �&       _                       �&      �&       x ���&      �&       { ���&      �&       ~ ���&      �&       y���                      �      �       U�             S             �U�                     �      �       U�             S             �U�                   �      �       u���      �       s��                  �      �       V                            %       U%      c       Qc      k       �U�                           %       U%      c       Qc      k       �U�                  (      c       T                 (      c       T                                        �(      �(       U�(      �(       V�(      �(       �U��(      }.       V}.      /       ��/      2       �U�2      �2       ���2      �2       �U��2      �2       ���2      5       �U�5      �5       V�5      �5       �U�                                        �(      �(       T�(      �(       S�(      �(       �T��(      1.       S1.      5       �T�5      05       S05      �5       ��~�5      �5       �T��5      �5       ��~�5      �5       �T��5      �5       ��~�5      �5       �T�                              �(      �(       Q�(      �(       \�(      �(       �Q��(      /*       \/*      },       �Q�},      �,       \�,      �5       �Q�                    �(      �(       R�(      �5       �R�                    �(      �(       X�(      �5       �X�                                        �(      �(       T�(      �(       S�(      �(       �T��(      1.       S1.      5       �T�5      05       S05      �5       ��~�5      �5       �T��5      �5       ��~�5      �5       �T��5      �5       ��~�5      �5       �T�                 �,      �,       8�                  �)      �)       Q�,      �,       0�                 &)      �)       �-}  },      �,       �-}                     &)      7)       s�7)      �)       ]},      �,       ]                 &)      �)       V},      �,       V                      T)      c)       q 
���c)      �)       R�)      �)       q 
���},      �,       q 
���                   &)      �)       0��)      �)       q 
���},      �,       0�                   T/      2       s���2      �2       s��                   n/      �/       0��/      �/       P                 �1      �1       0�                 �1      2       V                     �1      �1       Q�1      �1       q`��1      2       Q                      �1      �1       U�1      �1       uX��1      2       U                 �1      �1       s�#8                     H1      m1       0�m1      ~1       Q�2      �2       0�                        N1      b1       Qb1      m1       s��2      �2       Q�2      �2       s�                    U1      �1       P�2      �2       P                    �(      �(       U�(      �(       V�(      �(       V                    �(      �(       t���(      �(       s���(      �(       s��                       �(      �(       P�(      �(       P�(      �(       P�(      �(       0�                �(      &)       s��                �(      &)       1�                    �)      },       }  $0.��,      �,       }  $0.�                  �)      �)       s�                    �)      },       V�,      �,       V                    �)      },       s���,      �,       s��                  �)      *       q 
���                    !+      �+       u ���,      �,       u ��                    K*      f*       Tf*      p*       s�                        /*      [*       | 
���[*      p*       Pp*      },       | 
����,      �,       | 
���                                     �*      �*       Q�*      �*       q��*      �*       q��*      �*       q	��*      !+       q�!+      u+       Pu+      +       Y+      �+       P�+      �+       p��+      �+       P�+      �+       p��+      �+       P�+      �+       r�,      -,       P-,      B,       p�B,      l,       p�l,      p,       p�p,      },       Q�,      �,       P                    �*      },       T�,      �,       T                       !+      *+       0�*+      7+       1�7+      I+       RI+      S+       r�S+      \+       {�\+      _+       R                �+      ,       T                �+      ,       ���                  �+      ,       0�                �+      ,       T                �+      ,       ���                  �+      ,       0�                  �+      �+       P�+      �+       R�+      ,       P,      ,       p�,      ,       R,      ,       P                 �+      ,       Q                   ,      	,       p���	,      ,       r���                   ,      	,       p ���	,      ,       r~���                    �,      1.       \5      %5       \                        �,      �,       P�,      H/       ��2      �2       ���2      �5       ��                                �,      }.       V}.      /       ��/      H/       �U�2      �2       ���2      �2       ���2      5       �U�5      �5       V�5      �5       �U�                                      �,      1.       s��1.      H/       �T#��2      �2       �T#���2      5       �T#��5      05       s��05      �5       ��~#���5      �5       �T#���5      �5       ��~#���5      �5       �T#���5      �5       ��~#���5      �5       �T#��                        �,      �,       R�,      H/       w 2      �2       w �2      �5       w                           �-      .       q ��.      /      	 �����2      �2      	 ������2      
4      	 �����5      �5      	 �����                            U.      X.       q x !�����X.      �.      	 q ������.      �.       V�.      �.       v | ��.      /       V2      �2       V5      5      	 q �����                                                4-      =-       P=-      T-       p�T-      l-       p�l-      �-       p��-      �-       p��-      �-       p
��-      �-       p��-      �-       p��-      	.       ]	.      .       p�.      >.       ]>.      �.       P�2      �2       ^�2      3       ]3      3      
 q 1$~ "#�3      /3      
 q 1$~ "#�/3      G3      
 q 1$~ "#�G3      X3       }�X3      g3       }�g3      �3       }��3      �3       }��3      W4       \W4      ^4       p�^4      �4       P�4      �4       T�4      �4       \�4      5       P5      -5       ]-5      05       p��5      �5       ]�5      �5       T�5      �5       \�5      �5       P�5      �5       T                                 4-      �.       Z�.      /       ��~2      �2       ��~�2      �2       ��~5      05       Z05      �5       S�5      �5       S�5      �5       S�5      �5       Z                          a.      �.       P�.      �.       U�.      �.       S�.      �.       P�.      �.       p��.      /       U2      *2       U*2      *2       u
�*2      C2       u�C2      \2       u�\2      v2       u�v2      �2       U                      �.      �.       S�.      /       S2      �2       S                              �.      �.       Q�.      �.       | 
����.      /       Q/      /       | 
���2      !2       Q!2      v2       | 
���v2      �2       Q                      �.      �.       r 
����.      /       r 
���2      02       r 
���                      3      +3       Q+3      /3       q�/3      q3       Q                    �2      �2       [�2      �3       ��                    W4      5       R�5      �5       R                    �3      5       ]�5      �5       ]                   �3      �3       4��3      4       P                     W4      �4       Q�4      5       Q�5      �5       Q                 5      �5      
 @�F     ��5      �5      
 @�F     �                         5      05       s��05      �5       ��~#���5      �5       �T#���5      �5       ��~#���5      �5       �T#���5      �5       ��~#��                        5      05       Z05      �5       S�5      �5       S�5      �5       S�5      �5       Z                 5      �5       �q�  �5      �5       �q�                     5      �5       0��5      �5       P�5      �5       0�                       5      5       ]5      05       P05      >5       ]>5      >5       }�>5      m5       Um5      s5       ]s5      5       U�5      �5       ]                     5      �5       ^�5      �5       ^�5      �5       ^                      C5      m5       Qs5      {5       Q{5      5       u���                     >5      H5       } ���H5      m5       u~���s5      5       u~���                      P5      \5      
 @�F     �\5      m5       Ps5      x5      
 @�F     �                            �
      �
       U�
      s       Vs      x       �U�x      �       V�      �       �U��      �       V                      �
      �
       T�
      r       S�      �       S�      �       Q                            �
      �
       Q�
      w       ]w      x       �Q�x      �       ]�      �       �Q��      �       ]                            �
      �
       R�
      u       \u      x       �R�x      �       \�      �       �R��      �       \                             �
      H       0�H      L       PL      ]       Ri      x       Rx      �       0��      �       R�      �       0�                                    0�      )       P1      D       P�      �       0�                   5      x       1��      �       q  $0.��                              p      �       U�      �       S�      �       s��      �       s��      Y	       RY	      �	       s��	      
       R
      
       s�
      ,
       R,
      =
       s�                            p      |       T|      �	       \�	      �	       �T��	      �	       \�	      �	       �T��	      =
       \                            p      �       Q�      �	       V�	      �	       �Q��	      �	       V�	      �	       �Q��	      =
       V                             p      �       0��      �       P�      �	       T�	      �	       T�	      �	       0��	      
       T
      
       0�
      =
       T                 �	      �	       8�                     �      �	       ]�	      �	       ]�	      =
       ]                                U	      \	       u �8$y �!
���\	      w	       s��8$y �!
���w	      z	       q ��8$q��!
���z	      }	       r 8$q��!
���}	      �	       q ��8$q��!
����	      �	      @ t��1z ����s "#��8$t��1z ����s "#��!
���
      #
       u ��)
      ,
       q ���,
      3
       R3
      8
       t��1z ����s "#���                                 U	      Y	       s��8$s��!
���Y	      b	       r 8$s��!
���b	      w	       s��8$s��!
���w	      �	       q��8$q��!
����	      �	       u 8$q��!
����	      �	      & u 8$t��1z ����s "#��!
����	      �	      @ t��1z ����s "#��8$t��1z ����s "#��!
���
      )
       y ��)
      0
       q���0
      5
       Q5
      8
       t��1z ����s "#���                      U	      U	       RU	      U	       r�U	      Y	       r�Y	      w	       s�w	      w	       t��1t�����s "#�w	      w	       t��1t�����s "#�w	      �	       t��1t�����s "#�
      
       R
      
       r�
      )
       r�)
      )
       t��1t�����r "�)
      )
       t��1t�����r "#�)
      ,
       t��1t�����r "#�,
      =
       t��1t�����s "#�                                          U&      >       U>      Z       XZ      o       u�o      �       s��      �      
 q 1$s "#��      �      
 q 1$s "#��      �      
 q 1$s "#�                                      T      &       �T�&      {       T{      �       �T�                                      Q      &       �Q�&      v       Qv      �       V                              A      G       r ��G      K       | ��K      R       u ���R      �       ]�      �       q  } "��      �       } q ��      �       q  } "�                      K      O       | ��O      R       ]R      �       | ��                     K      W       RW      o      
 u ��4%�o            
 s ��4%�                                           0�&      �       0��      �       P�      �       U�      �      
 q 2$u "#��      �       q 2$u "��      �      
 q 2$u "#�                                  q &      v       q v             v                           @
      Y
       UY
      b
       �U�b
      |
       U|
      �
       \�
      �
       �U�                        @
      Y
       TY
      b
       �T�b
      
       T
      �
       �T�                          @
      Y
       QY
      b
       �Q�b
      s
       Qs
      �
       S�
      �
       �Q�                     W
      Y
       q b
      s
       q s
      �
       s                            W
      Y
       t u �Y
      b
       �T�U�b
      |
       t u �|
      
       t | �
      �
       �T| ��
      �
       �T�U�                                          �             U             u�             u�      �       S�      �       ^�      �       X�      �       x��             S      :       X:      o       So      �       ^�      �       X�      �       x��      �       S�      �       X�      �       S4      �       S                          �      8       T8             _      4       �T�4      F       TF      �       _                        �             Q             \      4       �Q�4      �       \                    �      8       P4      Y       P                               w      �       q ����(x "��      �      	 p (x "��      �       q ����(x "��      6       P6      N       pX�N      �       P�      �       pX��      �       P                          p       v ��4      �       v ��                  �      �       0�                                 ]4      �       ]                   8      Q       8�Q      {       P                        %       8�                    M      Y       ZY      �       ��                               3       U3      f       _f      g       �U�g      �       _                               .       T.      d       ^d      g       �T�g      �       ^                                                               J       QJ      R       ��~R      g       �Q�g      �       ��~�      �       �Q��      �       ��~�      �       �Q��      �       ��~�      �       �Q��      �       ��~�      �       �Q��      <       ��~<      l       �Q�l      �       ��~�      ,       �Q�,      �       ��~�      9       �Q�9      A       ��~A      �       �Q��      �       ��~                           J       RJ      �       �R�                                             J       XJ      R       ]R      g       �X�g      �       ]�      �       �X��      �       ]�      �       �X��             ]      z       �X�z      �       ]�      �       �X�                                                      N      R       Pg      z       Pz      ~       \~      �       P�             \�      �       \�      �       ���      �       \�      �       S�      -       0�-      E       P�      �       0��      C       \l      �       \e      p       Pp      z       0�z      �       \9      <       \�      �       \�      �       ���      �       S                                       �      �       P�             ~� �      �       P�      �       P�      �       ~� �      +       P+      �       ~� V      �       P*      4       P4      C       ~� �      �       ~� z      �       ~�                       �      �       V�      ,       Vz      �       V                 �             0�                                    �      �       T�      �       T�      �       �      V       ��~�             ��~�      *       ��~l      �       ��~z      �       T9      A       ��~�      �       ��~                     �      �       ���~���      �       P�             ���~��                     �      �       (�      �       (z      �       (                     �      �       (#��      �       (#�z      �       (#�                  o      �       0�,      N       0�                        (      �       V�      �      	 | 0$0&�,      p       Vp      u      	 | 0$0&�                          R      v       Rv      �       z v ��      �       z | 0$0&�,      e       Rp      u       z | 0$0&�                                    ,       YM      �       Q�      �       y } "��      �      	 y } " �,      C       QC      e       y } "�p      z      	 y } " �                      �      �       P�      �       pp��      �       P                   �      �       Q�      �      
 q v "#���                  �      �       q ?&��      �       V                  �      �       p �      �       pp                   �      �       Q�      �      
 q v "#���                  �      �       q ?&��      �       V                  N      e       P                              �      �       V�      V       V�      �       V�      *       Vl      �       Vz      �       V9      A       V�      �       V                                               �      �       P�      �       P�      +       p�+      a       ~� #�a             S             P      #       Y#      H       PH      N       YN      j       Pj      �       T�      �       S�      �       P�             P      6       U6      V       P�      �       P�      �       T�      �       S�             T      *       Sl      }       P}      �       Y�      �       P�      �       Yz      �       S9      A       S�      �       S                              �      �       _�      V       _�      �       _�      *       _l      �       _z      �       _9      A       _�      �       _                     �      �       (�      �       (z      �       (                     �      �       (�      �       (z      �       (                             �      �       Q�      �       q`��      V       Q�      �       Q�      *       Ql      �       Q�      �       Q                        �      �       q ���      +       p ���+      �      
 ~� ���z      �      
 ~� ���                  �             0��      �       0�                                        �       [�      �       ��~�      V      	 ��~����      �      	 ��~����      *      	 ��~���l      �      	 ��~���z      �       [9      A       ��~�      �      	 ��~���                            a      V       ��~�      �       ��~�      *       ��~l      �       ��~z      �       ��~9      A       ��~�      �       ��~                                �              0�       m       Um      �       q�      �       qp�      V       0��      �       U�      *       ql      �       0��      �       U                                    �      K       0�K      a       Ta      �       q�      �       qt�      V       0��      �       0��      �       T�      �       q�      *       ql      �       0��      �       T                   �      �       ]9      A       ]                 	      a       V                 	      a       �                   	      a       0�                 	      a       V                 	      a       �                   	      a       0�                            	             p�             S      '       p�'      '       p�'      .       S.      8       ~� #�8      M       SM      M       s�M      P       s�P      S       p s "#�S      \       s�\      a       S                          \       Q\      _       q�_      a       Q                         '      +       p���+      .       s p "#���.      P       s���P      S       p s "#���S      a       s���                         '      +       p���+      M       ~� #���M      P       s ���P      S       p s "���S      \       s ���\      a       ~� #���                                �       R�      V       R�      �       R�             Rl      �       R                             �      �       V�      �       VV      �       V*      l       V�      ,       V�      9       VA      �       V                                                                �      �       P�      �       p��      )       S)      =       Y=      d       Sd      j       Pj      y       Sy      �       P�      �       p��      �       S�      �       PV      m       p�m      �       S*      x       Sx      {       q s "�{      �       S�      �       q s "��      �       S�      �       P�      �       \�      �       Y�      �       \�      �       \�             Q             \      9       Q9      .       \3      �       \�      �       Q�      �       \�             Q             \      C       QC      V       \V      l       Q�      ,       S�      9       \A      u       \u      }       Q}      �       \                             �      �       _�      �       _V      �       _*      l       _�      ,       _�      9       _A      �       _                        �             (�      �       (V      �       (*      C       (�      �       (                          �      �       } ���      �       } ��V      �       } ��*      G       } ���      ,       } ��                              �      �       0��             [�      �       0�V      r       0�r      �       [*      C       0��      �       [�      ,       ��~                              �      �       0��      �       P�      �       ��~�      �       0��      �       S�      �       ��~V      �       0�*      C       0��      ,       ��~                     
             0�F      V       q�V      j       Q'      ,       0�                           �      �       p ���      �       { ���      �       ~� #����            	 { ��~�"�*      C       0��      �      	 { ��~�"��      ,       ��~���~�"�                     
             0�d      g       s ���g      j       TC      C       0�'      ,       0�                      
             0�      ,       R=      �       RC      C       0�'      ,       0�                  M      �       Vu      }       V                  M      �       ��  u      }       ��                    M      �       0�u      }       0�                  M      �       Vu      }       V                  M      �       ��  u      }       ��                    M      �       0�u      }       0�                         M      \       S\      t       s�t      t       s�t      �       Q�      �       S�      �       s��      �       s��      �       q s "#��      �       s��      �       Su      }       q�                     _      �       P�      �       p��      �       Pu      }       P                           t      x       s���x      {       q s "#���{      �       s����      �       s����      �       q s "#����      �       s����      �       s���                           t      x       s���x      {       q s "#���{      �       s����      �       s ����      �       q s "����      �       s ����      �       s���                       �      l       _�      9       _A      u       _}      �       _                       *      �       tp��      Z       tp�Z      c       T�      �       ����      l       tp�                              �      �       r ���      �       p ���      *       |���w      �       |����      �       |����      �       |����      �       |���                                           X      *       p ��w      �       X�      �       p ���      �       X�      �       p ���      �       X                             �             0�*      c       Xw      �       0��      �       
+��      �       0��      l       X�      �       0�                         *             Y�      �       3��      c       Y�      �       3��      �       0��      l       Y                      *      �       U�      Z       U�      �       0��      l       U                            �      �       z ���             p ��             q���&      3       z ��3      :       p ��:      >       q���                      �      �       | �8$8&��      �       q�8$8&�V      c       | �8$8&�c      g       q�8$8&�                       )       _                      3      �       ����      �       Q�      �       ���      9       ���                  3      �       _      9       _                 3      C       (                   �      �       P,      9       P                     �             _A      u       _}      �       _                     �             ���A      u       ���}      �       ���                     �             ���A      u       ���}      �       ���                     �             ���A      u       ���}      �       ���                    �      �       (A      T       (h      h       (                     �      �       (#`�A      T       (#`�h      u       (#`�                                  0�U      c       Ph      h       8�}      }       P                 �             T                �             R                    �      �       P�      ,       ��~                    �      �       U�      �       �U�                    �      �       T�      �       �T�                        �      �       U�      7       S7      A       �U�A      U       S                      �             T      A       �T�A      U       T                      �             Q      A       �Q�A      U       Q                        �             R      >       ]>      A       �R�A      U       R                        �             X      <       \<      A       �X�A      U       X                       �      �       U�      7       S7      A       �U�A      U       S                       �      �       u���      7       s��7      A       �U#��A      U       s��                       �             @<$�      #       P#      @       ^A      U       @<$�                     �      $       @<$�$      9       PA      U       @<$�                    �      :       VA      U       V                      �      �       T�      �       T�      �       �T1�                 �      �       U                 �      �       6��      �       0�                 �      �       u��                             �       A       0�A      E       PE      J       p�J      Y       PY      \       0�\      j       Qj      �       0��      �       P�      �       Q�      �       P                        �       9       Y9      U       0�U      {       Y{      �       0��      �       Y                         �       �        0��       J       PJ      Y       p�Y      �       P�      �       P                           �       �        u�              R      9       XY      \       Rj      p       Rp      {       X                                           Q      %       X%      )       R)      4       Q4      9       XY      \       Xj      p       X                                             q ����4$z "�      %       x ����4$z "�%      )       r ����4$z "�)      4       q ����4$z "�4      9       x ����4$z "�A      G       p ����4$u "�G      N      	 q 4$u "�N      Y       p����4$u "�Y      \       x ����4$z "�j      p       x ����4$z "�                   p       v        0�v       �        X                          s       �        Q�       �        R�       �        Q�       �        Q�       �        R                           �       �        p ����4$y "��       �        r ����4$y "��       �        q ����4$y "��       �        p ����4$y "��       �        r ����4$y "��       �        r ����4$y "��       �        r ����4$y "�                              �       �        P�       �        R�       �        Q�       �        P�       �        R�       �        R�       �        R                                    T       V        �T�                           P        0�P       V        8�                                   P       V        u                         3        1�                 `             U                 `             u� �                      }      �       R�      �       {��      �       R                     }      �       0��      �       Q�      �       Q                    �      �       X�      �       X                    �      �       Y�      �       Y                                          U       J       SJ      L       �U�L      l       Sl      n       �U�n      �       S                                  T       �       �T�                                  Q       �       �Q�                                          R       K       VK      L       �R�L      m       Vm      n       �R�n      �       V                                         U       J       SJ      L       �U�L      l       Sl      n       �U�n      �       S                                         u��       J       s��J      L       �U#��L      l       s��l      n       �U#��n      �       s��                      :      C       �T�L      n       �T�}      �       �T�                      :      C       �Q�L      n       �Q�}      �       �Q�                        :      C       VL      m       Vm      n       �R�}      �       V                        :      C       SL      l       Sl      n       �U�}      �       S                       �      �       U�      �       S�             S             U                       �      �       u� ��      �       s� ��             s� �             u� �                  �             P                 �      �       s� �0$0&�                        �&      "'       U"'      t(       St(      z(       �U�z(      �(       U                       �&      "'       U"'      t(       St(      z(       �U�z(      �(       U                      �&      "'       U"'      t(       St(      z(       �U�                  '      y(       ]                 '      b(       V                   '      "'       u��"'      b(       s��                    (      2(       T3(      3(       0�3(      ;(       \;(      J(       T                  +(      ;(       \                    �      �       U�      �       �U�                        �      �       T�      �       ^�      �       �T��      �       ^                       �      �       T�      �       ^�      �       �T��      �       ^                       �      �       t���      �       ~���      �       �T#���      �       ~��                       �      �       t���      �       ~���      �       �T#���      �       ~��                       �      �       t���      �       ~���      �       �T#���      �       ~��                      �      �       ]�      �       ]�      _       ]                                            p      {       P�      �       P�      �       P�      �       P�      �       P	             P5      K       P\      k       P�      �       P�      �       P�      �       P�      �       P�      �       PR      a       P                     �      �       _�      �       _�      _       _                                  �             _!      S       _      _       \_      x       _x      �       Q#      &       Q&      K       ���      �       _�      �       Q                      �      �       S�      �       S�      �       S                        �      �       ��_      �       ���      �       P�      �       ��                           �      �       0��      �       ���      �       0��      _       0�_      �       ��      �       ��                         �      �       0��      �       ���      �       0��      _       0�_      �       ��                   �             0�      _       V                              �      �       R�      #       ��B      Q       YQ      �       ���      �       P�      �       R�      �       P                  g      �       0�                                         U      �       V�      �       �U��      �       V�       	       �U� 	      /
       V                                  =       T=      �       S�      �       U�      
       �T�
      
       S
      /
       �T�                                 =       T=      �       S�      �       U�      
       �T�
      
       S
      /
       �T�                      /      3       P3      �       w 
      
       w                                     n      �       [�      �       [�      �       z �      �       {�	      @	       [@	      �	       ��
      
       [
      

       s 

      
       {�
      
       ��
      /
       [                        ;      =       P=      �       _�      �       ��
      
       _                              ;      �       0��      �       ���      �       ���      �       P�      7       ��7      
       ��
      
       0�
      /
       ��                                           `      �       0��      �       ]�      ,       ],      <       Q<      ]       ]]      m       Rm      �       ]�      �       P�      )       ])      V       QV      �       ] 	      
       ]
      
       0�
      /
       ]                              ?      p       [4      a       [a      e       {�e      �       [�      �       {��      �       [�              ��7      V       [�	      �	       [                                         `      �       0��      �       ^�      �       P�      �       ^�      �       ^ 	      	       ^	      	       p�	      m	       ^m	      p	       | 1&�p	      �	       \�	      �	       ^
      
       0�
      /
       ^                               `      �       0��      e       ��q      �       ��x              �� 	      �	       ���	      �	       \�	      �	       ��
      
       0�
      /
       ��                                   ;      �       0��      �       S�      �       0��      �       S�      �       _�       	       0� 	      �	       S�	      �	       P�	      �	       S�	      
       _
      
       0�
      "
       S"
      /
       _                                ;      �       0��      e       ��q      �       ���      �       0�x              ���      �       �� 	      �	       ���	      �	       1��	      �	       ��
      
       0�
      "
       ��"
      /
       1�                                     `      �       0��      e       _q      �       _�      �       _�      �       1��      x       2��      �       0��      C       1�F      �       1� 	      �	       _
      
       0�
      
       _
      
       _                      ?      �       \�      �       \�	      �	       \                    �      �       P�             ^                    �      �       0�V      �       0�                      i      �       Q�      �       q}��      �       Q                     b      �       v�#��      �       T�      �       tp��      �       v�#�                                              �      �       U�      D       VD      S       �U�S      �       V�      �       ���      �       V�      �       �U��             V      '       �U�'      :       V:      C       �U�C      o       Vo      3       ��3      E       �U�E      s       ��                                    �      �       T�      P       ^P      S       �T�S      �       ^�      �       �T��      $       ^$      '       �T�'      @       ^@      C       ����C      s       ^                                   �      �       T�      P       ^P      S       �T�S      �       ^�      �       �T��      $       ^$      '       �T�'      @       ^@      C       ����C      s       ^                                                 �      -       _S      �       _�      .       V.      N       ]N      �       V�      �       _'      B       _C      o       _o      w       Vw      |       ]|      �       V�             ]      +       V3      E       _E      P       VP      T       ]T      V       _V      s       ]                              �      D       SS      �       S�      �       w �      �       S�             S'      9       SC      o       S                           �      D       ]S      �       ]�      �       ]�      "       ]'      >       ]C      o       ]                               S      �       v���      �       ��#��'      :       v��:      C       �U#��C      o       v��o      3       ��#��3      E       �U#��E      s       ��#��                     w      �       P�      �       \C      o       
 �                                  �      �       0��      �       S�      �       T�      �       s��      �       S�      �       0��      �       w o              w       3       w E      s       w                        S      �       ~��'      @       ~��@      C       ��C      s       ~��                            `      n       Rn      �       w '      8       w 8      C       ��C      `       R`      o       w                    `      �       0�C      C       0�C      o       1�                              ;       \o      �       w �      �       RV      s       \                    �      �       P�             V                          0
      D
       UD
      J       SJ      N       �U�N      \       S\      `       �U�                          0
      =
       T=
      K       VK      N       �T�N      ]       V]      `       �T�                          8
      =
       T=
      K       VK      N       �T�N      ]       V]      `       �T�                          A
      D
       u��D
      J       s��J      N       �U#��N      \       s��\      `       �U#��                         A
      D
       u��D
      J       s��J      N       �U#��N      \       s��\      `       �U#��                  \
      �
       p �                  N
      \
       P                    �      �       U�      �       �U�                   �      �       U�      �       �U�                        �      �       U�      �       S�      �       �U��             U                       �      �       U�      �       S�      �       �U��             U                      �      �       P�             P             u                     �      �       P�             P             u                     �      �       0��      �       P�             0�                      �       �        U�               S       $       �U�                      �       �        T�       #       \#      $       �T�                     �       �        U�               S       $       �U�                  �       !       V                  �       $       P                      0      A       UA      �       S�      �       �U�                      0      E       TE      �       \�      �       �T�                     0      A       UA      �       S�      �       �U�                  =      �       V                  U      �       P                             8       U8      T       ST      V       �U�                            8       U8      T       ST      V       �U�                        !       u                         !       u                       D      L       PL      U       VU      V       P                          @      H       UH      a       Sa      b       �U�b      n       Sn      o       �U�                         @      H       UH      a       Sa      b       �U�b      n       Sn      o       �U�                    R      Z       Pb      m       P                        `      �       U�      /       S/      1       �U�1      9       U                       `      �       U�      /       S/      1       �U�1      9       U                     n      �       u���      /       s��/      1       �U#��                     n      �       u���      /       s��/      1       �U#��                  y      0       V                    �      �       U�      �%       �U�                                                          �      �       T�      @       S@      �       �T��      J       SJ      �       �T��             S      �       ��z�      �       �T��      ;        S;               �T�       J!       ��zJ!      w!       �T�w!      n"       ��zn"      R$       �T�R$      b$       ��zb$      �$       S�$      �$       �T��$      +%       S+%      N%       ��zN%      [%       �T�[%      �%       ��z                    �      �       Q�      �%       ��y                    �      �       R�      �       ��z                  �      �       X�      �       ��z                                                         �      �       T�      @       S@      �       �T��      J       SJ      �       �T��             S      �       ��z�      �       �T��      ;        S;               �T�       J!       ��zJ!      w!       �T�w!      n"       ��zn"      R$       �T�R$      b$       ��zb$      �$       S�$      �$       �T��$      +%       S+%      N%       ��zN%      [%       �T�[%      �%       ��z                                    �      �       ^~      %       ^%      4       P:      A       PA      Q       ^Q      �       0��      �       \�      �       ^�      �       P;               0��$      �$       ^                   �      �       P�      �%       ��z                                           �             P      @       ]�      J       ]�      �       P�             ]      �       ��z�      ;        ]       J!       ��zw!      n"       ��zR$      b$       ��zb$      �$       ]�$      +%       ]+%      N%       ��z[%      �%       ��z                                                         �      �       T�      @       S@      �       �T��      J       SJ      �       �T��             S      �       ��z�      �       �T��      ;        S;               �T�       J!       ��zJ!      w!       �T�w!      n"       ��zn"      R$       �T�R$      b$       ��zb$      �$       S�$      �$       �T��$      +%       S+%      N%       ��zN%      [%       �T�[%      �%       ��z                                                         �      �       t���      @       s��@      �       �T#���      J       s��J      �       �T#���             s��      �       ��z#���      �       �T#���      ;        s��;               �T#��       J!       ��z#��J!      w!       �T#��w!      n"       ��z#��n"      R$       �T#��R$      b$       ��z#��b$      �$       s���$      �$       �T#���$      +%       s��+%      N%       ��z#��N%      [%       �T#��[%      �%       ��z#��                                                         �      �       t���      @       s��@      �       �T#���      J       s��J      �       �T#���             s��      �       ��z#���      �       �T#���      ;        s��;               �T#��       J!       ��z#��J!      w!       �T#��w!      n"       ��z#��n"      R$       �T#��R$      b$       ��z#��b$      �$       s���$      �$       �T#���$      +%       s��+%      N%       ��z#��N%      [%       �T#��[%      �%       ��z#��                 �      �       U                    �      �       P�      �%       ��z                          I      �       T�      �       t��      �       T�      �       T�      �       t��      �       T�$      �$       T                     I      �       Q�      �       Q�$      �$       Q                          �       ];               ]                       d      �       0��      �       U�      �       0��      �       U;       \        0�\       a        Ua       z        0�z               U                                                           @       S@      �       �T��      J       SJ      ~       �T��             S      �       ��z�      ;        S       J!       ��zJ!      w!       �T�w!      n"       ��zn"      R$       �T�R$      b$       ��zb$      �$       S�$      �$       �T��$      �$       �T��$      +%       S+%      N%       ��zN%      [%       �T�[%      �%       ��z                             #      �       V�      �       V�      S"       VS"      Y"       UY"      [%       V[%      a%       Ua%      �%       V                                                             @       s��@      �       �T#���      J       s��J      �       �T#���             s��      �       ��z#���      �       �T#���      ;        s��;               �T#��       J!       ��z#��J!      w!       �T#��w!      n"       ��z#��n"      R$       �T#��R$      b$       ��z#��b$      �$       s���$      �$       �T#���$      +%       s��+%      N%       ��z#��N%      [%       �T#��[%      �%       ��z#��                                   @       ^�      J       ^�             ^�      ;        ^b$      �$       ^�$      +%       ^                                              @       ]�      J       ]�             ]      �       ��z�      ;        ]       J!       ��zw!      n"       ��zR$      b$       ��zb$      �$       ]�$      +%       ]+%      N%       ��z[%      �%       ��z                                                              @       S@      �       �T��      J       SJ      �       �T��             S      �       ��z�      �       �T��      ;        S;               �T�       J!       ��zJ!      w!       �T�w!      n"       ��zn"      R$       �T�R$      b$       ��zb$      �$       S�$      �$       �T��$      +%       S+%      N%       ��zN%      [%       �T�[%      �%       ��z                         #       U#      #       V                   @      �       VS      ~       V                   @      �       VS      ~       V                   �      �       VS      ~       V                   �      �       ��{S      l       ��{                                     �      J       ]�             ]      �       ��z�      ;        ]       J!       ��zw!      n"       ��zR$      b$       ��zb$      �$       ]�$      +%       ]+%      N%       ��z[%      �%       ��z                         �      �       R�      J       ^�      �       ^�               ^b$      �$       ^�$      +%       ^                       �      J       _�      �       _�               _b$      �$       _�$      +%       _                       �      J       V�      �       V�               Vb$      �$       V�$      +%       V                    m      �       \�$      &%       \                 �      �       ��|                 �      �       ��|                                �      �       V       Q!       Vw!      S"       VS"      Y"       UY"      n"       VR$      b$       V+%      N%       V[%      a%       Ua%      �%       V                              �             S      �       ��z       J!       ��zJ!      Q!       �T�w!      n"       ��zR$      b$       ��z+%      N%       ��z[%      �%       ��z                                 �      �       V       S"       VS"      Y"       UY"      b$       V�$      �$       V�$      �$       V+%      [%       V[%      a%       Ua%      �%       V                 �      �      
 ��|��|"�                	         �      �       D�       b$       D��$      �$       D��$      �$       D�+%      �%       D�                                           9       ]9      u       ^�      �       ]       �        ]�       �        ^�       �        Pw!      �!       ^�!      n"       ��zR$      b$       ��z+%      N%       ��z[%      �%       ��z                          c      u       _w!      n"       _R$      b$       _+%      N%       _[%      �%       _                        �!      n"       SR$      b$       S+%      N%       S[%      �%       S                                     �!      �!       s  $ &0��F     "��!      �!       s $ &0��F     "��!      �!       s  $ &0��F     "��!      7"       r 0��F     "�7"      n"       s  $ &0��F     "�R$      b$       s $ &0��F     "�+%      N%       r 0��F     "�[%      g%       s  $ &0��F     "�g%      q%       r 0��F     "�q%      ~%       s  $ &0��F     "�~%      �%       r 0��F     "�                           �!      �!       s  $ &0��F     "�!      �!       s $ &0��F     "�!      n"       s  $ &0��F     "R$      b$       s $ &0��F     "+%      N%       s  $ &0��F     "[%      �%       s  $ &0��F     "                            �!      7"       r 0��F     "�7"      Z"       s  $ &0��F     "�+%      N%       r 0��F     "�[%      g%       s  $ &0��F     "�g%      q%       r 0��F     "�q%      ~%       s  $ &0��F     "�~%      �%       r 0��F     "�                          �!      S"       VS"      Y"       UY"      Z"       V+%      N%       V[%      a%       Ua%      �%       V                    �!      Z"       ��z+%      N%       ��z[%      �%       ��z                     Z"      Z"       Pb%      g%       Py%      ~%       P                         E"      M"       ��z�M"      Y"       QY"      Z"       ��z�[%      a%       Qa%      g%       ��z�                     �!      n"       0�+%      N%       0�[%      �%       0�                  �       =!       ^                                #      u#       0�u#      �#       ��z�#      �#       _�#      �#       p��#      R$       ��z�1��$      �$       ��z�1��$      �$       ��zN%      [%       0�                        �#      �#       0��#      �#       ��#      $       _�$      �$       �                        #      R$       0��$      �$       0��$      �$       0�N%      [%       0�                          #      u#       0�u#      M$       ��z�$      �$       ��z�$      �$       ��zN%      [%       0�                        u#      �#       \�#      R$       \�$      �$       \�$      �$       \                      �#      �#       S�#      .$       S�$      �$       S                    `      e       Ue      j       �U�                    `      i       Ti      j       �T�                      �       �        U�       �        t�}��       �        �U�                        �       �        T�       �        P�       �        U�       �        �T�                            p      �       U�      �       ^�      �       �U��             ^      	       �U�	             U                            p      �       T�      �       ]�      �       �T��             ]      	       �T�	             T                   p      �       0�	             0�                  �      �       T                    p      �       U�      �       �U�                    p      �       T�      �       �T�                      p      y       Qy      �       P�      �       �Q�                      p      �       R�      �       Q�      �       �R�                 �      �       U                      �      �       U�      .       V.      7       �U�                      �      �       T�      4       ^4      7       �T�                      �      �       Q�      �       �Q��      2       ]                      �      �       R�      0       \0      7       �R�                  �      7       P                     �      �       U�      .       V.      7       �U�                     �      �       T�      4       ^4      7       �T�                 �      �       t                   �      6       _                 �      �       S                 �      (       ^                 �      (       \                 �      (       V                      @      R       UR      u       Su      v       �U�                     @      R       UR      u       Su      v       �U�                 @      A       u                  @      A       u                   ^      k       P                  c      t       S                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    `       r        Ur       |        �U�                        `       j        Tj       t        Pt       {        U{       |        �T�                       `       r        u�r       x        Tx       {        tx�{       |        �U#�                          �       �       U�      ?       V?      R       �U�R      �       U�      A       V                    �       �        T�       A       �T�                        �              Q      @       QR      �       Q�      �       Q                          �       �       R�      �       S�      R       �R�R      �       R�      A       �R�                          �       &       T&      �       �TR      k       Tk      �       �T�      �       T                      �       M       \R      �       \�      A       \                 ?      E       3�                          T      T       PT      z       p�z      �       p�      ?       s } "��      �       p��      �       p��      �       s } "��      8       Q                   ,      <       4�q      �       6�                         �       �       u���      ?       v��?      R       �U#��R      �       u���      A       v��                          3      T       P�      ?       ]�      �       P�      �       ]�      A       ]                  ,      <       0�                          ?       U�      �       U                             ?       ^�      !       ^!      8       ~�                  �      8       X                   �             X      !       R                  �      8       U                      �       �        U�       �        S�       �        �U�                    �       �        T�       �        �T�                  �       �        U                  �       �        v�                        @      �       U�      �       w �      �       ��}�      �       w                         @      �       T�      �       _�      �       �T��      �       _                                                  @      �       Q�      �       V�      �       �Q��      �       V�      �       �Q��      �       V�      
       �Q�
      �
       V�
      �
       �Q��
      �       V�      �       �Q��      �       ��}�      �       �Q��      �       V�      �       ��}�      �       V�             ��}      5       V5      �       ��}                    @      �       R�      �       �R�                    @      �       X�      �       �X�                       @      �       T�      �       _�      �       �T��      �       _                                      �      �       ]�      �       ]�      �       ]
      �
       ]�
      �       ]�      �       ��}�      �       ]�      �       ��}�      �       ]�             ��}      5       ]5      �       ��}                              �      i       ^i      �       �QO&�Q'�QO&
����      -	       ^-	      
       �QO&�Q'�QO&
���
      �
       ^�
      �
       �QO&�Q'�QO&
����
      �       ^                 Q      g       U                       �      Z       _             _-	      
       _�
      �
       _                       �      Z       S             S-	      
       S�
      �
       S                      b	      e	       Qe	      
       V�
      �
       V                   Z      Z       V-	      b	       V                 �      �       ^                                           �      �       Q�      �       V�      �       V�      �       �Q��      �       V�      	       �Q�
      �
       V�
      �
       �Q��
      �       V�      �       �Q��      �       ��}�      �       �Q��      �       V�      �       ��}�      �       V�             ��}      %       V5      �       ��}                               �      �       \�      �       \�      	       \
      
       \
      �
       U�
      �
       \�
      �
       U�
      �
       \�
      �       \�      %       \5      �       \                                    �      �       ]�      �       ]�      �       ]
      �
       ]�
      �       ]�      �       ��}�      �       ]�      �       ��}�      �       ]�             ��}      %       ]5      �       ��}                	                 �      �       S�      �       ^�      �       S�      �       ^�      �       S�      	       ^
      
       S
      �
       ^�
      }       S}      �       ^�      %       ^5      �       ^                 
      5
       ��}�
����}�
��" $ &�                        r
      
       P
      �
       ��}�      #       ��}�      �       ��}      %       ��}                     
      �
       0��             0�      #       ��}�      �       ��}      %       ��}                    
      �
       0��             0�             ��}                         
      �
       P�
      �
       S�
      �
       P�
      �
       S�      �       S                    �
      �
       P�             P                          �      �       ��}�      �       P�      �       ��}�             ��}5      �       ��}                               $       P$      �       ��}�      �       ��}5      �       ��}                        �             S      �       sp��      �       sp�5      �       sp�                                  a             0�      �       S�      �       ��}#      '       S,      ;       S�      �       0��      �       ��}�      �       ��}�             ��}5      �       ��}                      U      �       ]�      �       ]5      �       ]                            �       V�      �       V5      �       V                 k      �       _                 k      �       _                 k      �       _                  r      �       S                       0       M        0�M       R        PR       \        0�\       _        P                       0       J        0�J       O        QO       R        RR       \        0�\       _        R                          8       E        QE       M        PM       O        p�R       \        P\       ^        q u��                            #        T#       .        T                         -        0�                                  u                     
               P                u #�                      P      {       U{      �       S�      �       �U�                 P      R       u�                 P      R       u�                  [      �       V�      �       0�                      �      F       UF      G       �U�G      k       U                      �      B       TB      G       �T�G      k       T                    �      F       XG      k       X                   �      F       x�#�G      k       x�#�                   �      F       x� G      k       x�                               	       Q	             q`�      F       QG      k       Q                    @      B       TB      G       �T�                    @      F       UF      G       �U�                                p      �       U�      �       S�      �       �U��             S             q�~�             �U�      3       S3      5       �U�                                p             T      �       V�      �       �T��             V             U             �T�      4       V4      5       �T�                      �      �       P�      �       P�      �       P                               p      �       u��      �       s��      �       �U#��             s�             q�~�             �U#�      3       s�3      5       �U#�                    �      �       v�      )       ��                      �             V             U             �T�                      �             S             q�~�             �U�                  �             P                        �      �       U�      �       S�      �       �U��      �       U                       �      �       U�      �       S�      �       �U��      �       U                      �      �       U�      �       S�      �       �U�                  �      �       V                                                                              �             U      $       V$      ?       �U�?      �       V�      �       U�      �       V�      J       �U�J      T       UT      _       V_      �       �U��      �       V�      �       �U��      �       V�      �       U�      �       V�      m       ��~m      �       �U��      �       V�             �U�             U             V      �       �U��      �       V�      �       �U��              V       �        �U��       �        ��~�       �        �U��       !       ��~!      &!       �U�&!      /!       V                                                            �             T      $       S$      ?       �T�?      i       Si      �       ��~�      �       S�      J       �T�J      _       S_      �       �T��      �       S�      �       �T��      �       ��~�      �       �T��      �       S�      �       �T��      �       S�      �       �T��      �       ��~�      �       �T��              S       &!       �T�&!      /!       S                                        �             Q      $       \$      ?       �Q�?      �       \�      �       �Q��      �       \�      �       �Q��      �       \�      �       �Q��              \       &!       �Q�&!      /!       \                                                           �             T      $       S$      ?       �T�?      i       Si      �       ��~�      �       S�      J       �T�J      _       S_      �       �T��      �       S�      �       �T��      �       ��~�      �       �T��      �       S�      �       �T��      �       S�      �       �T��      �       ��~�      �       �T��              S       &!       �T�&!      /!       S                 $      *       3�                                     P      1       w 1      ?       ��~?      /!       w                   .      ]       0�                                   _      {       P7      D       Pz      �       P�      �       P�      	       PC      T       P�      �       P�      �       P�      �       PC       U        P                         �      �       P�      �       V      �       V�      �       V       m        V                                 �      /       0�>      �       ��~      O       0�O      l       ��~l      �       0��      �       ��~�      �       0�       C        ��~C       m        0�                                    �      q       0�q      �       
��      X       0�X      g       Pg      l       Xl      �       0��      �       0��      �       0�       3        P3       C        
��C       m        0�                      �             P      ;       Vm       �        V                           <       S;      f       S�      �       S                           9      f       S�      �       S�             S      �       S�      �       S       �        S                    @      �       \�      �       \                        n      �       P�      �       P�      	       P/      C       P                      e      �       V�      <       \;      f       \                           e      s       Vs      �       ^�      �       T�      �       ^�      <       V;      f       V                    �             P+      <       P                  �             T                  ;      P       0�                                  $       S?      :       S�      �       S�      �       S�      �       S�              S&!      /!       S                                           U      $       V?      :       V�      �       V�      �       V�      �       V�              V&!      /!       V                                  $       s��?      :       s���      �       s���      �       s���      �       s���              s��&!      /!       s��                             �      �       P�      :       ]�      �       ]�      �       ]�      �       P�              ]&!      /!       ]                                           P      $       w ?      :       w �      �       w �      �       w �      �       w �              w &!      /!       w                                            �      �       0��      �       _�             Q             _�      �       Q�      �       0��      Y       ��~]      f       Pj      �       0��      �       R�      �       P�      �       R�      �       ��~�      �       0�&!      /!       0�                      j      �       Q�              Q*!      /!       Q                    �      �       UA      z       U                       �      �       ['      +       1�+      �       [�      �       [                        �      �       [���             [�Z�T��             p �Z�T��      +       p �p�T��                                         ^      i       Si      �       ��~�      �       S�      �       �T�J      _       S�      �       ��~�      m       �T��      �       S�      �       �T�             �T��      �       ��~               �T��       &!       �T�                                                     ^      �       V�      �       U�      �       V�      �       �U�J      T       UT      _       V�      �       V�      �       U�      �       V�      m       ��~�      �       V             U             V�      �       V               V�       �        ��~�       �        �U��       !       ��~!      &!       �U�                                           ^      F       0�F      J       PJ      �       _�      �       0��      �       _�      �       0�J      _       0��      �       _�      m       ��~�      �       _             _�      �       _               _�       �        ��~�       !       ��~                               ^      �       0�J      _       0��      y       0�y      �       P�      �       0�             0��      �       0�               0�                                  >      B       RB      F       _F      �       ��~�      m       ��~�      �       ��~             ��~�      �       ��~               ��~�       &!       ��~                              �      �       ��~Z      _       P�      �       ��~�      �       ��~             ��~�      �       ��~               ��~                                      N      s       0�s      �       ]�      �       ]�      �       0��      m       S�      �       0��      �       4p ��      �       T�      �      	 4��~3��       �        S�       !       S
!      !       S                                �      �       \J      _       \�      m       \�      �       \             \�      �       \               \�       &!       \                            �             P      -       Q-      m       ��~             P               P�       &!       ��~                                     �      �       0��      �       ^�      �       0�J      _       0��      :       0�:      R       PR      m       ^�      �       0�             0��      �       0�               0��       &!       ^                  �      �       Q                    �      .       
 �;      J       
 �                    �      .       Q;      J       Q                    �      .       T;      J       T                   �             0�      .       P                     ]      #       S_      u       S�      )       S}      }       S                               ]      #       V_      l       Ul      u       V�             V             U             V              U       )       V}      }       V                      v      #       ^_      u       ^�      )       ^}      }       ^                       v      y       0�y      #       __      u       0��      )       0�}      }       _                 *      E      % r #���������
��#���������-( �                          �      E       Rp      u       P�             R             R$      )       P                  y      �       1��      #       \                      /      ;       Su      �       S)      �       Sf      }       S                                            /      �       V�      �       U�      �       V�      �       U�      4       V4      8       U8      ;       Vu      �       V)      N       VN      R       UR      �       Vf      j       Uj      p       Vp      t       Ut      }       V                       �      ;       \u      �       \)      �       \f      p       \                      �      ;       ^u      �       ^)      =       ^                      �      �       P�      �       _x      }       P                          �      �       1��      ;       _u      �       _=      _       4~ �_      c       5~ �c      �       4~ �f      p       4~ �                       /      ;       0�u      �       0�)      =       0�p      }       0�                      �             P9      ;       Pu      {       P                     �      �       S�      �       S�       �        S                               �      �       U�      �       V�      �       U�      �       V�      �       U�      �       V�      �       V�       �        V                    �      v       ^�       �        ^                         �      �       s���      �       Q�      �       s���      �       s���       �        s��                    u      �       _�       �        _                         �       ^�      �       ^                     �      �       U�             s��8%�             U                      �      �       t ���            	 s����      }       T�       �        T                    �      �       P�      �       P                    E      N       P�       �        P                         �       \�      �       \                      �      �       _�      �       _�      �       _                      .      5       R5      y      - s��
�� 
��#u  
��t "1$ $ &v� "��       �       - s��
�� 
��#u  
��t "1$ $ &v� "�                        
      =
       U=
      L
       VL
      O
       �U�O
      �       V                        
      (
       T(
      K
       SK
      O
       �T�O
      �       S                      
      /
       Q/
      =
       R=
      �       �Q�                  �      �       P                       
      (
       t��(
      K
       s��K
      O
       �T#��O
      �       s��                          0      k       Uk      x       �U�x      �       U�      �       �U��      �       U                        0      C       TC      N       SN      �       �T��      �       T                          0      k       Qk      x       �Q�x      �       Q�      �       �Q��      �       Q                          0      k       Rk      x       �R�x      �       R�      �       �R��      �       R                              0      k       Xk      x       �X�x      �       X�      �       �h�      �       �X��      �       �h�      �       X                                0      k       Yk      x       �Y�x      �       Y�      �       w �      �       �Y��      �       w �      �       �`�      �       Y                             0      k       3�k      x       Px      �       3��      �       P�      �       P�      �       3��      �       P                     0      N       0�N      k       T�      �       0�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  p      p       Rp      v       �R�                     	      4	       U4	      u	       �U�                       	      +	       T+	      ;	       P;	      u	       �T�                           	      7	       Q7	      `	       S`	      a	       �Q�a	      t	       St	      u	       �Q�                    ?	      D	       PD	      u	       Q                                 �       U�      "       S"      +       �U�+      ~       U~      -       S                               G       TG      k       �T�k      ~       T~      -       �T�                               9       Q9      k       �Q�k      ~       Q~      -       �Q�                                       b       Rb      =       ]=      +       �R�+      ;       ];      >       �R�>      k       ]k      ~       R~      -       �R�                                $       V+      7       V>      w       Vw      ~       t ~      -       V                       5      "       \+      9       \>      k       \~      -       \                                 _       0�_      r       Ps      �       P�      �       P+      ~       0�~      �       P                               �       u���      "       s��"      +       �U#��+      ~       u��~      -       s��                        =      "       ^+      =       ^>      k       ^~      -       ^                        W      �       ]�      �       }�~              ]              }�                    �      �       ]�      �       }�                      �             P             p|�             P                  �             Q                    �      �       ]�      �       }�                      �      �       T�      �       t��      �       T                                      �      �       Q�      �       R�      �       t����      �       R�      �       Q�      �       t��1%Ut��1$�!��      �       Q�      �       R�      �      > t��1%Ut��1$�!2%3t��1%Ut��1$�!2$�!��      �       r q !��      �       Q                    �              ]              }�                      �             P      !       p~�!      (       P                        -       Q                               �       U�      �       V�      �       �U��      �       U                             �       T�      �       �T��      �       T                                    m       Sm      o       u o      z       Sz      |       u |      �       S�      �       S�      �       u                                    m       s� m      o       u #@o      z       s� z      |       u #@|      �       s� �      �       s� �      �       u #@                        9      ?       Q?      C       q`�C      �       Q�      �       Q                �      �       0�                �      �       V                 �      �       s��                          0!      O!       UO!      �!       \�!      �!       U�!      �!       ^#      ,#       \F#      u#       \                                0!      O!       TO!      �"       S�"      �"       �T��"      #       S#      #       �T�#      >#       S>#      F#       �T�F#      u#       S                        0!      O!       QO!      �"       V�"      �"       ]�"      u#       �Q�                    0!      O!       RO!      u#       �R�                    0!      O!       XO!      u#       �X�                                G!      O!       TO!      �"       S�"      �"       �T��"      #       S#      #       �T�#      >#       S>#      F#       �T�F#      u#       S                              P!      k!       P!      �!       P�!      �!       P�!      �"       0��"      #       0�#      #       P#      ,#       PF#      b#       P                      w!      �!       P#      #       Pc#      k#       P                  #      ,#       P                      �!      "       P"      �"       s��"       #       s�                  �!      T"       X                    �!      �"       0��"      �"       1��"      �"       0�                 �!      ""       P                 T!      l!       S                       T!      �!       S#      >#       S>#      F#       �T�F#      u#       S                 �"      �"       S                 �"      �"       S                   '#      >#       S>#      F#       �T�                   '#      >#       S>#      F#       �T�                    �       �        U�       E       �U�                   �       �        U�       E       �U�                  �       E       R                        �       �        Z�       �        Q�       �        Z&      E       Z                    �              S              Z                 �              Q             r                      �       �        0��              P2      E       P                            .        U.       �        �U�                              _        T_       ~        �T�~       �        T                           .        U.       �        �U�                  $       �        R                     M       _        t 8%�_       ~        T~       �        t 8%�                      Q       t        Qt       ~        �T��~       �        Q                                U                                 U                                 u                       �      �       U�      �       S�      �       �U�                    �      �       T�      �       �T�                  �      �       v��                          �             U      b       Sb      h       u�~�h      �       S�      �       �U�                          g       ]h      �       ]                        D      R       0�R      _       V_      c       v�k      �       V                    R      k       \t      �       \                      �      �       U�      �       �U��      �       U                     �      �       U�      �       �U��      �       U                            �      �       Q�      �       \�      �       �Q��      	       \	      	       �Q�	      	       Q                       �      �       T�      �       ]�      	       ]	      	       T                   �      �       0��      	       1�	      	       0�                      �      �       0��      �       s��      	       s�	      	       0�                        �	      �	       U�	      �	       �U��	      �	       U�	      

       �U�                        �	      �	       T�	      �	       �T��	      �	       T�	      

       �T�                            �	      �	       Q�	      �	       S�	      �	       �Q��	      �	       Q�	      	
       S	
      

       �Q�                   �	      �	       0��	      �	       0��	      

       P                    �	      �	       T�	      �	      "  �F      �F     �T4 $0.( �                    �	      �	       T�	      

       �T�                      �	      �	       Q�	      	
       S	
      

       �Q�                    �	      �	       U�	      

       �U�                  �	      

       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                           '       U'      �       �U�                             X       TX      �       �T��      �       T                                               X       QX      y       Sy      z       �Q�z      �       S�      �       �Q��      �       S�      �       �Q��      �       S�      �       �Q��      �       S�      �       �Q��      �       Q                                \      s       Ps      �       Q�      �       P�      �       Q�      �       P�      �       Q�      �       P�      �       Q                      '      X       TX      \       �T��      �       T                    '      X       U�      �       U                            �      Z       UZ             S             �U�      7       S7      L       UL      l       S                        �      9       T9      7       �T�7      L       TL      l       �T�                      �      �       Q7      G       QG      L       P                        �             R      7       �R�7      L       RL      l       �R�                    �             ^      l       ^                   �             ^      l       ^                           �      Z       u��Z             s��             �U#��      7       s��7      L       u��L      l       s��                                  ,      1       �]�Q�p�� 1      5       �]�Q�p�\��5      A       �]�Q�p�\��V��A      P       �]�Q�P�\��V��P      Z       �]�Q�s��\��V��Z      �       �]��\��V���             �\��V��      7       �]��\��V��L      l       �]��\��V��                   �      Z       ~�#��
���7      L       ~�#��
���                      �      �       U�      �       S�      �       �U�                    �      �       T�      �       �T�                  �      �       V                                �      )       U)      2       ^2      D       ��~D      e       ^e      �       ��~�      �       ^�      �&       ��~�&      �&       ^                                                    �             T      2       S2      D       �T�D      e       Se      �       ��~�      $       �T�$      �       ��~�      �       S�      �       �T��      �       ��~�      �        �T��       !       ��~!      )#       �T�)#      ?#       ��~?#      %       �T�%      =%       ��~=%      �&       �T��&      �&       S                    �      )       Q)      �&       ��~                    �      )       R)      �&       �R�                    �      )       X)      �&       �X�                  j&      o&       P                                      %      2       _2      9       w 9      D       ��}D      �       _�      �       w �      <       V<      �       w �      �       V�      �&       w �&      �&       V�&      �&       w                                           %      2       0�D      �       0��      �       0��      �       8�      �       0��      �        V�       !       0�!      #       V)#      ?#       0�?#      �$       V�$      �$       0��$      %       V%      =%       0�=%      �%       Vo&      �&       V�&      �&       0�                                         U      �       0��      �       P�      �       P�      �       P�      �       P$      -       Pg      {       P�      �       P�!      �!       P�"      �"       0��#      �#       P$      %$       PC$      P$       0�                                           \@!      �!       \?#      �#       \�#      C$       \P$      �$       \�$      %       \o&      �&       \                                             �       0��      �        ]@!      �!       0��"      )#       ]?#      �#       ]�#      �#       ]�#      C$       0�P$      �$       0��$      �$       ]�$      �$       0��$      %       0�=%      �&       ]                                         �       0�@!      �!       0�?#      T#       0�T#      r#       
���#      C$       0�P$      �$       0��$      �$       Q�$      �$       0��$      %       0�o&      �&       
���&      �&       Q                                 t      �       Q�      �       P?#      {#       P�#      �#       P�#      �#       Q�$      �$       Po&      u&       Pu&      �&       q��~��&      �&       P                 �      �      
 F�F     �                 �      �       V                 �      �      
 ��F     �                 �      �       V                       $      
 ��F     �                       $       V                 J      g      
 w�F     �                 J      g       V                 �      �      
 ��F     �                 �      �       V                           �        \�"      �"       \                   +       N        0�N       �        Q                        �"      �"       P�"      �"       \=%      o&       \�&      �&       \                    �"      �"       P=%      p%       P                       �"      )#       0�=%      :&       0�:&      T&       1��&      �&       0�                   �%      o&       V�&      �&       V                 �"      �"      
 ��F     �                 �"      �"       V                 �"      �"      
 ��F     �                 �"      �"       V                     i      �      
 �F     ��"      �"      
 �F     �C$      P$      
 �F     �                     i      �       V�"      �"       VC$      P$       V                 �      �      
 k�F     �                 �      �       V                       �      �       S�       �        S!      @!       S�!      �"       S                                 �      �        S!      �!       S�!      �"       S�"      )#       S?#      �#       S�#      C$       SP$      �$       S�$      %       S=%      �&       S                            p       ]!      @!       ]�!      �"       ]                       ]       s�                                ^      m       P�      �       P�      �       P�      �       P!       !       P�!      �!       P"      "       PI"      T"       P                      �      x       \x      �       ]�       �        ]                         �      0       ^0      A       TA      M       ^�      �       ^�       �        ^                 9      ^      
 <�F     �                 9      ]       s�                 m      �      
 B�F     �                  �      �      
 N�F     ��      �      
 N�F     �                  �      �      
 \�F     ��      �      
 \�F     �                   x      �       U�      �       U                  |      �       T                  �       �        0�                            �      �       ��  �      )       ��  �       !       ��  )#      ?#       ��  �$      �$       ��  %      =%       ��  �&      �&       ��                                    �      �       ��~��      �       P�             �       �       ��~��      )       ��~��       !       ��~�)#      ?#       ��~��$      �$       ��~�%      =%       ��~��&      �&       ��~�                                    �      �       U�      <       V<      �       w �      �       V�      )       w �       !       w )#      ?#       w �$      �$       w %      =%       w �&      �&       V�&      �&       w                                 �      e       ^e      �       ��~�      �       ^�      )       ��~�       !       ��~)#      ?#       ��~�$      �$       ��~%      =%       ��~�&      �&       ^                            �      �       0��      )       0��       !       0�)#      ?#       0��$      �$       0�%      =%       0��&      �&       0�                                          �      �       0��      �       P�      e       _e      �       ��~�      $       ��~H�$      �       ��~�      �       _�      �       ��~�      �       ��~H�%      )       0��       !       ��~)#      ?#       ��~�$      �$       ��~H�%      =%       ��~�&      �&       _                                   �      �       U�      �       V�      �       0��      �       v�$      �       0��      �       V�      �       0��      �       w       )       w �       !       0�)#      ?#       0�%      =%       0��&      �&       V�&      �&       w                            �            
 �C     �$      �      
 �C     ��      �      
 �C     ��       !      
 �C     �)#      ?#      
 �C     �%      =%      
 �C     �                           �             ��(  $      �       ��(  �      �       ��(  �       !       ��(  )#      ?#       ��(  %      =%       ��(                                 �      e       _e      �       ��~�             ��~H�$      �       ��~�      �       ��~�       !       ��~)#      ?#       ��~%      =%       ��~                             �      e       ^e             ��~$      �       ��~�      �       ��~�       !       ��~)#      ?#       ��~%      =%       ��~                   H      T       1�T      ]       ��~e      �       ��~�      �       ��~                                   T       
 �T      �       ��}$      �       ��}�             ��}
      �       ��}�       !       ��})#      ?#       ��}%      =%       ��}                            T      T       1�e      �       1��      �       0�$      �       0��      �       0��       !       0�)#      ?#       0�%      =%       0�                           �      �       Y�      �      	 s 8$8&�
      @       Y@      a       ��~a      �      	 s 8$8&�)#      ?#       S                T      T       
 �T      �       V                 T      e       0�                  T      e       0�!      !       0�                               Z      h       Th      l       ^l      �       T�      �       ~�
             T      �       ~��       �        P4#      ?#       P                             T      e       0��      �       0��      �       ]$      �       0��      
       ]
      �       0��       !       0�)#      ?#       0�%      =%       0�                  T      e       0�!      !       0�                                          �      #       0�#      e       Pe      �       _�      �       P�      �       _�              [             0�$      �       _�      
       P
      �       _�       !       _)#      ?#       _%      -%       _-%      =%       [                                           U             ��~$      �       ��~�      �       ��~�       !       ��~)#      ?#       ��~%      =%       ��~                    �      �       S�      
       S                 �      �       V                 �      �       Q                 �      �       8                        �
      �
       U�
      �       S�      �       �U��      �       U                       �
      �
       U�
      �       S�      �       �U��      �       U                  �
      �       V                  �
      �
       U                    �      �       U�      Z       �U�                   �      �       U�      Z       �U�                  �      Z       Z                     �      �       0��             U*      O       U                       �      �       S�      �       R�      �       P�      O       R                                �      �       P�      �       u��      �       P�      �       R�             P*      4       P7      D       PO      U       P                     �             0�      *       u�#�*      9       0�9      O       q�#�O      Z       0�                        �      �      	 y ������             0�      #       [#      *       u *      O      	 y �����                      �      �       X�      *       X9      O       X                          *       U*      �       �U�                          k       Tk      �       �T�                         *       U*      �       �U�                        �       Y                           *       0�*      k       Xn      �       X                           `       R`      c       Pc      �       R                                    7       P7      :       x�:      c       Pc      f       Rf      m       Pn      t       Pw      �       P                         m       0�n      y       0�y      �       q�#�                      *      ?       UV      k       Uy      �       U                 �             U                 �      �       U                    �      �       P�      �       u                     �+      ,       U,      &,       P                                                        �+      $,       T$,      \,       Q\,      h,       qy�h,      s,       Q�,      �,       Q�,      �-       �T��-      �-       Q�-      �-       R�-      K.       �T�K.      �.       Q�.      �.       R�.      4/       �T�4/      �/       Q�/      �/       R�/      �0       �T��0      �0       qy��0      G1       QG1      P1       RP1      �1       �T��1      �1       Q�1      w4       �T�                    �+      �+       Q�+      w4       �Q�                                        �+      !,       R!,      v,       \v,      �,       �R��,      H-       \H-      �-       �R��-      z/       \z/      �0       �R��0      �2       \�2      �2       �R��2      23       \23      �3       �R��3      �3       \�3      w4       �R�                        �+      ,       X,      �,       ]�,      �,       �X��,      w4       ]                                       ,      !,       R!,      v,       \v,      �,       �R��,      H-       \H-      �-       �R��-      z/       \z/      �0       �R��0      �2       \�2      �2       �R��2      23       \23      �3       �R��3      �3       \�3      w4       �R�                        �,      �,       0��,      .-       P.-      �-       ~�~�23      �3       ~�~�                           \,      l,       p�l,      s,       T�/      �/       P�/      z0       \�0      �0       p��0      �0       T                              �+      ,       0�,      v,       V�,      �,       V�,      �,       }� �,      �-       _�-      0       V�0      23       V23      �3       _�3      �3       V                       v,      v,       PA.      K.       6��2      �2       P�2      �2       	���2      �2       3��3      �3       6�r4      w4       S                    L-      �-       V23      �3       V                    L-      �-       \23      �3       \                    �3      �3       P�3      �3       P                  .      .       U                  �.      �.       U                 �.      �.       U                 0      u0       }�                      0      �0       �Q��3      �3       �Q��3      w4       �Q�                   0      �0       V�3      �3       V�3      r4       V                  z0      �0       \�3      r4       \                  H0      u0       Q                              0      �0       0��0      �0       P�0      �0       S�0      �0       0��3      �3       6��3      �3       P�3      h4       Sh4      q4       Pq4      r4       S                 H0      n0       Q                 H0      n0       ��}�                  m1      {1       U                 �1      �1       U                 �1      �1       U                    �'      �'       U�'      �'       \                        �'      �'       T�'      �(       V�(      �(       �T��(      �+       V                    �'      (       Q(      �+       �Q�                                        �'      �'       R�'      {(       ^{(      �(       �R��(      !*       ^!*      +       �R�+      +       ^+      �+       �R��+      �+       ^�+      �+       �R��+      �+       ^�+      �+       �R��+      �+       ^�+      �+       �R�                                            �'      3(       X3(      �(       ]�(      �(       �X��(      	)       X	)      )       ])      ;)       X;)      �)       ]�)      *       X*      +       ]+      .+       X.+      �+       ]�+      �+       X�+      �+       ]�+      �+       X                                        �'      �'       R�'      {(       ^{(      �(       �R��(      !*       ^!*      +       �R�+      +       ^+      �+       �R��+      �+       ^�+      �+       �R��+      �+       ^�+      �+       �R��+      �+       ^�+      �+       �R�                                           �'      3(       X3(      �(       ]�(      �(       �X��(      	)       X	)      )       ])      ;)       X;)      �)       ]�)      *       X*      +       ]+      .+       X.+      �+       ]�+      �+       X�+      �+       ]�+      �+       X                              �(      )       \�)      �)       \�)      �)       S�)      �*       \�*      �*       [�*      �+       \�+      �+       S�+      �+       \                        �(      �(       |��(      	)       Q�*      �*       P�*      +       S�+      �+       S                                          �'      {(       0��(      )       0�)      )       P)      p)       0�p)      )       P)      �)       0��)      �)       P�)      u*       0�u*      �*       P�*      �*       S�*      �*       P�*      +       0�+      +       P+      �+       0�                  (      4(      
 �F     �                  (      3(       U                  A(      b(      
 �F     �                  A(      a(       U                        �)      \*       _�*      �*       _+      �+       _�+      �+       _                        �)      \*       ��;  �*      �*       ��;  +      �+       ��;  �+      �+       ��;                          �)      \*       �;  �*      �*       �;  +      �+       �;  �+      �+       �;                          �)      \*       V�*      �*       V+      �+       V�+      �+       V                                �)      �)       \�)      �)       S�)      \*       \�*      �*       \+      �+       \�+      �+       \�+      �+       S�+      �+       \                      �)      !*       	��+      +       	�� +      8+       ^�+      �+       	���+      �+       	��                                     �)      �)       \�)      �)       S�)      \*       \�*      �*       \�*      �*       S+      ;+       \;+      B+       SB+      I+       PI+      �+       S�+      �+       S�+      �+       \�+      �+       S�+      �+       \                                 �)      �)       \�)      \*       S�*      �*       S�*      �*       T+      ?+       S?+      �+       T�+      �+       t��+      �+       \�+      �+       T�+      �+       S                   H*      \*       R�+      �+       0�                   �)      H*       _+      8+       _�+      �+       _�+      �+       _                   �)      H*       \+      8+       \�+      �+       S�+      �+       \                    *      (*       P/+      8+       P                    �4      �4       U�4      �4       S                                �4      �4       T�4      '6       _76      D6       _D6      W6       Qz6      �6       _7      7       Q7      08       _<8      �@       _                        �4      �4       Q�4      76       �Q�76      D6       QD6      �@       �Q�                                                                      �4      �4       R�4      '6       ^'6      76       �R�76      _6       ^_6      z6       �R�z6      �6       ^�6      �6       �R��6      �6       ^�6       7       �R� 7      �7       ^�7      �7       �R��7      08       ^08      <8       �R�<8      m:       ^m:      ;       �R�;      ;       ^;      �<       �R��<      �<       ^�<      �=       �R��=      r>       ^r>      �?       �R��?      �?       ^�?      �?       �R��?      �?       ^�?      �?       �R��?      2@       ^2@      �@       �R��@      �@       ^                        �4      B5       XB5      q6       Vq6      z6       �X�z6      �@       V                        �;      �;      	 r 8$8&�<      3<      	 r 8$8&�r>      v>      	 r 8$8&��@      �@      	 r 8$8&�                    U<      ^<       r 
��v8#��
��7��>      �>       r 
��v8#��
��7�                          H6      W6       T7      7       T,9      :9       P:9      �9       S^>      r>       P                        �;      <       T<      <       t�<      �<       Tr>      �>       T}@      �@       T                             �;      �;       0��;      <       Z<      <       q�<      3<       Q3<      P<       Zr>      v>       Q}@      �@       0�                        �;      �;       y 1$��;      �<       Xr>      �>       X}@      �@       X                                                                   �4      '6       ^'6      76       �R�76      _6       ^_6      z6       �R�z6      �6       ^�6      �6       �R��6      �6       ^�6       7       �R� 7      �7       ^�7      �7       �R��7      08       ^08      <8       �R�<8      m:       ^m:      ;       �R�;      ;       ^;      �<       �R��<      �<       ^�<      �=       �R��=      r>       ^r>      �?       �R��?      �?       ^�?      �?       �R��?      �?       ^�?      �?       �R��?      2@       ^2@      �@       �R��@      �@       ^                       �4      B5       XB5      q6       Vq6      z6       �X�z6      �@       V                                   �7      �7       ^&:      5:       Pm:      ;       ^;      �<       ^�<      �=       ^F>      ^>       Qr>      �?       ^�?      �?       ^�?      �?       ^2@      �@       ^                               �4      '6       ]76      h6       ]z6      �6       ] 7      08       ]<8      �8       ]�8      �8       v8�9      ^>       ]r>      �@       ]                    �4      s6       \z6      �@       \                  �@      �@       P                    ,?      _?       R�?      �?       R                  W5      m5       U                   /=      E=       Uu@      }@       U                  �:      �:       U                  �;      �;       U                    =      "=       Um@      u@       U                      @      j       Uj      �       S�      �       �U�                      @      J       TJ      �       ]�      �       �T�                        @      c       Qc      �       V�      �       |��      �       �Q�                  �      �       R                  j      �       U                 �      �       U                 �      �       T                        �       1       U1      7       u�7      �       U�      �       u��      �       U                         �              0�      4       P7      a       Pk      �       P�      �       
��                       �       �        0��       b       Xk      �       X�      �       0��      �       1�                                d        Ud       h        u�h       �        U�       �        u��       �        U                           "       K        0�K       `        Ph       �        P�       �        q ��       �        P�       �       
 ��������                              "        0�"       �        Y�       �        Y�       �        0��       �        1�                        p      �       U�      �       S�      �       �U��      �       U                      p      �       T�      �       �T��      �       T                   �      �       Q�      �       Q                          �      �       V�      �      
 q 1%q "#��      �       V�      �       V�      �      
 q 1%q "#�                   �      �       �����      �       ����                     �      �       u�      �       s�      �       u                                    U      5       S5      6       �U�                               U                      �             U      0       u�0      Y       U                       �             0�      '       P0      W       PX      Y       0�                      `      �       U�      �       u��      �       U                       `      �       0��      �       P�      �       P�      �       0�                      �      F       UF      G       �U�G      k       U                      �      B       TB      G       �T�G      k       T                    �      F       XG      k       X                   �      F       x� G      k       x�                    �      F       x�G      k       x�                              	       Q	             q`�      F       QG      k       Q                    @      B       TB      G       �T�                    @      F       UF      G       �U�                      p      �       U�      �
       S�
      �
       �U�                  2
      �
       \                                   �      �       0��      "	       \"	      '	       |�'	      @	       \_	      a	       0�a	      s	       ]s	      �	       }��	      �	       ]�	      �	       0��	      �	       ]�	      �	       }��	      �	       ]2
      6
       0�6
      �
       ]                         _	      w	       \w	      �	       |H��	      �	       \�	      �	       |H��	      2
       \                  �      �
       V                            �             U      h       \h      o       �U�o             \      �       �U��      �       \                    �      6       T6      �       �T�                          �      �       Q�      �       V�      �       �Q��      �       V�      �       �Q�                      �      �       R�      y       ^y      �       �R�                      	      y       ^y      `       �R�o      n       �R��      �       �R�                          	      �       V�      `       �Q�o      n       �Q��      �       �Q��      �       V�      �       �Q�                      	      6       T6      `       �T�o      n       �T��      �       �T�                      	             U      `       \o      n       \�      �       \                       v             0�o      �       0��      n       0��      �       0�                         4      6       0�6      p       _p      v       Uv      `       _o      n       _�      �       _                                      4      6       T6      V       t�V      p       Tp      t       t�t      v       Tv      �       V�             So      �       S�      �       V�      -       S-      `       V`      n       S�      �       S�      �       V�      �       S                    y      `       ^o      n       ^�      �       ^                                       v      �       V�             So      w       Sw      �       V�      �       S�      -       V-      T       ST      `       V`      n       S�      �       S�      �       V�      �       S                            y              0�       )       P)      `       0�o      <       0�<      T       PT      n       0��      �       0�                          �      �       U�             S             �U�             S             �U�                      �      �       T�      �       U�             �T�                    �      �       P             P                                �             U      ,       S,      ]       �U�]      �       S�      �       �U��      �       S�             �U�      �       S                                  �      �       T�      J       V]      	       V�      �       V      !       V�             V             �T�      |       V�      �       V                            �             Q      V       \V      ]       �Q�]             \             �Q�      �       \                 �      �       ��]  �                                                 P]      q       Pu      �       P�      �       _�             P      �       _      9       P]      |       P|      �       _�      �       _                  �      �       P                               ,      J       S�      �       ^�      �       S/      E      
 s�Hq "�i      �       ^�             S|      �       ^�      �       ^                            X       ]]             ]      �       ]                 �      �       \                 �      �       \                        C       1��      �       1�                        C       S�      �       S                        C       V�      �       V                    3      F       [F      �       ���      �       s�#S�                         #       Z#      �       w                    -      C       _�      �       _                      �&      )'       Y)'      :'       y�:'      O'       Y                     '      %'       Q.'      :'       q�:'      ?'       Q                  �&      O'       P                  �&      '       X                        ��      '�       U'�      x�       Sx�      ��       �U���      ��       S                        ��      '�       T'�      ��       �T���      �       T�      ��       �T�                                ��      Ϋ       QΫ      '�       ]'�      ��       �Q���      ��       Q��      >�       ]>�      T�       �Q�T�      ��       ]��      ��       �Q�                          ��      '�       R'�      ��       �R���      ��       R��      �       ^�      ��       �R�                                      ��      '�       X'�      e�       \e�      o�       �X�o�      x�       \x�      ��       �X���      ��       \��      ��       X��      >�       �X�>�      J�       \J�      ��       �X���      ��       \                              ��      '�       Y'�      ��       �Y���      ��       Y��      >�       _>�      T�       �Y�T�      ��       _��      ��       �Y�                                     ��      x�       0�x�      ��       2���      ݮ       0�ݮ      �       P�      (�       V(�      8�       P8�      >�       V>�      O�       0�O�      T�       6�T�      ]�       P]�      ��       V��      ��       0�                ��      ��       �                    ��      ��       T��      �       t 2$s�
"�������      ��       �T2$s�
"������                ��      ��       S                ��      ��       ��~�                      ��      ��       ����      �       P�      ��       V��      ��       0�                    ��      ��       s���      �       \�      ��       ��~                   ��      ��       T��      ��       t���      ��       t���      ��       t���      ��       t.���      ��       | 1$| "4$s�
"#6�                    �      >�       \T�      ��       \                	ī      ī       Y                
ī      ī       r @B$ $0.�                         ī      e�       � o�      x�       � ��      ��       � >�      T�       � ��      ��       �                              ī      '�       X'�      e�       \o�      x�       \��      ��       \>�      J�       \J�      T�       �X���      ��       \                       ī      Ϋ       QΫ      2�       ]6�      e�       ]J�      T�       ]                     ī      Ϋ       TΫ      �       Q�      '�       t 2$u�
"������                           ī      '�       U'�      e�       So�      x�       S��      ��       S>�      T�       S��      ��       S                    �      �      H q2$u�
"��H$q2$u�
"#��@$!q2$u�
"#��8$!q2$u�
"#��!��      $�      � t 2$u�
"�����#2$u�
"��H$t 2$u�
"�����#2$u�
"#��@$!t 2$u�
"�����#2$u�
"#��8$!t 2$u�
"�����#2$u�
"#��!�                          q�      6�       ]o�      x�       ]��      ��       ]>�      J�       ]��      ��       ]                    |�      Ϭ       V��      ��       V                        �      .�       Po�      w�       P��      ��       P>�      J�       P                          ī      '�       0�'�      !�       5��~��;�      e�       5��~��o�      x�       5��~����      ��       5��~����      ��       5��~��                                      D�      X�       PX�      [�       V[�      j�       Pj�      |�       VϬ      �       P�      �       V�      �       P�      e�       Vo�      o�       Vo�      x�       2���      ��       V>�      E�       V                   ܫ      ܫ      
 q2$u�
"�ܫ      �       q2$u�
"#��      '�       t 2$u�
"�����#2$u�
"#�                                      �L      �M       U�M      DN       VDN      MN       �U�MN      nN       UnN      �N       V�N      O       UO      qQ       VqQ      �Q       U�Q      �R       V�R      �R       U�R      �S       V                                        �L      �L       T�L      �M       S�M      MN       �T�MN      ZN       SZN      dN       �T�dN      nN       TnN      P       SP      (Q       �T�(Q      �Q       S�Q      NR       �T�NR      �R       S�R      �S       �T�                              �L      !M       Q!M      HN       ]HN      MN       �Q�MN      _N       ]_N      dN       �Q�dN      nN       QnN      �S       ]                              �L      7M       R7M      JN       ^JN      MN       �R�MN      aN       ^aN      dN       �R�dN      nN       RnN      �S       ^                          �L      �M       X�M      FN       \FN      MN       �X�MN      nN       XnN      �S       \                                    �L      /N       Y/N      MN       �Y�MN      �N       Y�N      WO       �Y�WO      [P       Y[P      (Q       �Y�(Q      hQ       YhQ      NR       �Y�NR      �R       Y�R      �S       �Y�                   �L      �L       u� dN      nN       u�                        �L      �L       u� 7M      7M       T7M      HM       t�HM      M       TdN      nN       u�                                   M      RM       [`M      hM       { 
���hM      /N       [MN      dN       [nN      �N       [WO      �O       [P      [P       [(Q      �Q       [NR      QR       [                       M      M       p 8$z��!
���M      hM       z��8$z��!
���hM      nM       q 8$p��!
���nM      qM       r 8$p��!
���qM      M       p��8$p��!
���                          �M      N       q 
���nN      rN       q 
���WO      dO       q 
���P      /P       q 
���(Q      ,Q       q 
���                                        �M      /N       z �8$u �!
���nN      �N       z �8$u �!
����N      �N       z �8$����!
����N      WO       ����8$����!
���WO      �O       z �8$u �!
����O      P       z �8$����!
���P      [P       z �8$u �!
���(Q      ]Q       z �8$u �!
���]Q      hQ       z �8$����!
���hQ      �Q       ����8$����!
���NR      �R       z �8$����!
����R      �R       ����8$����!
���                                 �L      "N       0�"N      /N       QMN      JP       0�JP      dP       QvP      vP       Q(Q      �Q       0��Q      �Q       QNR      zR       0�zR      �R       Q�R      �R       0�                                    �L      &N       0�&N      /N       RMN      RP       0�RP      dP       RvP      vP       RvP      yP       r q �yP      �P       S(Q      �Q       0��Q      �Q       RNR      �R       0��R      �R       R�R      �R       0�                        �M      �M       P�M      �M      / ��4�H0H%�$!0)( 8/�������MN      YN       PYN      dN      / ��4�H0H%�$!0)( 8/�������                      �O      �O       0��O      P       PNR      VR       0�                            �O      �O       q ��8$p��!
����O      �O       u 8$p��!
����O      �O       u 8$��1��!
����O      �O       q ��8$��1��!
����O      �O       UNR      VR       q ��8$��1��!
���                      �N      O       0�O      WO       Q�R      �R       Q                    �N      WO       T�R      �R       T                             �N      O       p 8$q��!
���O      
O       q��8$q��!
���
O      O       ��2��8$��1��!
���.O      2O       { ��8${��!
���2O      5O       p 8${��!
���5O      IO       { ��8${��!
����R      �R       { ��8${��!
���                     vP      (Q       ���Q      NR       ���R      �S       ��                     vP      (Q       \�Q      NR       \�R      �S       \                     vP      (Q       ^�Q      NR       ^�R      �S       ^                     vP      (Q       ]�Q      NR       ]�R      �S       ]                   vP      yP       r q �yP      �P       S                         vP      (Q       V�Q      NR       V�R      �R       V�R      �R       U�R      �S       V                               �P      �P       P�P      �P       P�Q      �Q       P�Q      �Q       ���Q       R       0� R      R       P�R      �R       PtS      ~S       0�                	       vP      �P       v�P      (Q       _�Q      NR       _�R      �S       _                     �P      (Q       S�Q      NR       S�R      �S       S                        �Q      �Q       Z�R      gS       ZgS      ~S       ��~S      �S       Z                      R      !R       P!R      $R       qy�$R      FR       v#�
���                 R      FR       R                         R      !R      
 p r #3%�!R      $R      
 qyr #3%�$R      -R       v#�
��r #3%�-R      4R       P4R      FR       v#�
��r #3%�                  'R      FR       Q                   �R      gS       Y~S      �S       Y                  �R      tS       V~S      �S       V                      �R      hS       0�hS      tS       PtS      tS       0�~S      �S       0�                                      �R      #S       P-S      0S       P0S      gS       q~S      �S       P�S      �S       q�S      �S       P�S      �S       q�S      �S       P�S      �S       q�S      �S       P�S      �S       q                        S      S       t 
���S      #S      
 v�
���-S      gS      	 q �
���~S      �S      	 q �
���                     �R      -S       v-S      gS       Q~S      �S       Q                  ES      gS       T                        �S      �T       U�T      U       SU      'U       �U�'U      +U       S                      �S      T       TT      �T       _�T      �T       ��T      �T       ~��T      �T       ��T      �T       _'U      +U       _                    �S      /T       Q/T      +U       �Q�                        �S      �T       R�T      U       \U      'U       �R�'U      +U       R                        �S      T       XT      U       ]U      'U       �X�'U      +U       ]                        �S      �T       Y�T      �T       v��T      'U       �Y�'U      +U       Y                       �S      �T       0��T      �T       P�T      U       P'U      +U       0�                    T      �T       X'U      +U       X                    kT      �T       0�'U      +U       0�                 �S      �S       u#                 �S      �S       u#                 �S      �S       u#                 �S      �S       u#
                 �S      �S       u#                	 �S      �S       u#                  �T      �T       T                 �T      �T                               �%      �&       U�&      '(       �U�'(      @(       U@(      v(       �U�                            �%      d'       Td'      �'       T�'      (       T'(      P(       TP(      Z(       t�Z(      _(       T_(      g(       t�g(      v(       T                          �%      &       Q&      �&       S�&      '(       ��'(      1(       S1(      v(       ��                                �%      �&       R�&      �&       [�&      �&       �R��&      �&       R�&      �&       Z�&      �'       _�'      '(       _'(      @(       R@(      v(       _                        �%      �&       X�&      '(       �X�'(      @(       X@(      v(       �X�                    �%      �%       Y�%      v(       �Y�                             	&      �&       y�&      �'       [�'      (       [(      (       S(      '(       ['(      @(       y@(      v(       [                         	&      �&       y�&      �'       ���'      '(       ��'(      @(       y@(      v(       ��                        &      R&       QR&      �&       u#�
����&      �&       �U##�
���'(      @(       Q                                 &      9&      	 p �
���9&      �&      
 u�
����&      �&        
����&      �&       } 
����&      �'      	 w �
����'      '(      	 w �
���'(      6(      	 p �
���6(      @(      
 u�
���@(      v(      	 w �
���                       &      R&       u"��q �R&      �&       u"��u#�
����&      �&       �U#"���U##�
���'(      @(       u"��q �                         �&      �&       } 
����&      �'       ]�'      �'       }��'      �'       ]�'      '(       ]@(      v(       ]                              �&      �&       0��&      `'       X`'      �'       R�'      �'       X�'      (       X%(      '(       X@(      S(       XS(      _(       __(      v(       X                   	&      �&       y '(      @(       y                       	&      =&       Z=&      �&       y'(      @(       Z                    �%      �&       Y'(      @(       Y                                �&      �&       0��&      ,'       P,'      .'       Q9'      t'       Pt'      v'       Uz'      �'       P�'      �'       Y�'      �'       P�'      '(       P@(      v(       P                               �&      )'       [)'      `'       S`'      l'       Ql'      n'       q�n'      �'       Q�'      (       [(      (       S@(      n(       [n(      v(       S                          <'      E'      	 ~ �����'      �'       v 3$z "��'      (       ^(      (       Zn(      v(      	 ~ ����                            �#      $       U$      �$       �U��$      �$       U�$      �%       �U��%      �%       U�%      �%       �U�                          �#      �$       T�$      �$       T�$      �%       T�%      �%       Z�%      �%       T                            �#      ]$       Q]$      �$       �Q��$      �$       Q�$      �%       �Q��%      �%       Q�%      �%       �Q�                              �#      I$       RI$      L$       r 7�L$      w$       Rw$      �$       �R7��$      %%       R%%      �%       X�%      �%       R�%      �%       �R7�                            �#      ?$       X?$      �$       �X��$      �$       X�$      �%       �X��%      �%       X�%      �%       �X�                    �#      �#       Y�#      �%       �Y�                             �#      �#       zI$      �$       Y�$      �%       Y�%      �%       Q�%      �%       Y�%      �%       z�%      �%       P                   �#      �#       z�%      �%       z                      �#      7$       Y�$      �$       Y�%      �%       Y                     �#      �#      	 p �
����%      �%      	 p �
����%      �%      
 u�
���                   �#      �#       u"��y ��%      �%       u"��y �                              w$      �$       [�$      �$       {��$      �$       [�$      �%       [�%      �%       {��%      �%       [�%      �%       [                   �#      �#       z �%      �%       z                       �#      �#       [�$      �$       [�%      �%       [                      �#      n$       Z�$      %       Z�%      �%       Z                      w$      �$       Y�$      �$       P�%      �%       P                  �$      �$       y 3$p 3$s "�                         �$      %%       Y%%      R%       Q�%      �%       q��%      �%       Y�%      �%       Q                  %%      Z%       S                                    �$      %%       0�%%      5%       U5%      :%       P:%      <%       UE%      N%       PN%      Z%       Uv%      �%       U�%      �%       u 8$��%      �%       U�%      �%       0��%      �%       U                      #      h#       Qh#      �#       �Q��#      �#       Q                      #      V#       PV#      ^#       Y^#      {#       p�{#      �#       t #��#      �#       Y                 #      �#       u                        `Z      �Z       U�Z      [       S[      [       �U�[      �]       S                        `Z      �Z       T�Z      �Z       T[      V[       T�[      \       T                            `Z      �Z       Q�Z      [       V[      [       �Q�[      �[       V�[      \       Q\      �]       V                      4[      �[       Q\      �\       Qc]      �]       Q                       h[      ~[       q\      A\       qk\      }\       qc]      s]       q                          m[      ~[       Z\      7\       Z7\      A\       qk\      �\       Zc]      �]       Z                         �Z      �Z       u��Z      �Z       U�Z      [       ]�\      �\       ]�\      �\       U                  �\      c]       ^                    �\      �\       P�\      c]       _                 �\      c]       s��                 �\      c]        
���                          �Z      �Z       P�Z       [       \ [      [       P�\      �\       P�\      c]       \                		 �Z      �Z      
 t2$u�
"��Z      �Z       t2$u�
"#�                    �]      �]       U�]      �]       �U�                    �]      �]       T�]      �]       �T�                      �]      �]       Q�]      �]       R�]      �]       �Q�                      �*      �*       U�*      +       S+      +       �U�                 �*      �*       u�                        �]      �]       U�]      E^       SE^      O^       �U�O^      �a       S                          �]      �]       T�]      �]       Q�]      F^       VF^      O^       �T�O^      �a       V                                                   �]      �]       P�]      ^       0�O^      �^       0��^      �^       P_      2_       P3_      H_       PM_      e_       Pf_      j_       Pt_      �_       0��_      �_       P�_      �_       P�_      �_       P�_      �_       0��_      `       P�`      �`       0� a      a       Pa      3a       P4a      ?a       P                      [^      a^       Pa^      M_       ]�_      �a       ]                     `      `       Q`      `       q�`      `       | #�`      �`       | #��a      �a       | #�                      `      1`      	 p  $ &�1`      �`      , | �H0H%�$!0)( 8/�� $ &��a      �a      , | �H0H%�$!0)( 8/�� $ &�                      #`      q`      	 q �����q`      �`      . | #�H0H%�$!0)( 8/��������a      �a      	 q �����                  `      �`       Q                      �^      �^       P�^      M_       _�a      �a       _                      �^      �^       P�^      �^       \�a      �a       \                      �^      �^       P�^      �^       ^�a      �a       ^                   �^      �^       ^�^      M_       ^                         @      X@       UX@      d@       Sd@      j@       �U�j@      (A       S                  @      "@       u�                        @      X@       u��X@      d@       s��d@      j@       �U#��j@      (A       s��                     D@      X@       Pj@      ~@       P�@      A       P                 j@      �@       s��                     �@      �@       0��@      �@       V�@      �@       \�@      �@       V                 �@      (A       s��                                            ��      �       U�      "�       S"�      4�       �U�4�      �       S�      ��       �U���      8�       S8�      ��       ����      ��       �U���      �       S�      O�       �U�O�      ��       S��      ��       �U���      А       SА      ^�       �U�                              �      "�       V4�      �       V��      �       V�      �       VO�      ��       V��      ؐ       V:�      I�       V                                  �      "�       P"�      3�       _3�      ?�       P?�      _�       __�      �       P�      ��       _��      ��       P��      ��       _��      ��       P                      W�      �       ^��      ��       ^��      �       ^                              P�      [�       p } "�[�      �       | } "���      @�       | } "�@�      l�       ��} "���      �       | } "�ߏ      �       | } "�O�      ��       | } "�                       ��      @�       | } "�@�      l�       ��} "�ߏ      �       | } "�O�      ��       | } "�                           ��      ��       Vߏ      �       V�      �       VO�      ��       VА      ؐ       V:�      I�       V                               ��      8�       S8�      ��       ����      ��       �U�ߏ      �       S�      O�       �U�O�      ��       S��      ��       �U�А      ^�       �U�                      ��      ��       ^ߏ      ��       ^А      ^�       ^                        ��      ܌       p 
���܌      ��      
 ��~�
���ߏ      ��      
 ��~�
���А      ^�      
 ��~�
���                            q�      }�       0�}�      č       Tč      ��       ���      �       ��W�      ��       0�А      5�       ��:�      Y�       ��                           ��      �       0��      ��       P��      ��       ��ߏ      �       ���      �       0��      ��       ��А      ^�       ��                                               ��      ҍ       0�ҍ      �       P�      ��       _ߏ      �       0��      ��       ����      �       0��      �       _�      O�       ��O�      z�       0�z�      ��       P��      ��       ��А      �       _�      �       ���      :�       V:�      ?�       _?�      I�       ��I�      ^�       V                    �      @�       0�O�      ��       0�                  q�      }�       0�W�      ��       0�                    ��      ��       P��      ��       p�}���      ��       R                              ڍ      �       0��      y�       \��      ��       \�      �       \А      ސ       \ސ      :�       ]I�      ^�       ]                              �      �       p ���      )�      	 �����)�      ��       ]��      Ď       p ��Ď      ʎ       } ��ێ      ��       ]:�      I�       ]                    ώ      Ҏ       s p �Ҏ      ێ       ]                  �      *�       0�                 ��      ��       s��                 ��      �       | } "�                   ��      ߏ       V��      А       V                   ��      ߏ       S��      А       S                    �      ߏ       ]��      А       ]                      ��      �       p 
����      ߏ       ^��      А       ^                         �      N�       0�N�      R�       PR�      r�       Rr�      ʏ       ��~Տ      ߏ       0���      А       ��~                    ��      ��       0���      ��       P                      ��      ��       P��      ��       r �8$8&���      ��       r p "�8$8&p "���             Q                 ��      А       s��                        �0      �0       U�0      �1       S�1      �1       �U��1      53       S                    �0      �0       T�0      53       �T�                        �0      �0       Q�0      �1       _�1      �1       �Q��1      53       _                        �0      �0       R�0      �1       ]�1      �1       �R��1      53       ]                                �0       1       X 1      �1       \�1      �1       �X��1      �1       \�1      �1       X�1      m2       \m2      �2       X�2      53       \                 �0      �0       u�                  �0      �0       P                                   �0      �0       R�0       1       T�1      �1       T�1       2       X 2      T2       ��T2      a2       Ta2      m2        v 1$#������"�m2      �2       T�2       3       T 3      53        v 1$#������"�                   �0      �0       U�0      �0       Q                           �0      �0       t q "��0       1       Q�1       2       Q 2      a2       w m2      �2       Q�2      �2       w                         �0      1       P1       1       V�1      �1       P�1      53       V                    �0      �1       ^�1      53       ^                   31      �1       S�1      �1       S                          �f      �f       U�f      �f       s�|��f      �f       �U��f      g       Sg      g       s�|�                            �f      �f       T�f      �f       Q�f      �f       V�f      �f       �T��f      �f       Q�f      g       V                    �f      �f       Q�f      g       �Q�                      �f      �f       P�f      �f       P�f      g       P                   �f      �f       Sg      g       S                   �f      �f       u���f      �f       S                        0      B0       UB0      G0       PG0      p0       �U�p0      �0       P                          0      70       T70      k0       Vk0      p0       �T�p0      �0       T�0      �0       V                      0      ?0       Q?0      p0       �Q�p0      �0       Q                      J0      S0       PS0      j0       Sj0      p0       P                    $0      70       xtmv�70      G0       Tp0      �0       xtmh�                    +0      m0       \w0      �0       \                    20      o0       ]~0      �0       ]                              �;      �;       U�;      �;       V�;      �;       �U��;      9<       V9<      @<       �U�@<      �<       V�<      �<       �U�                              �;      �;       T�;      �;       Q�;      �;       S�;      �;       �T��;      8<       S8<      @<       �T�@<      �<       S                 .<      @<       8�                      �;      �;       \�;      ;<       \@<      �<       \                 �<      �<       0�                  H<      �<       } 
���                     �;      �;       0��;      �<       0��<      �<       V                            �a      �a       U�a      �a       S�a      �a       �U��a      �a       S�a      �a       q�x��a      �a       �U�                              �a      �a       T�a      �a       Q�a      �a       V�a      �a       �T��a      �a       V�a      �a       U�a      �a       �T�                  �a      �a       P                           �a      �a       u���a      �a       s���a      �a       �U#���a      �a       s���a      �a       Q�a      �a       �U#��                            Pe      ke       Uke      ue       Sue      we       �U�we      �e       S�e      �e       q�z��e      �e       �U�                              Pe      _e       T_e      ke       Qke      ve       Vve      we       �T�we      �e       V�e      �e       U�e      �e       �T�                  le      �e       P                           Pe      ke       u��ke      ue       s��ue      we       �U#��we      �e       s���e      �e       Q�e      �e       �U#��                      0A      gA       UgA      7B       \7B      :B       �U�                  OA      5B       V                     OA      gA       u��gA      7B       |��7B      :B       �U#��                     TA      {A       S{A      �A       s`��A      �A       S                  bA      �A       ]                     �A      �A       S�A      �A       sh��A      �A       S                  �A      B       ]                        �a      !b       U!b      6b       ^6b      9b       �U�9b      Je       ^                          �a      b       Tb      !b       Q!b      /b       S/b      9b       �T�9b      Je       S                    b      2b       \9b      Je       \                      Zb      ^b       P^b      �c       V�c      @e       V                    yb      d       ]d      qd        2$#����} "��d      Je       ]                          �b      �b       P�b      �b       T�b      �c       ���c      �c       T�c      Je       ��                       b      !b       u��!b      6b       ~��6b      9b       �U#��9b      Je       ~��                 td      �d       _                    �d      �d       P�d      �d       w                         �b      c       _c      c       Qc      �c       _�d      Je       _                             �b      c       Yc      fc       w fc      tc       y�tc      �c       Y�c      �c       w �1��d      >e       w >e      Je       Y                        �e      �e       U�e      �e       S�e      �e       �U��e      �f       S                          �e      �e       T�e      �e       Q�e      �e       \�e      �e       �T��e      �f       \                              �e      �e       P�e      �e       P�e      �e       V�e      ;f       P;f      <f       V<f      if       Pwf      �f       P                       �e      �e       u���e      �e       s���e      �e       �U#���e      �f       s��                    `�      f�       Uf�      g�       �U�                    `�      f�       Tf�      g�       �T�                    p�      v�       Uv�      w�       �U�                    p�      v�       Tv�      w�       �T�                         L      oL       UoL      wL       �U�wL      �L       U�L      �L       �U�                         L      rL       TrL      wL       �T�wL      �L       T�L      �L       �T�                       L      L       QL      vL       ZwL      �L       Z                           L      L       RL      vL       QvL      wL       �R�wL      �L       Q�L      �L       �R�                         L      vL       XvL      wL       �X�wL      �L       X�L      �L       �X�                   hL      oL       u�oL      vL       U                  �L      �L       P                         [L      hL       YhL      vL       RwL      �L       Y�L      �L       Y�L      �L       R                   L      IL       U�L      �L       U                  L      IL       T                   L      *L       P+L      IL       P                   L      IL       R                        @�      L�       UL�      ��       ]��      ��       �U���      �       ]                        @�      _�       T_�      ��       S��      ��       �T���      �       S                        [�      �       ^��      G�       ^�      ʗ       ^��      �       ^                      2�      G�       0�G�      �       _ʗ      ۗ       _                                 [�      �       0���      Ô       0�Ô      2�       \2�      G�       0�G�      �       V�      ��       v���      ��       q��      ��       0���      ��       \ʗ      ۗ       V��      �       0�                                      G�      j�       ^�w �\�P���      ��       P����      ��       ^����      ��       ^�P����      ��      	 ^�w ����      ��       ^�w �P����      ��       ^�w �\����      �       ^�w �\�P�ʗ      ӗ       ^�w �\�P�ӗ      ֗       ^�w �\��֗      ۗ       ^�w �\�P�                 ��      ؕ       0�                 ��      �       0�                   �      ʗ       �����      �       ���                   �      ��       ��  ��      ʗ       ��  ��      ��       ��                     �      ��       S��      ʗ       S��      ��       S                 ��      ʗ       2�                     <�      b�       0�b�      }�       V}�      ��       v���      ��       V                   �      b�       0�b�      ��       \��      ��       \                     �      b�       0�b�       �       ��~ �      l�       1�l�      ��       ��~��      ��       1�                       �      b�       0�b�      x�       ��~x�      }�       1�}�      ��       ��~��      ��       ��~                   �      b�       0�b�      ��       _��      ��       _                      +�      /�       P/�      ��       w ��      ʗ       w ��      ��       w                       +      V+       UV+      [+       �U�[+      f+       U                      +      S+       TS+      [+       �T�[+      f+       T                      +      Z+       QZ+      [+       �Q�[+      f+       Q                      +      Z+       RZ+      [+       �R�[+      f+       R                  G+      Z+       P                     +      V+       UV+      [+       �U�[+      f+       U                     +      V+       UV+      [+       �U�[+      f+       U                    +      G+       T[+      f+       T                   +      G+       P[+      e+       P                    &+      G+       X[+      f+       X                      �       F!       TF!      �"       �T��"      #       T                      �       F!       QF!      �"       �Q��"      #       Q                           �       F!       0�F!      A"       ]A"      F"       PF"      �"       ]�"      �"       ]�"      #       0�                       !      "       S"      &"       s�&"      9"       SF"       #       S #      #       u�
                     !      F!       1�F!      �"       [�"      #       1�                             �       !       P!      !       p�!      F!       RF!      F!       r�F!      F!       r�F!      z!       r�z!      �!       r��!      �!       T�!      �!       t��!      �!       T�!      "       t�"      "       T"      F"       XF"      �"       T�"      �"       T                    !      ="       VF"      #       V                        F!      "       RF"      S"       RS"      �"       tr��"      �"       R�"      �"       tr�                  j!      �"       X                        F!      "       r ��8$r��!
���F"      S"       r ��8$r��!
���S"      �"       tr��8$ts��!
����"      �"       r ��8$r��!
����"      �"       tr��8$ts��!
���                              F!      U!       r��8$r��!
���U!      ]!       x 8$r��!
���]!      `!       p 8$r��!
���`!      "       r��8$r��!
���F"      S"       r��8$r��!
���S"      �"       tt��8$tu��!
����"      �"       r��8$r��!
����"      �"       tt��8$tu��!
���                        F!      "       r��8$r��!
���F"      S"       r��8$r��!
���S"      �"       tv��8$tw��!
����"      �"       r��8$r��!
����"      �"       tv��8$tw��!
���                        �!      �!       q 
����!      �!       Q�!      �!       QF"      S"       Q                           F!      "       0�F"      �"       0��"      �"       P�"      �"       0��"      �"       P�"      �"       0�                   S"      �"       ^�"      �"       ^                        S"      w"       Qw"      �"       Y�"      �"       Q�"      �"       Y                          _"      �"       Y�"      �"       R�"      �"       Y�"      �"       Y�"      �"       R                        h"      h"       Ph"      �"       p��"      �"       t p "#��"      �"       P�"      �"       p��"      �"       p�                        n"      w"       R�"      �"       Q�"      �"       R�"      �"      + p �H0H%�$!0)( 8/�������                  �!      �!       Q                              �!      �!      	 p ������!      �!       P�!      "      + r�H0H%�$!0)( 8/�������"      "      	 p �����"      "       P"      "      + r�H0H%�$!0)( 8/��������"      �"       P                      �(      �(       U�(      �*       S�*      �*       �U�                            �(      �(       T�(      �(       Q�(      u)       Vu)      �*       �T��*      �*       V�*      �*       �T�                      �(      �(       P�(      )       P)      �*       Y                              
)      )       R)      )       r�)      B)       XB)      B)       x�B)      \)       x�\)      �)       x��)      �)       T�)      �)       t��)      �)       t��)      �)       t��)      *       x�*      *       x�*      *       ^*      E*       x�E*      M*       x�M*      Z*       ^Z*      p*       ~�p*      p*       ^p*      �*       ~��*      �*       ^                  )      �*       U                     ,)      �)       0��)      �*       R�*      �*       0�                     )      ,)       p 
���,)      �*       Z                     �(      �)       0��)      �*       V�*      �*       0�                     �(      �)       0��)      �*       \�*      �*       0�                      *      *       p 
���*      .*       P:*      d*       P                    \)      �)       p 
����)      *       p 
���                    `)      �)       ^�)      �)       ^                 �)      �)       ~ 8%�                       B)      �)       X�)      �)       T�)      �)       X�)      �*       T                     5)      �)       1��)      �)       ]�)      �*       ]                    V*      �*       Q�*      �*       q��*      �*       Q                    E*      S*       ��������p*      �*       P�*      �*       P                    a*      p*      & ~��@$~ ��H$!~��8$!~��!�v*      �*      & ~��H$~��@$!~��8$!~	��!�                        @       f        Tf       �        �T��       �        T�       �        �T�                    G       �        R�       �        R                    j       �        T�       �        �T1$����r"�                    �       �        P�       �        p��       �        p}��       �        p~��       �        p��       �        P                   �       �        Q�       �        q|��       �        Q                  �       �        T                       j       �        t ��8$t��!��       �        p �8$q �!��       �        �T1$����r"��8$q �!��       �       . �T1$����r"��8$�T1$����r"#��!�                      �?      �?       U�?      
@       �U�
@      @       U                 �?      �?       u�                 �?      �?       u�                        �?      @       S@      	@       T
@      @       S@      @       u�                        �G      �G       U�G      DH       SDH      NH       �U�NH      �K       S                          �G      �G       T�G      �G       Q�G      EH       VEH      NH       �T�NH      �K       V                    �G      KH       ^NH      �K       ^                                 �G      H       0�NH      �H       0��H      �H       _�H      �H       ��H      �H       ��H      �H       ��H      I       �I      cI       �cI      �I       _�I      �I       Q�I      �I       q��I      �I       q��I      �I       q��I      �I      	 }p "#�J      DJ       [�J      �J       _�K      �K       _                        �G      H       0�H      0H       ]0H      ?H       0�NH      �H       0��H      �H       P�H      �K       ]                  I      jI       Q                      �I      �I      	 { ������I      �I       [�I      DJ       w                        {I      �I       0��I      DJ       P�J      �J       P�K      �K       P                     J      DJ       X�J      �J       Q�K      �K       Q                         J      J       PJ      DJ       Q�J      �J       P�J      �J       R�K      �K       P�K      �K       R                            0U      �U       U�U      �W       _�W      Y       �U�Y      rY       _rY      �Y       U�Y      ]Z       _                            0U      �U       T�U      �W       ���W      Y       �T�Y      rY       ��rY      �Y       T�Y      ]Z       ��                    0U      hU       QhU      ]Z       ��                          0U      rU       RrU      �U       S�U      rY       ��~rY      �Y       S�Y      ]Z       ��~                      �W      �W       0��W      �X       ^�X      �X       ~��X      �X       ^                          �V      �V       0��V      �V       ^�V      �V       ~��V      �V       ^�W      �W       0��W      �X       ���X      �X       P                      [W      �W       U�W      �X       ��UY      rY       U                      `W      �W       T�W      �X       ��]Y      rY       T                      eW      �W       Q�W      �X       ��eY      rY       Q                      jW      �W       Y�W      �X       ��mY      rY       Y                      V       V       p | ����� V      $V       T$V      :W       ���| ������Y      �Y       S                      �W      �W       S�W      �X       ���X      �X       ��                  �W      �X       ]                        �U      �U       T�U      :W       ��0Z      9Z       ��9Z      LZ       u p u  $p  $,( �                        �U      �U       ^�U      V      ) ��~#��p "z ��~#��p " $z  $*( �V      $V      7 ��~#����~#��"z ��~#����~#��" $z  $*( �0Z      LZ       ^                      �U      V       \V      $V       r x { r x  ${  $,( �0Z      LZ       \                        �U      �U       S�U      :W       ��0Z      =Z       ��=Z      LZ       t r t  $r  $*( �                 �U      $V       �                    	V      �V       V�V      �V       ��                    V      $V       P$V      :W       ��                 V      :W       \                       V      -V       0�-V      1V       P1V      �V       U�V      :W       ��                  [V      �V       ]                   �V      �V       R�V      �V       R                     �W      X       ~ ������"���X      X       PX      pX       ~ ������"���                  >X      �X       P                    @X      eX       QeX      �X       �p �                   @X      GX       UGX      pX       | ���                   @X      JX       TJX      pX       v ���                   @X      ]X       R]X      pX       s ���                 @X      �X       _                            �              T       `       �T�`      j       Tj      �       �T��      )        T)       9        �T�                          �      :       R:      `       �R�`      �       R�      �       �R��      9        R                      �      V       V`      �       V�      9        V                             `      o       �y��8$y��!���o      r       �y��8$y��!��p t !��r      �       �y��8$y��!��P��      �      6 �z �8$s { O%s { "1&{ "31$ $ &| "#��!��P��      �       �z �8$y �!��P��      �       �z �8$y �!��x �)       9        �z �8$y �!��x �                    �      �       P)       4        P                  `      o       ���  �      )        ���                      `      j       Tj      o       �T��      )        T                  `      o      	 v�
����      )       	 v�
���                  `      o       \�      )        \                    `      o       [�      �       0��      )        [                   `      o       S�      )        S                       `      e       Pe      o       s { O%s { "1&{ "��      �       P�      )        P                     `      `       y�`      `       y�`      o       y��      �       y�               Y       )        y�                    `      o       y ��8$y��!��      �       y ��8$y��!�       )        y ��8$y��!�                      �?      �?       U�?      �?       �U��?      �?       U                 �?      �?       u�                 �?      �?       u�                        �?      �?       S�?      �?       T�?      �?       S�?      �?       u�                          �E      $F       U$F      gF       SgF      qF       �U�qF      �G       S�G      �G       U                            �E      F       TF      $F       Q$F      hF       VhF      qF       �T�qF      �G       V�G      �G       T                      �E      jF       \qF      �G       \�G      �G       u�                       F      @F       0�qF      �F       0��F      �F       _�F      �F       ��F      G       �G      1G       �1G      AG       �AG      �G       ��G      �G       0�                           F      @F       0�@F      ^F       ^^F      bF       0�qF      �F       0��F      �F       P�F      �G       ^�G      �G       0�                  G      G       Q                  AG      �G       R                      �      �       U�      �       �U��      �       U                      �      �       T�      �       �T��      �       T                     �      �       U�      �       �U��      �       U                   �      �       u�      �       u                          g      �g       U�g      �i       ��~�i      �i       �U��i      �i       U�i      j       ��~                          *g      7g       P7g      �g       u��g      �i       ��~�i      �i       u��i      j       ��~                          ;g      �g       T�g      �i       w �i      �i       ��~�i      �i       T�i      j       w                    ;g      �g       u�#�i      �i       u�#                    �h      �h       p q !��h      �h       P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                      �E      �E       U�E      �E       S�E      �E       �U�                 �E      �E       u                  �E      �E       u #�                        P      d       Ud      z       Tz      {       �U�{      �       T                    P      V       TV      �       �T�                    S      z       Y{      �       Y                    d      z       U{      �       U                     d      h       Ph      z       y�{      �       y�                      ��      ��       U��      ��       �U���      ��       U                      ��      ��       T��      ��       �T���      ��       T                     ��      ��       �h���      ��       Q��      ��       �h�                     ��      ��       T��      ��       �T���      ��       T                     ��      ��       U��      ��       �U���      ��       U                                      �6      �6       U�6      �7       _�7      o8       �U�o8      �8       _�8      �8       U�8      �8       �U��8      �8       _�8      �8       �U��8      �8       _�8      �8       U�8      �9       �U�                                      �6      �6       T�6      �6       [�6      7       Q7      ^7       [^7      o8       �T�o8      s8       Qs8      �8       [�8      �8       �T��8      �8       [�8      �8       Q�8      �9       �T�                      �6      �6       Q�6      �6       T�6      �9       �Q�                                    �6      �6       P�6      �6       p�7      7       T7      '7       t�'7      �7       ~��7      �7       ~��7      �7       u~��7      �7       U�7      �7       u��7      8       u~�8      o8       Uo8      s8       t��8      �8       ~��8      9       U~9      �9       U�9      �9       u��9      �9       u~��9      �9       U                                           �7      8       Y8      8       y�8      8       Y8      68       y��8      �8       Y�8      �8       y��8      �8       Y�8      �8       y��8      �8       Q�8      A9       XA9      K9       x�K9      K9       XK9      \9       x�\9      h9       X�9      �9       T�9      �9       Y�9      �9       Y                    �6      �6      	 } ������6      �6       ]                      �6      W7       Uo8      }8       U�8      �8       U                         7      �7       _�7      o8       �U�o8      s8       _�8      �8       _�8      �9       �U�                  @7      ^7      & } ��H$}��@$!}��8$!}��!�o8      s8       0�                        7      '7      & t ��H$t��@$!t��8$!t��!�'7      ^7      & ~ ��H$~��@$!~��8$!~��!�o8      s8      & t ��H$t��@$!t��8$!t��!��8      �8      & ~ ��H$~��@$!~��8$!~��!�                        �7      8       Qf8      o8       Q�8      �8       Q19      A9       T                         @7      Z7       Q�7      T8       ]f8      o8       ]o8      s8       0��8      9       ]19      h9       Y~9      �9       ]                          �7      �7       R8      o8       R�8      �8       R~9      �9       R�9      �9       R                      �7      ?8       Z?8      O8       z�O8      f8       z��8      9       Z9      9       z�9      19       z�19      �9       Z                 �7      �7       1�                      �7      �7       1��7      �7       {��7      8       [�8      9       [                                     8      8       1�8      8       0�8      o8       1��8      �8       1��8      �8       0��8      9       1�19      A9       0�A9      K9       1�K9      M9       0�M9      h9       1�~9      �9       1�                    t7      o8       P�8      �9       P                   7      77       P77      ;7       p|�;7      @7       Po8      o8       P                  7      )7      & } ��H$}��@$!}��8$!}��!�o8      o8      & } ��H$}��@$!}��8$!}��!�                   7      )7       0�)7      @7       Qo8      o8       0�                            6      %6       U%6      ~6       \~6      6       �U�6      �6       \�6      �6       �U��6      �6       \                               6      6       T6      !6       t�!6      :6       v�:6      E6       RE6      S6       r�S6      i6       r~�i6      t6       R6      �6       v��6      �6       �T#��6      �6       v�                    6      %6       Q%6      �6       �Q�                            6      %6       U%6      ~6       \~6      6       �U�6      �6       \�6      �6       �U��6      �6       \                   /6      E6       0��6      �6       0�                    /6      6       P�6      �6       P                              05      [5       U[5      �5       \�5      �5       �U��5      �5       \�5      �5       �U��5      �5       U�5      6       \                            05      [5       T[5      z5       Vz5      �5       S�5      �5       s��5      �5       s��5      �5       S�5      �5       T�5      �5       t��5      6       �T#�                        05      ~5       Q~5      �5       �Q��5      �5       Q�5      6       �Q�                             75      [5       U[5      �5       \�5      �5       �U��5      �5       \�5      �5       �U��5      �5       U�5      6       \                     z5      ~5      & v ��H$v��@$!v��8$!v��!��5      �5      & t ��H$t��@$!t��8$!t��!��5      �5      0 �T��H$�T#��@$!�T#��8$!�T#��!�                   p5      ~5       R�5      �5      
 s��#��5      6       0�                        �5      �5       P�5      �5       Q�5      �5       q|��5      �5       Q�5      6       T                  �5      �5       R                     75      75       T75      A5       t�A5      T5       t�T5      g5       Pg5      k5       p|�k5      p5       P�5      �5       t�                   A5      [5      & t ��H$t��@$!t��8$!t��!��5      �5      & t ��H$t��@$!t��8$!t��!�                   A5      [5       0�[5      p5       R�5      �5       0�                        �9      :       U:      �:       \�:      �:       �U��:      �:       \                      �9      :       T:      :       P:      �:       �T�                                �9      �9       Q�9      �:       ^�:      �:       T�:      �:       ^�:      �:       �Q��:      �:       ^�:      �:       T�:      �:       ^                       �9      :       U:      �:       \�:      �:       �U��:      �:       \                    :      <:       ]�:      �:       ]                           :      9:       v
�9:      Y:       SY:      Y:       s�Y:      `:       s�`:      e:       s|�e:      �:       S�:      �:       S�:      �:       v
�                         (:      J:       _J:      �:       ]�:      �:       }|��:      �:       ]�:      �:       ]�:      �:       _                   Y:      `:       s ��@$s��8$!s��!�`:      }:       su��@$sv��8$!sw��!�                      e:      m:      	 p �����m:      u:       Uu:      }:      	 p �����                    g:      }:      	 q �����}:      �:       ��������                             ;      ;       U;      u;       \u;      v;       �U�v;      �;       \�;      �;       �U��;      �;       \                       ;      ;       T;      ;       Q;      �;       �T�                            ;      ;       U;      u;       \u;      v;       �U�v;      �;       \�;      �;       �U��;      �;       \                      ;      k;       Vv;      �;       V�;      �;       V                           ;      .;       s
�.;      6;       R6;      O;       r�O;      `;       rx�`;      k;       Rv;      �;       s
��;      �;       s
�                    #;      v;       P�;      �;       P                   #;      6;       0��;      �;       0�                    �      �       U�      H       �U�                              �      �       T�             V             �T�      "       V"      .       T.      F       VF      H       T                          �      �       Q�      �       T�      .       �Q�.      4       T4      H       �Q�                    �      �       P�      �       p��      �       p�.      <       p�                    �      �      	 q �����.      <      	 q �����                      �            	 | �����      &      	 | �����.      H      	 | �����                    @      Y       UY      �       �U�                                @      I       TI      �       \�      �       �T��      �       \�      �       U�      �       �T��      �       \�      �       �T�                                @      ]       Q]             V      �       �Q��      �       V�      �       T�      �       �Q��      �       V�      �       T                          @      ]       R]      r       Tr      �       �R��      �       T�      �       �R�                    ^      c       Pc      r       p��      �       p�                    k      r      	 q ������      �      	 q �����                      n      w      	 } ������      �      	 } ������      �      	 } �����                  �      �       U�      <       u�                  �      <      & u ��H$u��@$!u��8$!u��!�                           �      �      & u ��H$u��@$!u��8$!u��!��      �       X�      �       R�             Y             R"      /       Y/      <       X                 �      �       0��      <       Z                          �      �       Y�      �       R�      �       Y�             R"      <       R                          �      �       P�      �       p��      �       P�      �       P�             p�"      ,       p�,      /       P                        �      �      	 q �����             q x !�����            	 q �����"      /      	 q �����                  �      �       U�      �       u�                  �      �      & u ��H$u��@$!u��8$!u��!�                       �      �      & u ��H$u��@$!u��8$!u��!��      )       X)      d       Yg      m       Xm      �       Y                 �      �       0��      �       Z                                6       Y6      _       Q_      d       Yg      m       Ym      �       Q                                     R      9       r�9      >       p u "#�>      >       R>      d       r�g      m       r�                        #      9       PU      X       p x !�X      d       Pg      �       P                  @      L       UL      �       u�                  L      �      & u ��H$u��@$!u��8$!u��!�                           L      L      & u ��H$u��@$!u��8$!u��!�L      �       [�      �       Q�      �       X�      �       Q�      �       X�      �       [                 L      L       0�L      �       Z                          X      �       X�      �       Q�      �       X�      �       Q�      �       Q                          e      e       Qe      z       q�z      �       q��      �       x 2$����u "#��      �       R�      �       r��      �       q 2$����u "#��      �       q 2$����u "#��      �       q 2$����u "#�                      z      �      	 p ������      �      	 p ������      �      	 p �����                    ~      �       q����      �       x 2$����u "#���                        0�      W�       UW�      *�       ��*�      8�       U8�      B�       ��                        0�      W�       TW�      ��       S��      ɉ       �T�ɉ      B�       S                            W�      W�       ��#�W�      z�       ��#�z�      ��       _��      �       ��      "�       x�"�      6�       |�6�      ɇ       _ɇ      S�       ��k�      ��       _��      ��       _��      *�       _                    z�      ��       T��      *�       ��                 z�      Ԇ       \                  ��      Ԇ       0�                              ��      Ԇ       1�Ԇ      �       ���      �       P�      k�       ��k�      }�       P}�      ��       ��ɉ      *�       ��                        Ԇ      �       \"�      ��       \k�      ��       \�      *�       \                        Ԇ      �       ]6�      y�       ]y�      ��       ^k�      ��       ]                            Ԇ      ��       ��;�      M�       PM�      ��       ��k�      |�       P|�      ��       ��ɉ      *�       ��                               y�      ��       ]��             ^      ·       }�·      ݇      
 ~ 2$v "#�݇      �      
 ~2$v "#��      �      
 ~ 2$v "#��      7�      
 ~ 2$v "#�7�      B�      
 ~2$v "#���      �       ^�      *�       ]                        ��      ��       U��      S�       w ��      �       U�      �       w                         ��      ·       0�·      7�       ^7�      <�       ~�<�      S�       ^�      �       0�                      y�      ·       0�·      3�       _<�      K�       _��      *�       0�                    ·      �       \�      S�       \                   ·      Շ       ~ 2$v "#����      !�       ~ 2$v "#���                          a�      n�       ]n�      ��       \��      
�       |�
�      (�       |~�(�      k�       \��      ��       \ɉ      �       \�      ��       ]                          ��      ��       T��      k�       w ��      ��       w ɉ      Չ       TՉ      �       w                             ��      ��       0���      k�       ^��      ��       ^��      ��       ~���      ��       ^݉      �       0�                       a�      ��       0���      k�       _��      ��       _ɉ      ��       0�                      ��      Ɉ       Q(�      @�       Q@�      O�       ��                   ��      ؈       } �8$v �!
���(�      k�       } �8$v �!
���                  �      �       T�      �       t�                        �4      �4       U�4      �4       �U��4      5       U5      (5       S                          �4      �4       T�4      �4       �T��4      5       T5      5       R5      (5       V                          �4      �4       Q�4      �4       �Q��4      5       Q5      5       Z5      (5       �Q�                    �4      �4       P�4      5       P                        pE      �E       U�E      �E       S�E      �E       �U��E      �E       U                    tE      �E       P�E      �E       P                    �      �       p��      �       u#�                    �      �       U�      �       �U�                    �      �       T�      �       t                               �             U      %       V%      +       U+      /       V/      6       �U�6      \       U\      |       V|      �       U                          �      �       T�      /       ]/      6       �T�6      O       TO      �       ]                      �             Q      6       �Q�6      `       Q`      �       �Q�                         �             0�+      /       P6      U       0�U      d      & t��H$t	��@$!t
��8$!t��!�n      |       P�      �       P                          �      �       s��      �       t��      �       T�      �       t��             t�6      O       s�O      |       t�                    �            & s��H$s��@$!s��8$!s��!�6      d      & s��H$s��@$!s��8$!s��!�                     �      �       t �             [6      |       [                      �      �      & t ��H$t��@$!t��8$!t��!��            & t ��H$t��@$!t��8$!t��!�O      d      & t ��H$t��@$!t��8$!t��!�                           �      �       	���      �      & t��H$t��@$!t��8$!t��!��      �       	���            & t��H$t��@$!t��8$!t��!�6      O       	��O      d      & t��H$t��@$!t��8$!t��!�                         �      �      & s��H$s��@$!s��8$!s��!��      �       Y�      �       R�             YO      |       Y                     �      �       0��             ZO      |       Z                          �      �      & s��H$s��@$!s��8$!s��!��      �       R�      �      & s��H$s��@$!s��8$!s��!��             R6      O      & s��H$s��@$!s��8$!s��!�O      |       R                  �             u `      |       Q                        �             U      %       V%      +       U+      /       V`      |       V|      �       U                 �      u       u                      !      0       r�0      5       r|�5      5       R5      @       r�@      m       r�                          !      0      + r �H0H%�$!0)( 8/�������0      5      + rt�H0H%�$!0)( 8/�������@      B      	 p �����B      P       PP      d      + r �H0H%�$!0)( 8/�������                      !      5       PD      P      	 q �����P      m       P                      !      0      , r��H$r	��@$!r
��8$!r��!�����0      5      , r|��H$r}��@$!r~��8$!r��!�����J      d      , r��H$r	��@$!r
��8$!r��!�����                  
      m       T                 
      m       Y                     !      0      & r��H$r	��@$!r
��8$!r��!�0      5      & r|��H$r}��@$!r~��8$!r��!�N      d      & r��H$r	��@$!r
��8$!r��!�                          ��      �       U�      o�       Vo�      �       �U��      �       U�      "�       V                          ��      �       T�      
�       _
�      �       �T��      �       T�      "�       _                    �      �       v��      %�       v�%�      %�       v�%�      ��       ]��      ��       }���      ��       }x���      ��       }|���      ��       ]                      %�      G�       PG�      J�       p�J�      _�      + v�H0H%�$!0)( 8/�������                      .�      _�       R_�      ��       w ��      �       ��                      `�      o�       0�o�      �       ^�      �       ~��      ��       ^                    o�      ��       V��      ��       V                    o�      ��       S��      ��       S                 ��      Յ      , }��H$}	��@$!}
��8$!}��!�����                        `�      o�       0���      ��       S��      Յ       QՅ      ݅       ���      ��       S                  �      �       T�      �       t�                    �      �       p��      �       u#�                    �      �       U�      �       �U�                    �      �       T�      �       t                               `      �       U�             V             U             V             �U�      3       U3      q       Vq      �       U                          `      �       T�             ]             �T�      /       T/      �       ]                      `      �       Q�             �Q�      U       QU      �       �Q�                        `      �       0�             P      J       0�J      q       P{      �       P                           l      �       s��      �       t��      �       T�      �       t��      �       t�      /       s�/      6       t�6      q       r 1$r "2$����s "#�                    s      �      & s��H$s��@$!s��8$!s��!�      Y      & s��H$s��@$!s��8$!s��!�                     s      �       t �      �       [      q       [                        �      �      & t ��H$t��@$!t��8$!t��!��      �      & t ��H$t��@$!t��8$!t��!�/      6      & t ��H$t��@$!t��8$!t��!�6      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                                   �       	���      �      & t��H$t��@$!t��8$!t��!��      �       	���      �      & t��H$t��@$!t��8$!t��!�      /       	��/      6      & t��H$t��@$!t��8$!t��!�6      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                  >      Y      n r 1$r "2$����s "#��H$r 1$r "2$����s "#��@$!r 1$r "2$����s "#��8$!r 1$r "2$����s "#��!�                         �      �      & s��H$s��@$!s��8$!s��!��      �       Y�      �       R�      �       Y/      q       Y                     �      �       0��      �       Z/      q       Z                                �      & s��H$s��@$!s��8$!s��!��      �       R�      �      & s��H$s��@$!s��8$!s��!��      �       R      /      & s��H$s��@$!s��8$!s��!�/      q       R                  �      �       u U      q       Q                        �      �       U�             V             U             VU      q       Vq      �       U                   P      d       u 4      =       u                      �      �       Y�      �       y��              y�       )       y|�=      Y       y�                    �      )       X=      Y       X                    �      )       R=      Y       R                    �      )       \=      N       \                         l      �       P�      �       P�      �       Q�             P             Q      4       P=      Y       P                   l      4       [=      Y       [                        �      �       q p "��      �       ]�      �       0��             ]             0�                          ��      ��       U��      ��       V��      ф       �U�ф      ��       U��      �       V                          ��      ��       T��      ΄       ^΄      ф       �T�ф      ݄       T݄      �       ^                    ��      ��       v���      ��       v���      ��       v���      k�       \k�      x�       |�x�      ��       |x���      ��       ||���      ��       \                      ��      ׃       P׃      ڃ       p�ڃ      �      + v�H0H%�$!0)( 8/�������                      ��      �       R�      Ą       w Ą      ф       ��                    ��      ��       0���      ��       ]                    ��      k�       _��      ��       _                      ��      k�      	 v �������      ��       X��      ��       ��                 ��      ��      , |��H$|	��@$!|
��8$!|��!�����                       ��      ��       0�^�      k�       Xk�      ��       Q��      ��       ��                     1�      9�       v s �9�      L�       TL�      ^�       v  �                  0      4       T4      F       t�                                 p�      )       u#�                    `      q       Uq             �U�                      d      w       Pw      �       yl��             �U#                    �      �       Q�             Q                                         d      �       0��      �      
 y z !
����      �       z 
����      �       0��      �      
 u p !
����      �       p 
����      �       0��      �       P�      �       p 
����      �       p 
����             P             0�             z 
���                             d      d       p�d      w       p�w      y       y|�y      �       Y�      �       R�      �       R�             R             Y             R                              �      �       Z�      �       q u ��      �      � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/����      �      � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/����            � �U##�H0H%�$!0)( 8/��t �#�U##�H0H%�$!0)( 8/������t �#����*( �U##�H0H%�$!0)( 8/���             Z             q u �                           1       T1      S       �T�                    $      A       RA      S       u                 $      R       0�                   $      $       r�$      +       r�+      A       r�A      R       R                    +      A      & r��H$r��@$!r��8$!r��!�A      S      2 u#��H$u#��@$!u#��8$!u#��!�                   +      A      & r��H$r��@$!r��8$!r��!�A      S      2 u#��H$u#��@$!u#��8$!u#��!�                      1      <       T<      A      ) �Tr�H0H%�$!0)( 8/���A      R      , �Tu#�H0H%�$!0)( 8/���                            ��      ς       Uς      #�       ]#�      &�       �U�&�      b�       ]b�      p�       Up�      z�       ]                            ��      ς       Tς      !�       \!�      &�       �T�&�      b�       \b�      m�       Tm�      z�       \                         ��      ς       u�ς      ς       }�ς      �       }��      �       }��      �       }�&�      b�       Sb�      p�       u�p�      z�       }�                      �      ��       P��      ��       p���      �      + }�H0H%�$!0)( 8/�������                        �      �       V&�      =�       V=�      A�       v�A�      b�       V                        &�      <�       s~��8$s��!
���G�      K�       s~��8$s��!
���K�      N�       p 8$s��!
���N�      b�       s~��8$s��!
���                                 p�             u#�                             I       UI      �       �U��      �       U                          1       u �      �       u                                   �       0��      �       Q�      �       0��      �       Q�      �       0��      �       Q                               i       Ql      �       Q�      �       Q�      �       Q�      �       t �#�                                          �       0��      �       r x "��      �       P�      �       0��      �       p u ��      �       P�      �       P�      �       0��      �       P�      �       0��      �       P                          I       X�      �       X                                      x�� �      $       x�� �$      I       YI      [       y�[      a       yx�a      f       y|�f      �       Y�      �       x�� ��      �       Y                          1      . x�� ��H$x�� ��@$!x�� ��8$!x�� ��!��      �      . x�� ��H$x�� ��@$!x�� ��8$!x�� ��!�                    l      �      & y��H$y	��@$!y
��8$!y��!��      �      & y��H$y	��@$!y
��8$!y��!�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       R�      �       �U#                       �      �       r�� ��      �       P�      �       p��      �       px��      �       p|��      �       P�      �       P                  �      �      . r�� ��H$r�� ��@$!r�� ��8$!r�� ��!�                     �      �      & p��H$p	��@$!p
��8$!p��!��      �      & p��H$p	��@$!p
��8$!p��!��      �      & p��H$p	��@$!p
��8$!p��!�                              �      8�       U8�      ��       S��      ��       vt���      ��       S��      ��       vt���      w�       �U�w�      ��       S                            �      8�       T8�      ��       ]��      Ł       �T�Ł      w�       ]w�      ��       T��      ��       ]                                �      8�       u�8�      8�       s�8�      j�       s�j�      j�       v�� �j�      ��       _��      ��       ���      ��       x���      ��       |���      ��       _��      ��       s���      ��       _Ł      w�       _w�      ��       s���      ��       _                          j�      ��       V��      ��       V��      Ł       �U#�Ł      w�       V��      ��       V                    D�      W�      & s��H$s��@$!s��8$!s��!���      ��      & s��H$s��@$!s��8$!s��!�                    u�      ��      . s�� ��H$s�� ��@$!s�� ��8$!s�� ��!���      ��      . s�� ��H$s�� ��@$!s�� ��8$!s�� ��!�                            ��      ��       0���      ��       w ��      ��       w ��      ��       PŁ      w�       w ��      ��       0�                              0�      Q�       SQ�      X�       QX�      ��       SŁ      ځ       S�      #�       S#�      .�       Q.�      [�       S                   ��      ��      & ��H$	��@$!
��8$!��!�ځ      ��      & ��H$	��@$!
��8$!��!�                        �      0�       R�      �       R[�      p�       Rp�      w�       ��                          ��      ��       0���      ��       Qځ      ��       Q��      �       ����      ��       0�                         0�      X�       s @%�X�      b�       s @%�b�      j�       Rj�      ��       s @%�Ł      ځ       s @%�                        0�      X�       s 
���X�      ��       s 
���Ł      ځ       s 
����      .�       s 
���.�      [�       s 
���                          ��      �       R�      �       ���      0�       ~ s ��      �       ~ s �[�      w�       ~ s �                  d      �       r�                    �      �       U�      X       �U�                         �      �       u�      �       Y�      N       �U#N      R       YR      X       �U#                         �      8       0�8      ;       Q;      K       0�K      N       QN      X       0�                          �      �       Q�      �       t �#��      8       Q;      P       QP      R      # t �#u t �#����u ����*( �R      X       Q                                         �      �       0��             
 z y !
���              y 
���             0�      "      
 u p !
���"      ,       p 
���,      8       0�8      ;       P;      B       p 
���C      K       p 
���K      N       PN      R       0�R      X       y 
���                               �      �       u#��      �       u#��      �       u#
��      �       y
��      �       Z�      8       R;      B       RC      N       RN      R       ZR      X       R                           �      �       u#��8$u#��!
����      �       y��8$y��!
����      :      " �U##��8$�U##��!
���;      M      " �U##��8$�U##��!
���N      R       y��8$y��!
���R      X      " �U##��8$�U##��!
���                           �      �       u#��8$u#	��!
����      �       y��8$y	��!
����      :      " �U##��8$�U##	��!
���;      M      " �U##��8$�U##	��!
���N      R       y��8$y	��!
���R      X      " �U##��8$�U##	��!
���                      �      8       [;      B       [C      X       [                    @      \       T\      �       �T�                    D      w       Rw      �       u                 D      �       0�                   D      D       r�D      D       r�D      w       r
�w      �       R                       D      H       r��8$r��!
���H      K       p 8$r��!
���K      w       r��8$r��!
���w      �       u#��8$u#��!
���                         D      W       r��8$r	��!
���W      b       q 8$r	��!
���b      e       p 8$r	��!
���e      w       r��8$r	��!
���w      �       u#��8$u#	��!
���                  \      r       T                                     ?       U?      �       \�      �       sv��      �       �U��      �       \�      �       U�      �       \                                   ?       T?      �       V�      �       �T��      �       V�      �       T�      �       V                     ?      ?       |�?      \       |�\      \       |�\      �       |
��      �       S�      �       |
�                    \      �       p 
����      �       P                    u      �       ^�      �       ^                        �      �       s~��8$s��!
����      �       s~��8$s��!
����      �       p 8$s��!
����      �       s~��8$s��!
���                        4       r�                        �      �       U�      �       �U��             U      
       �U�                      �      �       T�      �       t �             t                             �
      �
       U�
      �       ���      �       U�      �       ���             �U�      �       ��                            �
      �
       T�
      �       ���      �       T�      �       ���             �T�      �       ��                        �
      �
       Q�
      �       �Q��      �       Q�      �       �Q�                 �
      �
       u                  �
      �
       u #�u #�"�                  �
      �
      
 | 
��	��                                                       �
             Z<      K       Z�      �       Z      �       Z�             ZW      �       [�      �       { 
����      �       [�             ��R      �       Z�      �       [�      �       ���      N       ZN      �       [�      �       Q�      �       [             ��      !       Z:      d       Zz      �       Z                                                               �
      �
       
����
             [      )       
���)      V       [�      �       
����      �       [      �       [�             [      W       ]W      �       ^�             ^      E       ��E      �       [�      �       
���H      �       [�      �       ^N      �       ^�      �       ^�             ��             ^      !       [!      :       ]N      Y       [Y      d       
���d      z       ]                                             �      �       ��s      w       Vw      �       ���      �       0��             ��W      �       \�      �       z 
����             \�      �       0�H      d       ��d      �       0��      �       \N      �       \�      �       \             \N      d       0�                                               �      �       ��d      o       Vo      �       ���      �       1��             ��W      �       U�      �      	 u 0$0&��             Ud      h       Rh      �       ���      �       ��H      �       ���      �       UN      �       U�      �       U             UN      d       1�                           �
      �
       P�
      D       YD      I       T�      �       P             Y�             TH      d       T                      �
      �
       0��
      I       V�      �       0�      <       V                                                         �
      �
       P�
             T             ��~      q       T�      �       P�      �       T      �       T�             T      �       Y�      �       T�             Y      �       T�      �       Y�      G       XG      :       Y:      d       Td      z       Yz      �       X�      �       Y�      �       X�      �       Y                          �
      �
       P�
      �       ��~�      �       P�      �       ��~      �       ��~                          �
      �
       t �
      �       S�      �       S      C       SH      G       SI      �       S                                                  �
      I       0�K      �       V�      �       p,�      �       V�      �       0��      �       V      �       0��      �       V�      �       0��      �      
 p q !
����      �       p 
����      �      $ s z 1$r "������"#��q !
����      �       V�      �      * s z 1$r "������"#��q !���"
����      �       0��             V             0�      !       p 
���!      �       0��      �       V                                                                                          �
      �
       r��
             P             P      )       t 1$����r "#�)      I       P�      �       r��      �       ^      1       P1      9       t 1$����r "q "#�9      I       PI      d       t 1$����r "q " "#�d      �       ^�             ^      +       ��+      W       VW      j       Pj      �       V�      �       P�      �       v q "��      �       P�      �      	 v q " "��             P      ,       PR      k       Pp      �       R�      �       ���      �       P�      �       s z 1$r "������"��      �       ^�      H       ��H      �       ^�      �       V�      �       P�      �       ���      N       P�      �       P�      �       P�             P      !       s z 1$r "������"�!      N       ��N      d       ^d      z       ��z      �       P�      �       ��                                                                  W       TW      �       x��      �       X�      �       x��             x�      �       X�      �       x��      A       YA      N       UN      �       Z�      �       X�      �       Z�             X             x�!      :       Td      z       Tz      �       Y�      �       u��      �       x��      �       Y�      �       p��      �       x�                        B             ^      �       Z�             ^�      �       Z                           W       ��W      �       P�             ���      �       P                       �             ��N      }       ^}      �       R�      �       ^                                             u 
���              U       -       ^-      }       [}      �       Q�      �       [z      ~       U~      �       ^�      �       ��                  V      �       ���      �       ��                    �             U      |
       �U�                    �             T      |
       ��                            �      �       Q�      c	       _c	      d	       �Q�d	      t	       _t	      u	       �Q�u	      |
       _                 �      �       u                  �      �       u #�u #�"�                    d      Y	       Vu	      |
       V                    \      Y	       [u	      |
       [                       �      )	       t 
���K	      R	       t 
���u	      M
       t 
���b
      |
       t 
���                       �      )	      ( q 1$��"��8$q 1$��"#��!0$0&�K	      R	      ( q 1$��"��8$q 1$��"#��!0$0&�u	      M
      ( q 1$��"��8$q 1$��"#��!0$0&�b
      |
      ( q 1$��"��8$q 1$��"#��!0$0&�                             -      2       0�2      )	       Q)	      C	       q�K	      R	       Qu	      :
       Q:
      M
       q�b
      |
       Q                       �      �       q 1%��      �       P�             q 1%�      (       t 1%�                         �      �       t �      Y	       Rd	      
       R
      u
       Rw
      |
       R                                             �      �       0��      	       P	      R	       0�R	      Y	       Pd	      �	       0��	      �	      
 x } !
����	      �	       x 
����	      �	      " r v 1$| "����z "#��} !
����	      �	       P�	      �	       0��	      �	       P�	      
       0�
      "
       P'
      R
       0�R
      b
       Pb
      |
       0�                  �             ~�      2       ~�                  -      2       U                      �	      �	       P�	      �	       r v 1$| "����z "�
      '
       r v 1$| "����z "�                                    y      5y       U5y      �z       _�z      �}       ��~�}      �}       _�}      �}       �U��}      �}       ��~�}      R~       _R~      `~       U`~      j~       _j~      �~       ��~�~             _                                  y      5y       T5y      �z       ^�z      �}       �T��}      �}       ^�}      �}       �T��}      R~       ^R~      ]~       T]~      j~       ^j~      �~       �T��~             ^                                                5y      5y       �5y      ty       �ty      ty       �ty      �y       �Sz      kz       R�z      �z       v~��z      Q{       Sm{      {{       V{{      |       X|      %|       ��%|      i|       v~�i|      �|       S�|      I}       ^I}      �}       v~��}      �}       S�}      �}       R�}      �}       |����1$���� "#��}      �}       ��}      �}       ��}      $~       �j~      �~       v~��~             �                                 Jy      Py       s 
���Py      hy       Sky      �z       S�z      �}       ���}      �}       S�}      �}       ���}      R~       Sj~      �~       ���~             S                           z      �z       ��z      �}       ��~#��}      �}       ��}      �}       �U#��}      �}       ��~#��}      �}       �j~      �~       ��~#�                      'z      *z       Q*z      �}       ��~j~      �~       ��~                    3z      �z       V�}      �}       V�}      �}       V                      3z      [z       Q[z      �}       ��~j~      �~       ��~                      ;z      ?z       P?z      �}       ��j~      �~       ��                      �y      �y       V�y      �y       v 1%�~      6~       V6~      R~       \                              y      �z       0��z      U}       ��Z}      �}       ���}      �}       0��}      �}       ���}      j~       0�j~      �~       ���~             0�                            �y      �y       R�y      z       Q�~      �~       Q�~      �~       R�~      �~       ��~�~      �~       Q                     �y      �y       y �8$x �!
����~      �~       y �8$x �!
����~      �~       ��~��8$��~��!
���                    �y      �y       } 
����y      �y      	 } 
��1%��~      �~       } 
����~      �~      	 } 
��1%�                          �z      j{       ]j{      m{       [�{      �}       ]�}      �}       ]j~      �~       ]                                �z      '{        
����{      |       P|      %|       ��%|      E|        
���i|      {|        
���I}      �}        
����}      �}        
���j~      s~        
���                           �z      �z       s 
����{      |       R|      %|       ��%|      i|       s 
���I}      �}       s 
���j~      �~       s 
���                                   kz      �z       0��z      �z       \�z      �z       Y�z      Q{       \Q{      m{       |�m{      I}       \I}      �}       Y�}      �}       \�}      �}       0��}      �}       \j~      �~       \                        kz      �z       0�Q{      j{       ]j{      |       [|      %|       ���}      �}       0�                        kz      �z       0�Q{      m{       Pm{      |       Z|      %|       ���}      �}       0�                               �z      Q{       ��~��8$��~��!0$0&��{      �{       | 1$��~"��8$t �!0$0&��{      |      ( | 1$��~"��8$| 1$��~"#��!0$0&�|      Q|       ��~��8$��~��!0$0&�i|      �|       ��~��8$��~��!0$0&�I}      �}       ��~��8$��~��!0$0&��}      �}       ��~��8$��~��!0$0&�j~      �~       ��~��8$��~��!0$0&�                           kz      �z       ��~�z      m{       ��~#�m{      m{       ��~m{      �}       ��~#��}      �}       ��~�}      �}       ��~#�j~      �~       ��~#�                           kz      �z       ��z      m{       ��~#�m{      �{       ��~#��{      �}       ��~#��}      �}       ��}      �}       ��~#�j~      �~       ��~#�                           kz      �z       ��~�z      m{       ��~#�m{      �{       ��~�{      �}       ��~#��}      �}       ��~�}      �}       ��~#�j~      �~       ��~#�                             kz      Q{       VQ{      {{       V{{      �{       X�{      �|       V�|      I}       ��~I}      �}       V�}      �}       Vj~      �~       V                  �|      �|       ]                      }      }      
 p r !
���}      }       p 
���}      }       p 
��s "
���}      +}       ~��r !
��s "
���                                  @             U      �       _�      �       U�             _      	       �U�	      $       U$      �       _�      �       �U��      �       _                 @      B       u                  @      B       u #�u #�"�                                        �       S�             (      	       �U#($      W       SY      w       Sw      �       (�      �       �U#(�      �       S�      �       S                                       �       � �      �       u� �      �       Q�             �       	       �U#H$      2       Q2      �       � �      �       �U#H�      �       �                               �       T�      �       <�      	       T$      �       T                             �       � �      �       u� �      	       U$      �       U                  �      	       Q                        �      �      
 p r !
����      �       p 
����      �       q��r !
����      	       P                     2      2       Q2      Y       0�j      �       Q�      �       0�                          U       TU      7       T                        7       Y                                        B      ^       Pf      u       Pu      }       t 1$����y "#�}      �       P�      �       t 1$����y "{ "#��      �       P�      �       t 1$����y "r "{ "#��      �       P�      �       r 1$t 1$����"y "{ "#��             P             r 1$t 1$����"y "{ "#�             P      $       r 1$t1$����"y "{ "#�$      /       P/      1       r 1$t 1$����"y "{ "#�                       7       X                        B      ^       q 
����      �       q 
����      �       0��             q 
���      1       q 
���                 �      �       u                  �      �       u #�u #�"�                 �             t�                  �      �       r�                    P      j       Uj      �       �U�                    P      j       Tj      �       Z                  Y      �       Y                         Y             0�      	       P	      {       0�{             P      �       0�                     Y             0�      	       X	      �       0�                            ]      �       X�      �       X	             X      *       X^      �       X�      �       X                          {      �       P�      �       P�              P.      ^       P�      �       P                           �      �       P�      �       p��      �       p��      �       p��              p�.      B       p�B      �       U�      �       p��      �       U                      �      �       [�              [.      �       [                        �      �       Q�              Q.      U       Q�      �       Q                       �      �       p��8$p��!0$0&��              p��8$p��!0$0&�.      ^       p��8$p��!0$0&��      �       p��8$p��!0$0&�                       �      �       p��8$p��!
����              p��8$p��!
���.      ^       p��8$p��!
����      �       p��8$p��!
���                         �      �       T�              T.      :       T�      �       T�      �       x ��                  �      �       T                      q      t      
 p q !
���t      x       p 
���x      �       u��q !
���                    �      �       U�      C       �U�                      �      �       T�      �       X�      C       �T�                   �      �       u�      �       U                     �      <       0�<      =       P=      C       0�                      �      �       P�              Q=      B       Q                     �      �       Q�      �       q��      �       q��             q�      =       U=      B       q�                          �      )       X)      ,      
 q r !
���,      9       q 
���9      =       u��r !
���=      B       X                         �      �       q ��8$q��!
����      �       t 8$q��!
����      �       u 8$q��!
����              q ��8$q��!
���=      B       q ��8$q��!
���                         �      �       q��8$q��!
����      �       t 8$q��!
����      �       u 8$q��!
����              q��8$q��!
���=      B       q��8$q��!
���                     �              q��8$q��!0$0&�       5       t �8$y �!0$0&�=      B       q��8$q��!0$0&�                    �             R=      B       R                      P      g       Ug      �       u�{��      �       �U�                      P      n       Tn      �       �T��      �       T                     Z      n       t ��n      �       �T���      �       t ��                         Z      j       t 8%�j      x       Rx      �       �T8%��      �       R�      �       t 8%�                        `      q       Qq      �       T�      �       Q�      �       t 8%1$����u "
 �                  g      �       U                   l      �       U�      �       P                                    �v      �v       U�v      �v       ]�v      	w       }�{�	w      ;w       �U�;w      Jw       ]Jw      Rw       }�{�Rw      �x       �U��x      �x       U�x      �x       ]�x      y       �U�                            �v      �v       T�v      Rx       ^Rx      Ux       �T�Ux      �x       ^�x      �x       T�x      y       ^                               �v      �v       }��v      �v       }��v      ;w       S;w      Jw       }�Jw      pw       Spw      vw       ]vw      vw       Svw      vw       s�vw      �w       s��w      �w       s��w      Px       ]Ux      xx       ]xx      �x       V�x      y       S                        �v      �v       p 
����v      �v       | 
���;w      Gw       p 
���Gw      Jw       | 
���                           �v      �v       0�pw      vw       Pvw      ;x       _;x      Jx       PJx      Tx       �Ux      �x       _                         �v      �v       0��v      ;w       \Jw      Nx       \Ux      �x       \�x      y       \                          �v      �v       S�v      ;w       }�|�Jw      Rw       }�|�Rw      �x       �U#��x      y       �U#�                   Jw      pw       S�x      y       S                          ^w      bw       Pbw      kw       Rkw      �x       ���x       y       R y      y       ��                            �v      �v       V�v      �v       v 3%��v      	w       P#w      ;w       VJw      Vw       PVw      pw       v 3%��x      y       v 3%�                 vw      �w       s ��8$s��!
���                        �w      �w      
 t p !
����w      �w       p 
����w      7x       v 
���Ux      gx       v 
���                 �w      �w       s��8$s��!
���                     �w      �w       s��8$s��!0$0&��w      7x       ����8$w ��!0$0&�Ux      xx       ����8$w ��!0$0&�                  x      x       T                  ]x      xx       X                        �x      �x      
 p t !
����x      �x       p 
����x      �x       p 
��q "
����x      �x       v��t !
��q "
����x      �x       v��v~��8$!
��q "
���                  $      D       r�                 �      �       u�             u#�                      �      �       X�             R             0�                 �             0�                       �      �       0��      �       P�             0�             P                 �      �       u                            p+      �+       U�+      �,       ]�,      �,       �U��,      H-       ]H-      �-       U�-      �/       ]                            p+      �+       T�+      �,       V�,      �,       �T��,      H-       VH-      a-       Ta-      �/       V                            p+      �+       Q�+      �,       \�,      �,       �Q��,      H-       \H-      ~-       Q~-      �/       \                           p+      �+       u�
��+      �,       }�
��,      �,       �U#�
��,      H-       }�
�H-      �-       u�
��-      �/       }�
�                      �+      ~,       _�,      �,       _H-      /       _                           �+      �+       0��+      ~,       6��,      H-       6�H-      �.       0��.      /       8�/      /       6�/      /       0�/      g/       6�g/      l/       0�l/      }/       6�}/      �/       0�                         �+      �+       }�
#�,      ?,       Q?,      G,       q�G,      R,       q~�R,      x,       Q�,      H-       S/      �/       S                   �+      �+       }��,      �,       P                     �+      �+       r s "#��+      	,      
 s ��"#�?,      x,       S                        �+      �+       P�+      x,       ^�,      H-       ^/      �/       ^                       	,      ,       x 8$��#	��!
���,      R,       ��#��8$��#	��!
���R,      k,       r 
���k,      x,       ��#��8$��#	��!
���                      /,      ?,       Pf,      n,       P�,      �,       P                        �,      �,       y 
����,      +-      
 ���
���/      F/       y 
���l/      �/       y 
���                  �,      �,      & s ��H$s��@$!s��8$!s��!�                 �,      �,      & s��H$s��@$!s��8$!s	��!�                    �-      �-       P�-      �.       ���.      �.       ��                    �-      �-       U�-      �.       ]�.      �.       ]                 �-      �.       ^�.      �.       ^                     �-      �-       P�-      �-       P�.      �.       0��.      �.       8�                  �-      �-       R�-      �-       r��-      �-       r��-      m.       r�m.      �.       Q�.      �.       q|��.      �.       Q                 �-      P.       r ��8$r��!
���                   �-      B.       y 
���B.      �.       T                  .      v.       P                 m.      {.       T                m.      �.       U                       {.      �.       q��8$q��!
����.      �.       p 8$q��!
����.      �.       p 8$q��!
����.      �.       q~��8$q��!
���                 �      �       u                  �      �       t                   �      �       u #                 �      �       t #                      @E      HE       UHE      hE       ShE      iE       �U�                 @E      AE       u8                          @B      qB       UqB      �D       S�D      �D       �U��D      0E       S0E      1E       U                    ^B      �D       V�D      0E       V                   ^B      �D       \�D      0E       \                 0C      ;C       U                   �B      �B       S�D      �D       S                     �B      �D       s�
��D      �D       �U#�
��D      0E       s�
�                 �D      �D       s�                 �B      �B       S                 �B      �B       s�                                                               j      �j       U�j      �l       V�l      �l       T�l      n       �U�n      =n       V=n      On       �U�On      Xn       VXn      �n       �U��n      fo       Ufo      zo       Vzo      �o       U�o      �o       V�o      p       �U�p      (p       V(p      �r       �U��r      �r       U�r      s       Vs      _t       �U�_t      jt       Ujt      �u       �U��u      �u       V�u      wv       �U�wv      �v       V                                               j      �j       T�j      Nn       _Nn      On       �T�On      �n       _�n      fo       Tfo      zo       _zo      �o       T�o      �q       _�q      �q       P�q      �r       V�r      �r       _�r      �r       T�r      _t       __t      jt       Tjt      �v       _                         j      ]j       Q]j      _t       �Q�_t      jt       Qjt      �v       �Q�                         j      Tj       RTj      _t       �R�_t      jt       Rjt      �v       �R�                         j      _j       X_j      _t       �X�_t      jt       Xjt      �v       �X�                                 �k      �k       P�k      n       ��~Xn      �n       ��~�o      q       ��~�r      �r       ��~jt      �t       ��~�t      *u       ��~wu      v       ��~Iv      �v       ��~                       �j      �j       1�fo      zo       1��r      s       0�wv      �v       0�                          �j      �j       0��j      �j       1�n      (n       0�(n      =n       ��~fo      zo       0��r      s       0�                      �j      �j       p  $0)�fo      zo       p  $0)�s      s       ]                      k      $k       p  $0)�$k      �k       ��~�0)�On      Xn       ��~�0)�                    %k      Ck       p  $0)�On      Xn       p  $0)�                	        j      _j       0�_j      �j       \�j      �j       R_t      jt       0�                
      j      _j       0�_j      �j       ^_t      jt       0�                              >j      =n       SOn      �r       S�r      s       S_t      �t       S�t      @u       Swu      v       SIv      �v       S                   >j      _j       0�_t      jt       0�                                   m      n       _�o      p       _(p      �q       _�q      �q       P�q      �r       V�r      �r       _s      _t       _jt      �t       _*u      wu       _v      Iv       _                                    m      Km       PKm      n       T�o      p       T(p      3p       T3p      Np       0�Np      gp       Pjt      �t       0��t      �t       p ���t      �t       R�t      �t       p ���t      �t       ��
0$0.��                       hp      }p       0�}p      �p       T�p      �p       t��r      �r       T                     hp      }p       0�}p      �p       [�r      �r       [                    �p      �p       U�r      �r       U                  �p      �p       X                  �p      �p       R                   �p      �p      
  
G     ��p      �p       P                   �p      �p      
 �
G     ��r      �r      
 �
G     �                      �p      �q       \�q      �r       ��~*u      @u       \                      q      /q       P/q      �r       ��~*u      @u       P                           q      5q       V5q      >q       �>q      �q       V�q      �r       _*u      ;u       V;u      @u       �                       q      >q       �>q      �q       ]�q      �r       ��~*u      @u       �                           q      �q       0��q      �q       P�q      �r       ��~�r      �r       P�r      �r       v�
*u      @u       0�                      �q      �q       ~��q      zr       ^zr      �r       ~�                      �q      hr       ��~qr      zr       Pzr      �r       ��~                  �q      r       ��~�����5$} "�                     �m      n       _�o      p       _(p      /p       _                      �m      n       fylg��o      p       fylg�(p      /p       fylg�                   �m      �m       P�m      �m       Q                      �m      n       R�o      p       R(p      /p       R                  �m      n       Q                 n      n       _                 n      n       2FFC�                   n      n       P�o      p       P                 n      n       R                       �n      fo       Tzo      �o       T�r      �r       T�r      s       _                      �n      fo       fylg�zo      �o       fylg��r      s       fylg�                   �n      o       Ro      Ao       P                          o      fo       Qzo      �o       Q�r      �r       Q�r      �r       t��
��5$t�"��r      �r       ��
��5$�"�                    Co      fo       Pzo      �o       P                  zo      �o       R                                              ��      ��       U��      �       _�      �       �U�'�      ��       �U���      �       _�      ��       �U���      ��       }��      5�       }�5�      ��       _��      ��       �U�w�      1�       �U�A�      b�       �U�:�      J�       _J�      ��       �U���      ª       �U�ª      ˪       }�                                    ��      ��       T��      �       ]�      ��       �T���      ��       T��      �       ]�      5�       �T�5�      ��       ]��      :�       �T�:�      J�       ]J�      ˪       �T�                        ��      ��       Q��      ��       ��~��      ��       Q��      ˪       ��~                        ��      ��       R��      ��       �R���      ��       R��      ˪       �R�                        ��      ��       X��      ��       �X���      ��       X��      ˪       �X�                    �      �       8���      ��       :�                        ��      �       S��      �       S5�      ��       S:�      J�       S                                               ��      �       ^�      �       ��~'�      ��       ��~��      ��       ^��      Ӟ       PӞ      �       ^�      S�       ��~�      5�       ��~5�      ��       ^��      ��       ��~w�      1�       ��~A�      ��       ��~:�      E�       PE�      J�       ^J�      ��       ��~��      ˪       ��~                            ��      ͟       P͟      ޟ       Q�      0�       P0�      5�      	  
��1�ª      ƪ       Pƪ      ˪      	  
��1�                 ��      ę       }�                    ř      ڙ       P`�      l�       P                  m�      {�       P                  E�      S�       P                        3�      y�       \��      ��       \��      բ       ��~b�      +�       \                    ��      ��       P��      +�       _                      ��      ��       R��      ܤ       ��~��      +�       R                      �      �       P�      ��       ^��      +�       ^                      �      2�       P��      �       Y�      &�       Y                                    i�      y�       0�y�      �       V��      ��       V��      ġ       0��      r�       Vr�      բ       ��~1�      <�       V?�      `�       P`�      +�       V��      ��       V                      p�      |�       P|�      ��       ��~��      +�       ��~                                7�      S�       _S�      �       w ��      ��       w ��      w�       w 1�      A�       w b�      ��       _��      :�       w ��      ��       w                 	                   3�      y�       0�y�      ��       _��      �       0���      ��       0���      ��       0���      �       P�      ��       _��      ��       Z��      բ       ��~1�      A�       0�b�      :�       0�                
                 3�      y�       0�y�      ��       ^��      �       0���      ��       0���      �       0��      :�       P:�      w�       ^1�      A�       0�b�      :�       0���      ��       ^                    S�      ]�       pp�]�      �       ��~@�                     W�      ��       [��      ��       \��      ʢ       \                      �      %�       Y%�      m�       \��      ��       \                       W�      ��       _��      ��       Z��      ��       ]��      ��       }|���      բ       ]                      W�      ��       0��      %�       0�%�      r�       ]��      ��       ]                                �      �       ]�      �       �T�'�      ��       �T��      ��       �T���      ��       �T�w�       �       �T�A�      b�       �T�J�      ��       �T���      ª       �T�                                    �      w�       _��      �       _'�      s�       _�      ��       _��      ��       _w�       �       _A�      b�       _J�      '�       _'�      ��       ��~��      ˧       ��~��      ��       _                                 �      �       P�      �       ��~'�      ��       ��~�      ��       ��~��      ��       ��~w�       �       ��~A�      b�       ��~J�      ��       ��~��      ª       ��~                        ;�      ?�       P?�      ^�       Q��      �       Q�      U�       Q                         3�      7�       P7�      |�       S��      �       S�      ��       Sw�      �       S                           k�      w�       ]'�      ٝ       ]ٝ      s�       ��~��      ��       ]A�      b�       ]J�      d�       ��~                               k�      w�       _'�      s�       _��      ��       _A�      b�       _J�      '�       _'�      ��       ��~��      ˧       ��~��      ��       _                            |�      w�       S'�      ȝ       Sȝ      s�       ��~��      ��       SA�      b�       SJ�      d�       ��~                                 ��      w�       0�w�      ��       [��      ��       0�'�      :�       0�:�      >�       P>�      i�       [i�      Ý       ��~s�      ��       0���      ��       0�A�      b�       0�                                  ��      w�       0�w�      ��       w ��      ��       0�'�      x�       0�x�      ��       P��      s�       w s�      ��       0���      ��       0�A�      b�       0�J�      ��       w ��      ª       w                                   ��      ܦ       Pܦ      �       y 2$y "2$#,��      1�       ��~52$#,�1�      ��       U��      �       U�       �       U �      �       Q�      I�       U��      ��       P                                        ��      ]�       0�]�      a�       Pa�      ��       V'�      J�       0�J�      ѝ       Vѝ      s�       ��~s�      ��       V��      ��       0���      ��       VA�      b�       VJ�      d�       ��~r�      ��       P��      ��       V��      ª       V                                ��      w�       0�w�      ��       ^'�      e�       0�e�      i�       Pi�      ��       ^��      ��       0���      ��       ^A�      b�       ^J�      ��       ^��      ª       ^                                   q�      ��       V��             v�      Ϝ       v�Ϝ      ܜ       v�ܜ      �       v��      �       v��      �       v��      �       v��      �       v��      �       v	��      "�       v
�"�      "�       v�"�      ѝ       v�ѝ      s�       ��~#�A�      b�       VJ�      d�       ��~#���      ��       \��      ��       ]��      ��       }���      ��       }q�]�      4�       ]��      ��       ]��      ��       ]��      ��       ]                              ��      �       R�      1�       ��~1�      ��       R��      C�       RC�      ��       ��~��      �       P��      ��       R                                    ��      ��       0���      �       ]�      ��       }��      \�       ]��      1�       0���      ��       0���      �       ��~"�      4�       R��      ��       ��~��      ��       0���      ª       ��~                
             ��      w�       0�'�      ��       0���      ��       S��      �       P�      �       S�      R�       S��      ��       0�A�      b�       0�                       ��      �       \�      4�       |P���      ��       \��      ª       \                         {�      ��       0���      ��       T��      ��       R��      ��       TA�      b�       0�                 ��             ���
��4$p �                          {�      ��       P��      ��       P��      ��       p 1%���      ��       PA�      [�       P[�      b�       Q                         ��      ��       \��      �       }3$v "�      s�       \J�      Z�       }3$v "Z�      d�       }3$w "                    ˦      ��       T��      ˧       T                    �      �       0��      �       S                              �<      >       U>      ->       �U�->      K>       UK>      ^>       �U�^>      ?       U?      s?       �U�s?      }?       U                              �<      >       T>      ->       �T�->      K>       TK>      ^>       �T�^>      ?       T?      s?       �T�s?      }?       T                        �<      5=       Q5=      U>       VU>      ^>       �Q�^>      }?       V                    =      W>       \^>      }?       \                           =      '>       0�'>      +>       P+>      ->       Q->      K>       0�K>      ^>       Q^>      }?       0�                         =      K=       0�K=      K=       QK=      S=       q�a=      �=       Qh>      �>       Q�>      �>       Q                                          =      K=       ZK=      �=       P�=      	>       z { "�	>      ->       S->      7>       P7>      G>       S^>      h>       Sh>      �>       P�>      �>       z x "��>      �>       S�>      �>       P�>      s?       Ss?      }?       P                             =      �=       	���=      �=       ���=      �=       [h>      �>       	���>      �>       ���>      �>       	���>      �>       ��s?      }?       ��                       =      K=       	��K=      G>       ��^>      �>       ���>      }?       ��                           =      K=       	��K=      �=       [h>      �>       [�>      �>       Q�>      �>       [s?      x?       [                              =      K=       	��K=      �=       S�=      �=       Q�=       >       S->      4>       Sh>      �>       S�>      �>       Ss?      }?       S                               =      K=       	��K=      >       X->      G>       X^>      s>       Xs>      x>       Qx>      �>       X�>      �>       Xs?      }?       X                	         =      K=       0�K=      >       ^->      G>       ^^>      �>       ^s?      }?       ^                              �=      �=       0��=      >      
  �C     �>      ->       ]->      G>       0�^>      h>       0��>      �>       0��>      �>      
 ��C     ��>      �>       0��>      s?       ]s?      }?       0�                  �>      s?       ^                    @3      ^3       U^3      �3       �U�                      @3      O3       TO3      j3       Pj3      �3       �T�                     @3      k3       0�k3      �3       P�3      �3       P                     [3      �3       S�3      �3       S�3      �3       S                    3      �3       Q�3      �3       Q                          s3      �3       0��3      �3       r p ��3      �3       p  r "��3      �3       r p ��3      �3       0�                      [3      3       V3      �3       T�3      �3       V                    �3      4       U4      �4       �U�                      �3       4       T 4      %4       P%4      �4       �T�                     �3      &4       0�&4      �4       P�4      �4       P                      4      �4       \�4      �4       \�4      �4       \                    Q4      l4       Q�4      �4       Q                          24      l4       0�l4      |4       u p ��4      �4       p  u "��4      �4       u p ��4      �4       0�                      4      C4       VC4      �4       R�4      �4       V                    �(      �(       U�(      �(       �U�                    �(      �(       T�(      �(       �T�                            �/      �/       U�/      �/       S�/      �/       �U��/      �/       S�/      �/       �U��/      0       S                            �/      �/       T�/      �/       \�/      �/       �T��/      �/       \�/      �/       �T��/      0       \                            �/      �/       Q�/      �/       V�/      �/       �Q��/      �/       V�/      �/       �Q��/      0       V                        �/      �/       P�/      �/       P�/      �/       6��/      0       P                    �              U      �       �U�                      �       R       QR      h       �Q�h      �       Q                     �              0�      F       Uh      �       U                                      P             p`�      A       PA      F       p`�h      �       P                    �       �        U�       �        q0�                 �       �        U                        �      �       U�      W�       VW�      f�       �U�f�      z�       U                        �      �       T�      W�       ]W�      f�       �T�f�      z�       T                       �      �       U�      W�       VW�      f�       �U�f�      z�       U                   �      W�       Ss�      z�       0�                   �      �       	��f�      f�       	��f�      z�       P                  :�      J�       P                     �      0�       �H�0�      9�       Q9�      :�       �H�                 �      :�       S                 �      :�       V                            �        T�       �        �T�                                        P?       @        PG       H        Po       p        P                      P�      z�       Tz�      ��       �T���      ��       T                  t�      ��       X                  t�      ��       R                  t�      ��       Q                    t�      z�       Tz�      ��       �T�                  t�      ��       U                              ��      ͊       U͊      Ί       �U�Ί      ي       Uي      ڊ       �U�ڊ      �       U�      �       S�      �       �U�                              ��      ͊       T͊      Ί       �T�Ί      ي       Tي      ڊ       �T�ڊ      �       T�      �       V�      �       �T�                         ��      ͊       U͊      Ί       �U��      �       U�      �       S�      �       �U�                    ��      �       V�      �       �T�                    ��      �       S�      �       �U�                  ��      �       P                      �      '�       U'�      (�       �U�(�      O�       U                          �      '�       T'�      (�       �T�(�      9�       T9�      N�       VN�      O�       �T�                     �      '�       U'�      (�       �U�(�      O�       U                    4�      N�       VN�      O�       �T�                  4�      O�       U                  I�      L�       P                      P�      g�       Ug�      h�       �U�h�      ��       U                          P�      g�       Tg�      h�       �T�h�      y�       Ty�      ��       V��      ��       �T�                     P�      g�       Ug�      h�       �U�h�      ��       U                    t�      ��       V��      ��       �T�                  t�      ��       U                  ��      ��       P                          ��      ��       U��      ��       S��      ��       �U���      �       S�      �       �U�                            ��      ��       T��      ��       Q��      ��       V��      ��       �T���      �       V�      �       �T�                     ��      ��       P��      Ջ       Pڋ      �       P                    ��      �       V�      �       �T�                    ��      �       S�      �       �U�                  ֋      �       P                                    `�      ��       U��      ��       S��      ��       �U���      $�       S$�      *�       �U�*�      j�       Sj�      p�       �U�p�      ��       S��      ��       U��      ��       S                                    `�      ��       T��      ��       ]��      ��       �T���      )�       ])�      *�       �T�*�      o�       ]o�      p�       �T�p�      ��       ]��      ��       T��      ��       ]                                    `�      ��       Q��      ��       V��      ��       �Q���      %�       V%�      *�       �Q�*�      k�       Vk�      p�       �Q�p�      ��       V��      ��       Q��      ��       V                    x�      ��       P��      ��       P                                 ��      ��       u����      ��       s����      ��       �U#����      $�       s��$�      *�       �U#��*�      j�       s��j�      p�       �U#��p�      ��       s����      ��       s��                            ��      ��       P��      ͑       P�      �       P*�      9�       Pp�      w�       P��      ��       P                            q�      ��       \��      '�       \*�      m�       \p�      ��       \��      ��       u���      ��       \                   ��      �       s��p�      ��       s��                  �      �       U                   *�      Z�       s����      ��       s��                      ��      Ԓ       UԒ      Ւ       �U�Ւ      �       U                      ��      Ԓ       TԒ      Ւ       �T�Ւ      �       T                      ��      Ԓ       QԒ      Ւ       �Q�Ւ      �       Q                      ��      �       U�      �       �U��      2�       U                      ��      �       T�      �       �T��      2�       T                            ��      �       Q�      ��       V��       �       �Q� �      �       V�      �       �Q��      2�       Q                            ��      �       R�      ��       S��       �       �R� �      �       S�      �       �R��      2�       R                 ��      2�       �Np	                       ��      �       T�      �       �T��      2�       T                     ��      �       U�      �       �U��      2�       U                     �      �       R�      ��       S �      �       S                     �      �       Q�      ��       V �      �       V                     �      �       T�      ��       �T� �      �       �T�                     �      �       U�      ��       �U� �      �       �U�                     �      ��       P �      �       P�      �       \                          �      )�       U)�      3�       S3�      5�       �U�5�      L�       SL�      R�       �U�                            �      �       T�      4�       V4�      5�       �T�5�      M�       VM�      Q�       UQ�      R�       �T�                      �      �       Q�      )�       T)�      R�       �Q�                  *�      Q�       P                  5�      R�       �Q�                      5�      M�       VM�      Q�       UQ�      R�       �T�                      5�      L�       SL�      Q�       q�}�Q�      R�       �U�                     5�      C�       s��C�      Q�       QQ�      R�       �U#��                                ��      ��       U��      ��       S��      ��       �U���      j�       Sj�      o�       }�{�o�      s�       q�{�s�      t�       �U�t�      �       S                                ��      ��       T��      ��       Q��      ��       \��      ��       �T���      m�       \m�      s�       Us�      t�       �T�t�      �       \                        ��      ��       P��      Θ       PΘ      ј       Vt�      �       P                        ��      m�       \m�      s�       Us�      t�       �T�t�      �       \                          ��      j�       Sj�      o�       }�{�o�      s�       q�{�s�      t�       �U�t�      �       S                          ј      ژ       Pژ      &�       V&�      G�       PH�      s�       Pt�      �       P                        ��      o�       ]o�      s�       Qs�      t�       �U#��t�      �       ]                              Ъ      �       U�      &�       \&�      T�       |�}�T�      [�       �U�[�      o�       \o�      w�       Uw�      ��       \                            Ъ      �       T�      X�       VX�      [�       �T�[�      o�       Vo�      t�       Tt�      ��       V                       �      �       |��      &�       |�&�      T�       |�}�T�      [�       �U#�[�      o�       |�                    �      �       p 
���[�      l�       p 
���                  �      T�       V                    �      &�       \&�      T�       |�}�                  �      T�       S                     �      (�       0�(�      9�      	 s | #��O�      T�      	 s | #��                      (�      5�       P9�      =�       s���=�      N�       P                        ��      �       U�      ��       w ��      ��       ����      ɰ       w                           ��      ܯ       Tܯ      6�       _6�      ��       ����      ��       _��      ɰ       ��                        ��      د       Qد      ��       S��      ��       �Q���      ɰ       S                        ��      �       R�      ��       V��      ��       �R���      ɰ       V                         �      �       0��      �       P�      s�       \s�      z�       T{�      ��       0���      ɰ       \                    $�      =�       \=�      i�       _��      ��       \                       ,�      L�       ^L�      P�       ~�P�      i�       ^��      ɰ       ^                     ,�      3�       P3�      =�      	 s�
�����      ��       P                 ��      ɰ       �] �                        а      �       U�      ٱ       w ٱ      �       ���      �       w                           а      �       T�      i�       _i�      �       ���      �       _�      �       ��                        а      ��       Q��      ݱ       Sݱ      �       �Q��      �       S                        а      �       R�      ޱ       Vޱ      �       �R��      �       V                         �      �       0��      ,�       P,�      ��       ]��      ��       T��      ձ       0��      �       ]                     I�      p�       ]p�      ��       _�      �       ]                       Q�      }�       ^}�      ��       ~~���      ��       ^�      �       ^                    W�      p�       R�      �       R                 а      �       �� �                                �      *�       U*�      <�       �U�<�      w�       Uw�      �       V�      $�       U$�      �       V�      �       U�      W�       V                      e�      {�       U{�      ��       VͲ      �       V                  |�      ��       p ��                   ��      Ȳ       ]��      �       P                       �      $�       U$�      �       V�      �       U�      W�       V                  �      W�       ^                        �      m�       S�      c�       Sp�      ��       Sڻ      #�       S                        ��      ��       p ��ڻ      ��       p ����      �       p ���      #�       p ��                           ��      ٴ       0�ٴ      ��       T��      )�       T��      �       Tc�      p�       T��      ڻ       T                  �      @�       0�                                        �      $�       0��      �       P�      m�       \��      ��       P��      ��       ]K�      `�       _`�      ��       ]�      2�       0�2�      >�       P>�      c�       \��      ��       Pڻ      #�       0�#�      >�       ]                                                       �      �       P�      @�       T@�      F�       t�F�      X�       TX�      m�       S��      ��       P��      �       S�      �       s��      �       [�      '�       s�µ      е       s�е      ��       S��      �       s��      (�       S(�      3�       s�3�      W�       SW�      b�       s�b�      ��       S��      ��       S��      ��       s���      ��       S[�      `�       S��      ��       T��      ��       t���      ��       ti��      +�       P+�      /�       T/�      @�       t�                      d�      �       \)�      `�       \>�      W�       \                      ��      ��       T)�      3�       T3�      <�       p                 ��      ��       p                 �      g�       R                          x�      ��       \��      )�       \��      �       \c�      p�       \��      ڻ       \                            ܵ      �       Q�      6�       Q:�      d�       Qd�      z�       Pz�      ��       R��      ��       R                        ��      �       s��      �       [�      '�       s�µ      е       s�                          ��      �       R�      �       Z�      �       R�      �       Zµ      е       R                                               ��      �       s��      `�       [`�      h�       Rh�      l�       r�l�      z�       R��      ��       [��      µ       Rµ      µ       s�µ      е       s���      ��       Z��      ڷ       [ڷ      �       P�      �       S�      ��       P��      )�       [��      ��       R��      �       [c�      p�       [��      ڻ       [                                �      '�       U'�      `�       S`�      z�       Q�      µ       S��      ط       S��      )�       S��      Һ       Sc�      k�       S��      ڻ       S                     �      �       r @%��      �       R'�      C�       RK�      ^�       Q                                �      ��       Z��      ��       P��      ��       p 
�����      µ       P��      ̷       P��      )�       P��      ��       0�Һ      �       Z��      Ȼ       P                               ��      ��       0���      ��       s  { "���      µ       s  r "���      ÷       s  r "�÷      ̷       { s ���      )�       { s ���      ��       s  { "���      Ȼ       { s �                     ��      ��       �[�`�      ��       �[�#�      >�       �[�                      ��      �       ����      +�       U+�      <�       u|�<�      @�       U                       ��      ��       �[�`�      ��       �[�@�      ��       �[�#�      >�       �[�                         ��      ��       ���`�      й       ���й      ��       X@�      ��       ���#�      >�       ���                       ��      ��       S`�      '�       S@�      ��       S#�      >�       S                       ��      ��       ]`�      ��       ]@�      ��       ]#�      >�       ]                     ��      ��       ]`�      ��       ]#�      >�       ]                            ��      �       P�      �       q ��      ��       ss s  $0-( 4&�`�      '�       ss s  $0-( 4&�@�      ��       ss s  $0-( 4&�#�      >�       P                                ��      �       �[��      ?�       T?�      D�       t u "�D�      ��       T�      *�       T*�      B�       R��      ��       r p '���      ˹       R˹      ܹ       Pܹ      ��       x #�      >�       �[�                              ��      �       �[��      f�       Uf�      i�       u z "�i�      ��       U�      D�       U��      ҹ       Tҹ      Թ       t p "�Թ      �       T�      ��       ��#�      >�       �[�                           ��      �       �[��      q�       Z{�      ��       Z��      s�       Z��      ҹ       Uҹ      ܹ       u p "�ܹ      ��       P#�      >�       �[�                                ��      �       �[��      ��       [��      ��       P��      ��       t p "���      ��       P��      ��       [{�      '�       ['�      ��       S˹      ��       Q#�      >�       �[�                     ��      ��       ��#�`�      ��       ��#�#�      >�       ��#�                     ��      ��       ����`�      ��       ����#�      >�       ����                     ��      ��       �J�8�`�      ��       �J�8�#�      >�       �J�8�                     ��      ��       ����`�      ��       ����#�      >�       ����                        ж      ��       X`�      ��       X@�      ��       X#�      >�       X                   ж      �       Q#�      >�       Q                       �      �       r �      $�       P$�      *�      
 p ����z�*�      <�       P<�      ��      * rp���#?$��������# %!����z�                       �      �       r�      Q�       rtQ�      Q�       PQ�      Z�      	 p �J�8�Z�      c�       Pc�      ��      * rt�����z@$��������# %!�J�8�                  �      �       r�      {�       rx                  	

     �      �       r�      {�       r|{�      {�       P{�      ��      	 p ��#���      ��       P��      ��      * r|�����z># $��������%!��#�                     ��      ��       X`�      ��       X@�      ��       X                             ��      ��       0�`�      �       0��      ��       P��      �       Q�      �       P�      �      
 p ����z��      �       P@�      ��       0�                             ��      ��       0�`�      ��       0���      Ƹ       PƸ      ׸       Q׸      �       P�      �      	 p �J�8��      �       P@�      ��       0�                             ��      ��       0�`�      ��       0���      ��       P��      ��       Q��      ��       P��      ��      
 p ����z���      ��       P@�      ��       0�                                 ��      ��       0�`�      b�       0�b�      i�       Qi�      r�       Pr�      x�      	 p ��#�x�      {�       P@�      e�       0�e�      t�       Qt�      ��       0���      ��       Q                  8�      ��       R��      ��       r p '�                  ��      ��       Q��      ��       T                ��      ��       U                  ��      ��       S��      ˹       Q                      �      �       u �      �       Q�      �       R&�      >�       Q                    A�      F�       PF�      Q�       [�Q�      c�       Q                            �       Q�      �	       �Q��	      �	       Q                          �       R�      �	       �R�                          J       XJ      �	       �X�                            r	       Yr	      �	       �Y��	      �	       Y                        }      e	       Se	      o	      & u0�X�R"u �Xu "�Ru0-( | �o	      �	      ( u0�X�R"u �Xu "�Ru0-( u���	      �	       S                  �      �	       Z                            f      �       r p ��      �      	 ��}�p ��      o	      	 ��}�| �o	      �	       ��}�u���	      �	       ��}�u���	      �	      	 ��}�| �                           .       0��      �       0��	      �	       0�                         f      }       S}      �       u0x u } u0-( ��      �       u0�Xr "u } u0-( ��      �       u0�X�R"u } u0-( ��      �	      # u0�X�R"u �Xu "�Ru0-( �                           f      �       Z�      �       ~ u(v { +( ��      �       ~ u(v u8+( ��      �       ~ u(�Xu("�Ru8+( ��      �	      # u8�X�R"u(�Xu("�Ru8+( ��	      �	       ~ u(v u8+( �                     f      �       X�      �       �Xr ��      �	       �X�R�                   �      [	       v�0$0&v�0$0& $ &�[	      e	       v��0$0&v��0$0& $ &�                           	      	       p r "#��@&q "�	      %	       v �0$0& r "#��@&q "�%	      .	       X.	      1	       v �0$0& r "#��@&q "�1	      [	      * v �0$0& v �0$0& ?&"#��@&��}"�[	      e	      , v��0$0& v��0$0& ?&"#��@&��}"�                          .	      1	       X1	      N	      3 v �0$0& v �0$0& ?&"#��@&p "} "��}"s �N	      R	      ; v �0$0& v �0$0& ?&"#��@&s  $ &��}"p "} "#�R	      [	      9 v �0$0& v �0$0& ?&"#��@&s  $ &��}"p "} "�[	      e	      ; v��0$0& v��0$0& ?&"#��@&s  $ &��}"p "} "�                     .	      1	       S1	      N	       PN	      R	       p�                �      	       T                �      	       v �0$0&�                   	      	       P	      	      
 p r "#���                  	      	       p ?&�	      	       R                        w	      �	       S�	      �	       s��	      �	       S�	      �	       S                          w	      �	       P�	      �	       P�	      �	       s 2$� "
<�	      �	       s2$� "
<�	      �	       P                      w	      �	       R�	      �	       R�	      �	       R                                          �v      w       Uw      w       u�w      w       Uw      <w       u�<w      Bw       u�Tw      _w       U�w      �w       U�w      �w       R�w      �w       Ux      8x       u�8x      <x       u�<x      Ux       u�}x      �x       U�x      �x       u�                      �v      _x       T_x      }x       �T�}x      �x       T                            �v      w       Qw      �w       V�w      �w       �Q��w      zx       Vzx      }x       �Q�}x      �x       V                                  �v      Bw       RBw      �w       \�w      �w       �R��w      x       \x      (x       R(x      |x       \|x      }x       �R�}x      �x       \�x      �x       R                 �v      �v       t�                                 w      -w       Q-w      4w       p O��Bw      x       Qx      x       p ��x      8x       QBx      fx       Q}x      �x       Q�x      �x       p ���x      �x       Q                                           �v      Gw       0�Gw      �w       X�w      �w       p ���w      �w       X�w      �w       P�w      �w       X�w      �w       p O���w      �w      
 s �O���w      x      
 s~�O��x      x       Xx      Ux       0�Ux      fx       X}x      �x       p ���x      �x       X�x      �x       0�                            �v      w       Qw      �w       V�w      �w       �Q��w      zx       Vzx      }x       �Q�}x      �x       V                     -w      Bw       1�x      %x       3�+x      <x      
 u  s "x "��x      �x       2�                         �w      �w       2��w      �w      	 z r u "��w      �w      	 z r u "��w      x       1�x      x       0�}x      �x       3�                                  �I      J       UJ      fL       ���fL      �L       �U��L      KM       ���KM      )O       �U�)O      �O       ����O      
S       �U�
S      OS       ���OS      `V       �U�                    �I      jJ       TjJ      `V       �T�                    �I      J       QJ      `V       �Q�                    �I      (J       R(J      `V       ���                                    �I      K       XK      fL       ���fL      �L       �X��L      KM       ���KM      )O       �X�)O      DP       ���DP      
S       �X�
S      $S       X$S      OS       ���OS      `V       �X�                     
J      iL       0�iL      �L       ^�L      �L       P�L      `V       0�                      J      uJ       QuJ      K       ���#
S      $S       ���#                 J      \J       Q                   J      LJ       SLJ      \J       ���                \J      \J       ���                \J      \J       �Й�                                 \J      K       XK      fL       ����L      M       ���M      M       ����
(!�M      -M       ����	�
(!�-M      1M       Q1M      KM       ����	�
(!�)O      �O       ����O      DP       ����	�
(!�
S      $S       X$S      OS       ���                  \J      iL       ����L      `V       ���                         \J      �K       S�K      fL       ����L      �L       ���)O      OO       ���
S      OS       S                              \J      fL       ���fL      iL       �U��L      KM       ���KM      )O       �U�)O      �O       ����O      
S       �U�
S      OS       ���OS      `V       �U�                  \J      iL       �Й��L      `V       �Й�                                                    iL      iL       ^�L      �L       ����L      M       0�M      M       P5M      KM       PKM      �M       ^�M      )O       ^=O      OO       ���OO      �O       0��O      �O       P�O      S       ^JS      OS       0�OS      �S       ^�S      T       PT      �T       0��T      �U       ^�U      �U       0��U      V       ^V      >V       0�>V      `V       ^                      jJ      �J       T�J      K       s�
S      $S       s�                      uJ      K       Q
S      S       QS      $S       s�#P                         uJ      �K       V�K      fL       �Ș�L      �L       �Ș)O      OO       �Ș
S      OS       V                           zJ      }J       R}J      K       v�K      iL       ����L      
S       ���
S      $S       v�$S      `V       ���                           �J      �J       R�J      K       v�K      iL       ����L      
S       ���
S      $S       v�$S      `V       ���                                �J      K       ���K      iL       �Ț��L      M       �Ț�M      M       UM      
S       �Ț�
S      $S       ���$S      �S       �Ț��S      �S       T�S      `V       �Ț�                        �L      �L       ]�L      )O       _=O      OO       0�OO      
S       _OS      `V       _                   �L      �L        OO      �O                              �L      )O       ]OO      
S       ]OS      `V       ]                  K      K       ���
S      JS       S                  K      K       ���
S      JS       ���                  K      K       �Й�
S      JS       �Й�                    K      K       0�
S      (S       0�(S      JS       PJS      JS       0�                   K      fL       A��L      �L       A�)O      =O       A�                   K      fL       ��	  �L      �L       ��	  )O      =O       ��	                     K      fL       ����L      �L       ���)O      =O       ���                 K      �K       �ؙ                               K      wK       0�wK      �K       _�K      �K      	 y 3$| "# �K      �K       V�K      6L       0�6L      8L       |���"�
�?
��#3$| "8L      WL       0�WL      ^L       P^L      fL       V�L      �L       V�L      �L       ])O      =O       0�                               K      WK       A�WK      ^K       y 
�?
���^K      oK       u 1$p "�
�?
���oK      �K       u 1$|"�
�?
���L      L       } 
�?
���L      .L       q s "�
�?
���.L      6L       |s "�
�?
���6L      8L       |���"�
�?
���                          wK      �K       Z�K      L       S6L      fL       S�L      �L       S)O      5O       S                      fK      �K       [�K      fL       _�L      �L       _)O      =O       _                       �K      8L       ^LL      fL       ^�L      �L       ^)O      =O       ^                �M      �M                       �M      �M       v� �v� ��                   �M      �M       P�M      �M      
 p t "#���                  �M      �M       p ?&��M      �M       T                �M      �M                          �M      �M       R�M      �M      
 p r "#���                  �M      �M       r ?&��M      �M       P                     �N      �N       P�T      �T       P�T      U       �ؙ                   �N      �N       ����T      �T       ���                �N      
O                       �N      
O       v�                    �N      
O       Q
O      
O      
 q r "#���                  �N      
O       q ?&�
O      
O       R                U      <U                       U      <U       v�                    :U      <U       P<U      <U      
 p q "#���                  :U      <U       p ?&�<U      <U       Q                   �O      TR       _>V      `V       _                   �O      �Q       S>V      `V       S                   �O      TR       �Й�>V      `V       �Й�                   �O      OR       0�>V      `V       0�                      �O      �O       P�O      TR       ���>V      `V       ���                   �O      *P       Y*P      �P       ���                 nP      �P        #�����3$�.G     "                      P      P       p�P      �Q       ���#�>V      `V       ���#�                  P      P       | 0$����0$.�                      &P      *P       P*P      TR       �Ș>V      `V       �Ș                      DP      qP       PqP      TR       ���>V      `V       ���                  �P      �P       p @$�����                  Q      !Q       P                �P      �P       ���#                   �P      �P       p @$��P      �P       P                   �P      �P       P�P      �P      
 p q "#���                  �P      �P       p ?&��P      �P       Q                  �Q      �Q      	 q �����                  �Q      �Q       P                �Q      �Q       |                  �Q      �Q       Q                   �Q      �Q       P�Q      �Q      
 p q "#���                  �Q      �Q       p ?&��Q      �Q       Q                �S      �S       �К                �S      �S       v�                   �S      �S       Q�S      �S      
 p q "#���                  �S      �S       q ?&��S      �S       P                  T      �T       �����U      �U       ����                    9T      |T       R|T      �T       ���                      NT      hT       QhT      |T      & ���� $ &51$���� $ &"3$r "X�|T      �T      ) ���� $ &51$���� $ &"3$���"X�                  VT      �T       P                 VT      �T       Y                 VT      �T       Z                  \T      �T       U                  `T      �T       T                 �U      �U       T                �U      �U       ���                  (V      >V       T                 (V      >V       ���                 iL      �L       �Й�                 �      �       U                    `/      e/       Ue/      j/       �U�                    `/      i/       Ti/      j/       �T�                              �V      �V       U�V      �W       Y�W      �W       �U��W      �W       Y�W      X       �U�X      ?X       Y?X      QX       �U�QX      �X       Y                  �V      �V       T                                                    �V      �W       Q�W      �W       S�W      �W       Q�W      �W       S�W      �W       �Q��W      �W       Q�W      X       SX      X       �Q�X      X       QX      X       SX      X       �Q�X      %X       Q%X      )X       S)X      6X       Q6X      QX       SQX      \X       Q\X      �X       S�X      �X       Q                          �V      �W       0��W      �W       0��W      X       PX      @X       0�@X      QX       PQX      �X       0�                              �V      �V       U�V      �W       Y�W      �W       �U��W      �W       Y�W      X       �U�X      ?X       Y?X      QX       �U�QX      �X       Y                                 �V      �V       u�V      �W       y�W      �W       y�W      �W       yX      X       yX      'X       y)X      ?X       yQX      ^X       y�X      �X       y                                 �V      �V       u�V      �W       y�W      �W       y�W      �W       yX      X       yX      'X       y)X      ?X       yQX      ^X       y�X      �X       y                                 �V      �V       u �V      �W       y �W      �W       y �W      �W       y X      X       y X      'X       y )X      ?X       y QX      ^X       y �X      �X       y                      �W      �W       Q�W      X       SX      X       �Q�                  �W      �W       Q�W      �W       S                 �W      �W       y�����3$@*G     "                   X      X       SX      X       �Q�                   )X      6X       Q6X      QX       S                 %X      )X       S                 QX      �X       y$�                   QX      \X       Q\X      �X       S                  �W      �W       Q                 �W      �W       S                          `V      �V       U�V      �V       S�V      �V       �U��V      �V       S�V      �V       U                            `V      �V       T�V      �V       V�V      �V       �T��V      �V       T�V      �V       V�V      �V       T                          `V      �V       Q�V      �V       �Q��V      �V       Q�V      �V       �Q��V      �V       Q                      `V      �V       0��V      �V       0��V      �V       P�V      �V       0�                    7      67       U67      Y7       �U�                      7      ,7       T,7      M7       ZM7      Y7       �T�                    7      F7       QF7      Y7       �Q�                      7      07       R07      X7       VX7      Y7       �R�                      %7      07       rp �07      C7       r p �C7      M7       R                   %7      I7       s p �I7      M7       X                  O7      Y7       P                     $      _       R_      ~       t0~      �       R                     $      w       Pw      ~       u�(~      �       P                     $      -       0�-      :       q ��:      �       Q                  �      �       Z                 �      �       U                 �      
       T                            �#      K$       UK$      �$       _�$      �$       [�$      �(       �U��(      �(       U�(      )       _                          �#      F$       TF$      �$       w �$      �(       �T��(      �(       T�(      )       w                         $      $       S$      �$       ���$      �(       �T����
�	�U"#H��(      )       ��                       $      �%       0��%      �%       P!&      k(       0�z(      )       0�                              4$      C$       SC$      K$       u K$      O$        O$      �$       ���(      �(       S�(      �(       u �(      )       ��                     4$      F$       t ����
0Iv "#P�F$      �$       w �����
0Iv "#P��(      �(       t ����
0Iv "#P�                   4$      O$       R�(      �(       R                       4$      X$       0��(      �(       0��(      �(       S�(      �(       ��~                     4$      �$       \�$      �$       S�(      )       \                      7$      &'       ]z(      �(       ]�(      )       ]                                     �$      �$       \�$      K&       SK&      �&       \�&      '       R'      '       R'      &'       P4'      A'       [A'      i(       Pz(      �(       S�(      �(       P�(      )       \                    C$      X$       S�(      �(       u                              �$      �$       P�$      �$       U�$      �$       P�$      �&       Vz(      �(       V�(      �(       P�(      )       V                      X$      w(       ^z(      �(       ^�(      )       ^                      r$      z$       Pz$      �$       ���(      )       ��                   �$      .&       0�z(      �(       Q                  /%      O%       0�                     O%      y%       Qy%      ~%       q��z(      �(       Q                      Z%      ~%       Pz(      �(       P�(      �(       u u r  $0-( �                   �%      &      	 p 0$0&�&      &       q �0$0&�                      &      	&       P	&      &      
 p r "#���&      &       P                   &      	&       p ?&�	&      &       R                     K&      Y&       0�Y&      �&       0��&      �&       Q                  a&      �&       0�                     �&      �&       Q�&      �&       q���&      �&       Q                      �&      �&       P�&      �&       P�&      �&       u u r  $0-( �                 �&      �&       �T����
�	�U"#`                    �&      k(       V�(      �(       V                       �&      �&       �T����
�	�U"#`�&      &'       Q&'      i(       T�(      �(       T                     &'      A'       0�A'      i(       Z�(      �(       Z                     &'      A'       0�A'      i(       S�(      �(       S                      q'      �'       x � $0.�(      '(       0��(      �(       x � $0.�                        �'      �'       Q(      '(       Q�(      �(       Q�(      �(       Q                       �'      �'       p �'      �'       R(      '(       p �(      �(       R�(      �(       U                  �'      �'       X                  �'      �'       U                r$      �$       S                r$      �$       w �����
0Iv "#��                   �$      �$       P�$      �$      
 p q "#���                  �$      �$       p ?&��$      �$       Q                    0      �       U�      �       �U�                    0      �       T�      �       �T�                    0      �       Q�      �       �Q�                    0      �       R�      �       �R�                     0      �       r ����
�	u "#H��      �       �R����
�	u "#H��      �       �R����
�	�U"#H�                  M      �       X                  \      �       Z                      u      �       v 8&��      �       \�      �      / �U#�(#H�����8&1�U#�(#H�����8&0.( �                    �      �       V�      �       �U#�(#H�����
p;&�                  k      �       ]                     �      �       X�      �       T�      �       X                    �      �       R�      �       P                   �      �      	 u 0$0&��      �      	 u 0$0&�                        �      �       r�0$0&��      �       r��0$0&��      ,       P,      �       r�0$0&�                 �      �       t�0$0&��      �       t�0$r�0$+( 0$0&�                 �      �       t�0$0&��      �       t�0$r�0$-( 0$0&�                  $      �       Y                      /      8       P8      >       _>      �       r�0$0&u �                  g      �       _                  {      �       P                    I      ]       P]      g       r�0$0&u :$} 
 �                        P      {       U{      |       X|             �U�      @       X                      P      |       T|             �T�      @       T                 P      R       u�(                       P      {       t ����
�	u "#H�{      |       t ����
�	x "#H�|             �T����
�	�U"#H�      @       t ����
�	x "#H�                        t      x       Px      {       u {      |       x       @       x                             t      �       0��      �       ��~�      6       0�6      ;       Re      �       0��      �       ��~�      I       0��      %       0�%      %       ��~7      �       0��      �       R�      @       0�                                    t      |       0�|      `       [`      �       _�      �       [�             [6      �       [�             [I      }       [}      �       0��      %       [%      %       0�7      �       [�             Q"      >       [�             [      @       0�                                �      �       P�      �       U�      ;       x� ;      #       ��~a      {       P{      "       ��~�             ��~      @       x�                       �      �       P�      |       ��~      @       ��~                            C       UC      |       ��~      @       U                                            ;       U;      |       ��~|      �       ��}�      �       \�      I       ��}I      �       \�             ��}      %       \7      P       \P             ��}"      �       \�             ��}      @       U                      �      �       P�      |       ��~      @       ��~                           )       P)      6       p��6      ;       P                                x,� $ &Pp "�      ;       x,� $ &Px0"�                                    x0      )       P)      6       p��6      @       P                       @       x,� $ &Px0"�                                 �      �       P�      �       ��~�      #       ��}#      %       S7             S"      �       S�      �       ��~�             Q             P                       �      �       Q�      �       ��~#H�      #       ��}�      �       Q�             ��~#H                                        �      #       0�#      `       V`      d       0�d             V      �       1��      `       V`      �       1��      ;       V;      e       1�e      �       V�      }       1�}      �       0��             1�      %       V7             V"      �       V�             0�                              �      #       
 }��      �       PR      `       {� #0`      �       P;      e       P�      �       P<      <       P             P�             
 }�                                   �      #        ���      �       QV      `       {� #0`      �       P;      e       P�      I       QI      �       P�      �       Q<      <       Q             Q�              ��                            �      #       
 }�#      �       RV      �       R;      e       R�             RP      �       R�             
 }�                                     �      #        ��#      �       TV      �       R�      �       T;      e       Re      I       TI      �       R�      �       T�      %       T7      �       T"      :       T�              ��                            �      #       0�#      �       ^�      �       ^V      �       ^;      �       ^�      %       ^7             ^�             0�                                    �      #       0�#      �       ��}�      �       ��}V      �       ^�      �       ��};      e       ^e      I       ��}I      �       ^�      �       ��}�      %       ��}7             ��}�             0�                	                 �      #       
 }�#      �       X`      �       
 }��      �       X;      e       Re      I       XI      f       
 }��      �       R�      %       X7      �       X�             
 }�                
                   �      #        ��#      �       U`      �        ���      �       U;      e       Re      I       UI      f        ���      �       R�      %       U7      �       U"      0       U�              ��                                 �      #       0�/      `       ��}d      k       ��}{             ��}�      �       ��}�      ;       ��}e      I       ��}�      %       ��}7      P       ��}"      h       ��}                           �      #       0�#      =       _T      `       [`      %       _7             _"      �       _�             0�                        �      #       
 }�T      �       P*      /       p } -( �             P�             
 }�                        �      #        ��T      �       Q%      /       q { +( �             Q�              ��                                    �      #       
 }�#      `       ��}d             ��}�      T       ��}T      �       R�      �       ��}�      ;       ��}e      I       ��}�      �       ��}�      %       ��}7             ��}"      h       ��}�             
 }�                                    �      #        ��#      `       ��}d             ��}�      T       ��}T      �       T�      �       ��}�      ;       ��}e      I       ��}�      �       ��}�      %       ��}7             ��}"      h       ��}�              ��                                    �      #       0�#      `       ��~d             ��~�      T       ��~T      �       ^�      �       ��~�      ;       ��~e      I       ��~�      �       ��~�      %       ��~7             ��~"      h       ��~�             0�                                       �      #       0�#      `       ��~d             ��~�      T       ��~T      ]       _]      �       ��}�      �       ��~�      ;       ��~e      I       ��~�      �       ��~�             ��}      %       ��~7             ��~"      h       ��~�             0�                                    �      #       
 }�#      `       ��~d             ��~�      T       ��~T      �       X�      �       ��~�      ;       ��~e      I       ��~�      �       ��~�      %       ��~7             ��~"      h       ��~�             
 }�                      		              �      #        ��#      `       ��~d             ��~�      T       ��~T      �       U�      �       ��~�      ;       ��~e      I       ��~�      �       ��~�      %       ��~7             ��~"      h       ��~�              ��                            �      �       Y�      7       s0�      /       s0�             s0<      k       s0             s0                            �      �       Y�      7       s8�      /       s8�             s8<      k       s8             s8                      �      �       �4
  �      6       �4
  e      �       �4
        %       �4
  7      P       �4
  "      �       �4
                         �      �       ��~�      6       ��~e      �       ��~      %       ��~7      P       ��~"      h       ��~                      �      �       �T����
�	�U"#H��      6       �T����
�	�U"#H�e      �       �T����
�	�U"#H�      %       �T����
�	�U"#H�7      P       �T����
�	�U"#H�"      �       �T����
�	�U"#H�                              �      �       0��      �       [�      6       0�6      6       [e      �       0��      �       [      %       0�7      P       0�"      �       0��      �       [                        �             Q      %       Q7      P       Q"      5       Q5      >       ��~��~"#L                             �      �       Q�             Z      6       ��}      %       Q7      K       ZK      P       p q "#�"      >       Z>      h       ��}                      �      ;       ����      %       ����7      P       ����"      �       ����                  �      �       Q                  �             X                          �      �       q� �      �       qp�      �       T�             q�              qp                    �      �       U�             U                            �      �       R�      �       q� #8�      �       qp#8�      �       R�             q� #8             qp#8                      �      �       P�             P             u8                 �      �       q� #H�      �       u�                  �      �       q� #H�             u�                         p-      �-       U�-      �-       S�-      �-       U�-      �-       �U�                        p-      �-       T�-      �-       V�-      �-       T�-      �-       �T�                                )      w)       Uw)      Y*       SY*      h*       �U�h*      �*       S�*      
+       U
+      T,       ST,      �,       y��~��,      e-       S                        )      s)       Ts)      �*       �T��*      
+       T
+      e-       �T�                                )      �)       Q�)      Y*       ^Y*      h*       �Q�h*      �*       ^�*      
+       Q
+      T+       ^T+      �,       �Q��,      e-       ^                        5)      Y*       _h*      T+       _�,      L-       _L-      R-       PR-      e-       _                    5)      a*       \h*      e-       \                                     5)      w)       q ����
0Iu "#P�w)      �)       q ����
0Is "#P��)      Y*       ~ ����
0Is "#P�Y*      h*       �Q����
0I�U"#P�h*      �*       ~ ����
0Is "#P��*      
+       q ����
0Iu "#P�
+      T+       ~ ����
0Is "#P�T+      T,       �Q����
0Is "#P�T,      �,       �Q����
0Iy "
�J��,      �,       �Q����
0Is "#P��,      e-       ~ ����
0Is "#P�                              m)      �)       0��)      �)       P�)      �)       0��)      �)       Q�)      *       q�*      !*       Qh*      j*       0�
+      T+       0��,      �,       0�                         m)      Y*       s���h*      �*       s���
+      T,       s���T,      �,       y�|��,      e-       s���                   m)      �)       0�h*      j*       0�j*      t*       p ����Hs "#���                   �*      �*       Q�,      �,       Q                   �*      �*       (��*      �*       P                   �*      �*       P�,      �,       P                  �*      �*       R�,      �,       R                     �*      �*       P�*      �*       s#�#�
����,      �,       s#�#�
���                    �,      �,       T�,      -       r t +( �-      -       T                  C-      C-       TC-      e-       t 	��                  �,      e-       P                     -      -       p  �-      #-       Q#-      3-       p  �                 -       -       T                       -      '-       T'-      /-      
 q t "#���/-      3-       t ?&t "#���                  -      3-       t ?&�                	j*      �*       _                	 j*      t*       p ����Hs "#Ȗ�                   �*      �*       P�*      �*      
 p q "#���                  �*      �*       p ?&��*      �*       Q                  �)      !*       R                �)      *       r                    �)      *       P*      *      
 p x "#���                  �)      *       p ?&�*      *       X                 l+      �+       ^                     �+      �+       R�+      �+       P�+      �+       q                    �+      �+       P�+      �+      
 p t "#���                  �+      �+       p ?&��+      �+       T                �+      �+       T�+      �+      
 t  "#���                �+      �+       _                !*      8*       ~ ����
0Is "#��                   6*      8*       P8*      8*      
 p q "#���                  6*      8*       p ?&�8*      8*       Q                        �      D�       UD�      b�       Vb�      k�       �U�k�      _�       V                        �      >�       T>�      a�       Sa�      k�       �T�k�      _�       S                       �      M�       0�M�      d�       \d�      k�       Pk�      _�       0�                        2�      9�       P9�      ]�       w ]�      k�       ��k�      _�       w                  ��      T�       S                 ��      T�       V                       ��      Ӓ       0�Ӓ      1�       ]1�      @�       1�@�      T�       ]                     ��      G�       1�G�      O�       PO�      O�       1�O�      T�       0�                        Ò      Ӓ       0�Ӓ      1�       ��1�      B�       PB�      T�       ��                     Ò      �       ����      �       Q�      T�       ���                     Ò      ��       ^��      �       P�      T�       ^                   �      B�       _O�      T�       _                ��      �       0�                    ��      �       ����      �       R�      �       ���                ��      �       ���                ��      �       V                 ��      �       v�                  �      �       _                    @�      ��       U��      �       ��w                    @�      a�       Ta�      �       ��w                           ��      ͅ       0�ͅ      ��       ��w��      {�       ��w{�      ��       ��w�#���      �       ��w��      А       ��w!�      �       ��w                             ��      ͅ       0�ͅ      7�       ��w7�      J�       ��w�#�J�      N�       PN�      ��       ��w��      �       ��w��      А       ��w!�      �       ��w                     ̌      ،       ��w#�������H��w"#���،      �       { ����H��w"#���ȍ      ؍       ��w#�������H��w"#����      1�       { ����Hs "#���                  ��      ��       P                   ��      ��       u�����      �      	 ��w#���                                    ��      ��       v��v���v��v��v�����      Ї      ; ��w#�#����w#�#���X���w#�#����w#�#���Ї      �      E ��w#�#����w#�#�����w#�#����w#�#����w#�#�����      �      E ��w#�#����w#�#�����w#�#����w#�#����w#�#����      {�      ; ��w#�#����w#�#���X���w#�#����w#�#�����      ܋      ; ��w#�#����w#�#���X���w#�#����w#�#���܋      �       v��v���v��v��v���1�      �      ; ��w#�#����w#�#���X���w#�#����w#�#�����      А      ; ��w#�#����w#�#���X���w#�#����w#�#���!�      �      ; ��w#�#����w#�#���X���w#�#����w#�#���                        ��      ��       S��      |�       ��w��      ��       P��      �       ��w                    ��      ��       P��      �       ��x                     ��      �       ��x��      �       Q�      �       ��x�                                      ��      ͅ       Sͅ      �       [�      �       P�      R�       [R�      J�       ��wJ�      v�       [��      �       ��w�      �       [1�      �       ��w��      А       ��w!�      �       ��w                     ̌      ،       ��w#�������H��w"#���،      �       { ����H��w"#���ȍ      ؍       ��w#�������H��w"#����      1�       { ����Hs "#���                     ̌      ،       ��w#�������H��w"#Ȗ�،      �       { ����H��w"#Ȗ�ȍ      ؍       ��w#�������H��w"#Ȗ��      1�       { ����Hs "#Ȗ�                                   ��      ͅ       0�ͅ      Ї       S�      k�       Sk�      ��       \�      \�       S\�      �       ��w{�      ��       S��      ҋ       ��w܋      �       S�      1�       \                                   ��      ͅ       0�ͅ      Ї       ]�      v�       ]v�      ��       V�      T�       ]T�      �       ��w{�      ��       ]��      ȋ       ��w܋      �       ]�      1�       V                 r�      ��       T                             R�      j�       0�r�      V�       0���      ��       0���      �       0�1�      �       0���      А       0�!�      �       0�                                      ��      ��       	����      �       Z�      G�       RG�      X�       PX�      l�       Rl�      ~�       Z~�      ��       R��      ��       P��      Ї       Z�      �       Z��      ܋       Z܋      �       	��1�      Վ       Z                                ��      ��       0���      Ї       w �      {�       w ��      ܋       w ܋      �       0�1�      �       w ��      А       w !�      �       w                                   ��      ��       0���      e�       ��wl�      Ї       ��w�      {�       ��w��      ܋       ��w܋      �       0�1�      �       ��w��      А       ��w!�      �       ��w                           �      >�       ��wR�      V�       ��w��      �       ��w1�      �       ��w��      А       ��w!�      �       ��w                             �      R�       0�R�      �       ��w�      V�       ��w��      �       ��w1�      �       ��w��      А       ��w!�      �       ��w                               �      R�       0�\�      Ї       \�      V�       \�      _�       \_�      �       ��w{�      ��       \��      ܋       ��w܋      �       \                                    ��      ��       0���      G�       UG�      T�       p  $ &4$x "#T�      ��       U��      ��       p  $ &4$x "#��      �       U��      {�       U��      ܋       U܋      �       0�1�      �       U��      А       U!�      E�       U                               j�      Ї       0�Ї      �       P��      �       P�      {�       0���      �       0�1�      �       0���      А       0�!�      �       0�                    ��      ��       0�܋      �       0�                        ��      ��       0���      Ї       [�      a�       [܋      �       0�                      �      Ї       T�       �       T �      a�       {�                   ��      h�       Z~�      ��       Z                                    �      ,�       P,�      0�       p�0�      4�       �:�      T�       PT�      X�       p�X�      \�       �~�      ��       P��      ��       p���      ��       ���      ��       P                                Q�      a�       Qa�      �       ]�      �       ��w��      ��       ��w��             ]      ܋       ��w1�      Î       ��wÎ      Վ       z  $ &4$x "                                       Z�      a�       Ta�      o�       Ro�      x�       Tx�      ��       R��      ��       [��      �       t v  $t  $-( ��       �       t��w�v  $t  $-( ���      ċ       Rċ      ܋       [F�      V�       PV�      Y�       p�Y�      ��       P                                   Z�      a�       Ta�       �       Z �      (�       T(�      3�       [3�      ��       T��      Ǌ       {w �  ${  $+( ���      ��       T��      ��       {}   ${  $+( ���      ��       {w �  ${  $+( ���      ܋       Z                               Q�      a�       Ta�      o�       Ro�      É       TÉ      �       R�      �       ��w�      {�       R��      ��       ��w��      ܋       T1�      ��       ��w                                       Q�      a�       Ta�       �       Z �      (�       T(�      {�       [{�      P�       Te�      t�       T��      ��       [��      ܋       Z1�      ��       T��      Վ       VՎ      �       ��x��      А       ��x!�      �       ��x                                                Z�      a�       Ra�      ω       Sω      މ       Rމ      �       S�       �       ��w �      ��       R��      ��       T��      ��       R��      {�       ��w��      ��       R��      ��       ��w��      ͋       S͋      ܋       ��w1�      �       ��w��      А       ��w!�      ё       ��wۑ      ߑ       ��w                                                Z�      a�       Ra�      ى       \ى      މ       Rމ      ��       \��       �       ��w �      ��       \��      ��       T��      ��       \��      {�       ��w��      ��       \��      ��       ��w��      ׋       \׋      ܋       ��w1�      �       ��w��      А       ��w!�      Ƒ       ��wۑ      �       ��w                                                          a�      o�      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&���      ��       P��      ��       { 4$x "#u y 'y ���      ��      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&���      �      x t v  $t  $-(  $ &4$x "#u t v  $t  $-(  $ &4$x "#u ?&'t v  $t  $-(  $ &4$x "#u ?&��       �      � t��w�v  $t  $-(  $ &4$x "#u t��w�v  $t  $-(  $ &4$x "#u ?&'t��w�v  $t  $-(  $ &4$x "#u ?&� �      (�       yu yu ?&'yu ?&�O�      a�       Pa�      �       yu yu ?&'yu ?&��      �       t  $ &4$x "x q "��      �       t  $ &4$x "r  $ &4$x "���      ��       yu yu ?&'yu ?&���      ܋      0 { 4$x "#u { 4$x "#u ?&'{ 4$x "#u ?&�1�      D�       t  $ &4$x "r  $ &4$x "�D�      ��      " t  $ &4$x "��w� $ &4$x "���      ��      " v  $ &4$x "��w� $ &4$x "���      W�       PW�      [�      0  4$x "#y  4$x "#y ?&' 4$x "#y ?&���      ��       P!�      *�       P*�      M�      0  4$x "#y  4$x "#y ?&' 4$x "#y ?&�M�      ]�      6  4$x "#��w 4$x "#��w?&' 4$x "#��w?&�                            �      �       _1�      =�       _=�      �       ��w��      А       ��w!�      &�       ��w&�      �        ��w#H�������Q %3%�����                               w�      ��       T��      Վ       VՎ      b�       ]b�      ��       V��      Ϗ       ]��      ��       ]��      А       V!�      U�       ]U�      �       ��w                                   w�      ��       T��      ��       V��      ��       P��      �       V��      А       V!�      q�       Vq�      ȑ       Tȑ      ۑ       Vۑ      ��       T��      �       V                                 w�      Վ       0�Վ      W�       1�W�      b�       Pb�      ��       0���      ��       1���      �       P��      ��       1���      А       0�!�      �       1�                        ��      ��       	����      ��       VĐ      А       V]�      �       Q                       ��      ��       	����      А       V]�      ��       Z��      ۑ       Vۑ      �       Z                 w�      ��       ��w                     9�      [�       s { +�!�      /�       s { +�/�      ]�        4$x "{ +�                             q�      u�       p 4$x "#��w�u�      ȑ       t 4$x "#��w�ȑ      ۑ       v 4$x "#��w�ۑ      �       t 4$x "#��w��      ��       v 4$x "#��w���      ��       t 4$x "#��w���      �       v 4$x "#��w�                j�      r�       �$
                  j�      r�       0�                j�      r�       \                j�      r�       ��x�                j�      r�       ��w                j�      r�       ��w#@                 r�      r�       T                 �      T�       { ����H��w"#��                 �      T�       { ����H��w"#Ȗ                 �      3�       r q +�                      �      
�       1�
�      ;�       X;�      ?�       x�                 +�      /�       x ����x����3$p "                      L�      ��       1���      ��       X��      ��       x�                 ��      ��       x ����x����3$p "                      ِ      ��       R�      �       P�      �       R                  �      �       p��      �       P                        �      ,�       1�,�      ��       [��      ��       {���      ��       \                  ,�      F�       [                    S�      s�       U��      ��       U                    [�      s�       T��      ��       T                    ��      ��       Q��      �       ��w#@                    ��      ň       Pň      �      	 ��w#@#                 ��      ň       0�                         �      \�       U\�      �       S�      �       �U��      @�       S                       �      v�       Tv�      k�       \k�      @�       �T�                      ҂      �       PY�      k�       P~�      ��       P                 v�      ��       0���      т       T                            k�      *�       \*�      6�       |�;�      ��       0���      ڄ       1�ڄ      �       2��      ��       0���      �       1��      @�       \                 g�      @�       ���}�                	   g�      j�       Pj�      v�       s                 
   g�      j�       p�����3$ -G     "j�      v�       s #�����3$ -G     "                     g�      ��       ���|���      ��       Q��      @�       ���|�                    v�      ��       P��      т       P                ��      ��       0�                ��      ��       ���|�                ��      ��       S                ��      ��       s�                  ��      ��       T                   k�      6�       |  $ &
0Is "#P��      @�       |  $ &
0Is "#P�                   k�      6�       |  $ &
�	� "
���      @�       |  $ &
�	� "
��                    ��      	�       P�      @�       P                        ��       �       U �      �       }� � $ &54$}� "��      �       }�l� $ &54$}�l"��      @�       U                          ă      ��       Q��      �       p �      �       pP�      �       Q�      @�       p                   �      @�       Q                       ;�      ��       s� ���      �       s����      �       �U#����      ��       s� ���      �       s���                          Z�      ��       R��      ��       s���      ބ       R��      ��       R��      �       s�                   A�      ;�       V�      @�       V                 A�      T�       P                  C�      g�       Q                    C�      Y�       ���|�Y�      g�       V                    ph      th       Uth      uh       �U�                    ph      th       Tth      uh       �T�                    ph      th       Qth      uh       �Q�                    ph      th       Rth      uh       �R�                    �      �       T�      �       �T�                    �#      �#       U�#      �#       �U�                    �#      �#       T�#      �#       �T�                        ��      Ӂ       UӁ      ��       V��      ��       �U���      �       V                        ��      ́       T́      �       S�      ��       �T���      �       S                    ȁ      ��       \��      �       \                          �@      A       UA      `A       �U�`A      �A       U�A      �C       �U��C      �C       U                          �@      A       TA      `A       ��`A      �A       T�A      �C       ���C      �C       T                        �@      A       X`A      �A       X�C      �C       P�C      �C       X                      �@      A       Z`A      �A       Z�C      �C       Z                         �@      A       Y$A      B       Y�B      �B       Y�C      �C       Y�C      �C       Y                    �@      _A       _`A      �C       _                              A      A       8�A      :A       ]�A      �A       4��A      �A       ]�A      �C       ]�C      �C       8��C      �C       4�                                                                  �@      �@       X�@      �@       P�@      �@       p���@      A       PA      A       ^5A      HA       XHA      LA       x��LA      lA       XlA      xA       PxA      �A       p���A      �A       P�A      �A       ^�A      �A       S�A      �A       X�A      �A       x���A      �A       X�A      B       SB      %B       P%B      ;B       p� �@B      PB       VPB      TB       TTB      �B       V�B      �B       p� �:C      :C       P:C      IC       p� ��C      �C       P�C      �C       X                      A      :A       \�A      �A       \�A      �C       \                          A      A       ^�A      �A       ^�A      �A       S�A      �A       ^�A      gC       ^�C      �C       ^                        %B      �B       P�B      �B       ���B      "C       P:C      \C       P�C      �C       P                   �B      :C       V�C      �C       V                   �B      "C       P�C      �C       P                   �B      :C       v���C      �C       v��                 bB      �B       S                   bB      �B       P�B      �B       ��                 bB      �B       \                  �B      �B       S                  �B      �B       P                    �B      �B       T�B      �B       s��                  �B      �B       ^                   XC      �C       S�C      �C       s��                 XC      �C       \                 XC      gC       ^                            gC      xC       ^xC      C       ~��C      �C       ^�C      �C       S�C      �C       s���C      �C       S                    \C      `C       p s8�`C      �C       P                    �      >       U>      s!       �U�                        �      >       T>      /        ^/       >        �T�>       s!       ^                 �      �       u0                 �      �       u,� $ &Pu0"�                       �      >       t ����
�	u "#H�>      /        ~ ����
�	�U"#H�/       >        �T����
�	�U"#H�>       s!       ~ ����
�	�U"#H�                    �      5        V>       s!       V                  �      >       X                            9        ]9       >        	�0�T $0)( 	�#�>       s!       ]                    >      /        S>       s!       S                               i      w       Vw      �       x��F       Z        Vn       �        x���       �        Z�       �        y 3$v "��       �        Z�       	!       Zi!      s!       x��                                    i      �       \       "        P>       F        PF       X        \X       Z        Pi       x        \x       z        Pz       d!       \d!      i!       Pi!      s!       \                        i      �       PF       T        Pi       t        Pz       �        Pi!      n!       P                     i      �       \F       Z        \n       s!       \                        n      w       t | �w      �       | x��0$0&�F       Z        t | �n       7!       | x��0$0&�\!      s!       | x��0$0&�                       �      �       0�z       �        0��       	!       Ui!      s!       0�                             �      �       q X�z       �        q X��       �        [�       �        T�       �        [�       	!       Ti!      s!       q X�                          �       �        T�       �        P�       �        T�       �        T�       	!       P                       �       �        Y�       �        z �0$0&��       �        Y�       	!       Y                      �      �       0��      �       Ui!      s!       0�                      �      �       [	!      7!       [7!      \!       ��                 �      �       P                 �      �       | u 0$0&�                   �              P              
 p t "#���                  �              p ?&�               T                                �	      s
       Us
             S      �       ���      h       Sh      {       �U�{      �       ���      �       �U��      M       S                                    �	      s
       Ts
      x       ^x      �       ���      �       T�      `       ^`      {       �T�{      �       ���      �       �T��      &       T&      M       ^                       �
             s0      �       ��M      h       _{      �       ��                         L
      h
       u8h
      s
       u(�      �       s8�      �       s(�      �       s8             s(      &       s8                                             L
      e
       Pe
      h
       t �0$0&�h
      ~
       Q�      �       P�      �       p}��      �       ~ �0$0&��      �       _�             Q.      2       R2      M       _�      �       P�             t �0$0&�             Q      &       P&      =       Q                       
      h       \h             s�      h       \�      M       \                       
      e       ]e             s�      h       ]�      M       ]                              
      
       P
      s
       us
      m       ���      �       s�      h       ���      &       s&      M       ��                              '
      *
       P*
      s
       u s
      �       ���      �       s �      �       ���      &       s &      M       ��                     '
      P       V�      Y       V�      M       V                                      C             s0      �       PM      h       _{      �       P3      �       S�      �       R�      �       R             Q3      �       P�      �       p���      �       P�      "       _Q      �       _�      �       S                                  N       RN      �       w M      h       R{      �       w "      Q       w �      �       w                            "       p#��
���"             s�(##��
���M      h       s�(##��
���                          C      X       PX      �       ��M      U       PU      h       ��{      �       ��                     C      �       [M      h       [{      .       [                     C      �       YM      h       Y{      .       Y                         C      ]       x ]      x       ~x             ��#M      h       x �      �       q 1$s "                           C      �       UM      c       Uc      h       z 2$z "4$ "�{      �       U�      �       T�      �       U                             C             U      �       T�      �       t� �      �       TM      c       Uc      h       z 2$z "4$ "�{      �       P�      �       U�      �       T                       C             0�      �       _M      h       0�{      �       _                 �      �       p�0$0&t�0$0& $ &�                 �      �       p�0$0&t�0$0& $ &�                        $       R$      $      
 r s "#���                        $       r ?&�$      $       S                  >      E       QE      E      
 q r "#���                  >      E       q ?&�E      E       R                        Q      h       Q�      �       Q�             qx�      .       Q                              c      h       P�      �       P�      �       U�      .       R.             _"      Q       _�      �       _                      c      h       X�      �       X�             x~�      .       X                      c      h       0��      �       0��      �       P             P                      +              \"      Q       \�      �       \                     +              ^"      Q       ^�      �       ^                     +             _"      Q       _�      �       _                      3      �       S�              R"      Q       R�      �       S                     �      �       R�              Q"      Q       Q                            7      �       R�      �       T�      �       R�      �       T�      �       R�      �       s�                       �      �       R�      �       P�              P"      Q       P                                                  I      X       s�0$0&u  $ &�X      ]       P]      �       s�0$0&u  $ &��      �        s�0$0&s� #�0$0& $ &��      �       u t�0$0& $ &��      �       P�      �       u t�0$0& $ &��      �        s�0$0&s� #�0$0& $ &��      �       0��             Y              y u "�       �       Y�      �       z ��             0�"      6       Y6      ;       z �;      L       YL      Q       T�      �       s�0$0&u  $ &��      �        s�0$0&s� #�0$0& $ &�                                             I      i       s�0$0&x  $ &�i      s       Qs      �       s�0$0&x  $ &��      �        s�0$0&s� #�0$0& $ &��      �       x t�0$0& $ &��      �       Q�      �       x t�0$0& $ &��      �        s�0$0&s� #�0$0& $ &��      �       0��      �       T�      �       0��              T"      0       T0      ;       t �;      C       T�      �       s�0$0&x  $ &��      �        s�0$0&s� #�0$0& $ &�                       o      �       T"      0       T0      ;       t �;      C       T                          o      �       Y�      �       z �"      6       Y6      ;       z �;      L       YL      Q       T                    �      �       T0      ;       T                   0      6       Y6      ;       z �                   �      �       Y-      ;       	��                     {      �       s {�0$0& $ &��      �       p�0$0&{�0$0& $ &��      �       pH�0$0&{�0$0& $ &�                   {      �       p�0$0&{�0$0& $ &��      �       pJ�0$0&{�0$0& $ &�                     {      �       z�0$0&s  $ &��      �       z�0$0&p�0$0& $ &��      �       z�0$0&pH�0$0& $ &�                   {      �       z�0$0&p�0$0& $ &��      �       z�0$0&pJ�0$0& $ &�                  {      �       Z                 {      �       [                  s      �       ]                  �      �       ^                      �-      �-       U�-      �.       S�.      �.       �U�                      �-      .       0�.      t.       1�t.      �.       2�                   �-      �-       u� ��-      .       s� �.      �.       s��                                @             U      a       \a      h       �U�h      }       \}      �       U�             \      3       U3      �       \                        @             T      ^       S^      h       �T�h      �       S                                @             Q      c       ]c      h       �Q�h      }       ]}      �       Q�             ]      '       Q'      �       ]                                @             R      _       V_      h       �R�h      }       V}      �       R�             V      3       R3      �       V                                    @      s       Xs      }       �X�}      �       X�      �       �X��      �       X�      �       U�      '       �X�'      3       X3      [       U[      �       �X�                                    @      v       Yv      e       ^e      h       �Y�h      }       ^}      �       Y�      �       ^�      �       Y�      '       ^'      J       YJ      �       ^                         f      �       0��      �       Q�      %       q� �%      }       Q}      �       0�                       �       |                         �      �       Q'      .       Q.      3       u3      E       QE      [       |                             �      �       Q�             _'      .       Q.      3       u3      >       _>      C       p q "#�C      �       _                   �             ]t�'      �       ]t�                          �.      �.       U�.      U/       VU/      [/       T[/      \/       �U�\/      ]/       U                    �.      W/       \W/      [/       U                 
/      @/       s @*G     "                 
/      )/      # s @*G     "#�����3$�.G     "                        �F      �F       U�F      �F       V�F      G       �U�G      �I       V                        �F      �F       T�F      �F       w �F      G       ��G      �I       w                           �F      �F       Q�F      �F       \�F      G       �Q�G      �G       \�G      �I       �Q�                 �F      �F       u�                         �F      �F       0��F      �F       P�F      G       _G      G       r G      �I       _                uG      �I       _                   �G      �G       P�I      �I       0�                  uG      ~G        ~G      �I       V                     zG      �G       P�G      �G       v��G      �I       ��                  zG      �I       S�I      �I       ��                      �G      �G       |�H      =I       \=I      AI       |�                     zG      �G       0�`I      }I       \}I      �I       |�                 zG      �G       	��                 H       H       P                 H       H       p�����3$ -G     "                        H      �H       ^�H      �H       X�H      �H       ��1I      JI       X                            H      /H       X/H      AH       ��AH      QH       XpH      H       X�H      �H       P�H      �H       X                           �H      �H       T�H      I       ^I      I       TI      %I       ^%I      )I       P)I      4I       ^                  kI      }I       P                  �I      �I       0�                 �      �       U                 �      �       T                        @1      �1       U�1      �2       �U��2      �2       U�2      �3       �U�                              @1      �1       T�1      �2       ]�2      �2       �T��2      �2       T�2      I3       ]I3      N3       �T�N3      �3       ]                            @1      d1       Qd1      �2       _�2      �2       �Q��2      M3       _M3      N3       �Q�N3      �3       _                              @1      �1       R�1      Z2       ^Z2      �2       �R��2      �2       R�2      3       ^3      N3       �R�N3      �3       ^                        @1      �1       X�1      �2       �X��2      �2       X�2      �3       �X�                          �1      �1       | v ��1      �1       R�1      �2       | v ��2      E3       | v �N3      �3       | v �                      �1      �1       P�1      �2       Q�2      �3       Q                         �1      Z2       | v "2~ "�Z2      �2       | v "2�R"��2      3       | v "2~ "�3      E3       | v "2�R"�N3      �3       | v "2~ "�                              �1      �2       R�2      �2       rr��2      �2        | v "?%v "| "1&q ?%q "1&�R"��2      �2       p r "��2      .3       R.3      23        | v "?%v "| "1&q ?%q "1&�R"�23      73       p r "�N3      �3       R�3      �3       | v "?%v "| "1&q ?%q "1&~ "�                                  �1      `2       T`2      �2       q r "��2      �2       q r ">��2      �2      # | v "?%v "| "1&q ?%q "1&q "�R"��2      3       T3      .3       q r "�.3      E3      # | v "?%v "| "1&q ?%q "1&q "�R"�N3      �3       T�3      �3      " | v "?%v "| "1&q ?%q "1&q "~ "�                                 �1      �1       r ?��1      B2       PB2      T2       r ?�T2      f2       s x �f2      �2       ^�2      3       P3      3       r ?�N3      R3       PR3      �3       r ?��3      �3      " | v "?%v "| "1&q ?%q "1&~ "?�                                 �1      	2      	 @r ?�	2      c2       Xc2      �2       P�2      3       X3      3      	 @r ?�N3      W3      	 @r ?�W3      �3       X�3      �3      	 @r ?��3      �3      % @| v "?%v "| "1&q ?%q "1&~ "?�                        �1      l2       Ul2      �2       [�2      3       UN3      �3       U                           �1      -2       @u �-2      ?2       Z?2      i2       @u �i2      �2       T�2      3       @u �N3      �3       @u �                               �1      �2       0��2      �2       P�2      �2       P�2      3       0�3      +3       P23      N3       PN3      �3       0��3      �3       P                     ?2      T2       q ?�T2      y2       ZW3      ~3       q ?�                         @1      �1       @��1      �2       S�2      �2       @��2      D3       SN3      �3       S                      0      M       UM      �       �U��      �       U�      �       �U�                      0      M       TM      �       �T��      �       T�      �       �T�                  0      M       0��      �       0�                    0      M       b�M      �       Y�      �       b�                      0      M       QM      k       Pn      �       P�      �       Q                              �       R�      �       r/��      �       R�      �       rQ�                  S      �       T                     S      _       q t �_      {       R{      �       u q t q t 0-( �                      �      �       T�             u�(      #       T                       �      �       Q�      �       t0�             u�(#0      #       Q                       �      �       R�             r 4!�             R             Q      #       R                         �      �       0��      �       p ���             P             u�(      #       P                 �      #       U                 �      �       T                    �             U      ~       �U�                    �      p       Tp      ~       �T�                    �             Q      ~       �Q�                     �             q ����
�	u "#H�             q ����
�	�U"#H�      ~       �Q����
�	�U"#H�                  
      ~       Y                    .      �       S�      ~       ��                   .      p       �Q����
P9t "#P�p      ~       �Q����
P9�T"#P�                   .      p       �Q����
P9t "#Pp      �       �Q����
P9�T"#P                      L      Y       PY      �       Q�      ~       ��                  �      �       0�                    �      �       0��      d       _                      �      �       ���      K       ]N      d       ]                   �      R       PR      d       pH�                   �      �      
 q 2 $0.��      N       p0�2 $0.�                 �      N      ' y�8$8& $�Q����
�	�U"#h� $)�                           $       t { �$      '       QC      N       Q                        N       [                 $      -       Q                   -      4       Q4      4      
 q r "#���                  -      4       q ?&�4      4       R                .      9       �Q����
P9t "#P�                .      9       t� ��-(�-� �                   7      9       P9      9      
 p q "#���                  7      9       p ?&�9      9       Q                        `#      �#       U�#      �#       S�#      �#       U�#      �#       �U�                        `#      �#       T�#      �#       V�#      �#       T�#      �#       �T�                        �!      �!       U�!      !#       �U�!#      5#       U5#      U#       �U�                        �!      �!       T�!      !#       �T�!#      5#       T5#      U#       �T�                    �!      �!       Q�!      U#       �Q�                    �!      C#       _D#      U#       _                    �!      ?#       ]D#      U#       ]                         �!      �!       q ����
P9u "#P��!      �!       �Q����
P9u "#P��!      !#       �Q����
P9�U"#P�!#      5#       �Q����
P9u "#P�5#      U#       �Q����
P9�U"#P�                     �!      �!       0��!      !#       \D#      U#       \                       �!      "      ! | ����8�Q����
P9"�U"#��"      "      ! |����8�Q����
P9"�U"#��"      !#      ! | ����8�Q����
P9"�U"#��D#      U#      ! | ����8�Q����
P9"�U"#��                   z"      �"       p q "#��@& $ &��"      �"        s �r  $ &v q "#��@& $ &�                      �"      �"       p q ��"      !#       RD#      U#       R                                       �"      �"       p q ��"      �"       R�"      �"       Q�"      �"       P�"      �"       R�"      �"       q p ��"      �"       Q�"      #       sp �#      #       PD#      L#       PL#      P#       p 	��P#      S#       PS#      U#       p �                �"      �"       _�"      	#       _                 �"      �"       R�"      �"       q p �                      �"      �"       P�"      �"      
 p q "#���#      	#       Q	#      	#      
 p q "#���                    �"      �"       p ?&��"      �"       Q#      	#       q ?&�	#      	#       P                 "      *"       _                 "      *"       P                   #"      *"       Q*"      *"      
 q r "#���                  #"      *"       q ?&�*"      *"       R                W"      ^"       _                W"      ^"       R                  W"      ^"       Q^"      ^"      
 q t "#���                  W"      ^"       q ?&�^"      ^"       T                x"      z"       _                  x"      z"       Pz"      z"      
 p q "#���                  x"      z"       p ?&�z"      z"       Q                        P�      s�       Us�      ��       V��      ��       �U���      ��       V                        P�      m�       Tm�      ��       S��      ��       �T���      ��       S                    h�      ��       \��      ��       \                        �{      �{       U�{      �}       ]�}      �}       �U��}      i�       ]                    �{      �{       T�{      i�       ��x                         0|      0|       0�0|      p}       Vp}      u}       v�u}      �}       V�}      c       V�      �       VB�      i�       V                     0|      0|       0�0|      �}       ��x�}      �       ��x�      �       ��x�#��      i�       ��x                         0|      0|       1�0|      �}       \�}      �}       \�}      �}       0��}      �~       \�      �       \b�      i�       \                           (       ��x#������8��x"#��(      c       s ����8��x"#���      �       ��x#������8��x"#��B�      b�       s ����8u "#��                  �|      �|       P                    0|      0|       P0|      �}       ��x�}      i�       ��x                              �|      �|       q��q���q���q����|      �|       ~�#��~�#���Y��T���|      g}      0 ��x#�#����x#�#���Y����x#�#���g}      �}      : ��x#�#����x#�#�����x#�#�����x#�#����}      :~      0 ��x#�#����x#�#���Y����x#�#����      �      : ��x#�#����x#�#�����x#�#�����x#�#���b�      i�       q��q���q���q���                 �{      �{       u                     �{      �{       p�{      �{       u #                    �{      �}       _�}      i�       _                     �{      `|       ��y�`|      g|       Qg|      i�       ��y�                            |      p|       Sp|      �|       P�|      �}       S�}      �~       S�      �       Sb�      i�       S                           (       ��x#������8��x"#��(      c       s ����8��x"#���      �       ��x#������8��x"#��B�      b�       s ����8u "#��                           (       ��x#������8��x"#��(      c       s ����8��x"#���      �       ��x#������8��x"#��B�      b�       s ����8u "#��                 w|      �|       T                        �|      �|       0��|      g}       R�}      :~       Rb�      i�       0�                                �|      �|       	���|      }       Q!}      N}       QQ}      g}       Q�}      �}       Q�}      '~       Q*~      :~       Qb�      i�       	��                    �|      �|       0�b�      i�       0�                        �|      �|       0��|      }       P�}      �}       Pb�      i�       0�                        �|      �|       T�|      ,}       u�=}      g}       u��}      :~       T                            }      ,}       P=}      _}       P�}      �}       P�}      �}       p�~      *~       P*~      .~       p�                r|      w|       0�                r|      w|       ��y�                r|      w|       ]                r|      w|       }�                  w|      w|       T                 p      �       s ����8��x"#�                 p      �       s ����8��x"#�                 p      �       p r -�                      :~      X~       1�X~      �~       X�~      �~       x�                 {~      ~       x ����x����3$p "                      �~      �~       1��~             X             x�                 �~      �~       x ����x����3$p "                        �x      �x       U�x      g{       Sg{      o{       �U�o{      �{       S                      �x      �x       T�x      �y       \�y      �{       �T�                      Ry      �y       P�y      �y       P�y      z       P                 �x      @y       0�@y      Qy       T                            �y      �z       \�z      �z       |��z      {       0�{      Z{       1�Z{      o{       2�o{      x{       0�x{      �{       1��{      �{       \                 �x      �{       ��~�                	   �x      �x       P�x      �x       s                 
   �x      �x       p�����3$ -G     "�x      �x       s #�����3$ -G     "                     �x      &y       ��}�&y      0y       Q0y      �{       ��}�                    �x      0y       P1y      Qy       P                ;y      @y       0�                ;y      @y       ��}�                ;y      @y       S                ;y      @y       s�                  @y      @y       T                   �y      �z       |  $ &
P9s "#P��{      �{       |  $ &
P9s "#P�                   �y      �z       |  $ &
�	� "
P���{      �{       |  $ &
�	� "
P��                    z      �z       P�{      �{       P                        (z      �z       U�z      �z       }� � $ &54$}� "��z      �z       }�l� $ &54$}�l"��{      �{       U                          Dz      `z       Q`z      dz       p dz      sz       pP�{      �{       Q�{      �{       p                   �{      �{       Q                       �z      {       s� �{      g{       s�� �g{      o{       �U#�s�o{      x{       s� �x{      �{       s�� �                          �z      !{       R!{      %{       s�%{      ^{       Rx{      {       R{      �{       s�                   �y      �z       V�{      �{       V                 �y      �y       P                  �x      �x       Q                    �x      �x       ��}��x      �x       V                                  9        U9       �       w �      �       �@�      �       w �      �       U                                    9        Q9       z       ^z      �       �Q��      �       ^�      �       Q�      �       �Q�                                9        1��       �        1��      �       y��      �       U�      �       1�                  �       �        V�      �       V                            �       �        0��       '       V8      =       U=      E       VE      N       QN      V       q�V      z       Q�      �       V                    �       z       \�      �       \                    �       �        0��              P�      �       0�                      M       S       	 �Y�p�g       �        �Y�U��       �       	 �Y�p�                                p/      �/       Q�/      �/       �Q��/      �/       Q�/      0       �Q�0      E0       QE0      �0       �Q��0      �0       Q�0      51       �Q�                              p/      �/       R�/      0       �R�0      0       R0      +0       r �+0      �0       �R��0      �0       R�0      51       �R�                 p/      51       ���  �                 p/      51       ���  �                           p/      �/       T�/      �/       uȌ��/      �/       T0      �0       T�0      
1       T1      51       T                                     p/      �/       q ����
P9t "#P��/      �/       �Q����
P9t "#P��/      �/       �Q����
P9u "
h9��/      �/       q ����
P9t "#P��/      �/       �Q����
P9t "#P�0      E0       q ����
P9t "#P�E0      �0       �Q����
P9t "#P��0      �0       q ����
P9t "#P��0      �0       �Q����
P9t "#P��0      
1       �Q����
P9t "#P�1      51       �Q����
P9t "#P�                                                                     p/      �/       R�/      �/       Q�/      �/       P�/      �/       q ��/      �/       R�/      �/       Q�/      0       P0      0       Q0      0       P0      z0       Rz0      �0       r 	���0      �0       R�0      �0       P�0      �0       R�0      �0       P�0      �0       q ��0      �0       P�0      �0       pp��0      �0       P�0      �0       Q�0      �0       P�0      �0       R�0      1       P1      
1       �Q����
P9t "#p
1      1       P1      1       Q1      1       P1      (1       R(1      51       rJ�                           p/      �/       0��/      0       [0      0       0�0      !0       1�!0      �0       [�0      �0       0��0      51       [                               p/      �/      
 q  $@L$)��/      �/       �Q $@L$)��/      �/      
 q  $@L$)��/      0       �Q $@L$)�0      E0      
 q  $@L$)�E0      �0       �Q $@L$)��0      �0      
 q  $@L$)��0      51       �Q $@L$)�                      z0      �0       Q1      $1       Q$1      51       q*�                 �3      �3       T                  �3      �3       U                 �3      �3       Q                 �3      �3       R                                     4      H4       QH4      ~4       P~4      �4       �Q��4      5       Q5      5       P5      75       �Q�75      i5       Qi5      q5       Pq5      �5       Q�5      7       �Q�                                                   4      �4       R�4      �4       �R��4      5       R5      75       �R�75      l5       Rl5      q5       �R�q5      �5       R�5      �5       �R��5      �5       R�5      6       �R�6      &6       R&6      L6       �R�L6      Y6       RY6      b6       �R�b6      �6       R�6      �6       �R��6      �6       R�6      7       �R�                                           4      �4       X�4      �4       �X��4      5       X5      75       �X�75      �5       X�5      �5       �X��5      �5       X�5      6       �X�6      �6       X�6      �6       �X��6      �6       X�6      �6       �X��6      7       X                                 4      [4       Y[4      �4       �Y��4      5       Y5      75       �Y�75      i5       Yi5      q5       �Y�q5      �5       Y�5      7       �Y�                            4      �4       T�4      5       T75      �5       T�5      �5       u��~��5      �5       T6      7       T                                        4      H4       q ����
0It "#P�H4      ~4       p ����
0It "#P�~4      �4       �Q����
0It "#P��4      5       q ����
0It "#P�5      5       p ����
0It "#P�75      i5       q ����
0It "#P�i5      q5       p ����
0It "#P�q5      �5       q ����
0It "#P��5      �5       �Q����
0It "#P��5      �5       �Q����
0Iu "
HI��5      �5       �Q����
0It "#P�6      7       �Q����
0It "#P�                                                    4      34       R34      84       S�4      �4       R�4      �4       p ��4      5       R5      55       P55      75       R�5      �5       P�5      �5       R�5      �5       S�5      �5       P�5      �5       R6      6       P6      6       RG6      L6       RL6      b6       P�6      �6       s x "��6      �6       S�6      �6       s x ��6      �6       S                        4      34       0�34      84       1�84      �4       V�4      5       0�5      7       V                                    4      H4       q  $@L$)��H4      ~4       p  $@L$)��~4      �4       �Q $@L$)���4      5       q  $@L$)��5      5       p  $@L$)��5      75       �Q $@L$)��75      i5       q  $@L$)��i5      q5       p  $@L$)��q5      �5       q  $@L$)���5      7       �Q $@L$)��                                  �4      �4       q p ��4      �4       Q6      )6       Q)6      L6       PL6      �6       Q�6      �6      6 u s �Q����
0It "#ps �Q����
0It "#p0-( ��6      �6       Q�6      �6      6 u s �Q����
0It "#ps �Q����
0It "#p0-( ��6      7       P                           �4      �4       0�b6      �6       0��6      �6       Q�6      �6       X�6      �6       x ��6      �6       0��6      �6       Q�6      �6       X                         �4      �4       P�6      �6       P�6      �6       t#�#�
����6      �6       P�6      �6       t#�#�
���                     �5      �5       r q ��5      �5       r s ��5      6       P                    `7      n7       Un7      �7       �U�                          `7      k7       Tk7      �7       S�7      �7       �T��7      �7       S�7      �7       �T�                          `7      v7       Qv7      �7       V�7      �7       �Q��7      �7       V�7      �7       �Q�                    `7      v7       Rv7      �7       �R�                    w7      �7       P�7      �7       �\                  �7      �7       �U�                  �7      �7       �R�                    �7      �7       V�7      �7       �Q�                    �7      �7       S�7      �7       �T�                        �7      �7       U�7      �:       _�:      �:       �U��:      }?       _                        �7      �7       T�7      �7       P�7      �:       \�:      }?       �T�                    U8      �:       0��:      }?       0�                    �7      �7       P�7      U8       \                   �7      �7       U�7      U8       _                               �7      �7       p ����
�	u "#H��7      �7       | ����
�	u "#H��7      �:       | ����
�	 "#H��:      �:       �T����
�	 "#H��:      �:       �T����
�	�U"#H��:      �;       | ����
�	 "#H��;      ?       �T����
�	 "#H�?      }?       | ����
�	 "#H�                  �7      �7       S                    �7      �7       v  $ &Ps "��7      �7      	 p Ps "�                  �7      �7       P                  �7      U8       S                    8      /8       Q/8      48       q� 48      L8       Q                  8      U8       Y                    8      $8      	 r 3
���?8      B8       R                    (8      /8      	 u 3
���:8      =8       R                         U8      �:       \�:      �:       �T��:      �;       \�;      ?       �T�?      }?       \                   U8      �:       _�:      }?       _                       U8      �:       \�:      3;       \?      !?       \c?      }?       \                       U8      �:       _�:      3;       _?      !?       _c?      }?       _                         U8      �:       | ����
�	 "#H��:      �:       �T����
�	 "#H��:      �;       | ����
�	 "#H��;      ?       �T����
�	 "#H�?      }?       | ����
�	 "#H�                   U8      �8       | ����
�	 "#P�:      �:       | ����
�	 "#P                   U8      �8      0 | ����
�	 "#H� $ &P| ����
�	 "#P"��:      �:      0 | ����
�	 "#H� $ &P| ����
�	 "#P"�                   U8      �8       | ����
�	 "#h�:      �:       | ����
�	 "#h                          �8      �9       Q�9      �:       R�:      3;       S?      !?       Rc?      }?       R                          �8      �9       R:      �:       Q�:      &;       Q?      !?       Qc?      }?       Q                   U8      �8       �(#H�����8&��:      �:       �(#H�����8&�                          �8      �8       T�8      �:       P�:      3;       P?      !?       Pc?      }?       P                    �8      �8       x t  $ &��8      �9      	 x  $ &�                  9       9       q�0$0&� 9      ^9       q�0$r�0$+( 0$0&�                  9       9       q�0$0&� 9      ^9       q�0$r�0$-( 0$0&�                  %9      �9       T                          �9      �9       X�9      �:       X�:      3;       X?      !?       Xc?      }?       X                      $:      �:       U?      !?       Uc?      }?       U                    c:      �:       T?      !?       T                      c:      z:       [~:      �:       [?      !?       [                       �:      �:       �T�3;      �;       \�;      ?       �T�!?      c?       \                     �:      �:       _3;      ?       _!?      c?       _                      P;      W;       SW;      �;       ��!?      c?       ��                       �:      �:       0�P;      �>       0��>      �>       P!?      c?       0�                          g;      k;       Sk;      �;        �;      �;       ��!?      A?        A?      c?       ��                     g;      �;       | ����
P9r "#P��;      �;       | ����
P9�("#P�!?      A?       | ����
P9r "#P�                    k;      �;       S!?      c?       S                        x;      �;       U�;      �;       ��!?      1?       U1?      c?       ��                                �:      �:       R�;      E=       SE=      Q=       TU=      ]=       T]=      v=       R�=      �=       S�=      X>       Ri>      ?       SS?      c?       S                    �;      �;       T1?      A?       T                                 �:      �:       ^�;      �;       p q "#��@& $ &��;      �;       ~  $ &u q "#��@& $ &��;      ?       ^1?      =?       ~  $ &u q "#��@& $ &�=?      A?       ~  $ &��q "#��@& $ &�A?      E?      + ~  $ &��~  $ &��?&"#��@& $ &�E?      N?       PN?      c?       ^                  4=      v=       P                    �:      �:       V8=      i>       V                       �:      �:       P8=      E=       PE=      v=       Qv=      i>       P                       �:      �:       Xv=      �=       0��=      X>       XX>      i>       0�                       �:      �:       [v=      �=       0��=      X>       [X>      i>       0�                    �=      �=       1�%>      7>       0�                     �=      �=       p0�=      >       Q2>      X>       Q                  �=      >       T2>      X>       T                    �=      �=       YF>      X>       Y                  �=      �=       U                 �;      �;       T                 �;      �;       ^                   �;      �;       P�;      �;      
 p q "#���                  �;      �;       p ?&��;      �;       Q                      �;      <       0�<      �<       Q�<      =       Q                      �;      <       
���<      #<       U&<      =       U                  �;      <       0�                   <      3<       TB<      �<       T                    <      &<       RT<      �<       R                    <      &<       [s<      �<       [                    |<      �<       Z�<      �<       Y                     |<      �<       0��<      �<       P�<      �<       P                      �<      �<       y �<      �<       Z�<      �<       y                    �>      �>      	 p 0$0&��>      �>       q �0$0&�                      �>      �>       P�>      �>      
 p r "#����>      �>       P                   �>      �>       p ?&��>      �>       R                          �?      �?       U�?      �?       S�?      #@       �U�#@      I@       SI@      �@       �U�                          �?      @       T@      @       \@      #@       �T�#@      +@       T+@      �@       \                    �?      �?       Q�?      �?       R                        �?      �?       R�?      �?       P�?      �?       Q#@      :@       Q                           �?      �?       S�?      �?       s���?      @       S@      @       s��@      @       S;@      �@       S                                �?      �?       P�?      @       P@      @       s8@      @       PI@      `@       Qd@      z@       Qz@      �@       s8�@      �@       Q                 �?      �?       r8                   �?      �?       q8#@      :@       q8                    �?       @       ^#@      �@       ^                      �?      @       U#@      .@       U.@      :@       q0                    �?      "@       _#@      �@       _                      �?      @       R#@      :@       R:@      �@       ��                  ;@      B@       P                   x@      z@       q v �z@      �@       Q                   �@      �@       Q�@      �@      
 q t "#���                  �@      �@       q ?&��@      �@       T                          �C      D       RD      CD       \CD      iE       �R�iE      {E       \{E      �F       �R�                        D      �D       V3E      JE       ViE      �E       V�E      F       V                    D      xD      ' s 
��@$����@>$����+( �����iE      �E      ' s 
��@$����@>$����+( �����                      D      D       PD      dE       ]iE      �F       ]                   ?D      CD       | @$�����CD      uD       �R@$�����                      hD      uD       U�D      �D       U�E      F       U                        �D      �D       T3E      ?E       TF      F       T-F      6F       T                          1E      3E       UJE      QE       U�E      �E       U(F      -F       P�F      �F       U                      �D      �D       r t #��D      �D       R�E      �E       R                          .D      �D       P3E      FE       PiE      �E       P�E      F       P-F      SF       P                              2D      �D       X3E      <E       X<E      FE       v(iE      �E       X�E      F       X-F      SF       XSF      �F       ��                       2D      �D       v,3E      FE       v,iE      �E       v,�E      F       v,                       2D      �D       v03E      FE       v0iE      �E       v0�E      F       v0                       2D      �D       v43E      FE       v4iE      �E       v4�E      F       v4                       2D      �D       v83E      FE       v8iE      �E       v8�E      F       v8                          6D      �D       _3E      JE       _iE      �E       _�E      F       _-F      yF       _                       6D      �D       v� 3E      FE       v� iE      �E       v� �E      F       v�                  ?D      eD       ]                     ?D      CD       | @$�CD      RD       \RD      eD       �R@$�                      RD      YD       \YD      aD      
 r | "#���aD      eD       R                     RD      YD       | ?&�YD      aD       RaD      eD       | ?&�                  �D      3E       _                  �D      E       | p �                    �E      �E       Q�E      �E       ��                  �E      �E       | p �                �E      �E       S                �E      �E       U                   �E      �E       R�E      �E      
 r t "#���                  �E      �E       r ?&��E      �E       T                    OF      SF       QSF      �F       ��                  TF      |F       | p �                            �X      �X       U�X      MY       VMY      TY       �U�TY      �Y       V�Y      �Y       �U��Y      �[       V                  �X      �X       T                                �X      �X       Q�X      @Y       \@Y      TY       �Q�TY      �Y       \�Y      �Y       �Q��Y      1Z       \1Z      Q[       �Q�Q[      �[       \                    �X      �X       R�X      �[       �R�                            �X      �X       U�X      MY       VMY      TY       �U�TY      �Y       V�Y      �Y       �U��Y      �[       V                    �X      �X       q�Y      Y       Q                   �X      Y       PY      Y       P                   �Y      �Y       \�Y      �Y       �Q�                            TY      �Y       Q�Y      �Y       Q�Y      1Z       QQ[      �[       Q�[      �[       Q�[      �[       Q                        TY      �Y       \�Y      1Z       \1Z      Q[       �Q�Q[      �[       \                                            TY      �Y       P�Y      �Y       �T��Y      �Y       P�Y      �Y       �T��Y      1Z       P1Z      Q[       �T�Q[      }[       P}[      �[       �T��[      �[       P�[      �[       �T��[      �[       P�[      �[       �T��[      �[       P�[      �[       �T�                    TY      �Y       V�Y      �[       V                    �Y      �Y       P�Y      �Y       S                   �Z      �Z       ~d��Z      [       \                  �Z      Q[       Q                   �Z      [       |[      Q[       Z                  �Z      Q[       P                   �Z      [       |[      Q[       Y                   �Z      [       |[      Q[       R                   �Z      [       |[      Q[       X                   �Z      [       |[      Q[       T                 �Z      [       |                  1Z      �Z       \                 �Y      �Y       \                 �Y      �Y       \                 x[      �[       \                   �[      �[       \�[      �[       \                    �[      �[       P�[      �[       P                 �[      �[       \                  �[      �[       P                            �[      �]       U�]      �^       S�^      �^       U�^      6_       �U�6_      N_       SN_      �_       U                          �[      �]       T�]      '_       ��'_      6_       �T�6_      N_       ��N_      �_       T                            �[      \       Q\      �]       S�]      '_       ��'_      6_       �Q�6_      N_       ��N_      �_       S                        �[      K\       RK\      �]       ���]      N_       �R�N_      �_       ��                         +\      �]       t� ��]      '_       ��#H�'_      6_       �T#H�6_      N_       ��#H�N_      �_       t� �                     8\      o\       Qo\      �]       t0N_      �_       t0                    
\      /_       \6_      �_       \                  \      �\       P                 K\      o\       1�                     8\      Y\       YY\      �]       t,N_      �_       t,                      8\      �]       ^�]      N_       ��N_      �_       ^                          K\      v\       Ry\      �]       R�]      '_       ��6_      N_       ��N_      �_       R                            K\      o\       Ro\      {\       V~\      �]       V�]      '_       ��6_      N_       ��N_      �_       V                      �]      0^       _�^      �^       _6_      N_       _                    '^      '^       ^'^      �^       ~ :�I_      N_       ^                            /\      3\       Q3\      p^       w p^      {^       ��{^      +_       w +_      6_       ��6_      �_       w                     t\      �\       Q�\      �\       x��0$0&�                 �\      �\       \                 �\      �\       R                          �\      �\       Q�\      �\      
 q y "#����\      �\       [�\      �\       q ?&q "#����\      �\      # |  $ &��|  $ &��?&"#���                       �\      �\       q ?&��\      �\       Y�\      �\       q ?&��\      �\       |  $ &��?&�                �\      �\       \                �\      �\       V                 Y]      Y]       @�Y]      Y]       8�|_      �_       @��_      �_       8�                  C^      �^       T                         Y^      a^       q p r "#��@&�a^      d^       q t  $ &��r "#��@&�d^      k^      ( q t  $ &��t  $ &��?&"#��@&�k^      x^       Qx^      �^      ( v t  $ &��t  $ &��?&"#��@&�                     �]      �]       s �]      	^       s  s� "�	^      �^       V�^      �^       s �^      �^       s  s� "��^      �^       T6_      N_       V                         �]      	^       s	^      �^       ]�^      �^       s�^      �^       ]6_      N_       ]                C^      Y^       T                C^      Y^       ��                   R^      Y^       PY^      Y^      
 p r "#���                  R^      Y^       p ?&�Y^      Y^       R                  �^      '_       R                  �^      '_       T                    �^      �^       r | ��^      �^       P�^      �^       U                �^      �^       ��                   �^      �^       P�^      �^      
 p q "#���                  �^      �^       p ?&��^      �^       Q                �^      _       U                �^      _       ��                  �^      _       P_      _      
 p q "#���                  �^      _       p ?&�_      _       Q                    �_      �_       U�_      ch       �U�                            �_      �_       T�_      `       _`      $a       �T�$a      :a       _:a      Pa       �T�Pa      �a       _�a      ch       �T�                    �_      �_       Q�_      ch       ��}                    �_      �_       R�_      �_       ��}                          �_      �_       P�_      �_       ��}$a      2a       ��}2a      6a       Pa      �a       P                      �_      $a       �U�Pa      a       �U��a      ch       �U�                      �_      $a       ��}Pa      a       ��}�a      ch       ��}                      �_      $a       ��}Pa      a       ��}�a      ch       ��}                          �_      `       _`      $a       �T�Pa      a       _�a      �a       _�a      ch       �T�                        �_      �_       0�Pa      ]a       0�]a      ra       P�a      �a       0�                                  	`      `       Z`      `       \*`      /`       \/`      {`       0��c      ?d       \�d      �d       |��d      e       2�[e      �e       0��f      �f       0�                          D`      �`       \�`      $a       ��~�a      �a       ��~d      ?d       \�f      �f       \�g      �g       ��~                                           D`      �`       [�`      $a       ^�a      �a       ^�a      �b       _�b      kc       [kc      �c       _d      ?d       [�e      �e       _�e      �e       [f      tf       _tf      �f       [�f      hg       [mg      �g       _�g      �g       ^�g      �g       _�g      ch       [                    D`      {`       | ����
�	{ "#H�d      ?d       | ����
�	{ "#H��f      �f       | ����
�	{ "#H�                               U`      �`       S�`      $a       ��~�a      �c       ��~d      ?d       S�e      �e       ��~f      �f       ��~�f      �f       S�f      hg       ��~mg      ch       ��~                                       m`      $a       V�a      �a       V�a      �b       \�b      �c       V�c      �c       \�c      �c       V1d      ?d       V�e      �e       Vf      tf       \tf      �f       V�f      hg       Vmg      ch       V                 �f      �f       p X�                                        m`      $a       S�a      �a       S�a      �b       S�b      �b       ��~�b      c       S c      kc       Pkc      �c       S1d      ?d       S�e      �e       Sf      �f       S�f      �f       S%g      5g       ��~5g      ;g       Smg      �g       S                                 m`      �`       0��`      $a       _�a      �a       _�a      �b       ��~�b      �b       S�b      c       ��~�c      �c       ��~1d      ?d       0�f      �f       ��~�f      �f       0��g      �g       _                               m`      $a       0��a      �a       0��a      c       ��~�c      �c       ��~1d      ?d       0�f      �f       ��~�f      �f       0��g      �g       0�h      ch       Q                                   m`      $a       0��a      �a       0��a      c       ��~ c      Ac       YAc      Lc       y�Lc      kc       Y�c      �c       ��~1d      ?d       0�f      �f       ��~�f      �f       0�%g      5g       Y�g      �g       0�                                m`      $a       0��a      �a       0��a      �b       V�b      �b       1��b      �b       V�c      �c       V1d      ?d       0�f      Of       Vof      tf       1��f      �f       0��g      �g       0�                                           m`      $a       0��a      �a       0��a      b       Zb      b       ��~b      �b       Z�b      �b       ��~�b      c       Z�c      �c       Z1d      ?d       0�f      /f       Z/f      5f       ��~5f      _f       Z_f      of       ��~of      tf       Ptf      �f       Z�f      �f       0��g      �g       0�                     �`      �`       R�`      �`       R�`      �`       P                       �`      �`       S�`      �`       0��`      a       Q�g      �g       S                          �`      �`       Q�`      �`       Q�`      �`       S�`      $a       \�g      �g       Q�g      �g       s0                 �`      a       Q                 �`      $a       \                �`      "a       ��~                �`      "a       ^                   �`      a       |q�a      a       R                 a      "a       P                        �a      b       ]0b      �b       ]�c      �c       ]f      tf       ]                 �a      b       ]                 �a      b       S                �a      b       ��~                �a      b       _                   �a      �a       s}��a      b       R                  b      b       P                 5f      tf       ]                 5f      tf       S                5f      of       ��~                5f      of       _                   5f      [f       s}�[f      _f       R                  `f      df       P                    �f       g       R5g      Ng       ��~�g      h       R                        �f       g       UBg      Ng       U�g      %h       UAh      ch       U                      �f      5g       XLg      Ng       X�g      ch       X                        	g      g       Qg       g       p r��g      �g       p r��g      h       ur�                   	g      5g       Z�g      ch       Z                       	g      g       q z �g       g       Q�g      �g       Q�g      h       } uz ruz r0-( �                2c      Lc       [                2c      Lc       T                2c      Lc       P                          �c      �c       S�c      �c       P�c      �c       Pmg      g       P�g      �g       P                        �c      �c       R�c      �c       Rmg      �g       R�g      �g       R                 �c      �c       _                 �c      �c       P                 �c      �c       S                 �c      �c       _                 �c      �c       R                 �c      �c       S                       ?d      �d       \e      [e       \�e      f       \�f      �f       \hg      mg       \                       ?d      �d       [e      [e       [�e      f       [�f      �f       [hg      mg       [                    ?d      Ld       | ����
�	{ "#H��e      f       | ����
�	{ "#H��f      �f       | ����
�	{ "#H�hg      mg       | ����
�	{ "#H�                      ?d      Qd       S�e      f       S�f      �f       | ����
�	{ "#`hg      mg       | ����
�	{ "#`                        ?d      �d       Ve      [e       V�e      f       V�f      �f      0 | ����
�	{ "#X� $ &X| ����
�	{ "#`"�hg      mg      0 | ����
�	{ "#X� $ &X| ����
�	{ "#`"�                   Ld      �d       Se      [e       S                 Ld      Ld       u  $0.�                    \d      �d       Pe      [e       P                  ld      �d       R                  td      �d       Q                    e      e       Q"e      [e       Q                 �e      �e       0�                 �e      �e       [                  �e      �e       X                  �e      �e       ��~                   �e      �e       Q�e      �e       {0                  �e      �e       T                     �e      �e       Q�e      �e       q���e      �e       Q                  �e      �e       q�0$0&��e      �e       qH�0$0&�                   �e      �e       P�e      �e      
 p r "#���                  �e      �e       p ?&��e      �e       R                      �h      �h       U�h      �h       S�h      �v       �U�                                              �h      �h       T�h      ki       _ki      �j       ]�j      ck       _ck      dk       �T�dk      �n       _�n      p       ]p      3p       _3p      �p       ]�p      �s       _�s      t       ]t       u       _ u      )u       ])u      �v       _�v      �v       ]                                  �h      �h       Q�h      �h       ��~�h      dk       �Q�dk      �m       ��~�m      �n       �Q��n      �n       ��~�n      �u       �Q��u      �u       ��~�u      �v       �Q�                                  �h      �h       R�h      �h       ��}�h      dk       �R�dk      �m       ��}�m      �n       �R��n      �n       ��}�n      �u       �R��u      �u       ��}�u      �v       �R�                            �h      �h       P�h      �h       ��}dk      �k       ��}�k      �m       ��}�n      �n       ��}�u      �u       ��}                        �h      �h       ��}dk      �m       ��}�n      �n       ��}�u      �u       ��}                        �h      �h       ��~dk      �m       ��~�n      �n       ��~�u      �u       ��~                                          �h      ki       _ki      �j       ]�j      Nk       _dk      �n       _�n      p       ]p      3p       _3p      �p       ]�p      �s       _�s      t       ]t       u       _ u      )u       ])u      �v       _�v      �v       ]                            �h      �h       S�h      Nk       �U�dk      Fl       SFl      �n       �U��n      �n       S�n      �v       �U�                       �h      �h       0��k      �k       0��k      �k       P�n      �n       P�n      �n       0�                                        �h      �h       ^�h      �h       ~��h      �h       ^�h      Ni       0�*k      4k       ~�4k      Nk       2��m      �n       ^p      3p       ^�p      �p       0�+t      8t       ^)u      Gu       ^�u      av       0�                      dk      �k       ��}#P��k      �m      	 ��}#����n      �n       ��}#P��u      �u      	 ��}#���                   �k      �m       ��}�u      �u       ��}                   �k      �m       _�u      �u       _                   �k      �m       ���u      �u       ��                    �k      �m       U�u      �u       U                      l      "l       P"l      �m       ��}�u      �u       ��}                   l      �m      	 ��}#����u      �u      	 ��}#���                   l      *l       V*l      ql       ��}#��                 ql      �l       0�                     ql      �l       0��l      �m       \�u      �u       \                       ql      �l       0��l      m       ]m      m       ]m      �m       Y�u      �u       ]                      �l      m       [m      {m       [{m      �m       P�u      �u       [                       �l      �l       R�l      �l       r���l      �m       R�u      �u       r��                  �l      �m       Z                  �l      �m       Y                 �l      �m       u�8$8& $�� $)�                                    �l      �l       t x ��l      �l       Q�l      �l       ~ t x t x 0-( ��l      m       x t t x t x 0-( �m      Im       QIm      Rm       t p �Rm      Ym       T]m      `m      $ q u �0$0&p u �0$0&p 0-( �`m      rm      & q u �0$0&ru �0$0&r0-( �rm      �m       P                   6m      Rm       t x -�Rm      �m       u �0$0&x -�                    Vm      ]m       T]m      `m      $ q u �0$0&p u �0$0&p 0-( �`m      dm      & q u �0$0&ru �0$0&r0-( �                   ]m      dm       Tdm      dm      
 p t "#���                  ]m      dm       t ?&�dm      dm       P                    �l      �l       Q�l      �l       ~ t x t x 0-( ��l      �l       x t t x t x 0-( �                   �l      �l       Q�l      �l      
 q ~ "#���                  �l      �l       q ?&��l      �l       ^                            )i      Ni       0��m      �n       1�p      3p       1��p      �p       0�+t      8t       1�)u      Gu       1�                                                )i      ki       _ki      �j       ]�j      �j       _�m      �n       _�n      p       ]p      3p       _3p      �p       ]�p      �q       _r      �s       _�s      t       ]t      8t       _Xt       u       _ u      )u       ])u      �u       _av      �v       _�v      �v       ]                          )i      Ni       � ��m      �n       ��p      3p       ���p      �p       � �+t      8t       ��)u      Gu       ��                      5i      Ni       U�m      n       T�p      �p       U                                        @i      hi       ]hi      �j       ��~�m      �n       ]�n      p       ��~p      3p       ]3p      �p       ��~�p      �p       ]�s      t       ��~+t      8t       ]u      )u       ��~)u      Gu       ]�v      �v       ��~                             �j      �j       ��~X��p      �p       ��~X�8t      Xt       ��~X�Xt      tt       p X�tt       u       ��~X��u      �u       p X�av      �v       ��~X�                
                                      @i      Ni       Uki      �j       S�m      n       Tn      �n       S�n      �p       S�p      �p       U�p      �p       ��~�p      Eq       QEq      �q       s��r      )r       q� �1r      �r       Q�r      +s       s��+s      �s       Q�s      t       St      +t       s��+t      8t       Su       u       ��~ u      Gu       SGu      �u       s���v      �v       S                                                         @i      Ni       0�ki      ~j       _~j      �j       [�m      n       0�n      �n       \�n      �o       _�o      p       Sp      3p       \3p      �p       _�p      �p       0��p      �q       [r      Hr       [Xr      ]r       Q]r      �s       [�s      t       _t      +t       [+t      8t       \u       u       [ u      )u       _)u      Gu       \Gu      wu       [wu      �u       ��~�v      �v       _                                        @i      ki       0�ki      �j       ��~�m      �n       0��n      �o       ��~�o      p       ��~p      3p       0�3p      �p       ��~�p      �p       0��s      t       ��~+t      8t       0�u      )u       ��~)u      Gu       0��v      �v       ��~                 �m      n       �(                 �m      n       �(#�����3$ -G     "                      @i      Ni       0��m      �m       0��m      n       P�p      �p       0�                            �i      Wj       V�n      p       V3p      �p       V�s      t       V u      )u       V�v      �v       V                   �i       j       ~ "�o      'o       ~ "�                     �i       j       vs�o      �o       vs�Cp      �p       vs�                   �i       j       ��~1&~ ""�o      'o       z 1&~ ""�                          So      {o       R{o      �o       q 	���o      �o       z 1&~ "# 	���o      �o       T\p      �p       X                    yp      �p       Y�p      �p       z ~ "# 	�p �                            eo      no       q u �no      to       q t �to      �o       U`p      cp       t u �cp      fp       t { �fp      �p       T                            {o      �o       q r ��o      �o       Q�o      �o       x z 1&r ~ "z 1&r ~ "0-( �|p      p       r { �p      �p       r q ��p      �p       R                    _o      ho       Tho      �o        &p A-( �                    _o      ~o       X~o      �o        Jp A-( �                     �o      �o       vs��s      t       vs��v      �v       vs�                  �s      �s       ^                      �s      �s       R�s      �s       ~ 	���s      t       Q                      �s      �s       ~ t ��s      �s       ~ q ��s      t       T                    �s      �s       ~ r ��s      t       ^                     �o      �o       &��s      �s       Q�v      �v       &�                     �o      �o       J��s      �s       U�v      �v       J�                         7n      Gn       Q�n      �n       0��n      �n       P p      $p       Q$p      .p       s(>u      Gu       s(                                 n      @n       0�@n      Qn       SQn      `n       Q�n      �n       0��n      �n       V�n      �n       Sp       p       0� p      3p       S)u      Gu       0�                          n      en       V�n      �n       V�n      �n       Sp      3p       V)u      Gu       V                       n      @n       p 8�p       p       p 8�)u      3u       p 8�3u      >u       s�8�                        n      (n       r 8�(n      3n       v�8�p       p       r 8�)u      Gu       r 8�                   xt      �t       U�u      �u       ��~                      t      u       X�u      �u       Xav      �v       X                      �t      u       T�u      �u       Tav      �v       T                      �t      �t       P�t      �t       r u��t      �t       xu�                     �t      �t       S�t      �t       tx�av      �v       S                       �t      �t       p s ��t      �t       P�t      �t       y r s ur s u0-( ��t      �t       y xs uxs u0-( �                    �t      u       Rav      �v       R                     q      q       
��q       q       p u � q      9q       P                 .q      9q       _                 .q      9q       R                 .q      9q       Q                      ]r      �r       P7s      �s       PGu      Tu       P                   _s      rs       q� �rs      �s       R                    �j      k       ��}�q      �q       ��}8t      Xt       0��v      �v       ��}                    �j      k       _�q      r       _8t      Xt       _�v      �v       _                   �j      �j       ��}�����
�	 "#H��q      �q       ��}�����
�	 "#H�8t      Xt       � ��v      �v       ��}�����
�	 "#H�                        �j      �j       P�q      �q       PHt      Xt       P�v      �v       P                        �j      k       R�q      r       RSt      Xt       R�v      �v       R                   �j      k       P�q      r       P                      �j      �j       U�j      k       pk      k       p@                 �j      	k       Q                    �j      �j       Q�j      	k       p�                   �j      	k       T                      �q      �q       U�q      r       pr      r       p@                 �q      	r       Q                    �q      �q       Q�q      	r       p�                   �q      	r       T                   uk      �k       0��n      �n       0�                   uk      �k       ��}#h��n      �n       ��}#h�                   uk      �k       V�n      �n       V                     uk      yk       Uyk      �k       _�n      �n       _                    zk      �k       P�n      �n       P�n      �n       P                 �n      �n       0�                 �n      �n       ��}#h�                 �n      �n       V                 �n      �n       _                 �n      �n       P                 �k      �k       1�                 �k      �k      	 ��}#���                 �k      �k       V                   �k      �k       U�k      �k       _                  �k      �k       P�k      �k       P                 �k      �k       1�                 �k      �k      	 ��}#���                 �k      �k       V                 �k      �k       _                 �k      �k       P                 v      av       0�                 v      av       _                  v      av       X                  v      -v       ��~                   v      -v       Q-v      av       0                  $v      av       T                     $v      9v       Q9v      Wv       q��Wv      av       Q                  -v      9v       q�0$0&�9v      Dv       qH�0$0&�                   =v      Dv       PDv      Dv      
 p r "#���                  =v      Dv       p ?&�Dv      Dv       R                  �v      �v       R�v      �v       �R�                          p�      ��       U��      2�       V2�      9�       �U�9�      D�       VD�      K�       �U�                 p�      K�       ���  �                         p�      ��       0���      �       ]�      "�       1�"�      6�       ]9�      H�       ]                       p�      )�       1�)�      9�       P9�      9�       1�9�      ;�       0�;�      K�       P                          ��      ��       0���      �       ^�      $�       P$�      8�       ^9�      J�       ^                     ��      Ҁ       ���Ҁ      ـ       Qـ      K�       ���                       ��      �       S�      �       P�      1�       S9�      C�       S                   �      $�       \9�      F�       \                �      �       0�                    �      �       ����      �       R�      �       ���                �      �       ���                �      �       V                 �      �       v�                  �      �       \                    `�      �       U�      ��       �U�                    `�      |�       T|�      ��       �T�                    `�      z�       Qz�      ��       �Q�                    `�      ��       R��      ��       �R�                      `�      ��       X��      ��       S��      ��       �X�                 `�      a�       u�                     l�      ��       V��      ��       P                      �      �       U�      b       w b      m       ��}                    �      �       T�      m       ��}                     �      �       Q�      �       ]�      [       ^                      �      �       R�      [       V[      m       �R�                     �      �       0��      �       _�      �       _                   �      �       Q�      [       ]                       �      �       0��      �       |��      �       \�             |�                     0      D       ��}�D      N       RN      O       ��}�                 0      O       ^                 0      O       ��}                 0      O       w                  �      �       2�                 �      �       U                 �      �       u�                 �      �       u� �                      0      D       UD      �       V�      �       �U�                      0      H       TH      �       \�      �       �T�                      0      H       QH      �       S�      �       �Q�                 c      }       W                 c      }       1�                 c      }       \                 c      }       V                 p      �       1�                 p      �       U                 ~      �       u�                 �      �       u� �                                        }       U}      �       ]�      �       �U��      �       U�             ]             �U�      O       UO      �       ]�      �       U                                    7       T7      �       V�             V      +       T+      �       V�      �       T�      �       V                                    7       Q7      �       \�             \      +       Q+      �       \�      �       Q�      �       \                                          G       RG      }       [}      �       �R��      �       [�             �R�      +       R+      a       [a      �       ���      �       R�      �       [                                        K       XK      �       ^�      �       �X��             ^             �X�      +       X+      �       ^�      �       X�      �       ^                           �       0��      �       P�      �       0��             P      �       0�                                     7       0�7      }       Z�      �       Z             0�      +       1�+      a       Za      �       ���      �       1��      �       3��      �       Z                   �      �       U�             U                       K      Z       0�Z      }       S�      �       S�      �       0�                                G      }       R�      �       R�      �       �+      =       R=      O       u O      a       } a      �       ��      �       R                           K      Z       XZ      }       Q�      �       Q�      �       P�      �       } �����32$x "<��      �       X                u      �       ��
  �      �       ��
                    u      �       [�      �       [�      �       ��                  u      }       u��      �       }�                  u      �       0��      �       0��      �       P                    y      �       P�      �       P                  �      �       ���
  +      �       ���
                        �      �       [�      �       �R�+      a       [a      �       ��                      �      �       U�      �       ]+      O       UO      �       ]                  �      �       0�+      �       0�                    �      �       R�      �       _+      �       _                    �      �       0��      �       P+      �       0�                   +      O       UO      �       ]                   +      a       [a      �       ��                 +      �       _                 +      a       P                   +      T       _T      a       Ra      �       ��                                    @;      �;       U�;      �;       V�;      �;       p��;      �;       �U��;      �;       V�;      A<       p�A<      B<       �U�B<      ]<       V]<      s<       p�s<      t<       �U�                              @;      ;       T;      �;       ]�;      �;       �T��;      �;       ]�;      B<       �T�B<      o<       ]o<      t<       �T�                              @;      g;       Qg;      �;       \�;      �;       �Q��;      ;<       \;<      B<       �Q�B<      m<       \m<      t<       �Q�                              @;      �;       R�;      �;       S�;      �;       �R��;      �;       S�;      B<       �R�B<      j<       Sj<      t<       �R�                    @;      �;       X�;      t<       �X�                              @;      �;       Y�;      �;       ^�;      �;       �Y��;      ?<       ^?<      B<       �Y�B<      q<       ^q<      t<       �Y�                    �;      �;       P�;      �;       P                    G;      �;       Y�;      �;       ^                   @;      �;       X�;      �;       �X�                   @;      �;       U�;      �;       V                                   _;      �;       U�;      �;       V�;      �;       p��;      �;       �U��;      �;       V�;      A<       p�A<      B<       �U�B<      ]<       V]<      s<       p�s<      t<       �U�                                   _;      �;       U�;      �;       V�;      �;       p��;      �;       �U��;      �;       V�;      A<       p�A<      B<       �U�B<      ]<       V]<      s<       p�s<      t<       �U�                  _;      s;       X                   _;      k;       Pk;      s;       u                   c;      k;       p ����Hu"H�k;      s;       u�����Hu"H�                       �;      ?<       ^?<      B<       �Y�B<      q<       ^q<      t<       �Y�                         �;      .<       S.<      1<       s�1<      8<       SB<      j<       Sj<      t<       �R�                       �;      ;<       \;<      B<       �Q�B<      m<       \m<      t<       �Q�                       �;      �;       ]�;      B<       �T�B<      o<       ]o<      t<       �T�                       �;      A<       _A<      B<       �U#�B<      s<       _s<      t<       �U#�                   �;      �;       0��;      B<       P]<      t<       P                     �;      9<       V]<      k<       Vk<      t<       ��                 �;      �;       ���
  B<      ]<       ���
                   �;      �;       ^B<      ]<       ^                 �;      �;       _B<      ]<       _                   �;      �;       0�B<      X<       0�X<      ]<       P                       �;      �;       P�;      �;       v�;      �;        B<      W<       P                  �;      =<       ]                    �;      <       U<      !<       ��!<      B<       U                 �;      B<       T                       �;      �;       ���;      !<       R!<      #<       r 1&�#<      )<       R)<      .<       ��.<      B<       R                          �;      <       r  q �<      	<       q x �	<      <       r  q �<      <       r  t ���<      B<       Q                          �      
       U
      �       ^�      �       �U��      N       ^N      Q       U                      �      
       T
      N       ��N      Q       T                                �      �       Z�      �       ]�      �       Z�      �       Z�      �       }��      �       ]�      �       Z�      N       }�N      Q       Z                              .       ].      �       U�              U�      �       U                     .      �       ^�      �       �U��      N       ^                  .      u       U�      �       U                  .      u       Z�      �       Z                  .      u       { | "#��      �       { | "#�                  .      u       Q�      �       Q                     .      T       { | "# T      q       T�      �       { | "#                    =      u       P�      �       P                  =      u       { | "#�      �       { | "#                  =      u       q �      �       q                       =      d       Rd      l       r�l      u       R�      �       R                   �      �       ^�      N       ^                  �      �       ���      N       ��                     �      �       Z�      P       _�      N       _                   �      �       U�      �       P                    �      �       0��      �       0��             P                 �      �       p ����H{ "�                      �              X�      �       X�      N       ��                 �      �       p ����H{ "                      �              Y�      �       Y�      N       ��                    P      i       Ui      �       _                                      y 3%�             Y      #       p  y "�#      *       y p �*      3       p  y "�      N       Z                                   T      #       t p "#�#      *       t p "�*      3       t p "#�                          #       q p "#�#      *       q p "�*      3       q p "#�                       @       Z                  3      @       q p "�                      u      z       �Y��z      ~      
 �Y�R��~      �       ��������                        �             U      5       S5      ;       �U�;      |       S                          �             T      ;       �T�;      Q       TQ      d       Ud      |       �T�                        �             Q      :       ]:      ;       �Q�;      |       ]                                   R      6       V;      |       V                     �      ,       0�,      ;       P;      |       0�                     �             0�      ;       Q;      |       0�                 G      |       S                  G      d       Ud      z       �T�                G      z       V                 G      d       Q                G      ]       V]      z       \                      P      w       Uw      �       ]�      �       �U�                      P      w       Tw      �       V�      �       �T�                    c      n       Pn      w       u                      g      �       S�      �       sh��      �       S                 w      �       V                   w      �       S�      �       sh�                          �      �       U�      �       V�      �       �U��      �       U�             V                        �      �       T�      �       S�      �       �T��             S                          �      �       Q�      �       �Q��      �       Q�      �       R�             �Q�                    �      �       0��      �       0��             P                  �      �       P                    �             U      �       Q                  �      �       X                        �       T                       ,       X                       ,       T                 ,      M       q��                 M      �       q��                 �      �       q��                      �:      �:       U�:      /;       S/;      1;       �U�                 �:      *;       V                 �:      �:       V                 �:      �:       V                 �:      ;       V                 �:      ;       s� �                 �:      ;       V                 �:      ;       s� �                    p      �       U�      7       [                      p      �       T�      �       u��      7       �T�                          p      �       Q�      �       S�      �       �Q��      �       S�      7       �Q�                    p      �       R�      7       �R�                          p      �       X�      �       V�      �       �X��      �       V�      7       �X�                   u      �       u��      �       {��      7       {��                      �      �       V�      �       V�      7       �X�                      �      �       S�      �       S�      7       �Q�                        �      �       U�      �       {���      �       U�      7       {��                   �      �       Q�      �       u                            z      �       0�g      �       R�      �       R�      �       0��      �       P�             0�                       �      �       0��      �       {���      �       0��      7       {��                              n       Qn      q       q�q      �       Q�      �       {��      7       {�                  !      2       SP      ]       S                  !      2       QP      ]       Q                       +      2       P2      2      
 p r "#���V      Y       PY      ]       R                      +      2       p ?&�2      2       RV      Y       p ?&�Y      ]       r ?&�]      ]       R                        �      �       P�      [       pP�[      �       P�      �       P                �      �       S                  �      �       p�      �       pX                   �      �       Q�      �      
 q | "#���                  �      �       q ?&��      �       \                �      �       S                   �      �       Q�      �      
 q | "#���                  �      �       q ?&��      �       \                      %       S                        %       \%      %      
 | } "#���                        %       | ?&�%      %       ]                %      ,       S                  %      ,       Q,      ,      
 q ~ "#���                  %      ,       q ?&�,      ,       ^                            �       R�             R      ,       rP�,      7       R                   @      �       u��      �       ^                               P�             P                 @      �       u                   �             {���             {��                    	      �       U�      7       U                          P      P       PP      Z       p �Z      �       y u� $ &��      �       P�      �       p ��      �       y ~ � $ &��      �       y u� $ &�                P      j       �Q��      �       �Q�                    P      Z       p �Z      j      	 y u���      �       p ��      �      	 y ~ ��                      c      j       Pj      j      
 p ~ "#����      �       P�      �      
 p  "#���                    c      j       p ?&�j      j       ^�      �       p ?&��      �       _                        0      U       UU      /       ]/      L       | L      �       �U�                      0      D       TD      �       V�      �       �T�                      0      Q       QQ      �       S�      �       �Q�                       0      Y       0�Y      ]       P]      �       \�      �       �Q                  �      �       U�      �       U                        �      �       P�      �       p~��      �       P�      �       P�      �       p~��      7       P                 p      �       |��                   p      �       |���      �       Q�      �       qh��      �       Q                 �      �       |�                   �      �       |��      �       Q�      �       qh��      "       Q                  K      T       P                    s      �       1��      �       T�      �       T             T=      J       T                    x      �       1��      �       T                   x      �       ���      �       Z                 x      �       X                   x      �       0��      �       Q                     �      �       r �q ����1$��"���      �       r �u 1$��"���      �       r|�u 1$��"��                 �      �       T                 �      �       _                 �      �       X                   �      �       0��      �       Q                     �      �       r �q ����1$ "���      �       r �u 1$ "���      �       r|�u 1$ "��                 �             T                 �             ^                 �             X                   �      �       0��             Q                     �      �       r �q ����1$~ "���             r �u 1$~ "��             r|�u 1$~ "��                       =       T                       =       ]                       =       X                                0�      =       Q                           "       r �q ����1$} "��"      8       r �u 1$} "��8      =       r|�u 1$} "��                        P      �       U�             �U�             U      %       �U�                                      P      �       T�      �       �T��      �       X�              X              x�      4       Y8      R       YR      W       y�W      b       Zb      }       T}      �       Z�      �       z��             T      #       z�                        P      �       Q�             �Q�             Q      %       �Q�                          P      �       R�             ]             �R�             R      %       ]                          P      �       X�             ^             �X�             X      %       ^                        P      �       Y�      �       S�             �Y�      %       S                      P             �              P      %       �                     t      {       u��             U                               u��                  �      b       Z                    �             T      %       T                        �      �       pP��      �       P�              pP�              p0�                    �      �       [�      �       [                              4       pP�8      B       PB      R       pP�R      W       p0�                        4       [                       W      ]       1�]      b       {�b      r       {~�x      }       {��      �       {~�                    �      �       Q      %       Q                        �      �       Y�      �       Y�      �       r<�      �       r                     �      �       X�      �       y q ��      �       X                         ]      b       Rx      �       R�      �       rP��      �       R�      �       rP��      �       R      %       R                    �              U      b       �U�                    �       �        T�       b       �T�                     �       �        t ����
�u "#��              �T����
�u "#�      b       �T����
��U"#�                     �       �        t ����
�u "#��              �T����
�u "#�      b       �T����
��U"#�                  �       �        P�       �        p�                       �       �        �T����
�u "#��       L       QL      \       qh�\      a       Q                   �              �T����
�u "#�      b       �T����
��U"#�                 �       �        �T����
�u "#�                                   qp3      T       PT      a       qp                                  T3      <       p r �<      a       T                      %       q                          %       P%      %      
 p t "#���                        %       p ?&�%      %       T                �       �        x                    �       �        Q�       �       
 q r "#���                  �       �        q ?&��       �        R                                �      �       U�      0       S0      :       �U�:       !       S !      !       U!      8!       S8!      B!       �U�B!      :#       S                                �      �       T�      3       \3      :       �T�:       !       \ !      !       T!      ;!       \;!      B!       �T�B!      :#       \                                                �      �       Q�      :       ��:      �        Q�        !       �� !      B!       QB!      �!       ���!      �!       Q�!      �!       ���!      �!       Q�!      �!       ���!      �!       Q�!      "       ��"      �"       Q�"      �"       ���"      �"       Q�"      :#       ��                                      �      �       R�      �       [�      /       w /      :       ��:      �       [�       !       w  !      !       R!      B!       [B!      �!       w �!      �!       [�!      :#       w                                                        �      �       q  $ &
�t "#��      �       q  $ &
�| "#��      3       ��� $ &
�| "#�3      :       ��� $ &
��T"#�:      �        q  $ &
�| "#��        !       ��� $ &
�| "#� !      !       q  $ &
�t "#�!      ;!       q  $ &
�| "#�;!      B!       q  $ &
��T"#�B!      �!       ��� $ &
�| "#��!      �!       q  $ &
�| "#��!      �!       ��� $ &
�| "#��!      �!       q  $ &
�| "#��!      �!       ��� $ &
�| "#��!      �!       q  $ &
�| "#��!      "       ��� $ &
�| "#�"      �"       q  $ &
�| "#��"      �"       ��� $ &
�| "#��"      �"       q  $ &
�| "#��"      :#       ��� $ &
�| "#�                   �      �       q  $ &
�t "#� !      !       q  $ &
�t "#�                   �      �       q  $ &
�t "#� !      !       q  $ &
�t "#�                                                  -      1       R1      �       ���             R             s      !       R:       !       ��!      B!       ��B!      w!       Rw!      !       s!      �!       R�!      �!       ���!      "       R"      �"       ���"      �"       Q�"      #       ��#      #       ��$#      :#       ��                                             O      /       Vl      �       V�      �       Q�      �       s�      
       T
             s:       !       V!      9!       V9!      B!       �U#B!      w!       @��!      �!       V�!      �!       @�
"      "       @�"      �"       V�"      �"       @��"      $#       V                                v      �       1�k      w       1�w       !       ��!      !       0��!      �!       0��!      �!       ��"      �"       ���"      �"       ��                        v      /       Vk       !       V!      !       V�!      �!       V"      �"       V�"      $#       V                                                  z      z       0���z      �       0���0��0���      �       0��������      :      	 �����o      o       0���o      G        0���0��0��G       �        Z�����0���        !       Z�����U�!      !       0���!      !       0���0��0��B!      �!      	 ������!      �!       0����!      �!       0���0��0���!      �!       0��������!      �!       Z�����U��!      "      	 �����"      ?"       Z�����0��?"      C"       Z�����0��C"      H"       Z�����U�H"      �"       0���0��0���"      �"       0��������"      �"       0���0��0���"      �"       1���0��0���"      �"       1���R�0���"      :#       0�������                       �      �       ]�!      �!       ]�"      �"       ]�"      :#       ]                 �      �       }�1&} �" $ &�                       �      �      
 }1&}"��      �       Q�      �       R�      �      
 }1&}"�                 �      �       ���1&t " $ &�                 �      �       t u "#��@& $ &�                 �      �       ���1&}�1&t "} ��                   �      �       T�      �      
 t u "#���                  �      �       t ?&��      �       U                   �"      �"       z 	���"      #      
 ��# 	��                    �"      #       R#      #       ��v "# 	��                   �"      �"       q z ��"      #       U                     �"      #       r t �#      	#       Z	#      #       T                         l       0�$#      :#       0�                                     *       V*      8       Q8      K       VK      X       v 	��X      l       R$#      (#       V(#      ,#       v`�,#      1#       V1#      5#       R5#      :#       V                         l       ��� $ &
�| "#�$#      :#       ��� $ &
�| "#�                                        v q �       K       RK      l       Q$#      1#       R1#      :#       Q                 l      �       V                 l      �       ��                      �      �       r ����      �       T�      �       r ���                    �      �       Q�      �       ��v "# 	�v ���                     �      �       q  $ &
�| "#���              | x "#�              q  $ &
�| "#��                 �             T                                R            
 r y "#���                               r ?&�             Y                 5      @       q  $ &
�| "#��                   5      9       R9      @       ��                   9      @       R@      @      
 r x "#���                  9      @       r ?&�@      @       X                        �       !       ��  �!      �!       ��  "      �"       ��  �"      �"       ��                          �       !       T�!      �!       T"      �"       T�"      �"       T                            �      R        [R        !      	 t ���"��!      �!      	 t ���"�"      H"      	 t ���"�H"      �"       [�"      �"       [                        �       !       |���!      �!       |��"      �"       |���"      �"       |��                         �      G        |��G        !       |���!      �!       |��"      H"       |��H"      �"       |���"      �"       |��                         �              Y               |�R       V        RV       �        [�       �        |�                                        �      �       X�      �       ���              ~ |�� $ &�               ~ p �       .        Xy       �        X�       �        r� $ &u ��       �        x u ��       �        X"      Y"       XY"      r"       ���"      �"       ��                          �      G        Rb        !       R�!      �!       R"      �"       R�"      �"       R                          �      �       R�       !       ���!      �!       ��"      �"       ���"      �"       ��                            Q        TQ       �        �T�                             
        t ����0u"�
       &       
 t 0u"�z       �        �T����0u"�                    .       Q        SQ       g        Q�       �        Q                 .       Q        X                   T       g        T�       �        T                  V       g        T�       �        T                      �      �       U�      K       SK      M       �U�                      �      �       T�      L       VL      M       �T�                      �      �       U�      	       �U�	      #	       U                         �      9       0�9      E       T�      �       T�      �       0��      �       ��	      #	       0�                      �      9       0��      �       q ����      �       Y	      #	       0�                     �      �       Q�      �       q��      �       Q	      #	       Q                          9       0�	      #	       0�                   �      7       T	      #	       T                         �      9       0�9      h       Vh      n       v�n      	       V	      	       �U#	      #	       0�                     �      �       U�      	       �U�	      #	       U                     �      �       U�      	       �U�	      #	       U                 �      �       [                       �             P             pP�             P	      #	       P                  Q      r       Z                 [      r       0�                      �      �       1��      �       z��      	       z�"	      #	       1�                 �      �       Z                  �      	       T                  �      	       Q                    �      �       u�      	       �U#"	      #	       u                      0	      �	       Q�	      1
       Q1
      4
       q��4
      �       Q                    0	      �	       R�      �       R                 0	      �       T                 0	      �       U                                   �	      �	       0��	      �	       [�	      �	       0�D
      O
       [O
      �
       q!�8$8&��
      �
       [�
             q!�8$8&�k      �       q!�8$8&��      �       [�      �       q!�8$8&�                             �	      �	       P�	      �	       q0�	      �	       qh�	      �	       q0�	      9
       PD
      �       P�      �       P                      D
      O
       0��
      �
       0��      �       0�                       �	      �	       w D
             w k      �       w �      �       w                        �	      �	       �DD
             �Dk      �       �D�      �       �D                    S
      �
       Vk      �       V                      Z
      ]
       ~ s �]
      �
       ^k      �       ^                    �
      �
       S�
      �
       S                    �
             V�      �       V                      �
      �
       ~ s ��
             _�      �       _                 �	      �	       0�                    �	      	
       V
      9
       V                      �	      	
       ^
      
       ~ s �
      9
       ^                        %       0�                    %      5       V8      k       V                      %      5       _F      L       ~ s �L      k       _                            �      �       U�      
       S
             �U�      �       S�      �       �U��      �       S                            �      �       R�             ^             �R�             ^      �       �R��      �       ^                            �      �       X�             \             �X�             \      �       �X��      �       \                 �      �       ��q  �                            �      �       T�             V      �       V�      �       s �      �       V�      �       P�      �       V�      �       P�      �       ~                        �      �       Q�      �       qP��             Q�      �       Q                       �      �       R�      �       rt��             R�      �       R                      �      |       _�      �       _�      �       _                           j       _j      |       h��      �       h�                        f       S                                      0�      $       V$      (       P1      5       V5      :       0�:      L       ��                                 0�5      :       } ���:      L       Q                         5       ]5      C       }�C      f       ]                                    0�      V       \V      ]       T]      a       |�a      f       \                       f       ^                          x      |       0��      �       \�      �       T�      �       |��      �       \                            �      �       U�      �       S�      �       �U��             S             �U�      !       U                              �      �       T�      �       V�      �       �T��      �       T�             V             �T�      !       T                            �      �       T�      �       V�      �       �T��      �       T�             V             �T�                          �      �       U�      �       S�      �       �U��             S             �U�                      �      �       P�      �       P             P                   �      �       u �      �       s                  �      �       s                    �      �       T�      �       V                 �      �       s�                     �      �       s��             s� �             �U#H�                     �      �       s��             s� �             �U#H�                 �      �       T                   �      �       P�      �       s(                   �      �       p ����Hs0"H��      �       s(�����Hs0"H�                 �             V                 �             s� �                   �             s� �             �U#H�                   �             s� �             �U#H�                  �      �       V                   �      �       P�      �       s�                    �      �       p ����Hs� "H��      �       s� �����Hs� "H�                      0      5       Q5      9       qy�9      �       �Q�                          0      W       RW      `       �R�`      |       R|      �       P�      �       �R�                      R      W       X`      l       Xl      �       Q                         R      W       Q`      i       Qi      o       sy�o      u       �Q#3%�u      �       S�      �       �Q#3%#	��                          �      �       U�             \             �U�      -       \-      0       �U�                    �      �       T�      �       t ����1����-( ��      0       �T����1����-( �                  �      �       Q                      �      �       R�             S      *       S                        �             ]            " �T1�T $0)( ����34$�U"#�      /       ]/      0      " �T1�T $0)( ����34$�U"#�                        0       P                 �             |                         p      {       U{      �       T�      �       �U��      �       T                      x      {       U{      �       T�      �       �U�                  {      �       U                            `      �       U�      �       S�      �       u���      �       �U��      �       S�      �       �U�                          `      �       T�      �       V�      �       �T��      �       V�      �       �T�                  c      w       P                          p      �       T�      �       V�      �       �T��      �       V�      �       �T�                            p      �       U�      �       S�      �       u���      �       �U��      �       S�      �       �U�                    �      �       P�      �       P                      z      �       \�      �       T�      �       \                           z      �       u��      �       s��      �       u���      �       �U#��      �       s��      �       �U#�                 z      �       \                   z      �       T�      �       V                   z      �       u��      �       s�                             z      �       u��      �       s��      �       s� ��      �       u`��      �       �U#H��      �       s��      �       �U#�                             z      �       u��      �       s��      �       s� ��      �       u`��      �       �U#H��      �       s��      �       �U#�                 z      �       T                   z      �       P�      �       u(                   ~      �       p ����Hu0"H��      �       u(�����Hu0"H�                   �      �       \�      �       T                   �      �       V�      �       �T�                     �      �       s� ��      �       u`��      �       �U#H�                     �      �       s� ��      �       u`��      �       �U#H�                     �      �       s� ��      �       u`��      �       �U#H�                  �      �       V                   �      �       P�      �       s�                    �      �       p ����Hs� "H��      �       s� �����Hs� "H�                        �             U      �       ]�      �       �U��      F       ]                      �      �       T�              t�              �T�                    �      �       Q�      F       Q                    �      �       V�      F       V                          �      �       S�      �       x �             S             P      F       S                   �             1�/      �       0��      F       0�                �      �       ��^  �                      !      8       q�0$0&��             q �0$0&�             q�0$0&�>      F       q �0$0&�                    /      �       U�      F       U                            /      8       S8      F       PF      M       p�M      �       P�      �       Z�             V      $       P                    /      8       Y�             Y>      F       Y                  /      �       Y�      F       Y                             8       0��      �       0��             1�             0�>      F       1�                  $      >       P                                              @#      i#       Ui#      �#       ��|�#      $       �U�$      �*       ��|�*      d-       �U�d-      �-       ��|�-      �.       �U��.      �.       ��|�.      4       �U�4      74       ��|74      g5       �U�g5      o5       ��|o5      �7       �U��7      8       ��|8      B8       �U�                                  @#      �#       T�#      �#       _�#      $       �T�$      �'       _�'      g5       �T�g5      o5       _o5      �7       �T��7      8       _8      B8       �T�                    @#      �#       Q�#      B8       ��|                                              @#      w#       Rw#      �#       ��|�#      $       �R�$      �*       ��|�*      d-       �R�d-      �-       ��|�-      �.       �R��.      �.       ��|�.      4       �R�4      74       ��|74      g5       �R�g5      o5       ��|o5      �7       �R��7      8       ��|8      B8       �R�                         �)      �)       P�)      4       ��{74      g5       ��{o5      �7       ��{8      B8       ��{                                   l*      �*       0��*      �*       ��|�*      *+       [*+      d-       ��|�-      �.       ��|�.      �3       ��|�3      4       ��|�#�74      g5       ��|o5      �7       ��|8      B8       ��|                          a#      �#       Q�#      �#       ��|$      �)       ��|4      74       ��|g5      o5       ��|�7      8       ��|                          a#      i#       Ui#      �#       ��|$      �)       ��|4      74       ��|g5      o5       ��|�7      8       ��|                            a#      �#       T�#      �#       _$      �'       _�'      �)       �T�4      74       �T�g5      o5       _�7      8       _                            a#      i#       ��}�i#      z#       Uz#      �#       ��}�$      �)       ��}�4      74       ��}�g5      o5       ��}��7      8       ��}�                                �#      �#       S$      �$       S�$      �*       ��|d-      �-       ��|�.      �.       ��|4      74       ��|g5      o5       ��|�7      8       ��|                     s$      �$       0��$      �$       T�$      �$       R%      %       T                      �$      �$       T�$      %       Tg5      o5       T                 s$      �$       0�                           s$      ,%       \,%      9%       S9%      �'       ��|g5      o5       \�7      �7       S�7      8       ��|                   s$      %       Pg5      o5       P                          �$      �$       Q�$      �$       px�$      �$       Q�$      �$       pg5      o5       Q                     �$      �$       Z�$      �$       Q�$      %       Rg5      o5       Z                         %      ,%       \,%      9%       S9%      �'       ��|�7      �7       S�7      8       ��|                     %      ,%       \,%      �'       S�7      8       S                          %      9%       P9%      �'       \�7      �7       P�7      �7       �7      8       \                       %      9%       0�9%      �'       V�7      �7       0��7      8       V                            9%      \%       Q\%      &       s ��|3&9��8�`&      �&       Q�&      �&       s ��|3&9��8��&      $'       s ��|3&9��8��7      8       s ��|3&9��8�                              9%      �%       P�%      &       s��|3&9��8�d&      �&       P�&      �&       s��|3&9��8��&       '       s��|3&9��8� '      $'       P�7      8       s��|3&9��8�                        s%      &       U�&      �&       U�&      $'       U�7      8       U                       s%      &       T�&      �&       T�&      $'       T�7      8       T                        �%      &       Q�&      �&       Q�&       '       Q�7      8       Q                        �%      &       R�&      �&       R�&       '       R�7      8       R                  s%      �%       T '      $'       T                  s%      �%       U '      $'       U                       �%      �%       X�%      �%       u ?&u 'u ?&� '      
'       X
'      $'       u ?&u 'u ?&�                  �%      �%       R '      $'       R                   s%      �%       4� '      $'       4�                    �%      �%       R�&      �&       R�&      �&       R�7      �7       R�7      �7       R                    �%      �%       Q�&      �&       Q�&      �&       Q�7      �7       Q�7      �7       Q                       �%      �%       Y�&      �&       q ?&q 'q ?&��&      �&       Y�&      �&       q ?&q 'q ?&��7      �7       Y�7      �7       q ?&q 'q ?&�                     �%      �%       P�&      �&       P�&      �&       P�7      �7       P�7      �7       P                   �%      �%       4��&      �&       4�                      H'      g5       0�o5      �7       0��7      �7       0�8      B8       0�                          H'      �+       ��}��+      �+       R�+      g5       ��}�o5      �7       ��}��7      �7       ��}�8      B8       ��}�                      H'      o'       Qo'      �'       qp��'      �'       Q�7      �7                              P'      s'       Ps'      �'       p���'      �'       P�7      �7       ��}                  P'      b'       R�7      �7       0�                          �'      �'       0��'      �'       ��|�'      �'       P�'      0)       ��|4      74       ��|                    �'      (       Y(      `(       S                             �'      (       Y(      (       V(      v(       Vv(      )       ��|)      )       S)      0)       ��|4      4       ��|4      74       ^                                �'      �'       Y�'      (       S(      v(       ��|v(      �(       S�(      �(       ^�(      )       ^)      )       S)      +)       V+)      0)       S4      74       S                      (      (       \(      (       V(      X(       \                           v(      �(       S�(      �(       V�(      �(       ^�(      +)       V+)      0)       S4      74       V                           �'      	(       V	(      q(       ��{v(      �(       U�(      �(       ])      +)       ]+)      0)       U                      �'      v(       ^v(      )       ��|)      0)       \4      74       ��|                                  (      (       ]-(      [(       ][(      v(       \v(      �(       U�(      �(       _�(       )       _ )      +)       ]+)      0)       U4      74       ]                              (      (       _9(      v(       _v(      �(       ��|�(      �(       S�(      )       S)      0)       \4      74       \                     Q(      v(       Pv(      )       ��|)      0)       P                      �(      �(       P�(      0)       P4      74       P                       �'      �(       0��(      )       \)      0)       _4      74       _                �#      $       ��}�                 �#      $       S                                          �)      !*       |�!*      )*       ��~#�)*      �+       |��+      �+       q��+      �+       |��,      �-       |��.      �.       |��.      c/       ��~#�c/      i/       |��0      �0       ��~#��0      41       |�4      4       ��~#�05      g5       |�o5      �5       |�                                         �)      !*       |��!*      )*       ��~#��)*      �+       |���+      �+       q���+      �+       |���,      �-       |���.      �.       |���.      c/       ��~#��c/      i/       |���0      �0       ��~#���0      41       |��4      4       ��~#��05      g5       |��o5      �5       |��                            �)      *       ^*      *       Td-      r-       ^�.      �.       T�.      �.       ^�.      �.       T                               �)      �)       U�)      �)       ��|�)      *       P*      *       U*      *       Qd-      r-       U�.      �.       P�.      �.       U                                   �)      �*       ^�*      d-       ��|d-      �-       ^�-      �.       ��|�.      �.       T�.      �.       ^�.      4       ��|74      g5       ��|o5      �7       ��|8      B8       ��|                             �)      �)       U�)      d-       ��|d-      r-       Ur-      4       ��|74      g5       ��|o5      �7       ��|8      B8       ��|                      �)      �*       Sd-      �-       S�.      �.       S                            �)      �)       t 	���)      �)       T�)      �*       Vd-      r-       Tr-      �-       V�.      �.       V                                 �)      �)       0��)      )*       1�)*      d-       ��|d-      r-       0�r-      �.       ��|�.      �.       1��.      4       ��|74      g5       ��|o5      �7       ��|8      B8       ��|                �)      �)       U                �)      �)       ��|#�                
  �)      �)       P�)      �)      
 p q "#���                  �)      �)       p ?&��)      �)       Q                    k6      �6       P7      �7       Q                         d6      �6       Q�6      �6       x�7      7       P7      <7       [<7      T7       x�                  *6      �7       U                  d6      �7       T                    �6      �6       R�6      �6       R                    )7      \7       R_7      �7       R                               �*      �*       ��|�*      *+       [*+      d-       ��|�-      �.       ��|�.      4       ��|74      g5       ��|o5      �7       ��|8      B8       ��|                               �*      �+       ��}��+      �+       R�+      d-       ��}��-      �.       ��}��.      4       ��}�74      g5       ��}�o5      �7       ��}�8      B8       ��}�                            �*      �*       Q�*      �*       qp��*      +       Q+       +       qp� +      5+       Q�5      �5       Q                             �*      �*       Z�*      �*       P�*      �*       p���*      +       P+       +       p�� +      *+       P�5      �5       Z                   �*      �*       Y�5      �5       Y                                %+      5+       0�5+      M+       [P+      y+       [�,      d-       [�-      �-       [05      g5       [o5      �5       [�5      �5       0�                     5+      @+       s �,      -       s -      d-       V                      -      -       V-      8-       U8-      =-       Q=-      d-       U                  �,      d-       P                   -      
-       U
-      d-       Q                        `+      m+       Q�-      �-       Q05      g5       Qo5      �5       Q                       `+      m+       Q�-      �-       Q�-      �-       P05      35       P                         `+      m+       Q�-      �-       Q05      55       Q55      g5       Po5      �5       P                             �+      �+       U�+      �,       ��|�-      �.       ��|�.      �3       ��|74      05       ��|�5      �7       ��|8      B8       ��|                      �+      �+       ��}��+      �+       R�+      �+       ��}�                  �+      �+       ��|                      �+      �+       \�+      �+       Q�+      �+       \                       �+      �+       S�+      �+       U�+      �+       sP��+      �+       S                   �+      �+       P�+      �+       u                      �+      �,       ��|�-      .       ��|�4      5       ��|                     �+      �,       ��}��-      .       ��}��4      5       ��}�                     �+      �,       ��|�-      .       ��|�4      5       ��|                        �+      P,       \P,      �,       V�-      �-       \�4      �4       V                  �+      U,       _                          �+      K,       0�K,      _,       Q_,      p,       \p,      �,       Q�-      �-       0��4      �4       Q                                          �+      ],       ]],      �,       ��|�-      �-       ]�-      �.       ��|�#��.      41       ��|�#�41      4       ��|�#�74      �4       ��|�#��4      �4       ��|�#��4      �4       ��|�4      05       ��|�#��5      �7       ��|�#�8      78       ��|�#�78      B8       ��|�#�                   �+      �+       p  $ &
���~"#��+      �+       } $ &
���~"#�                   �+      �+       p  $ &
�q "#��+      �+       } $ &
�q "#�                            �+      ,       P,      4,       P4,      �,       ��|�-      �-       P�-      .       ��|�4      5       ��|                      _,      p,       \|,      �,       \�4      �4       Q                  �,      �,       ^                  �,      �,       S                 �-      �-       ��}                   �-      �-       ��}�-      .       P                 �4      �4       ��}                 �4      �4       ��}                      7.      �.       S74      i4       S5      05       S                          7.      H.       R_.      �.       R�.      �.       s(74      i4       R5       5       R                              .      �.       U�.      �.       s0r � $ &��.      �.       s0s(� $ &�74      C4       UC4      J4       s0q �J4      i4       s0r � $ &�5       5       U                  �.      �.       u q ��.      �.       U                   �.      �.       Q�.      �.      
 q r "#���                  �.      �.       q ?&��.      �.       R                 74      G4       U                   G4      N4       UN4      N4      
 q u "#���                  G4      N4       u ?&�N4      N4       Q                      �.      �0       ��|i4      �4       ��|�5      6       ��|8      78       ��|                      �.      �0       ��}�i4      �4       ��}��5      6       ��}�8      78       ��}�                      �.      c/       ��|� $ &
���~"#�c/      i/       ��|� $ &
�| "#��5      �5       ��|� $ &
�| "#�                      /      /      
 ��~p "#�/      c/       ��|
���~"#��5      �5       ��|
�| "#�                   /      c/       ��~�5      �5       ��~                            /      c/       0�c/      �0       Vi4      �4       V�5      �5       0��5      �5       P�5      6       V8      78       V                             /      ./       0�./      c/       Rc/      k/       0�k/      �0       \i4      �4       \�5      �5       R�5      6       \8      78       \                   /      �/       S�5      �5       S                        /      �0       ^i4      �4       ^�5      6       ^8      78       ^                                    /      ./       S./      c/       Pc/      k/       Sk/      �/       R�/      �/       p �/      �/       R�/      �0       Si4      �4       S�5      �5       P�5      6       S8      78       S                  �/      �/       P                    g0      �0       r ����3$v "�5      �5       r ����3$v "6      6       r ����3$v "                 i4      �4       v                                (0      L0       0�L0      _0       Q_0      b0       Rb0      g0       Qg0      �0       \�0      �0       Pi4      �4       0��5      �5       P6      6       P                       �0      �0       U�5      6       U8      8       U8      8       s0                   i4      k4       u p �k4      u4       U                   u4      |4       U|4      |4      
 p u "#���                  u4      |4       u ?&�|4      |4       P                  �5      �5       u z ��5      �5       U                   �5      �5       P�5      �5      
 p q "#���                  �5      �5       p ?&��5      �5       Q                     �0      �1       ��|*2      �3       ��|78      B8       ��|                     �0      �1       ��}�*2      �3       ��}�78      B8       ��}�                 �0      41       ��|� $ &
���~"#�                 �0      41       ��|� $ &
���~"#�                      1      ~1       Yl3      z3       Y�3      �3       Y                     1      �1       _*2      �3       _78      B8       _                  1      41       P                      ?1      ~1       Ql3      �3       Q�3      �3                                G1      S1       0�S1      ~1       S�1      �1       R.3      ?3       Vl3      �3       S                              G1      ~1       T~1      �1       R�1      �1       R*2      32       R32      l3       Vl3      �3       T78      B8       V                         G1      S1       QS1      ~1       P�2      I3       Rl3      v3       P�3      �3       Q                     G1      S1       0�S1      ~1       Rl3      �3       R                      ]2      �2       X�2      �2       ��|I3      l3       T78      B8       T                            f2      i2       T�2      �2       T�2      �2       ^I3      Y3       x t �Y3      l3       X78      =8       X=8      B8       ^                    ]2      i2       [�2      �2       [�2      �2       ��|                          i2      �2       Q�2      �2       U�2      �2       ��|V3      l3       Q78      B8       Q                     �2      �2       r0�2      )3       r0?3      I3       r0                            �2      �2       Q�2      �2       r0t ��2      3       Q3      )3       r0t �?3      C3       QC3      I3       r0t �                    �2      �2       Q!3      ?3       Q                      i2      �2       @<$��2      �2       PV3      l3       @<$�78      B8       @<$�                   �2      �2       q ~ ��2      �2       Q                   �2      �2       Q�2      �2      
 q { "#���                  �2      �2       q ?&��2      �2       [                 ?3      G3       Q                  3      3       Q3      3      
 q { "#���                  3      3       q ?&�3      3       [                  3      3       Q3      3       r0�t �                 3      3       Q                3      3       q ?&�                r3      �3       s0                   ~3      �3       P�3      �3      
 p r "#���                  ~3      �3       p ?&��3      �3       R                �3      �3       q0                   �3      �3       P�3      �3      
 p r "#���                  �3      �3       p ?&��3      �3       R                   �1      �1       ��|�1      *2       [                 �1      *2       ��}�                   �1      �1       0��1      *2       P                  �1      *2       Q                  �1      *2       Y                  �1      *2       Z                    P8      d8       Ud8      e8       �U�                    P8      d8       Td8      e8       �T�                    P8      d8       Qd8      e8       �Q�                    P8      d8       Rd8      e8       �R�                          p8      �8       U�8      -:       S-:      7:       �U�7:      A:       UA:      �:       S                            p8      �8       T�8      :       �T�:      %:       T%:      7:       �T�7:      A:       TA:      �:       �T�                            p8      �8       Q�8      :       �Q�:      %:       Q%:      7:       �Q�7:      A:       QA:      �:       �Q�                      �8      �8       Q�8      9       _:      %:       Q                          �8      �8       T�8      �8       t ����1����-( ��8      :       �T����1����-( �:      %:       t ����1����-( �%:      7:       �T����1����-( �A:      �:       �T����1����-( �                        �8      �8       U�8      -:       S-:      7:       �U�A:      �:       S                     �8       9       P%:      (:       Pa:      g:       P                             �8      �8      ' t ����1����-( ����0u "#��8      �8      ( �T����1����-( ����0u "#��8      :      ( �T����1����-( ����0s "#�:      %:      ' t ����1����-( ����0s "#�%:      -:      ( �T����1����-( ����0s "#�-:      7:      ) �T����1����-( ����0�U"#�A:      �:      ( �T����1����-( ����0s "#�                   �8      �8       u :      %:       s                      9      :       ^A:      a:       ^g:      �:       ^                     9      :       \A:      a:       \g:      �:       \                     9      :       VA:      a:       Vg:      �:       V                     9      :      ( �T����1����-( ����0s "#�A:      a:      ( �T����1����-( ����0s "#�g:      �:      ( �T����1����-( ����0s "#�                                9      �9       0��9      �9       P�9      :       0�:      :       P:      :       0�A:      a:       0�a:      a:       Pg:      �:       0��:      �:       P                    '9      V9       PV9      �9      	 s ��"#8                   �9      �9       ��A:      V:       ��                 �9      �9       V                 �9      �9       V                 �9      �9       ��                 �9      �9       \                 �9      �9       \                 �9      �9       ��                 �9      �9       ^                 �9      �9       ^                          �<      �<       U�<      �<       �U��<      �<       U�<      �<       S�<      =       �U�                        �<      �<       T�<      �<       �T��<      �<       T�<      =       �T�                          �<      �<       Q�<      �<       �Q��<      �<       Q�<      �<       V�<      =       �Q�                          �<      �<       Q�<      �<       �Q��<      �<       Q�<      �<       V�<      =       �Q�                        �<      �<       T�<      �<       �T��<      �<       T�<      =       �T�                          �<      �<       U�<      �<       �U��<      �<       U�<      �<       S�<      =       �U�                    �<      �<       P�<      =       P                         �<      �<       u��<      �<       �U#��<      �<       u��<      �<       s��<      =       �U#�                 �<      �<       u                     �<      �<       \�<      �<       \                    �<      �<       ]�<      =       ]                          =      /=       U/=      8=       �U�8=      Z=       UZ=      �=       S�=      �=       �U�                          =      /=       T/=      8=       �T�8=      e=       Te=      �=       V�=      �=       �T�                        =      /=       Q/=      8=       �Q�8=      _=       Q_=      �=       �Q�                          =      /=       R/=      8=       �R�8=      \=       R\=      �=       ]�=      �=       �R�                          =      /=       R/=      8=       �R�A=      \=       R\=      �=       ]�=      �=       �R�                        =      /=       Q/=      8=       �Q�A=      _=       Q_=      �=       �Q�                          =      /=       T/=      8=       �T�A=      e=       Te=      �=       V�=      �=       �T�                          =      /=       U/=      8=       �U�A=      Z=       UZ=      �=       S�=      �=       �U�                    j=      �=       P�=      �=       P                         =      /=       u�/=      8=       �U#�A=      Z=       u�Z=      �=       s��=      �=       �U#�                 =      =       u                     "=      /=       PA=      i=       P                    &=      3=       \A=      �=       \                                �&      
'       U
'      E'       �U�E'      i'       Ui'      �'       V�'      �'       �U��'      x(       Vx(      �(       �U��(      �(       U�(      �(       V                        �&      
'       T
'      ;'       S;'      B'       ~�~�B'      E'       �T�E'      �(       S                          �&      
'       Q
'      E'       �Q�E'      i'       Qi'      �(       �Q��(      �(       Q�(      �(       �Q�                                  �&      
'       R
'      E'       �R�E'      i'       Ri'      �'       \�'      �'       �R��'      /(       \/(      �(       �R��(      �(       R�(      �(       \�(      �(       �R�                     �&      B'       ^B'      E'       �T#��E'      �(       ^                       �&      
'       t��
'      ;'       s��;'      B'       ~P�B'      E'       �T#��E'      �(       s��                   �&      D'       _E'      �(       _                                   �&      '       0�'      3'       ��~E'      �'       0��'      �'       ��~�'      (       0�(      %(       P%(      *(       ��~*(      *(       P*(      �(       ��~�(      �(       0��(      �(       ��~                               �&      '       0�'      3'       ]E'      �'       0��'      �'       ]�'      (       0�(      "(       ]"(      *(       s��s��6$ $ &�*(      �(       ]�(      �(       0��(      �(       ]                    �&      �&       U�&      �&       �U�                      �&      �&       T�&      �&       u�~��&      �&       �T�                    �&      �&       Q�&      �&       �Q�                      �      �       U�      �       P�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                      p      }       U}      �       P�      �       �U�                        #      7#       U7#      �%       �U��%      �%       U�%      J&       �U�                        #      �#       T�#      �%       �T��%      �%       T�%      J&       �T�                        #      �#       Q�#      3%       �T#�%      �%       Q�%      J&       �T#                           #      �#       t �#      !$       P!$      3%       �T�%      �%       �T�%      �%       t �%      J&       �T                         C$      �%       W�%      �%       w��~��%      �%       W�%      �%       w��~��%      J&       W                      4%      Z%       P�%      �%       P�%      �%       P                    E$      $       p 
 �&      J&       p 
 �                    E$      $       W&      J&       W                      �      �       U�      �       T�      �       �U�                   �      �       u �      �       U                      P&      q&       Uq&      �&       V�&      �&       �U�                      P&      h&       Th&      �&       S�&      �&       �T�                   P&      r&       0�r&      �&       P                                            �      �       U�      *       ^*      -       �U�-      q       ^q      t       �U�t      T       ^T      w       Uw      �       ^�      �       U�      >       ^>      �       U�      i"       ^i"      l"       �U�l"      #       ^                    �      �       T�      #       ��~                      �      �       Q�             U�"      �"       U                        �      �       Q�             r�             q��"      �"       Q                         -      �       ��~�8$8&�-      e       ��~�8$8&�t      >       ��~�8$8&�      3       ��~�8$8&�2"      M"       ��~�8$8&�l"      �"       ��~�8$8&�                                   -      �       ^-      e       ^t      T       ^T      w       Uw      �       ^�      �       U�      >       ^>      >       U      3       ^2"      M"       ^l"      �"       ^                               =      N       0�N      �       ��-      e       ��t      d       ��d      j       ���#�      >       ��2"      M"       ��l"      �"       ��                       =      N       0�N      _       S�      �       S      >       S                          K       ~�      >       ~�                    @      K       T9      >       T                          �      �       ��~�8$8&�-      `       ��~�8$8&�t      (       ��~�8$8&�R      �"       ��~�8$8&��"      #       ��~�8$8&�                        �      �      	 u 1$~�"�             ��1$~�"      i       Tt      �       T                                          �      �       ^-      `       ^t      T       ^T      w       Uw      �       ^�      �       U�      >       ^>      �       U�      (       ^R      i"       ^i"      l"       �U�l"      �"       ^�"      #       ^                            �      �       U���      �       U�Q��      �       R�Q��      2       U�Q�2      i       U��t      �       U�Q�                                             �      )       V�\�)      ,       �\��      �       T���      �       T�Q��      �       P�Q��      "       T�Q�'      ;       V�S�;      >       V�Q�>      �       T�Q�t             V�\�      �       V���      �       V�S��      �       Z�S��      �       �S�2"      M"       T�Q�                                                �      �       V���      �       V�\��      �       R�\��      �       R�V��      �       \�V��      )       V�\�)      ,       �\�C      F       V��F      i       V�\�i      �      
 �������      �      
 ������-      T      
 ������t      t       V�\�t      �       U�Q��      �      
 ������2"      M"      
 ������l"      �"      
 ������                      �      �       P�      i       ~�t      �       ~�                               �      q       Pq      �       _�      �       _-      T       _t      �       P�      �       _2"      M"       _l"      �"       _                              �      �       ]�      �       \-      T       ]t      �       ]�      �       \2"      M"       ]l"      �"       ]                                          �      u       Su      �       V�      �       S�      �       V�             s�      �       S�      �       V�      �       ]�      �       V-      T       s�t      �       S�      �       ]2"      ="       Vl"      �"       s�                                                     	 r 8$8&�u      x       q 38$8&�x      �       v �38$8&��      j       v �38$8&��      �       v �38$8&��      �      	 p 8$8&�U      �      	 p 8$8&�-      T       v �38$8&�2"      ="       v �38$8&�l"      x"       v �38$8&�x"      �"       s�38$8&��"      �"       v �38$8&��"      �"       s�38$8&�                      �      �       T�      �       P�      �       T                  �      �       Q                                      0       T0      [       Q[      n       T-      T       Tl"      �"       T�"      �"       [�"      �"       Q�"      �"       [                                          0       Q0      U       TU      a       Pa      n       Q-      T       Ql"      {"       Q{"      �"       [�"      �"       P�"      �"       T�"      �"       Q�"      �"       T                                "      0       R0      O       XO      n       R-      T       Rl"      �"       R�"      �"       Q�"      �"       R�"      �"       X                                    %      0       X0      L       RL      R       PR      n       X-      T       Xl"      �"       X�"      �"       Q�"      �"       X�"      �"       R�"      �"       Q                    X      a       [a      n       YI      T       Y                    a      a       Ya      n       [O      T       U                            �      >       V]      m       Vm      p       Rp      �       V�      �       Z�      �       V                        �      ;       S;      >       Q`      �       S�      �       S                                       �       ^�      �       U�             ^>      �       U�      3       ^R      2"       ^M"      i"       ^i"      l"       �U��"      #       ^                                �      �       \�      �       |��             \>      (       \R      �       \�!      �!       \M"      e"       \�"      #       \                            �             S>      (       SR      �       S�!      �!       SM"      b"       S�"      #       S                     �      �       s(�      �       T             T                             �      �       ]             Q>             ]R      �       ]�!      �!       ]M"      g"       ]�"      #       ]                        ^      �       U�             ^R      2"       ^M"      X"       ^�"      #       ^                                     �      �       ���      �       V�      �       _�              v��       !       V!      !       v�!      $!       �$!      �!       _�!      �!       V�!      �!       V�!      "       V""      2"       V                      �      �        \!      �!       \"      ""       \                         �      �       0��      �       ���      �       P�      �!       ���!      2"       ��                                                          �      
       Q
             UR      �       U�      �       P�             P             T      �       P�      �       T�      �       P               Q                U        X        QX       `        p `       o        Qo       |        U|       �        Q�       !       P�!      �!       P�!      �!       Q�!      "       P"      ""       Q""      2"       PM"      X"       U�"      #       P                                             �             UR      �       U             T$      �       T                U)       `        Uo       |        U�       �        U�       !       T�!      �!       T�!      �!       U�!      "       T"      ""       U""      2"       TM"      X"       U                                  S!      �!       S                          �       ]�              ]!      �!       ]                    �      �       R�!      �!       R                      �             TR      �       T�!      �!       TM"      X"       T                        �             0�      F       PK      �       P�      �       P$!      <!       P                              F       Qd      s       Qs      v       Tv      �       Q                          F       Rh      �       R                            :       x  $ &q �:      F       ~� $ &q ��      �       x  $ &q �                             :       r x "1x  $ &�:      F       ~� $ &r "1~� $ &��      �       r t "1x  $ &��      �       r x "1x  $ &�                	 ^      t       ���                 t      }       ���                 }      �       ���                   �      
       Q�!      �!       Q                     �      
       ����!      �!       ����!      �!       R                           �      �       ����      �       R�      �       ����      
       R�!      �!       ����!      �!       R                       �      �       ���             P�!      �!       ���!      �!       r                    �      
       0��!      �!       0�                   �       �        Q"      "       Q                     �       �        ���"      "       ���"      "       P                         �       �        ����       �        p��       �        ����       �        p�"      "       ���"      "       P                            �       �        P�       �        T�       �        P�       �        T"      "       P"      "       p                      &      U       P�!      �!       P""      2"       P                       &      U       ����!      �!       ���""      -"       ���-"      2"       Q                           &      :       ���:      L       q�L      L       ���L      U       q��!      �!       q�""      -"       ���-"      2"       Q                              +      :       Q:      L       RL      P       QP      U       R�!      �!       R""      -"       Q-"      2"       q                    b      �       P�!      �!       P                     b      �       ����!      �!       ����!      �!       U                           b      z       ���z      �       U�      �       ����      �       U�!      �!       ����!      �!       U                    g      �       Q�!      �!       Q                   g      �       R�!      �!       R                   �       !       P�!      "       P                     �       !       ����!      �!       ����!      "       U                           �       �        ����       �        U�       �        ����       !       U�!      �!       ����!      "       U                    �       !       Q�!      "       Q                   �       !       p �!      "       p                  �      �       s�7
���                   +       [        Q"      ""       Q                     +       `        ���"      "       ���"      ""       P                         +       ?        ���?       C        p�C       C        ���C       U        p�"      "       ���"      ""       P                            0       ?        P?       C        TC       G        PG       U        T"      "       P"      ""       p                         P      �       T�      �       Q�      �       �T��      <       T                              P      x       Qx      �       �Q��      *       Q*      �       �Q��      �       Q�      �       �Q��      <       Q                              P      x       Rx      �       �R��      J       RJ      �       �R��      �       R�      �       �R��      <       R                                P      x       Xx      �       �X��             X      �       �X��      �       X�      �       �X��      +       X+      <       �X�                                P      x       Yx      �       �Y��             Y      �       �Y��      �       Y�      �       �Y��      '       Y'      <       �Y�                               n      x       Z�      �       P�      �       Z�      g       Zg      �       S�      �       Z�      �       S�      <       Z                          q      x       S�      d       Sd      g       Q�      �       S�      <       S                           q      }       Z�      A       ZA      �       X�      �       Z�      �       X�      <       Z                    �      �       Pl      �       t 3&0$0&u�� $ &s u� "��      �       q 0$0&u�� $ &s u� "�                 l      �       �t 70$0&&�                             �             x�7
���      �       �X#�7
����      �      	 | 7
����      �       �X#�7
����            	 | 7
���      +       x�7
���+      <       �X#�7
���                      �      1       T1      5       P5      P       �T�                    �      �       Q�      P       �Q�                        �             R             �R�             R      P       �R�                    �      �       X�      P       �X�                    �      �       Y�      P       �Y�                      �             Q      9       Q9      O       x �Q"1x  $ &u ��&�                       �             p r �             P              P       P       x  $ &�R�                  K      P       P                                       &       T&      a       �T�a      �       T�      =       �T�=      C       TC      U       �T�U      �       T�      �       �T�                                     &       Q&      a       �Q�a      �       Q�      =       �Q�=      E       QE      U       �Q�U      �       Q                                     &       R&      a       �R�a      �       R�      =       �R�=      E       RE      U       �R�U      �       R                                       &       X&      a       �X�a      �       X�      =       �X�=      E       XE      U       �X�U      �       X�      �       �X�                                         &       Z.      B       RB      K       PK      Z       Za      �       Z�             [             Q=      S       ZS      U       [U      �       Z                                      &       [&      Z       u� $ &�R�a      �       [�      �       Q�      =       u� $ &�R�=      P       [P      U       u� $ &�R�U      �       [                                 +       Za      �       Z�      )       T=      E       ZE      U       TU      �       Z                         <      B       r 3&�B      K       p 3&�K      Z       z 3&��             { 3&�             q 3&�             Q                   <      Z       z 7��             { 7�             q 7�                             a      �       x�7
����      =       �X#�7
���=      E      	 v 7
���E      U       �X#�7
���U      �      	 v 7
����      �       x�7
����      �       �X#�7
���                      �
      �       U�      �       �U��      �       U                  �
      �
       T�
      �       �T�                    �
      {       Q{      �       �Q�                    �
      4       R4      �       �R�                    �
             X      �       �X�                    �
             Y      �       �Y�                                        4       Y4      G       y r ����&�G      J       q z "1z  $ &r ����&�J      `       q z "1z  $ &u �����&�`      x       Rx      �       Y�      �      > z �Q"1z  $ &u ��&x z �Q"1z  $ &u ��&0*( ��      �      = z �Q"1z  $ &u ��&0z �Q"1z  $ &u ��&0*( ��      �      = z �Q"1z  $ &u ��&0z �Q"1z  $ &u ��&0*( �                          h       Pm      �       P                    �      �       R�      �       P�      �       R                     �
             x�7
���      �       �X#�7
����      �       �X#�7
���                 �      �       Y                  �      �       Q�      �       P�      �       p��      �       P                   �      �       X�      �       X                  �      �       T                    �
      �
       Q�
      �
       �Q�                  �
      �
      	 q  $ &�                      
      _
       U_
      a
       Ra
      �
       U                      S
      _
       U_
      �
       R�
      �
       R�
      �
       R                    
      
       Q
      S
       PS
      �
       Q                    W
      �
       P�
      �
       P                              �      S       US      �	       S�	      �	       v�}��	      �	       �U��	      �	       S�	      �	       v�}��	      
       �U�                    �      X       TX      
       �T�                    �      X       QX      
       �Q�                    �      X       RX      
       �R�                    �      X       XX      
       �X�                    �      X       YX      
       �Y�                       X      �       s� #8E	      d	       s� #8�	      �	       s� #8�	      �	       s� #8                       X      �       s� #(E	      d	       s� #(�	      �	       s� #(�	      �	       s� #(                       X      �       s� #E	      d	       s� #�	      �	       s� #�	      �	       s� #                       X      �       s� #E	      d	       s� #�	      �	       s� #�	      �	       s� #                       X      �       s� E	      d	       s� �	      �	       s� �	      �	       s�                       f      �       RY	      d	       R�	      �	       R                      f      �       TY	      d	       T�	      �	       T                      t      �       QY	      d	       Q�	      �	       Q                      t      �       XY	      v	       X�	      �	       X                    �      �       1��	      �	       2�                    �      �       Y�      	       Q                                     E       UE      K       SK      N       |�}�N      Q       �U�Q      �       S�      �       |�}��      �       �U�                           U       TU      �       �T�                           U       QU      �       �Q�                           U       RU      �       �R�                           U       XU      �       �X�                       U      {       s� #(�      �       s� #(Q      \       s� #(n      �       s� #(                       U      {       s� #�      �       s� #Q      \       s� #n      �       s� #                       U      {       s� #�      �       s� #Q      \       s� #n      �       s� #                       U      {       s� �      �       s� Q      \       s� n      �       s�                      U      {       s� #(�      �       s� #n      �       s� #(                     U      {       s� #�      �       s� #(n      �       s� #                    �      �       2�|      �       1�                    �             Y             Q                            �      �       U�             S             �U�      Z       SZ      `       �U�`      �       S                                        �      �       T�             \             �U#X      &       T&      ]       \]      `       �T�`      {       T{      �       \�      �       T�             \      >       T>      �       \                                      �      �       Q�             V             �U#`      [       V[      `       �Q�`      u       Qu      �       V�      �       Q�             V      '       Q'      �       V                   �      �       u� �      �       y �                   �      �       u� �      �       p �                �              V                �              \                 �      �       u�                    �      �       u� �      �       T                  �      �       U�              S                 �              P                 �              ]                      �      �       U�      �       V�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                        �      �       R�      �       P�      �       p ��      �       �R�                      �      �       X�      �       r ��      �       �X�                  �      �       S                  �      �       P                  �      �       \                            �      �       U�      �       S�      �       �U��      }       S}      �       �U��      �       S                    �      �       T�      �       �T�                            �      �       Q�      �       _�      �       �Q��      �       _�      �       �Q��      �       _                            �      �       R�      �       P�      �       �R��      �       P�      �       V�      �       �R�                        �      �       X�      �       �X��      �       X�      �       �X�                          �      �       QH      l       Z�             Q,      b       Z�      �       Q                               �      �       ^�      �       |<      K       PK      l       u�      �       P�             |,      <       u�      �       |                        �      �       P�      �       V�             P      ~       V�      �       P                      �      �       ^�      �       ^�      �       ^                       �             P�      �       P�      �       V�      ,       P�      �       P                                �      7       \7      l       Um             ��      �       U�      �       \�      ,       \,      <       UV      �       U�      �       \                             �      l       Tl             ��      �       T�      �       t��             T             R             r�      ,       T,      C       t�C      �       T�      �       R                                �      <       U<      x       \x      �       �U��      �       \�      �       U�      .       \.      5       �U�5      �       \                                �      <       T<      x       V�      �       V�      �       T�      �       X�             ��      ,       V5      �       V                                  �      <       Q<      =       S=      �       �Q��      �       S�      �       Q�      +       S+      5       �Q�5      u       Su      �       �Q�                            �      (       R(      <       Z<      �       �R��      �       R�             ��      �       �R�                            �             X      x       ^x      �       �X��      2       ^2      5       �X�5      �       ^                          �      <       Y<      �       �Y��      �       Y�      
       ]
      �       �Y�                                 �             r t �      <       [<      5       �R�T�5      :       1�:      x       P�      �       �R�T��      �       [�             ��      i       �R�T�i      u       	��u      �       P                          �      �       _�      �       �X�Q��      4       _4      5       �X�Q�5      �       _                          4      7       P7      �       ]�      �       }��      �       ]�      �       ]
             ]                        T      T       UT      �       Y�      �       ���      �       U�      �       Y                     <      �       P�      �       P
             0�                     T      �       R�      �       ���      �       R                          �             Y      E       ��E      S       Y      J       YJ      u       ��u      �       Y                        '      ,       P,      x       U[      `       P`      �       U                    5      x       Qi      �       Q                      E      c       Rc      f       r q "�f      x       Ru      �       R                   E      x       Xu      �       X                             �             Q              T       3       u u"�Q      r       Qr      {       T{      �       uu"��      �       Q                        �      #       R#      3       uu "�T      u       Ru      �       uu("�                            �             P      	       u0u "�	             P      #       u0r "u "�#      3       u 1$u0"u"�T      ]       P]      a       u8u("�a      x       Px      �       u(1$u8"u"�                        �      �       Q�      �       u u"��      �       Q�      �       uu"�                              �      �       P�      �       R�      �       u u"��      �      	 u� u"��      �       P�      �       R�      �       u(u"��      �      	 u� u"�                         �      �       T      -       T-      6       p 6      F       QF      Q       T                  �      e       Y                                  �      �       p��      �       z��      �       r��      �       R�      �       P�      �       R�      �       p��      �       P             RF      Q       R                    -      6       p ?      F       Q                      �              T      u       �T�u      �       T                        �             	 p q8�      
       r 8�
      I      	 p q8�u      �       r 8�                 .      U       Q                     )      ')       U')      S)       �U�                     )      *)       T*)      K)       SK)      S)       �T�                     )      .)       Q.)      S)       �Q�                     )      .)       R.)      K)       VK)      S)       �R�                 7)      K)       �U�                 7)      K)       �Q�                 7)      K)       V                 7)      K)       S                 K)      K)       0�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                    �      �       R�      �       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                    �      �       R�      �       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       Q�      �       Q�      �       �Q0�Q $@L$.( �                    �      �       R�      �       �R�                                      0      d       Ud      �       V�      �       �U��      �       V�             �U�      |       V|      �       �U��             V      "       �U�"      z       Vz      �       �U�                                      0      �       T�      �       �T��      �       S�             �T�      |       S|      �       �T��             S      "       �T�"      �       S�      r       ��~r      �       �T�                                            0      �       Q�      �       �Q��      �       Q�             �Q�      +       Q+      |       _|      �       �Q��      �       Q�             _      "       �Q�"      1       _1      �       �Q��      �       _�      �       �Q�                                  0      |       R|      �       �R��      �       R�             �R�      +       R+      �       �R��      �       R�      �       ��~�      �       �R�                                0      �       X�      �       �X��      �       X�             �X�      +       X+      �       �X��      �       X�      �       �X�                                     a      �       ^�      �       �T#���      �       ^�             �T#��      |       ^|      �       �T#���             ^      "       �T#��"      �       ^�      r       ��~r      �       �T#��                                     a      �       t���      �       �T#���      �       s���             �T#��      |       s��|      �       �T#���             s��      "       �T#��"      �       s���      r       ��~#��r      �       �T#��                         a      �       Z�      �       Z      +       Z�      �       Z�      �       ��}                                   a      �       0��      �       \�      �       0��      �       R�             \      �       0��      �       \�      �       0��      �       \�      r       ��~                                   a      �       0��      �       ]�      �       0��      �       R�             ]      �       0��             R      �       ]�      �       0��      �       ]�      r       ��~                                           a      �       q  $HM$)���      �       �Q $HM$)���      �       q  $HM$)���             �Q $HM$)��      +       q  $HM$)��+      |         $HM$)��|      �       �Q $HM$)���      �       q  $HM$)���               $HM$)��      "       �Q $HM$)��"      1         $HM$)��1      �       �Q $HM$)���      �         $HM$)���      �       �Q $HM$)��                                           a      �       q  $@N$)���      �       �Q $@N$)���      �       q  $@N$)���             �Q $@N$)��      +       q  $@N$)��+      |         $@N$)��|      �       �Q $@N$)���      �       q  $@N$)���               $@N$)��      "       �Q $@N$)��"      1         $@N$)��1      �       �Q $@N$)���      �         $@N$)���      �       �Q $@N$)��                  �      G       U                       >      �       0�;      z       0�z      �       P�      �       V�      �       0�                        �      �       0��      C       ]C      H       }�H      c       ]                   �             0�      )       P                        B      H       PH      n       s�n      �       ��~;      �       ��~                      Z      `       P`      j       ��}j      �       ��}��-3�-� �;      �       ��}��-3�-� �                      j      n       Pn      �       ��~;      [       ��~                   j      �       ��;      �       ��                   �      �       Y�      L       ��}                 �      ;       ��                    �      '       U'      /       �U�                      �      *       T*      .       u�~�.      /       �T�                    �      .       Q.      /       �Q�                      �       �        U�       �        P�       �        �U�                    �       �        T�       �        �T�                    �       �        Q�       �        �Q�                              1        U1       y        Qy       �        �U�                      (       w        p��w       y        q#��y              
 �U##��                      �       �        U�       �        T�       �        �U�                   �       �        u �       �        U                      �      �       U�      �       V�      �       �U�                      �      �       T�      �       S�      �       �T�                   �      �       0��      �       P                                     c       Uc      +       �U�+      2       U2      3       �U�3      >       U>      �       �U��      �       U                                        T      +       �T�+      N       TN      �       �T��      �       T                                             t      #       �T#+      2       Q2      3       t3      >       Q>      N       tN      �       �T#�      �       t                                       t       #       �T+      N       t N      �       �T�      �       t                           0      �       U�      �       _�      �       P�      �       ^�      �       �U�                  H      �       ^                          O      l       Pl      �       u� �      �       � �      �       p� �      �       ���~                  U      �       X                         U      {       U�{      }       Q}      �       T�      �       Q�      �      ! w #�;�4�4��������@�4%�;� 4%�                       �      �       ^�             _             ]      �       ���~                         A       VA      Q       v�Q      �       V                         U      �       0��      (       \(      /       _/      o       1�o      �       _�      �       1�                          /      9       S9      ;       s 1&�;      D       SD      ]       } | 1&�{      �       S�      �       S                      /      M       P�      �       P�      �       P                 �      �       ^                  �      �       \                    �      �       S      �       S                     �      �       ~�       $       T)      I       T                     �      �       0��      J       _�      �       _                     �      �        s���      �       R�      �       R                          �      �       U�      �       w �      �       �`�             w       !       �`                    �      �       T�      !       �l                          �      �       P�      �       S�             P              S       !       P                                �       -       U-      .       �U�.      G       UG      L       y�~�L      X       SX      Y       �U�Y      �       U�             �U�                            �       -       T-      .       �T�.      E       TE      Y       �T�Y      �       T�             �T�                              �       -       Q-      .       �Q�.      @       Q@      L       PL      Y       �Q�Y      �       Q�             �Q�                                �       �        R�       �        Y�       3       PY      }       Y}      �       P�      �       P�      �       P�             P                            �       -       X-      .       �X�.      L       XL      Y       �X�Y             X             �X�                          -       R.      =       R                                  �      �       T�      �       t��      �       U�      �       u��      �       U�      �       P�      �       U�      �       P�      �       U�      �       T�             U                       �      �       P�      �       P�      �       P�             P                    �      �       U�      �       �U�                    �      �       T�      �       �T�                    �      �       Q�      �       �Q�                      �      �       R�      �       P�      �       �R�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                      �      �       Q�      �       P�      �       �Q�                    0      A       UA      Y       �U�                      0      >       T>      Q       PQ      Y       �T�                    `      q       Uq      �       �U�                        `      �       T�      �       U�      �       \�      �       �T�                      y      �       V�      �       |��      �       �T#�                      }      �       S�      �       |��      �       �T#�                        p      �       U�      
       ^
      �
       �U��
      +       ^                    p      �       T�      +       ��                                  p      �       Q�      s	       \s	      
       ��
      G
       \G
      �
       �Q��
      �
       \�
      �
       ���
      �       ���      +       \                          �      �       R�      g	       [6
      G
       ��q ��
      �
       [�      �       ��q ��      �       [�      �       [                          �      k	       Z6
      G
       | p ��
      �
       Z�      �       | p ��      �       Z�      �       Z                                �      �	       S�	      �	       Q�	      
       S6
      Y
       S�
             S             
 �      [       Sg      l       Ul      �       S�      �       s�~��      �       0��      +       S                                        �      �	       X�	      �	       V�	      �	       
 ��	      
       V6
      `
       X�
      �
       X�
      �
       0��
             V             U      B       Vg      l       0�l      �       V�      �       Q�      �       X�      �       X�      	       x �      +       
 �                      �	      �	       QG
      `
      	 ������
             0�Y      l       U~      �       
 �                        �	      �	       0�G
      `
       | ���
      �
       
 ��
             UY      l       
 ��      �       Q�      +       0�                                �      {	       V{	      
       \6
      G
       V�
      �
       V�
      �
       \�
             |�      �       \�      �       |��      �       \�      +       V                                            �      �	       T�	      �	       ]�	      �	       }��	      
       ]
      G
       T�
      �
       T�
      �
       \�
      �
       |��
      �
       \�
      =       ]=      g       }�g      �       ]�      �       T�      �       ]�      �       T�             ]             }�      +       ]                             �      �       X�      �       ��8&��      
       ��6
      G
       ZG
      `
       ���
      �       ���      �       Z�      +       ��                                     �      �       Q�      �	       U�	      
       ��
      G
       UG
      �
       ���
      �
       U�
      �       ���      �       U�      �       ���      �       U�      +       ��                        (	      �	       _�	      
       _�
      �
       _�
      .       _.      l       Ql      ~       _~      �       U                    B	      
       ���
      �       ��                    c	      
       ���
      �       ��                            �             U      6       S6      7       �U�7      P       SP      Q       �U�Q      o       S                        �             T      Q       �T�Q      d       Td      o       �h                        �             Q      Q       �Q�Q      d       Qd      o       �l                          �       U�      �       �U�                      #      2       Q2      6       p�6      �       Q�      �       Q                      &      g       Pg      }       T}      �       P                            l       Rl      }       u� }      �       R                      �      �       U�      D       ]D      t       Ut      �       �U�                               �       W�      }       S}      �       sP��      �       S�      ?       sP�?      D       SD      t       W                   �      �       S�      ?       sP�                 /      ?       P                          �      �       U�      \       V\      _       �U�_             V      �       U                                �      �       W�      �       S�      �       P�      ?       S?      H       PH      I       s �_      n       Sn      s       s �      �       W�      �       ��{�                     `      c       p t 3${ "�c      g       w t 3${ "��      �       P                 `      t       x q 3$y "�                            �      �       1��      �       \�      I       \I      M       |�M      ^       \_      s       \s      w       |�w             \                          �      �       X�      �       x 1&��      �       X_      r       Xr      w      	 | | 1&�w            	 ||  1&�                �      ?       S                   �             P      (       P                      �      �       T�             U      "       Q"      %       R                    �      �       U�      #       �U�                    �      �       T�             S      #       �T�                    �      �       Q�      #       �Q�                    �      �       R�             V      #       �R�                              �U�                              �Q�                              V                              S                              0�                          �/      0       U0      00       �@00      �0       �U��0      �0       U�0      �0       �U�                          �/      0       T0      00       ��00      �0       �T��0      �0       T�0      �0       �T�                                    �/      00       Q00      o0       So0      q0       �Q�q0      �0       S�0      �0       �Q��0      �0       S�0      �0       �Q��0      �0       S�0      �0       Q�0      �0       S                        �/      00       R00      �0       �R��0      �0       R�0      �0       �R�                        �/      00       X00      �0       �X��0      �0       X�0      �0       �X�                                  10      A0       PD0      P0       PP0      p0       Vq0      }0       P�0      �0       V�0      �0       P�0      �0       V�0      �0       P�0      �0       V                          �,      �,       U�,      ;.       S;.      E.       �U�E.      N.       UN.      �/       S                                              �,      �,       T�,      .       V.      E.       �T�E.      N.       TN.      n.       Vn.      r.       Ur.      �.       V�.      �.       �T��.      �.       V�.      �.       U�.      �.       V�.      /       �T�/      /       V/      �/       �T��/      �/       V                  �.      �.       0�	/      /       0�                    �,      >.       \N.      �/       \                             �,      C-       0�C-      Y-       PY-      6.       ]E.      N.       0�N.      �.       ]�.      �.       0��.      ~/       ]~/      �/       0��/      �/       ]                       	.      .       0�s.      �.       _�.      �.       0��.      /       _/      �/       _                         �.      �.       0��.      �.       P�.      �.       V�.      	/       V	/      /       0�/      �/       V                        �.      �.       P�.      /       ^/      "/       P"/      �/       ^                 /      y/       ]                     /      /       }�/      "/       U"/      y/       }�                        �-      	.       VN.      n.       Vn.      r.       Ur.      s.       V�.      �.       U�.      �.       V                         �-      	.       ^N.      n.       ^n.      r.       Tr.      s.       ^�.      �.       T�.      �.       ^                      �-      	.       0�N.      j.       0�j.      r.       Pr.      s.       _�.      �.       P�.      �.       0�                  K-      �-       V�.      �.       V/      /       V                  K-      }-       S}-      �-       V�.      �.       V/      /       V                    K-      Y-       PY-      �-       ]�.      �.       ]/      /       ]                        K-      Y-       p�Y-      �-       }��-      �-       U�-      �-       }��.      �.       }�/      /       }�                     K-      �-       0��-      �-       P�-      �-       0��.      �.       P/      /       3�                    �,      �,       U�,      �,       �U�                    �,      �,       T�,      �,       �T�                    �,      �,       Q�,      �,       �Q�                    �,      �,       R�,      �,       �R�                   �,      �,       u�,      �,       U                          p	      �	       U�	      �	       V�	      �	       �U��	      
       V
      
       �U�                  {	      �	       S�	      �	       0�                    	      �	       \�	      
       \                 �	      �	       S                     �	      �	       s��	      �	       U�	      �	       s�                                    P)      �)       U�)      P*       SP*      S*       |�~�S*      U*       }h�U*      V*       �U�V*      �*       S�*      �*       |�~��*      �*       }h��*      �*       �U��*      �*       S                          ])      U*       ]U*      V*       �U#�V*      �*       ]�*      �*       �U#��*      �*       ]                       ])      F*       0�F*      V*       U�V*      �*       0��*      �*       U��*      �*       0�                    �)      �)       P�*      �*       P                        �)      �)       S�)      5*       SV*      �*       S�*      �*       S�*      �*       S                        �)      �)       s��)      5*       s�V*      �*       s��*      �*       s��*      �*       s�                         �)      �)       V�)      5*       VV*      �*       V�*      �*       V�*      �*       V                               �)      �)       P�)      �)       P�)      *       vt �*      *       vv�V*      g*       vv��*      �*       P�*      �*       vt ��*      �*       vv�                        �
      �
       U�
      �
       S�
      �
       �U��
      �       S                  �      �       P                  r      �       t 
���                                 p ��             q ��                    =      A       p ��A      R       q ��                    0
      4
       U4
      5
       �U�                    0
      4
       T4
      5
       �T�                   0
      4
       T4
      5
       �T�                   0
      4
       U4
      5
       �U�                    `
      u
       Uu
      {
       �U�                    `
      l
       Tl
      {
       �T�                    `
      q
       Qq
      {
       �Q�                  `
      q
       Qq
      v
       �Q�                  `
      l
       Tl
      v
       �T�                  `
      u
       Uu
      v
       �U�                    `
      l
       q ����t �����l
      u
       Tu
      v
       �Q�����T�����                  `
      v
       0�v
      v
       P                    0      :       U:      b	       �U�                            0      ^       T^      �       Z�      \       zp�\      �       Z	      %	       Z%	      C	       PR	      b	       T                              0      v       Qv      �       U�      �       ���      	       Q	      	       U	      R	       ��R	      b	       Q                                                        6      �       _�      �       P�      �       ^�      �       ]�      �       \�      �       V�             S             T             ��      0       R0      8       [8      >       Y>      D       XD      J       UJ      P       TP      V       RV      \       Q\      �       _	      a	       _a	      b	       �U
���                                   J      ^       P^      �       ���      �       ��p "��      �       ��p "~ "��      �       ��p "} "~ "��      �       zp��} "��"~ " "��      �       zp��| "~ " "��"} "�\      g       ���      �       ���      �       U	      	       ��%	      R	       RR	      X	       PX	      b	       ��                        p      �       P�      �       p��      �       �D�#�	      	       P                                                                        �      C       UC      
       S
             �U�      )       S)      �       �U��      o       So      y       Uy      �       S�      �       �U��      %       S%      r       �U�r      �       S�      �       �U��      �       S�      �       �U��      �       S�      �       �U��      �       S�              �U�               S       `        �U�`       f        Uf       \"       �U�\"      f"       Uf"      �#       �U��#      �#       S�#      �$       �U��$      �$       S�$      B)       �U�                        �      '       T#      )       	��`       f        T\"      f"       T                                            '      H       	��H      P       Py      �       P�      �       P�      �       P      )       	���      �       	���      �       	���      �       P@      �       	���      �       P�      �       P�      %       	��%      0       P�      �       P�      �       	��-      C       Pi      t       P�      �       	���#      �#       	��                                
       p ��
      @       x ��r      |       x ��|      �       s 1����$      �$       s 1���                                                                                                                     �      �       Q�      �       Z�      �       Q             P      g       0�g      z       Zz      �       0��      �       Z�      	       0�	      )       0�r      w       Qw      z       Z~      �       	���             Z             0�      8       0��      �       Z�      �       0��      �       Z�      X       ��X      [       Z_      �       1��      �       ���             Z.      E       ZE      Q       0�Q      q       0��      �       Z�      -       Z.      b       Pb      �       0��      �       Z�      �       Q�             P�      �       0�'       *        ZC       `        	��f       s        Zs       �        0��       �        Z�       �        Q�       !       Z!      �!       ���"      �"       Z�"      �"       0��"      �"       0�Q#      f#       0��#      $       Z$      $       Z�$      �$       Z�$      �$       	���$      �$       P�$      %       Z%      8%       ��8%      Y%       	���%      �%       Z�%      �%       P�%      &       Z&      2&       ���&      �&       P�&      *'       	��@'      E'       	��w'      �'       	���'      �'       P�'      �'       	���'      �(       ��)      )       	��                                        �      �       S�      �       �U��      �       S�      �       �U��      �       �U��      -       �U��              �U�       `        �U�f       \"       �U�f"      �#       �U��#      �$       �U��$      B)       �U�                    �      �       Z�      �       Z                                                               �      �        7��      �       R�      �       Q�      �       P�      �       |�      S       TS      �       X)      X       ��#      #       0�      *        7�|      �       P�      �       |g      �       R�      �       ��~�       !       |�!      �!       Ps"      �"       X�"      0#       |$      -$       X-$      i$        7��$      �$        7�"%      Y%       	��$&      2&       	��*'      1'       |1'      E'       zE'      R'       |R'      X'       ��~#�'      �'       	���(      )        7�                                                                    �      �       _:      O       _d      q       _z      H       _H      w       0�w      �       _�      �       _�      �       _�             _      �       _�             0��             _�      �       _'       `        _f       �        _�       �        _�       �!       _s"      �"       _�"      �"       P�"      Q#       _$      $       0�$      i$       _�$      �$       _�$      Y%       _�%      �%       _&      2&       _�&      �'       _�'      �(       _�(      )       _                                                                                                            �      �       ]?      O       ]d      q       ]z      �       ]�      �       }x��      �       ]�      �       }��      �       ]�             R             rx�      )       R)      C       ]H      w       0�w      �       ]�             ]      +       R+      .       rx�.      8       R8      k       ]s      �       ]�      �       R�      �       rx��      �       R�      �       r��      I       RI      �       ]�             ]      E       ]E      c       Rc      f       rx�f      q       Rq      �       ]�      �       }��      �       ]�             0��             ]�      �       R'       `        ]f       �        ]�       �        R�       �!       ]s"      �"       ]�"      �"       R�"      �"       rx��"      �"       R�"      �"       ]�"      Q#       ]$      $       0�$      m$       ]m$      �$       }��$      �$       ]�$      �$       }��$      %       R%      Y%       ]�%      �%       ]&      2&       ]�&      �'       ]�'      �(       ]�(      )       ]                                                                                           �      �       V1      �       V�      �       Y�             V             v�      �       V�             V      %       v�%      �       V�             Q      �       V�             V      1       Y1      U       VU      ]       v�]             V�              V'       `        Vf       �        V�       �        Q�       "       Vs"      �"       V�"      �"       v��"      f#       V�#      -$       V-$      L$       YL$      �$       ��~�$      �$       V�$      �$       Y�$      �$       V�$      %       Q%      Y%       V�%      �%       V�%      �%       V�%      2&       V�&      '       V*'      �'       V�'      �(       V�(      )       ��~)      &)       V                                                    �      �       ^5      �       ^�      �       ^�             ^             ^�              ^'       `        ^f       �        ^�       "       ^s"      f#       ^�#      �$       ^�$      Y%       ^�%      �%       ^�%      �%       ^�%      2&       ^�&      �'       ^�'      �(       ^�(      &)       ^                                                                    �      �       [?      �       [�      �       [�      �       [X      �       [      �       [�      �       ��~�      -       [3      �       [�      �       [�             ['       Z        [s       �        [Q#      f#       [�#      �#       [�#      $       P$      $       [-$      L$       [L$      �$       ��~�$      �$       [�$      �$       [�%      �%       [�%      �%       [�%      �%       |� �%      �%       [�%      &       P*'      E'       [�'      �'       |� �'      �'       [�(      )       ��~                               K      O       x�L      P       x��      �       x r ��      �       Xs       �       	 |� �{ ��#      �#       q��$      �$       q { ��%      &       { p �                                                                                       �      �       Z�             	���             Z             0�H      q       Zr      �       P�      �       0��      �       Z�      �       0��             0�      0       Z0      9       0�9      Z       0��      �       Z�      �       0��      �       0�      u       Zv      �       P�      �       0��      �       Z�      -       1�-      b       Zc      �       P�      �       Z�      �       0��      �       0�%      -       Z       '        0�f       s        Z�       �        Z"      &"       0�f"      s"       Pf#      p#       Zp#      �#       P�#      �#       Z�#      �#       	��Y%      �%       P�%      �%       P�%      �%       Z2&      a&       P�&      �&       Z�'      �'       P�(      �(       	���(      �(       P=)      B)       	��                   �             Sf       s        S                   �             \f       s        \                                             H       |�             |!      �       |�             Q�      �       |�      �       Q�             |�%      �%       |g&      p&       |�&      �&       |�&      �&       u�(      �(       u&)      /)       |/)      B)       p                                   H       Qp      �       Q�      �       Q�%      �%       Qg&      �&       Q�&      �&       Q�(      �(       Q&)      B)       Q                                          -      8       P8      C       RC      H       q ���      �       p ���      �       q ����      �       P�      �       R�%      �%       p ���%      �%       |���g&      s&       Ps&      �&       R�&      �&       P�(      �(       P&)      ))       p ��))      B)       q ���                                                     �             _�             _      �       _
             _       -       _       '        _f       s        _�       �        _"      \"       _f"      s"       _f#      �#       _�#      �#       _Y%      �%       _�%      �%       _�%      �%       _2&      �&       _�&      �&       _�'      �'       _�(      �(       _&)      B)       _                                                               �             ]�             ]      %       ](             ]             }x�      H       ]H      R       }x�R      y       ]      �       ]�      �       }x��      �       ]
      �       ]�      �       }x��      �       ]       -       ]       '        ]f       s        ]�       �        ]"      \"       ]f"      s"       ]f#      �#       ]�#      �#       ]Y%      �%       ]�%      �%       ]�%      �%       ]2&      �&       ]�&      �&       ]�'      �'       ]�(      �(       ]&)      B)       ]                                                                   �             V�             V      �       V�             v�      =       V=      L       v�L      �       V�      �       v��      �       V�      �       v��      -       V       '        Vf       s        V�       �        V"      \"       Vf"      s"       Vf#      �#       V�#      �#       VY%      �%       V�%      �%       V�%      �%       V2&      �&       V�&      �&       V�'      �'       V�(      �(       V&)      B)       V                                                   �             ^�             ^      -       ^       '        ^f       s        ^�       �        ^"      \"       ^f"      s"       ^f#      �#       ^�#      �#       ^Y%      �%       ^�%      �%       ^�%      �%       ^2&      �&       ^�&      �&       ^�'      �'       ^�(      �(       ^&)      B)       ^                                                                                 �             [�             [      H       [H      q       R�      �       R�      u       [�      �       U�      '       [-      b       [h      -       [       '        [f       s        [�       �        [�       �        U"      V"       [f"      s"       Uf#      t#       Ut#      }#       x� }#      �#       U�#      �#       [Y%      b%       Ub%      �%       [�%      �%       [�%      �%       x� �%      �%       [2&      ]&       U]&      a&       u� g&      �&       [�&      �&       [�&      �&       R�&      �&       P�'      �'       R�'      �'       U�'      �'       R�(      �(       [�(      �(       U�(      �(       R&)      B)       [                                          �      �       t��      �       t��       �        p�j"      s"       r u �f#      p#       { u ��#      �#       q��#      �#       TY%      b%       r u ��'      �'       q��'      �'       T�'      �'       u r ��(      �(       r u ��(      �(      	 x� �u �                                        �       S�      �       s��      �       S       '        S�       �        Sf"      s"       Sf#      �#       SY%      b%       S�%      �%       S2&      I&       S                                                                             �      �       \�             X             |             \      �       \-      6       \6      9       P9      b       Xb      �       ��~�      -       \       '        \f       s        X�       �        \"       "       \f"      s"       \f#      �#       \�#      �#       \Y%      b%       \b%      �%       ��~�%      �%       \�%      �%       \2&      F&       \g&      �&       \�&      �&       \�&      �&       U�&      �&       \�'      �'       \�(      �(       U�(      �(       \&)      /)       \/)      B)       P                         O       Ss       �        S                       #       |                              K      a       Pa      h      	 r 3$| "�h      s         t 2$�lG     "�����3$| "�s"      "       P"      �"      	 r 3$| "��"      �"      (  |�����2$�lG     "�����3$| "�$      -$       P                          �"      �"       P�"      0#       |0#      8#       P<#      Q#       PE'      R'       |R'      X'       ��~#                 �"      �"       ��~�"      #        x ����2$�lG     "�p ��~�"�                         S      �       Us"      .#       U.#      0#       Q$      -$       UE'      N'       U                   ~      )       S%      "%       S&      $&       S                     ~      �       X�      )       ��%      "%       ��&      $&       ��                           ~      �       Y�      �       ���      )       | �%      %       | �%      "%       ��~# �&      &       | �&      $&       ��~# �                           ~      �       R�      �       ��~�      )       |�%      %       |�%      "%       ��~#�&      &       |�&      $&       ��~#�                        ~      �       P�      '       ��~%      %       ��~&      &       ��~                     �      (       P(      )       ��%       %       P %      "%       	��&      !&       P!&      $&       	��                     �      �       P�      )       ��~%      "%       ��~&      $&       ��~                 �      �       P�&      '       0�                    �      #       S!      �!       S�'      �(       S                      �      #       ��~!      �!       ��~�'      @(       ��~b(      �(       ��~                        �      �       ����      �       Y�      #       ���!      �!       ����'      �(       ���                        �      #       ���!      ^!       ���^!      b!       Yb!      �!       ����'      �(       ���                        �      �       ����      �       P�      #       ���!      �!       ����'      �(       ���                        �      #       ���!      O!       ���O!      b!       Pb!      �!       ����'      �(       ���                    �      #       ��!      �!       ���'      �(       ��                     �      !       ���#�!      �!       ���#��'      �(       ���#�                 !      !       ��~                                    �      �       P�      "       Pc!      �!       P�!      �!       	���!      �!       P�!      �!       ��~�'      1(       P1(      <(       	��N(      O(       PO(      b(       ��~b(      q(       Pq(      x(       	��x(      �(       P                       �      #       ��~)!      O!       PO!      �!       ��~�'      �(       ��~                 T      �       S                  T      Y       ��~                   T      [       R[      �       ��                    T      [       X[      �       ��~                    T      [       Y[      �       ��~                 \      �       P                  E$      �$       9��(      )       9�                	  E$      �$       5��(      )       5�                
  E$      �$      
 �mG     ��(      )      
 �mG     �                  E$      �$      
 �lG     ��(      )      
 �lG     �                   E$      �$       S�(      )       S                 E$      �$      
 �lG     ��(      �(      
 �lG     �                 E$      �$      
 �mG     ��(      �(      
 �mG     �                 E$      �$       5��(      �(       5�                 E$      �$       9��(      �(       9�                   M$      �$       P�(      �(       P                   E$      �$       S�(      )       S                E$      E$       ��                  E$      E$       ��                  E$      E$       ��                  E$      E$       ��                          �      �       U�      #       S#      %       �U�%      .       U                   �      �       U�             S                 �             V                        P      �       U�      �       T�      �       �U��      �       U                      �      �       U�      N       SN      P       �U�                      �      �       T�      O       VO      P       �T�                    �      �       Q�      P       �Q�                             V                              s                        �      	       U	      B       SB      L       �U�L      �       S                          �             T      C       VC      L       �T�L      U       TU      �       V                          �      �       Q�      G       ]G      L       PL      U       QU      �       ]                         �             P      ,       ^L      U       Pk      �       Q�      �       0�                      �      $       \$      (       UL      U       \                               �      ,       _,      I       ^I      L       �U#PL      U       _U      `       ^`      �       R�      �       w �      �       R                                  �       U�             �U�      )       U)      �       �U��      �       U                                      �        T�       L       XL      ]       T]      J       XJ      �       P      )       T�      �       X                            t        Qt       �       ��}                            �        R�       �       ��}                            |        X|       �       ��}                            �        Y�       �       ��}                              �       �      )       ��      �       �                            �      �       U�      �       ��}4�      �       ��}�1�             ��}�1�)      ]       ��}�1�]      v       r�                            A      V       PV      [      	 p ��}���      �      	 p ��}���      �       | r �$��}���      �       Pt      �       U�      �       | ��|�{ �$�                                L       0�d      j       ��}j      �       T�      �       ��}�      �       T�      �       ��}                                   R      �       	���      �       Q�      )       Z)      =       Q=      �       Z      �       Q�      �       q��      �       T�      �       Q)      v       Q                                           h       �        T�       �        ?��              T             t�      /       T7      L       	��]      �       T�      �       ��}      &       P&      *       p�J      �       0��      �       S             S)      v       S�      �       T�      �       t��      �       T                                                   �       �        1��       �        P�       �        p��       �        r�)      L       0�L      Y       PY      ]       R�      �       0��             Q      v       Q�              T              R=      o       Uo      �       T�      �       T�      �       t��      �       T}      �       R�      �      
 1��|�1$��      �       R�      �       0�                        �      �       ��|             ��|)      b       ��|f      v       U                           �       �        P�       �        q �              Y      L       0�L      ]       q ]      �       Y�      �       Y                 �      �       1{ $1��      �       1r $1�                 		

                                       ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               ��}�               W               ��}�               ��}�               ��}�               ��~�               ��~�               ��~�               ��~�       h        ��~�h       �        U�       �        P7      L       ��}��      �       ��}��      �       p 2$� "
(��      �       p 2$� "
,��             p 2$� "
(�             p 2$u "�      *      
 p 2$u "#�*      4      
 p2$u "#�R      �       �      >       �a             �             PL      ]       �#�]      �       ��      �       ��}�                         R      �       0��      P       ^      �       ^             ^)      v       ^                                                       �       �0���      �       ���}��      �       �Y����}��             T�Y����}�             T�Y��_�      �       ���}�      #       ���}�#      D       �X����}�D      a       �X��a      �       T�X����}��      �       T�X��V��            
 �X��V�      )       �0��)      L       �X��L      X       T�X��X      ]       T�X��U�]      v       ���}��      �       �0��                              R      �       [�      )       X)      =       [=      �       X      �       [�      �       R�      �       R�             [)      �       [                                    7      L       ��~��      �       ��~��      �       p 2$� "���      �       p 2$� "���             p 2$� "��V      [       ��}4��      �       ��}4��      �       ��}�      �       _�      �       |��      �       _�      �       ��~�                                               p z �      L       S�      �       p q 2$� "
0���      �       P�      �       p 1$��      �       P�      �       p q 2$� "
0���      �       S�      �       p q 2$� "
0���      �       S                            R      �       0��      �       P)      7       P=      =      	 ��}�x �=      [      # ��}�x ������}�����-( �[      o       1u $��      �      # ��}�x ������}�����-( ��      �       1t $�             P)      v       P                     
      $
       U$
      %
       �U�                     
      $
       T$
      %
       �T�                    @
      U
       UU
      [
       �U�                    @
      L
       TL
      [
       �T�                    @
      Q
       QQ
      [
       �Q�                     @
      L
       q ����t �����L
      U
       TU
      [
       �Q�����T�����                   @
      V
       0�V
      [
       P                                   /       U/      %       S%      -       �U�-      �       S�      �       U�      �       S                                     D       TD      �       V-      >       V>      l       T�      �       V�      �       T�      �       V                   �             ]l      v       ]�      �       ]                   �             ^l      v       ^�      �       ^                   �             Sl      v       S�      �       S                     �      �       P�             Vl      v       V�      �       V                                �*      +       U+      f+       Sf+      n+       �U�n+      �+       S�+      �+       �U��+      �+       S�+      �+       �U��+      �,       S                                  �*      +       T+      +       V+      �+       �T��+      �+       T�+      �+       V�+      �+       �T��+      �+       V�+      O,       �T�O,      �,       V                              �*      +       Q+      )+       ])+      �+       �Q��+      �+       Q�+      �+       ]�+      �+       �Q��+      �,       ]                              �*      +       R+      )+       \)+      �+       �R��+      �+       R�+      �+       \�+      �+       �R��+      �,       \                     )+      e+       \e+      n+       0�n+      �+       \�+      �+       \                          )+      I+       ^T+      m+       ^m+      n+       Pn+      |+       ^�+      �+       ^�+      �+       P                  �+      �+       P                    A+      F+       VF+      i+       \n+      �+       V                  �+      �+       SO,      �,       S                 �+      �+       s                     �+      �+       PO,      X,       P                    O,      T,       s�T,      X,       UX,      �,       s�                       �+      ,       V,      ,       0�,      1,       V1,      4,       v q �4,      O,       V                  �+      O,       S                    �+      B,       0�B,      M,       P                    �+      ,       Q,      ,       V,      A,       Q                        �             U      *       S*      4       �U�4      �	       S                          �             T      4       �T�4      �       _�      �       T�      �	       _                          �             Q      4       �Q�4      �       \�      �       Q�      �	       \                                 �             0�      +       V+      4       P4      �       V�      �       0��      �       1��      �       0��      �	       V�	      �	       1��	      �	       V                                         �      1       ^1      4       �U#L4      X       ^_      _       0�_      ~       ^~      �       P�      �       ^�      �       Q�      W	       ^W	      k	       Qk	      	       ��	      �	       ^�	      �	       ���	      �	       ^�	      �	       P�	      �	       ^                                   �      /       ]/      4       �U#H4      [       ]_      _       0�_      �       ]�      �       w �      ~       ]~      �       P�      R	       ]R	      W	       QW	      �	       ]�	      �	       P�	      �	       ]                                        �      �       P�      &       w &      )       P)      4       ��4      g       w g      �       0��      �       w �      �       P�             
 ��      	       w 	      %	       P	      �	       w �	      �	       0��	      �	       P                           4      _       Pg      k       P�      �       P�             P	      %	       P�	      �	       P                                       4      _       P�      �       P�      �       Q�             P      #       QM      |       Q|      �       ��	      %	       PB	      R	       ]R	      k	       Qk	      	       ���	      �	       ���	      �	       P                   �      	       S	      �	       S                    �      �       [�      	       ��	      �	       [                    �      �       [�      	       ��	      �	       [                    �      �       U	      �	       U                      �      ,       U,      d       Sd      w       �U�                  �      v       V                 �      $       U                                  U      �       Q                 p      �       Q                                 h       Uh      �       S�      �       �U��      �       U�      �       �U�                    4      l       Z�      �       Z                   4      X       Q�      �       Q�      �       0�                       4      4       Q4      E       VE      X       @<$�[      �       V�      �       V�      �      
 q 1%q "#�                        p       �        U�       �       S�      �       �U��      �       S                          �       J       VR      e       Re      s       vx�s      �       R�      �       V�      �       9��      �       V                            �       �        u�       �        U�       �        ss      �       T�      �       s�      �       U�      �       s                    M      M       QM      V       q�V      �       X                  O      �       P                   �       >       S�      �       S                    �       >       P�      �       P                          �      �       U�      M       SM      U       �U�U      ^       U^      �       S                          �      �       T�      N       VN      U       �T�U      ^       T^      �       V                    �      P       \^      �       \                           �             0�             P      H       ]U      ^       0�^      �       ]�      �       0��      �       ]                 ^      �       V�      �       V                 ^      �       S�      �       S                 ^      �       ]�      �       ]                  o      �       ^�      �       ^                    �      �       P�      �       P�      �       ��                    �	      
       U
      �       �U�                        �	      
       T
      1
       V1
      �
       �T��
             V      �       �T�                        �	      
       Q
      �
       ]�
      �
       �Q��
      �       ]                            �	      
       R
      R
       \R
      �
       �R��
      �       \�      �       �R��      �       \                    �	      �
       S�
      �       S                     �	      
       R
      |
       \|
      |
       0��
      �       \�      �       \                       �	      
       Q
      �
       ]�
      �
       �Q��
      �       ]                       �	      
       T
      1
       V1
      �
       �T��
             V      �       �T�                   �	      �
       S�
      �       S                          �	      R
       0�R
      i
       _n
      |
       _�
      �       0��      �       _�      �       _�      �       0�                 �
      �
       0�                   U
      c
       Vc
      |
       \�      �       V                 �      �       S                     �      �       s��      �       U�      �       s�                  �      �       P                 �      �       0�                �
      �
       S                 �
      �
       s                   �
      �
       P                 �
      �
       s�                              0       V0      3       v q �3      r       Vr      y       v�`�y      �       V�      �       V�      �       0�                          �       S�      �       S                         �       0��      �       0�                        I       Q                       I             
 �      �       
 ��      �       ^�      �       ^                      _             P�      �       P�      �       P                      �      �       U�      �       V�      �       �U�                  �      �       S�      �       0�                   �      �       u8�      �       \                 �      �       S                                              U               S               �U�       G        SG       H        �U�H       b        Sb       c        �U�                             1        P2       F        PH       ]        P                                                        �n      �n       U�n      �s       ^�s      �t       ���~�t      Hv       ��~8�Hv      cv       ^cv      �|       ���~�|      �|       ��~8��|      ��       ���~��      Ǆ       ^Ǆ      I�       ���~I�      i�       ^i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      {�       ���~{�      ��       ��~8���      �       ���~�      �       ��~8��      #�       ���~                                  �n      �n       T�n      �s       S�s      Hv       �T�Hv      cv       Scv      ��       �T���      Ǆ       SǄ      I�       �T�I�      i�       Si�      #�       �T�                            �n      �n       Q�n      %�       �з~%�      1�       qз~1�      s�       �з~s�      w�       qз~w�      #�       �з~                            �n      o       Ro      %�       �ط~%�      1�       qط~1�      s�       �ط~s�      w�       qط~w�      #�       �ط~                    �n      �p       X�p      #�       �X�                  �n      �p       Y                  �n      �p       �                           �n      %�       �%�      1�       q1�      s�       �s�      w�       qw�      #�       �                                 �n      �t       0��t      �t       ]Hv      ||       0�||      �|       P�|      �|       0��|      �|       ]�|      ��       0���      ��       P��      #�       0�                                    �n      o       Po      �p       ~��p      �t       ���~Hv      �|       ���~�|      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      p�       ���~�      #�       ���~                                  Ho      �o       T�o      �r       _�r      Hv       ��~Hv      cv       _cv      %�       ��~%�      1�       q�~1�      s�       ��~s�      w�       q�~w�      #�       ��~                       Ho      �s       \Hv      cv       \��      Ǆ       \I�      i�       \                           Ho      �p       ~8�p      %�       �̷~%�      1�       q̷~1�      s�       �̷~s�      w�       q̷~w�      #�       �̷~                       Ho      �s       v @$�Hv      cv       v @$���      Ǆ       v @$�I�      i�       v @$�                	                                             Ho      �s       0��s      �t       ���~Hv      cv       0�cv      �y       ���~z      �|       ���~�|      ��       ���~��      Ǆ       0�Ǆ      I�       ���~I�      i�       0�i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      S�       ���~S�      S�       PS�      O�       ���~O�      ��       0���      ֐       1�֐      Ǔ       0�Ǔ      �       Y�      ӕ       0�ӕ      �       2��      ��       ���~��      �       0��      �       ���~�      >�       0�>�      #�       ���~                
                                   Ho      �s       0��s      �t       ���~Hv      cv       0�cv      �|       ���~�|      ��       ���~��      Ǆ       0�Ǆ      I�       ���~I�      i�       0�i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      O�       ���~O�      S�       PS�      �       ���~��      F�       ���~�      k�       ���~k�      r�       0�r�      #�       ���~                                           Ho      �s       0��s      �t       ���~Hv      cv       0�cv      �|       ���~�|      ,}       ���~,}      E~       1�E~      ��       ���~��      Ǆ       0�Ǆ      I�       ���~I�      i�       0�i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      #�       ���~                                                                Ho      �s       0��s      �t       ���~Hv      cv       0�cv      �y       ���~z      �|       ���~�|      �       ���~7�      ��       ���~��      Ǆ       0�Ǆ      I�       ���~I�      i�       0�i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      ω       ���~߉      g�       ���~t�      �       ���~#�      /�       P/�      O�       ���~O�      �       0��      '�       ���~��      ݘ       0�ݘ      �       P�      �       ���~�      �       0��      +�       ���~�      #�       ���~                       Ho      �r       ]�r      �r       ��~Hv      Vv       ]Vv      cv       ��~                                                                                                                                                                                                                     Ho      Ps       0�Ps      �t       _Hv      cv       0�cv      �|       _�|      �|       _�|      �|       U�|      l~       _l~      �~       U�~      �~       _�~      �~       U�~      �       _�      �       U�      �       _�      �       Q�      +�       _+�      A�       UA�      ہ       _ہ      �       U�      a�       _a�      t�       Ut�      Æ       _Æ      �       U�      �       _�      ?�       U?�      I�       _I�      i�       0�i�      ��       _��      ��       U��      w�       _w�      Ŋ       UŊ      ۊ       _ۊ      �       U�      #�       _#�      b�       Ub�      w�       _w�      ��       U��      H�       _H�      `�       U`�      �       _�      &�       U&�      C�       _C�      ��       U��      ؏       _؏      ��       U��      Y�       _Y�      ��       U��      ֐       _֐      ��       U��      ґ       _ґ      ��       U��       �       _ �      ǒ       Uǒ      ђ       _ђ      �       U�      2�       _2�      ?�       U?�      f�       _f�      ��       U��      �       _�      9�       U9�      �       _�      �       U�      0�       _0�      o�       Uo�      ��       _��             U      w�       _w�      ��       U��      ��       _��      ��       U��      �       _�      3�       U3�      ��       _��      ��       U��      ��       _��      ��       U��      �       _�      �       U�      �       _�      �       U�      4�       _4�      W�       UW�      �       _�      5�       U5�      ��       _��      ��       U��      �       _�      ��       U��      �       _�      $�       U$�      ,�       _,�      2�       U2�      T�       _T�      r�       Ur�      ��       _��      ��       U��      '�       _'�      /�       U/�      J�       _J�      W�       UW�      #�       _                            �r      Hv       ��~cv      %�       ��~%�      1�       q�~1�      s�       ��~s�      w�       q�~w�      #�       ��~                                                                                                  �s      �t       S�t      �t       S�t      �t       r �t      �t       Scv      �v       S�w      �w       S�x      �x       S�y      �y       Sz      "z       S�z      {       S|      3|       S�|      �|       S�|      5}       SE~      _~       S�~      �~       SJ      t       S�      �       SI�      n�       S��      р       S�      ��       S�      k�       Sk�      �       �ȷ~7�      u�       SǄ      !�       Sv�      ��       S��      �       Si�      ��       S��      ��       Pχ      ��       S��      ��       Sn�      p�       Sp�      u�       Pu�      ��       S߉      �       SO�      w�       S��      ��       S�      ,�       St�      �       S�      .�       S{�      ��       S��      ��       S                                               Ho      �s        -1��s      bt       ���~bt      gt      	 ���~�1�gt      �t       ���~Hv      cv        -1�cv      �|       ���~�|      ��       ���~��      Ǆ        -1�Ǆ      I�       ���~I�      i�        -1�i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      ��       ���~��      S�       ���~�      #�       ���~                                           Ho      bs       0�bs      �s       �й~�s      �s       R�s      �s       PHv      cv       0�A�      L�      	 �й~p "�L�      U�       PU�      �       ���~��      Ǆ       0�i�      q�      	 �й~p "�q�      ��       P!�      v�       ���~I�      i�       0���      χ       ���~��      Ӌ       ���~                                                     Ho      �s       	���s      �s       0��s      �t       ���~Hv      cv       	��cv      �|       ���~�|      �}       ���~�}      �}       S�}      �}       p��}      ~       PE~      ��       ���~��      Ǆ       	��Ǆ      '�       ���~'�      )�       P)�      i�       ���~v�      I�       ���~I�      i�       	��i�      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      "�       ���~�      #�       ���~                    �|      �|       P�|      �|       q�                          �|      �|       Pw�      |�       P|�      ��       S��      \�       �ȷ~w�      ��       �ȷ~                       w�      ��       ���~#`���      \�       ~� �\�      w�       ���~#`�w�      ��       ~� �                       w�      |�       P|�      ��       S��      \�       �ȷ~w�      ��       �ȷ~                               w�      Ŋ       UŊ      ۊ       _ۊ      �       U�      #�       _#�      b�       Ub�      i�       _w�      ��       U��      ��       _                            ��      ��       V��      �       Y�      �       T�      �       Z�      &�       TK�      \�       Y                  ��      ��       [                     ��      K�       0�K�      \�       1�w�      ��       0�                   ي      �       1�#�      &�       1�                    ��      i�       ]w�      ��       ]                               ��      Ŋ       UŊ      ۊ       _ۊ      �       U�      #�       _#�      b�       Ub�      w�       _w�      ��       U��      ��       _                        Ɋ      �       S�      ��       s|���      \�       Sw�      ��       S                      ي      �       P�      �       x p "��      &�       X                  ��      �       P                 ��      �       s|                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                   &�      K�       [w�      ��       [                     &�      K�       Uw�      ��       U��      ��       _                     *�      \�       Uw�      ��       U��      ��       _                       �~      �~       0��~      �~       V�~             v~�             V                    �~      �~       P�~             S                 �~             _                        _~      l~       0�l~      �~       \�~      �~       |��~      �~       \                    \~      l~       Pl~      �~       V                  _~      �~       S                    l~      t~       P�~      �~       P                       L~      l~       _l~      �~       U�~      �~       _�~      �~       U                 8      J       _                        T�      k�       Pk�      �       ]u�      |�       P�      O�       ]                           T�      k�       0�k�      r�       Vr�      x�       vz�x�      |�       T|�      ��       vz���      �       Vu�      |�       0�                    ��      ��       P��      �       Z                    ��      ��       P��      �       [                  ��      ��       ^                  ��      �       X                    k�      r�       \��      �       \                    k�      r�       SЃ      �       S                     H�      �       _u�      |�       _�      O�       _                 J�      O�       _                      V�      x�       P��      Ȃ       P!�      3�       P                    |�      ��       P��      ��       Q                      
�      �       P�      1�       ���~� $ &#�1�      A�       P                 
�      Q�       ���~�                 Q�      Q�       P                  �      1�       ��                  �      1�       Q                    ��      �       ���~��      ʇ       ���~��      Ӌ       ���~                 ��      Ȃ       P                      ��      �       ���~��      ��       U��      ʇ       ���~��      Ӌ       ���~                        Ȃ      �       P��      ��       P��      ��       T��      ��       P                !�      _�       ���~                 !�      3�       P                !�      _�       ���~                    3�      K�       PK�      O�       R                      Ԏ      ؎       P؎      �       [�      ��       [                      �      �       P�      ��       Z؏      ��       Z                      �      �       P�      F�       Y�      ��       Y                         ]�       x �1)��      ��       x �1)�                    �      �      	 z p { ��      �      	 z p { �                   �      �       2��      ��       2�                   �      �       U�      ��       U                         ��      &�       U&�      /�       _/�      ��       U��      ��       _؏      ��       U                    +�      F�      	 y z p ��      �      	 y z p �                   +�      T�       4��      �       4�                   +�      T�       U�      �       U                     /�      ��       U��      ��       _؏      �       U                  �      �       P                    �      �       P�      �       T                  �      ��       P                    �      �       P�      �       T                  Ȝ      Ԝ       P                            �      "�       P"�      ��       ]��      ��       P��      ��       ][�      h�       Ph�      �       ]                        ��      ��       V'�      +�       P+�      4�       VW�      ��       V                      ��      ��       \/�      4�       PW�      �       \                       "�      &�       R��&�      +�       ���~��+�      .�      	 ���~�R�.�      �       ���~����~�                   S�      W�      	 R����~�W�      �       ���~����~�                      M�      ��       X�      �       X4�      W�       X                        U�      Y�       PY�      ��       \�      /�       \4�      W�       \                        \�      `�       P`�      ��       V�      '�       V4�      W�       V                      e�      i�      	 p  $ &�i�      ��       ���~� $ &��      �       ���~� $ &�                          m�      ��      	 s  $ &���      1�       S�      4�       S4�      R�      	 s  $ &�R�      �       S                      {�      ��      	 p  $ &���      l�       ���~� $ &��      �       ���~� $ &�                    ��       �       R �      ,�       ���~                    ��       �       Q �      Q�       ���~                    ,�      B�       TB�      U�       t0�U�      ��       ���~#0�                       ϙ      [�       ][�      ��       ���~��      ��       P��      �       ���~                         ϙ      N�       �ػ~�N�      W�       QW�      ��       �ػ~���      ��       T��      �       �ػ~�                   ϙ      ��       U��      �       }                 ��      �       ���~                 ��      �       �ػ~�                   ��      Ě       QĚ      ߚ       ���~#                  �      3�       P                    ߖ      �       P�      3�       T                 ��      3�       ���~                  z�      ��       P                  M�      T�       P                    H�      L�       PL�      O�       T                  �      �       P                    ��      �       P�      �       T                    ,�      6�       Pk�      r�       P                        '�      +�       P+�      6�       Xf�      j�       Pj�      r�       X                    �      �       P�      ��       p �                  v�      ��       P                    q�      u�       Pu�      |�       T                                         C�      G�       PG�      ��       Y֐      �       Y�      ��       Yґ      ��       Y �      |�       Y|�      ��       Qђ      ��       Y�      =�       Y�      �       Y0�      �       Y��      �       Y�      >�       Y                                             K�      ��       X֐      �       X�      �       XS�      ��       Xґ      ��       X �      u�       Xђ      =�       X�      �       X0�      4�       X��      �       X��      ݘ       Xݘ      �       P�      �       ���~�      �       X�      >�       ���~                                                                O�      q�      	 up 8�q�      ��      
 uu8�֐      �      	 up 8��      '�      	 up 8�S�      t�      	 up 8�ґ      ��      	 up 8� �      �      	 up 8�0�      >�      	 up 8�O�      ]�      	 up 8�l�      ��      	 up 8�ђ      �      	 up 8��      �      	 up 8��      �      	 up 8��      9�      
 uu8�9�      =�      
 8��      �      	 up 8��      �      	 p 8�0�      O�      	 up 8�O�      o�      
 uu8�o�      ��      
 8���      ��      	 up 8���            
 uu8�      ƕ      
 8���      И      	 up 8�И      �      
 uu8�                                                            8�      O�       0�O�      q�       up 8x �q�      ��       uu8x �֐      �       up 8x ��      �       up 8x �S�      t�       up 8x �ґ      ��       up 8x � �      �       up 8x �0�      >�       up 8x �O�      ]�       up 8x �l�      u�       up 8x �ђ      �       up 8x ��      �       up 8x ��      �       up 8x ��      9�       uu8x �9�      =�       8x ��      �       up 8x ��      �       p 8x �0�      4�       up 8x ���      ��       up 8x ���             uu8x �      ƕ       8x ���      И       up 8x �И      �       uu8x �                 �      ��       S                    R�      \�       P\�      ��       p�                   +�      =�       Q=�      �       ���~                 +�      >�       1�                    ݒ      �       S�      �       S                    ��      �       Y�      �       Y                     �      ��       0���      �       1��      �       0�                         0�      2�       1�2�      Q�       [Q�      f�       {�j�      �       [�      �       [                                �      �       \�      2�       V2�      C�       TC�      Q�       { ~ "#�Q�      f�       { ~ "�j�      ��       T��      �       V�      �       T                       �      �       up 8x ��      o�       Zo�      ��       z���      �       Z�      �       z�                    0�      2�       Pc�      f�       } p "�                 H�      W�       V                  H�      U�       P                   U�      W�       PW�      W�      
 p q "#���                  U�      W�       p ?&�W�      W�       Q                   o�      ��       Z�      �       Z                     o�      ��       U�      �       U�      �       _                       s�      ��       U��      �       _�      �       U�      �       _                  ��      ˒       P                  |�      ˒       Y                  e�      l�       P                    `�      d�       Pd�      g�       T                  F�      H�       P                    A�      E�       PE�      J�       T                  �      �       P                  �      '�       T                �      �       T                 �      �       P                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                  �      ��       P                  �      ��       T                  x�      ��       T                 S�      t�       ���~#�	                  (�      S�       P                 �      '�       ���~#�	                  ��      �       P                    ��      ��       P��      �       T                    �      ��       P��      �       X                    �      �       P�      �       Y                    ~�      ��      	 q 
��#���      ��       r�	�
��#�                    ~�      ��       Q��      ��       P��      ��       p t '�                     ݘ      �       1��      �       T�      >�       T                                                                     O�      ��       U��      ֐       _֐      ��       U��      ґ       _ґ      ��       U��       �       _ �      ǒ       Uǒ      ђ       _ђ      �       U�      2�       _2�      ?�       U?�      f�       _f�      ��       U��      �       _�      9�       U9�      �       _�      �       U�      0�       _0�      o�       Uo�      ��       _��             U      �       _��      ��       U��      �       _�      �       U�      �       _�      5�       U5�      >�       _                 �      �       U                 �      0�       ���~                 �      �       6�                 E�      `�       ���~�`�      ��       �ع~�                 l�      ��       ��~                 l�      ��       ���~�                 `�      ��       �ع~�                  ��      ��       P                  ��      ��       T                  n�      ��       P                  Y�      _�       P                    T�      X�       PX�      a�       T                    M�      Q�       PQ�      f�       X                    E�      I�       PI�      f�       Y                    �      �      	 q 
��#��      5�       r�	�
��#�                    �      �       Q�      *�       P*�      *�       p t '�                  N�      T�       P                  I�      ^�       T                N�      V�       T                 N�      T�       P                   T�      V�       PV�      V�      
 p q "#���                  T�      V�       p ?&�V�      V�       Q                        ��      ��       P��      ��       S��      ؛       V؛      ݛ       S                  ��      ��       P                    ��      ��       Pћ      ݛ       P                    ��      ��       P��      ��       T                    ��      ��       P��      ��       X                    ��      ��       P��      ��       T                    4�      d�       P'�      /�       P                          @�      Y�       QY�      [�       q�[�      `�      
 uu3&�`�      d�      
 3&�'�      /�       Q                    ]�      d�       T*�      /�       T                     4�      `�       U`�      g�       _'�      /�       U                            :�      >�       P>�      v�       Xv�      y�       Py�      ��       X�      �       P�      �       X                    A�      O�       PO�      #�       T                               A�      v�       Xv�      y�       Py�      �       Q�      �       P�      ��       X��      ��       Q��      �       X�      #�       Q                   A�      O�       PO�      #�       T                   A�      W�       UW�      #�       _                          A�      ��       0��2����      ŝ       V�S�؝      ۝       x ��۝      ߝ       x �x��      �       0��2���      #�       V�S�                        ��      Ν       ]Ν      ߝ       Pߝ      �       ]�      #�       ]                              ��      ��       P��      ��       p t ���      ŝ       Pʝ      Ν       }�Ν      ߝ       Pߝ      �       p q "��      �       P�      �       p t "��      �       P�      !�       P                      ��      ��       ^��      ��       ~���      �       ^�      #�       ^                   S�      W�       UW�      #�       _                   ��      ��       V����      ��       V�S�                  ��      �       ��                    ��      �       P�      �                         ��      چ       P                 v�      چ       ���~                    �      
�       P
�      6�       X                    �      �       P�      �       V                        :�      \�       P\�      ��       ]��      �       P�      �       ]                 ��      �       ���~                 ��      ��       �ػ~�                 �      �       ���~                 �      �       �ػ~�                 {      �{       �̷~                   {      �{       ��}��{      �{       P                     {      �{       ��L��{      �{       P�{      �{       ��~                 {      �{       ���~                     {      !{       �ػ~�!{      ${       U${      �{       �ػ~�                �{      �{       ��~                �{      �{       U                      �x      !y       V!y      �y       \n�      u�       V                       �x      �x       0��x      y       ]y      qy       Sqy      �y       sz��y      �y       Sn�      u�       0�                    <y      @y       P@y      �y       Z                    Ny      Ry       PRy      �y       [                  Zy      �y       ^                  fy      �y       X                  uy      �y       ]                  �y      �y       V                   �x      �y       _n�      u�       _                �      �       _                  �w      �x       S                      �w      �w       V�w      �w      	 p 3&��w      �w      
 3&�                       �w      �w       0��w      5x       V5x      qx       v|�qx      �x       V�x      �x       v��x      �x       p�                      x      `x       [�x      �x       P�x      �x       [                    x      #x       P#x      `x       Z                  *x      �x       \                  9x      `x       X                 9x      �x       \                  Lx      �x       ]                 �w      �x       _                    �v      �v       Sw      �w       S                    �v      �v       V�v      �v      	 p 3&�                           �v      �v       0��v      �v       Vw      'w       V'w      -w       v�-w      0w       Y0w      [w       V[w      �w       v|��w      �w       V                    Dw      Hw       PHw      �w       Z                            w      $w       \$w      'w       ^'w      *w       P*w      ^w       \^w      �w       ^�w      �w       ^                  Pw      �w       [                  ^w      �w       \                  sw      �w       ]                 sw      �w       \                   �v      �v       _w      �w       _                      À      р       Rр      �       �ȷ~�      0�       �ȷ~                    ��      ��       Z��      р      	 p 3&�                     ��      À       0�À      +�       Zd�      �       Z�      �       z��      +�       Z+�      0�       z�                    ��      �       ^+�      ��       ^                        ��      ��       P��      E�       [��      �       [�      0�       [                            �      �       R�      +�       ��~+�      E�       R��      ��       R��      �       ��~�      0�       ��~                      +�      d�       Vс      �       V+�      0�       V                       ��      d�       ]��      ��       P��      �       ]�      0�       ]                          �      E�       X      ہ       Xہ      �       S�      �       X�      0�       X                      �      d�       S�      �       S�      0�       S                  �v      w       _��      ��       _                         ��      +�       _+�      A�       UA�      ہ       _ہ      �       U�      0�       U                 �v      �v       t 8$p !0$0&�                      �v      �v       T�      �       P�      ��       T                  �v      �v       P                   ��      �       p�~��      �       T                       �      �       s ���      
�       R
�      
�       r p "�
�      �       p r "#l�7�      G�       R                       y�      �       s ���      ��       R��      ��       	�r ���      ��       T��      ��       R                  &�      n�       T                    ��      �       RӋ      �       R                    ݈      �       TӋ      ��       T                    ��      !�       XӋ      �       X                  �      6�       P                         �p      %�       �ط~%�      1�       qط~1�      s�       �ط~s�      w�       qط~w�      #�       �ط~                    �p      �q       ~���q      �q       P�q      �r       ��~                �p      �r       ]                    �p      0r       ���~�0r      Br       QBr      �r       ��~                    �p      r       ���~�r      0r       Q0r      �r       ��}                    �p       r       �ع~� r      r       Qr      �r       ��}                  �p      �p       ~8�p      �r       �̷~                �p      �r       �з~                �p      �r       ^                    �p      �p       U�p      �p       ���~��p      �r       T                �q      �q       U                �q      �q       ��}�                �q      �q       ��L                �q      �q       ^                �q      �q       U                �q      �q       ��}�                �q      �q       ��L                �q      �q       ^                �q      �q       ����                �q      �q       U                �q      �q       ��}�                �q      �q       ��L                �q      �q       ^                �q      �q       ���~�                "q      �q       @�                "q      �q       _                "q      �q       \                "q      �q       ��}�                 �o      �o        �                   �o      �o       T�o      �o       _                 �o      �o       \                 �o      �o       ���~�                 �o      Ep       D�                 �o      Ep       _                 �o      Ep       \                 �o      Ep       �ع~�                 Ep      �p       D�                 Ep      �p       _                 Ep      �p       \                 Ep      �p       ���~�                �p      �p       _                �p      �p       ���~�                                   �r      �r       R�r      �t       ���~Hv      cv       Rcv      �|       ���~�|      %�       ���~%�      1�       q��~1�      s�       ���~s�      w�       q��~w�      p�       ���~�      #�       ���~                 �r      �r       R                 �r      Ps       ��~I�      d�       ��~                   �r      �r       _�r      Ps       ��~I�      d�       ��~                 �r      Ps       \I�      d�       \                        �r      �r       0��r      s       Ps      Ps       _I�      Y�       _Y�      c�       Td�      d�       0�                   Ps      bs       A���      Ǆ       A�                       Ps      bs       ���~���      ��       ���~���      ��       U��      Ǆ       ���~�                                A�      L�      	 �й~p "�L�      U�       PU�      �       ���~i�      q�      	 �й~p "�q�      ��       P!�      v�       ���~��      χ       ���~��      Ӌ       ���~                 �t      �t       _                   �t      �t       ]�|      �|       ]                   �t      �t       ��~�|      �|       ��~                 �t      Pu       ���~�                 �t      Pu       ��}�                	 �t      3u       ��}                 Pu      �u       ���~�                 Pu      xu       U                 �u      �u       �ع~�                 �u      �u       U                 �u      v       ���~�                 �u      v       U                v      6v       _                 v      6v       S                 qv      �v       _                   �y      �y       _�      	�       _                  z      Bz       _��      ��       _                   �z      |       _߉      �       _                 ,}      M}       ���~�M}      E~       �ع~�                 Y}      �}       ��~                 Y}      �}       ���~�                 M}      E~       �ع~�                 �}      �}       P                �}      �}       ���~�                 �}      �}       ��                 �}      �}       ���~                       J      �       _�      �       U�      �       _χ      �       _                       �      '�       ���~�O�      W�       ���~�W�      [�       U[�      w�       ���~�                      )�      =�       P=�      [�       ���~� $ &�[�      i�       P                 )�      ~�       ���~�                 ~�      ~�       P                  ;�      [�       ��                  ;�      [�       R                     ��      �       _{�      ��       _��      ��       _                       ��      ƌ       ���~�{�      ��       ���~���      ��       U��      ��       ���~�                 Ռ      �       _                        @[      �[       U�[      {\       S{\      �\       �U��\      !]       S                        @[      z[       Tz[      ~\       \~\      �\       �T��\      !]       \                        @[      �[       Q�[      |\       V|\      �\       �Q��\      !]       V                        @[      �[       R�[      \       w \      �\       ��~�\      !]       w                       @[      +\       X+\      �\       �X��\      !]       X                          @[      \       Y\      �\       �Y��\      �\       Y�\      �\       �Y��\      �\       Y�\      !]       �Y�                               ~[      �[       0��[      �[       T�[      �[       ^�[      \       T�\      �\       T�\      �\       T�\      �\       Y�\      	]       T                   ~[      �[       0��[      �[       p�                     \      A\       0�A\      b\       1�b\      �\       2�                   \      \       0��\      �\       1�                   \      \       P�\      �\       P                   b\      {\       S{\      �\       �U�                   b\      {\       S{\      �\       �U�                        �X      �Y       U�Y      qZ       SqZ      {Z       �U�{Z      6[       S                          �X      !Y       T!Y      0Y       R0Y      ^Z       ]^Z      {Z       �T�{Z      6[       ]                        �X      Y       QY      0Y       X0Y      �Y       _�Y      6[       �Q�                        �X      Y       RY      wY       \wY      }Y       Q}Y      6[       �R�                      �X      Y       XY      �Y       V�Y      6[       �X�                        �X      ,Y       Y,Y      xZ       ^xZ      {Z       �U#Ȓ{Z      6[       ^                         �Y      �Y       Z���Y      �Y       Z�_��Y      lZ       �_�{Z      �Z       Z�_��Z      �Z       ���_��Z      6[       �_�                   �Y      �Y       \���Y      lZ       \�V�{Z      6[       \�V�                     �Y      �Y       [���Y      �Y       [�P�{Z      �Z       [�P��Z      �Z      
 ������                 cY      cY       V                 cY      cY       \                 cY      cY       _                 cY      cY       ]                          @W      �W       U�W      =X       S=X      LX       �U�LX      gX       UgX      �X       S                        @W      oW       ToW      �W       \�W      GX       ]GX      �X       �T�                        @W      hW       QhW      �W       V�W      IX       ^IX      �X       �Q�                   �W      �W       \���W      =X       \�V�gX      �X       \�V�                  LX      gX       0�                        �U      V       UV      |V       S|V      �V       �U��V      �V       S                          �U      V       TV      V       \V      �V       �T��V      �V       T�V      �V       \                              �U      V       QV      CV       VCV      PV       QPV      hV       s�hV      �V       �Q��V      �V       Q�V      �V       V                   �U      V       U�V      �V       S                        �             T      �       �T��      �       T�      �       �T�                        �      &       Q&      �       �Q��      �       Q�      �       �Q�                        �      �       R�      �       �R��      �       R�      �       �R�                        �             X      �       �X��      �       X�      �       �X�                    �      �       � �      �       Z                                  �      �       S�      P       R�      �       S�      �       R�      �       r �
              R       -       r �I      ]       Ru      �       r �                                �             P      g       X�      �       P�      �       X       #       X#      9       x �I      S       XS      u       x ��      �       x �                 #      #       �X�                 #      #       �R�                 #      #       Q                `      g       u��                `      g       
3��                 g      g       P                g      g       p ?&�                 i      u       u��                 i      u       Ι}�                  g      i       Pi      i      
 p q "#���                  g      i       p ?&�i      i       Q                x      �       u��                x      �       
�L�                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       u��                �      �       
3��                 �      �       P                �      �       p ?&�                 �      �       u��                  �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                �      �       u��                �      �       3� �                   �      �       P�      �      
 p q "#���                  �      �       p ?&��      �       Q                        �V      �V       U�V      W       SW      W       �U�W      3W       S                      �V      �V       T�Q��V      W       T�V�W      3W       \�V�                            �O      �O       U�O      5Q       S5Q      ?Q       �U�?Q      R       SR      R       �U�R      U       S                    �O      9P       T9P      U       ��~                            �O      �O       Q�O      :Q       ]:Q      ?Q       �Q�?Q      R       ]R      R       �Q�R      U       ]                  �O      �O       R�X�                    �O      �O       Y�O      U       �Y�                        �O      �O       u����O      �O       \�O      �O       u����O      gP       \R      �R       \                        �O      �P       _R      �S       _�S      �S       _�T      U       _                                     �O      iP       0��0��iP      6Q       V�\�6Q      8Q       �\�?Q      R       V�\�R      �R       0��0���R      �R       V�0���R      �R       V�\��R      �R       V�\��R      S       V�\�S      <S       V�\�<S      U       V�\�                           �O      �P       0�?Q      IQ       0�R      �S       0��S      �S       1��S      �S       0��T      U       1�                     �O      dP       SR      �S       S�T      U       S                   �O      dP       \R      �R       \                     �O      dP       _R      �S       _�T      U       _                     �O      dP       ]R      �S       ]�T      U       ]                     �O      dP       �O�  R      �S       �O�  �T      U       �O�                       �O      dP       ��  R      �S       ��  �T      U       ��                        \P      ^P       t p �^P      dP       TR      iR       T                  jR      �R       P                .P      @P       Y                 .P      2P       P                   2P      @P       P@P      @P      
 p t "#���                  2P      @P       p ?&�@P      @P       T                @P      DP       X                  @P      DP       QDP      DP      
 q ~ "#���                  @P      DP       q ?&�DP      DP       ^                 R      6R       Y                 R      R      
 r v #5&�                   6R      DR       YDR      DR      
 p y "#���                  6R      DR       y ?&�DR      DR       P                  DR      HR       QHR      HR      
 q x "#���                  DR      HR       q ?&�HR      HR       Q                      qR      }R       t x �}R      �R       Q�R      �R       t x �                  mR      �R       P                      �R      �R       Q�R      �R      
 q r "#����R      �R       U                   �R      �R       q ?&��R      �R       R                   �R      �R       R�R      �R       q y �                 �R      �R       P                      �R      �R       R�R      �R      
 p r "#����R      �R       P                     �R      �R       r ?&��R      �R       P�R      �R       r ?&�                         @      Y@       UY@      B       SB      B       �U�B      �J       S                                     @      c@       Tc@      ?A       w ?A      �A       ��~�A      B       w B      B       ��~B      B       w B      �B       ��~�B      I       w I      tI       TtI      �J       w                                      @      c@       Qc@      v@       Vv@      �A       �Q��A      �A       V�A      �G       �Q��G      �G       V�G      I       �Q�I      I       QI      zI       VzI      �J       �Q�                                                     @      c@       Rc@      A       ^A      �A       ��~�A      �A       ^�A      B       �R�B      �B       ��~�B      �F       �R��F      �G       ��~�G      �G       ^�G      H       ��~H      �H       �R��H      �H       ��~�H      I       ^I      )I       R)I      zI       ^zI      �I       �R��I      �I       ^�I      �J       ��~                                         @      c@       Xc@      �A       ��~�A      B       �X�B      �C       ��~�C      �F       �X��F      H       ��~H      �H       �X��H      I       ��~I      tI       XtI      zI       ��~zI      �I       �X��I      �J       ��~                         @      c@       Yc@      I       �Y�I      !I       Y!I      �J       �Y�                                         �@      �@       ����@      A       _#A      �A       _B      8B       _HB      �B       ^�B      �B       _�F      �F       _�F      �G       ��~�G      H       ^�H      �H       ��~�H      I       ����I      �I       ����I      �J       ��~                        P@      c@       Pc@      I       ��~I      tI       PtI      �J       ��~                   �@      �@       w #(�H      �H       w #(                                          �@      A       0�A      �A       VB      0B       VHB      �B       V�F      �G       V�G      H       VH      9H       0�9H      GH       r�GH      ]H       R]H      �H       r��H      �H       V�I      �I       0��I      �J       V                                          �@      A       	��A      A       \#A      )A       	��)A      �A       \B      &B       \HB      VB       ]cB      iB       	��iB      �B       ]�B      �B       \�F      �G       \�G      H       ]�H      �H       \�I      �I       	���I      �J       \                   �H      �H       ��~��H      �H       Q                           �A      �A       ��~��A      �A       U�F      �F       U�F      �G       ��~��H      �H       ��~��I      �J       ��~�                         �A      �A       U�F      �F       U�F      �G       ��~��H      �H       ��~��I      �J       ��~�                       �F      �F       U�F      �G       ��~��H      �H       ��~��I      �J       ��~�                     �F      �G       ��~��H      �H       ��~��I      �J       ��~�                     �F      �G       ~���H      �H       ~���I      �J       ~��                            �F      nG       TnG      {G       ~��H      �H       T�I      J       T$J      ^J       T^J      �J       ~�                        nG      {G       P�I      J       PXJ      ZJ       P�J      �J       P                             �F      rG       0�rG      {G       Q�H      �H       0��I      
J       0�
J      J       Q$J      �J       0��J      �J       Q                        �F      rG       0�rG      �G       1��H      �H       0��I      
J       0�
J      $J       1�$J      �J       0��J      �J       1�                           �F      �F       0��F      nG       Q�H      �H       Q�I      �I       Q$J      EJ       QZJ      }J       Q                     �F      G       ��~��I      J       ��~�$J      ZJ       ��~�                   %G      {G       ��~�ZJ      �J       ��~�                 G      �G       ��~�                	  
J      $J       ��~��J      �J       ��~�                   C      C       ��~�C      GC       T                 OC      sC       Q                   9H      GH       P�H      �H       P                      gH      sH       PsH      �H       q�H      �H       P                 gH      �H       U                 �H      �H       P                  qH      �H       ��                  qH      �H       X                   9H      GH       Q�H      �H       Q                �@      �@       ���                    �A      �A       R�G      �G       R                    �A      �A       ^�G      �G       ^                        �G      �G       0��G      �G      	 p ~  ��G      �G       p ~ O��G      �G      	 p ~  �                     �A      �A      
 1r 7$1��A      �A       1�Q#(} 7$1��G      �G      
 1r 7$1�                  �A      �A       R�G      �G       R                  �A      �A       ^�G      �G       ^                    �A      �A       R�A      �A      
 } �Q#("�                  �A      �A       ^                  �A      �A       B�                  �A      �A       P                       �B      C       S{C      �E       S�E      �F       SH      H       SzI      �I       S                                  	C      C       0��C      �C       0��C      �D       V	E      (E       [(E      4E       T4E      �E       t��E      �E       T�E      �E       VF      �F       VH      H       0�zI      �I       V                    cE      �E       R�E      �E       r�                	 	   	 �B      C       s{C      �C       s�C      �C       PH      H       s                           �C      �C      
 p < $0.��C      �D       v5$s "#�< $0.��E      �E      
 p < $0.�F      UF       v5$s "#�< $0.�nF      }F       v5$s "#�< $0.�zI      �I       v5$s "#�< $0.�                            �C      %D       U%D      �D       x 
���F      LF       x 
���LF      nF       t 
���nF      }F       x 
���zI      �I       x 
���                              D       D       P D      YD       y 
���YD      �D       | 5$s "#<�
���F      2F       y 
���2F      UF       | 5$s "#<�
���nF      }F       | 5$s "#<�
���zI      �I       | 5$s "#<�
���                           D      %D       u �%D      �D       x 
���F      LF       x 
���LF      nF       t 
���nF      }F       x 
���zI      �I       x 
���                             D       D       p � D      YD       y 
���YD      �D       | 5$s "#<�
���F      2F       y 
���2F      UF       | 5$s "#<�
���nF      }F       | 5$s "#<�
���zI      �I       | 5$s "#<�
���                           D      3D       Z3D      �D       @<$x 
��{ x 
�� $0.( �F      LF       @<$x 
��{ x 
�� $0.( �LF      nF       @<$t 
��{ t 
�� $0.( �nF      }F       @<$x 
��{ x 
�� $0.( �zI      �I       @<$x 
��{ x 
�� $0.( �                                D      D       QD       D       @<$p { p  $0.( � D      YD       @<$y 
��{ y 
�� $0.( �YD      �D      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( �F      2F       @<$y 
��{ y 
�� $0.( �2F      UF      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( �nF      }F      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( �zI      �I      / @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( �                          D      �D       QF      uF       QuF      }F      � @<$x 
��{ x 
�� $0.( @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( @<$x 
��{ x 
�� $0.(  $@<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.(  $,( �zI      �I       Q�I      �I      � @<$x 
��{ x 
�� $0.( @<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.( @<$x 
��{ x 
�� $0.(  $@<$| 5$s "#<�
��{ | 5$s "#<�
�� $0.(  $,( �                          'D      �D       U�D      �D       p �F      }F       UzI      �I       U�I      �I       p �                 nD      �D       U                     'D      �D       
 ��F      �F       
 ��zI      �I       
 ��                     'D      �D       
 ��F      �F       
 ��zI      �I       
 ��                     'D      �D       0�F      �F       0�zI      �I       0�                  uD      �D       s t "#(��I      �I       s t "#(�                           �C      �C       s t "#��C      �C       s t "H��C      �D      
 v5$s "#��E      �E      
 v5$s "#�F      �F      
 v5$s "#�zI      �I      
 v5$s "#�                
           �C      uD      
 v5$s "#�uD      �D       s t "#(��E      �E      
 v5$s "#�F      }F      
 v5$s "#�zI      �I      
 v5$s "#��I      �I       s t "#(�                  4E      VE       T                 4E      VE       ]                  @E      VE       ��                  @E      VE       P                 �E      �E       0�                 �E      �E       �R�                     9H      NH       QNH      WH       q`�]H      �H       Q                   I      LI       QLI      pI       r                    I      )I       ���)I      pI       R                            �             U      �       Y�      �       U�      �       Y�      �       U�      �       Y                                �             T      �       �T��      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T�                                      �      S       QS      �       �Q��      �       Q�      �       �Q��             Q      c       w c      �       �Q��      �       Q�      �       w �      �       Q�      �       �Q�                        �      %       0�%      S       P�      �       0��      �       0�                   �      �       T�      �       T                                     �      S       QS      �       �Q��      �       Q�      �       �Q��             Q      c       w c      �       �Q��      �       Q�      �       w �      �       Q�      �       �Q�                          W       PW      Y       T                     G      O       r t "#��@&�O      Q      8 w #�z�O%w #�z�"1& $ &y� $ &t "#��@&�Q      c      g w #�z�O%w #�z�"1& $ &y� $ &w #�z�O%w #�z�"1& $ &y� $ &?&"#��@&�                      G       y                      G       w #�z�2�                   @      G       RG      G      
 r t "#���                  @      G       r ?&�G      G       T                      �      �       x��      �       T�      �       t��      �       T                 �      �       X                        �      �       x { ��      �       {  x "��      �       | { ��      �       {  | "��      �       p�                     I      S       Z�      c       Z�      �       Z�      �       Z                       �      �       p ����#5$y "#��      �      
 r5$y "#��      �      
 r 5$y "#��             p ����#5$y "#�                                �      W       TW      z       �T�z      �       T�      �       �T��      �       T�      �       �T��      �       T�      �       �T�                                   �      �       P�      �       R�             P      !       R#      8       P8      >       Q>      C       PU      W       0��      �       P�      �       u$                   d      k       Pk      k      
 p r "#���                  d      k       p ?&�k      k       R                 �      �       u                   �      �       t r ��      �       �Tr �                 z      �       u                   z      �       T�      �       �T�                      �      �       T�      �      
 p t "#����      �       P                     �      �       t ?&��      �       P�      �       t ?&�                        p.      �.       T�.      �/       �T��/      �/       T�/      �/       �T�                        p.      /       R/      ,/       �R�,/      N/       RN/      p/       �R�p/      �/       R                              p.      /       X/      ,/       �X�,/      </       X</      p/       �X�p/      �/       X�/      �/       �X��/      �/       X                      p.      T/       YT/      p/       �Y�p/      �/       Y                                          �.      /       T/      "/       { p��,/      N/       TN/      \/      
 p�p��p/      /       T/      �/       p�z ��/      �/       T�/      �/       p�z ��/      �/       T�/      �/       { z ��/      �/       T�/      �/       { z ��/      �/       T�/      �/       { z �                       �.      "/       P,/      \/       Pp/      �/       P�/      �/       P                     �.      �.       Q�.      �.       P�/      �/       Q                  �.      �.       T�/      �/       T                 �.      �.       P                    �.      �.       ���/      �/       ��                    �.      �.       Z�/      �/       Z                 (/      ,/       U                N/      `/       Y                 N/      Y/       X                   Y/      `/       X`/      `/      
 p x "#���                  Y/      `/       x ?&�`/      `/       P                        �-      �-       U�-      �-       V�-      �-       �U��-      m.       V                        �-      �-       T�-      �-       �T��-      .       T.      m.       �T�                          �-      �-       Q�-      �-       S�-      �-       �Q��-      .       Q.      m.       S                 X.      d.       T                 �-      �-       P                     �-      .       T.      Q.       �T�X.      X.       �T�                   �-      Q.       \X.      X.       \                    .      <.       0�<.      Q.       TX.      X.       T                   .      Q.       PX.      X.       P                 .      .       |�&                                              0�      }�       U}�      ޟ       _ޟ      ţ       �U�ţ      �       _�      ��       �U���      ��       U��      ]�       _]�      �       �U��      S�       _S�      ��       �U���      ��       _��      �       �U��      ��       U��      w�       �U�w�      ��       _                                              0�      }�       T}�      ��       V��      �       ���      ţ       �T�ţ      �       ���      ��       �T���      ��       T��      ]�       V]�      �       �T��      +�       ��+�      :�       �T�:�      K�       ��K�      �       �T��      ��       T��      ��       �T�                                              0�      }�       Q}�      �       ]�      ţ       �Q�ţ      �       ]�      ��       �Q���      ��       Q��      ]�       ]]�      �       �Q��      S�       ]S�      ��       �Q���      ��       ]��      �       �Q��      ��       Q��      w�       �Q�w�      ��       ]                     j�      }�       u ��      ��       u ��      ��                                  t�      ��       S˦      Χ       SΧ      �       p �      �       S��      ��       S                         W�      ��       \ţ      �       \��      ]�       \�      S�       \�      ��       \                                         ��      ��       s���      ޟ       _ޟ      ţ       �U�ţ      �       _�      ��       �U�˦      ��       �U�]�      �       �U��      S�       _S�      ��       �U���      ��       _��      �       �U���      w�       �U�w�      ��       _                      ��      z�       Pţ      �       P�      S�       P                        Ğ      ş       Yţ      �       Y�      S�       Yw�      ��       Y                       Ğ      ş       Xţ      �       X�      S�       Xw�      ��       X                          Ğ      ��       0���      ��       s˦      ��       0�]�      �       0���      �       0��      *�       s*�      ��       0�                     ��      ��       Q��      ��       | �      *�       ��~                           ��      �       q�ţ      �       q��      �       #��      '�       q�'�      +�       #�:�      K�       #�                       ��      ş       Rţ      �       R�      S�       Rw�      ��       R                                         ��      ��       s���      ޟ       _ޟ      ţ       �U�ţ      �       _�      ��       �U�˦      ��       �U�]�      �       �U��      S�       _S�      ��       �U���      ��       _��      �       �U���      w�       �U�w�      ��       _                   ��      �       �1   ţ      ��       �1                      ��      �       �   ţ      ��       �                      ��      �       ���ţ      ��       ���                   ��      �       ���ţ      ��       ���                                   ��      ޟ       _ޟ      ţ       �U��      ��       �U�˦      ��       �U�]�      �       �U�S�      ��       �U���      ��       _��      �       �U���      w�       �U�w�      ��       _                     ��      �       �����      ��       ���w�      ��       ���                     ��      ��       T��      ş       s�w�      ��       T                  Ɵ      �       P                              �      ţ       �   �      ��       �   ˦      ��       �   ]�      �       �   S�      ��       �   ��      �       �   ��      �       �   *�      w�       �                                 �      ţ       ����      ��       ���˦      ��       ���]�      �       ���S�      ��       �����      �       �����      �       ���*�      w�       ���                                  �      ţ       ����      C�       ���C�      L�       TL�      ��       ���˦      ��       ���]�      �       ���S�      ��       �����      �       �����      �       ���*�      w�       ���                              �      ţ       S�      ��       S˦      ��       S]�      �       SS�      ��       S��      �       S��      �       S*�      w�       S                             �      ţ       0��      ��       0�˦      ��       0�]�      �       0�S�      ��       0���      �       0���      w�       0�                    �      t�       VS�      _�       V_�      f�       0�                               �      ţ       ����      �       ���˦      ��       ���]�      �       ���f�      ��       �����      �       �����      �       ���*�      w�       ���                               �      ţ       S�      �       S˦      ��       S]�      �       Sf�      ��       S��      �       S��      �       S*�      w�       S                   �      _�       s�ԩ      ��       s�                              �      <�       0�<�      B�       1�B�      u�       \u�      {�       1�{�      �       \�      ��       1���      ��       1�l�      ��       \ �      �       \ԩ      =�       \E�      I�       1�I�      ��       \                     H�      _�       �#�'�ԩ      ߩ       p�'�ߩ      ��       �#�'�                   �      H�       0�H�      _�       �#�'�0.�ԩ      ��       �#�'�0.�                         �      _�       [Ĩ      ��       [ԩ      ��       [��      ��       w ª      ͪ       P                	           �      �       ]l�      ��       ]]�      �       ]ԩ      ��       ]��      ͪ       ]*�      w�       ]                         ,�      *�       ^l�      ��       ^]�      c�       ^ �      �       ^ԩ      ��       ^                            m�      ~�       P~�      ��       u�#�
��@$�A�      j�       V|�       �       V��      ͪ       V*�      w�       V                     A�      Y�       �B$x �*�      G�       �B$x �G�      ]�       �B$��~��                    ʡ      �       Q]�      i�       Q                          �      Y�       X]�      w�       Xw�      |�       s�*�      G�       XG�      ]�       ��~                  ��      ��       s��                  ��      ��       Y                  ��      ��       0�                  ��      ��       s��                  ��      ��       Q                  ��      ��       V                  ��      6�       s��                  ��      1�       Y                  ��      6�       ]                  ��      6�       s��                  ��      �       s�                  ��      6�       V                           ��      ţ       S�      �       S˦      l�       Sf�      ԩ       Sͪ      �       S��      �       S                           ��      ţ       s���      �       s��˦      l�       s��f�      ԩ       s��ͪ      �       s����      �       s��                 ��      â       V                            #�      g�       Z��      ��       q t ���      ţ       Zh�      j�       p r �j�      ��       P��      ��       p r ���      ��      	 q��r �                             ��      #�       0�#�      ţ       \�      K�       \˦      l�       \f�      ��       \ͪ      �       \��      �       0�                      ��      K�       P˦      l�       Pf�      �       P                     ��      ţ       Y�      ��       Y��      �       Y                       ��      ţ       X�      )�       X)�      3�       x���      �       X                           �      ţ       ]�      �       ]˦      l�       ]f�      ԩ       ]ͪ      �       ]��      �       ]                           �      ţ       ^�      �       ^˦      l�       ^f�      ԩ       ^ͪ      �       ^��      �       ^                      ��      ţ       v���      B�       v��˦      l�       v����      �       v��                      ��      ţ       v���      B�       v��˦      l�       v����      �       v��                      �      ţ       v���      B�       v��˦      l�       v����      �       v��                      �      ţ       v���      B�       v��˦      l�       v����      �       v��                               �      #�       0�#�      ţ       R�      ?�       0���      ��       0���      ;�       [m�      ��       0���      �       R˦      l�       [                           �      ţ       NB$��      �       NB$�˦      l�       NB$�f�      ԩ       NB$�ͪ      �       NB$���      �       NB$�                           �      ţ       �B$��      �       �B$�˦      l�       �B$�f�      ԩ       �B$�ͪ      �       �B$���      �       �B$�                 ��      â       V                 ��      �       s��                 ��      �       s��                 ��      �       s��                �      ��       �U%                  �      ��       �!%                  ��      ��       �b%                  ��      ��       �.%                  ��      �       �o%                  ��      �       �;%                  �      �       �|%                  �      �       �H%                            Ԥ      �       2��      -�       X˦      ݦ       0�ݦ      �       Ya�      l�       Y                              Ԥ      �       �����      �       Y�      $�       U$�      -�       Y˦      ݦ       ����ݦ      �       R�      �       X�      @�       Ra�      l�       X                      ��      -�       R�      �       U/�      l�       U                        �      -�       U��      �       X;�      a�       Qa�      l�       X                      Τ      -�       Q˦      7�       Qa�      l�       Q                y�      ��       T                y�      ��       ���|�                   ��      ��       Q��      ��      
 p q "#���                  ��      ��       q ?&���      ��       P                �      ��       T                  �      ��       Q��      ��       s�                   ��      ��       P��      ��      
 p q "#���                  ��      ��       p ?&���      ��       Q                   Ԩ      Ԩ       s��Ԩ       �       ��~ª      ͪ       s��                   Ԩ       �       0�ª      ͪ       0�                   Ԩ      ��       [ª      ͪ       P                   Ԩ      Ԩ       s��Ԩ      ��       Rª      ͪ       s��                   Ԩ      ��       Qª      ͪ       Q                   Ԩ       �       Vª      ͪ       V                  �      ��       V                 �      ��       s�                     �      ��       ��~���      ��       R��      ��       ��~�                     �      ��       ��~���      ��       T��      ��       ��~�                 �      ��       s�#                 �      ��       P                   �      ��       s��S�      f�       s��                 �      *�       P                 t�      ��       s��                 t�      ��       V                 ��      ��       s��                    ��      ��       Q��      ��       |                    ��      ��       R��      ��       s�                 �      ]�       s�                 �      ]�       s��                            �_      �_       U�_      �_       \�_      �_       �U��_      �`       \�`      �`       �U��`      �`       \                            �_      �_       T�_      �_       V�_      �_       �T��_      �`       V�`      �`       �T��`      �`       V                     �_      �_       P�_      �_       P�`      �`       P                           �_      �_       U�_      �_       \�_      �_       �U��_      �`       \�`      �`       �U��`      �`       \                   �_      �_       t�_      �_       v                   �_      �_       t �_      �_       v                   �_      �_       0��_      �_       P                 �_      �_       3�                   �_      �_       0��_      &`       0�                   �_      �_       v�_      `       v                   �_      �_       v�_      `       v                    �_      �_       P�_      &`       P                  `      `       R                 `      !`       Q                    �_      �_       0�&`      i`       0��`      �`       0�                    �_      �_       v(&`      Y`       v(�`      �`       v(                    �_      �_       v &`      U`       v �`      �`       v                   R`      ``       R                 R`      d`       P                  �_      �_       1�i`      �`       1�                 �_      �_       v8i`      �`       v8                 �_      �_       v0i`      �`       v0                  �`      �`       R                 �`      �`       Q                          �m      n       Un      <n       \<n      ?n       �U�?n      Qn       \Qn      Xn       �U�                      �m      n       Tn      n       Vn      Xn       �T�                  	n      n       P'n      ?n       P                         �m      n       Un      <n       \<n      ?n       �U�?n      Qn       \Qn      Xn       �U�                      �m      9n       S?n      Nn       SNn      Wn       U                   �m      n       tn      n       Q                   �m      n       t n      n       T                �m      	n       S                  �m      	n       0�	n      	n       P                      n      'n       ]?n      Sn       ]Sn      Wn       Q                      n      'n       V?n      On       VOn      Wn       T                      n      'n       S?n      Nn       SNn      Wn       U                    #n      'n       P?n      Wn       P                     n      'n       S?n      Nn       SNn      Wn       U                 n      #n       1�                    �=      �=       U�=      >       �U�                    �=      �=       T�=      >       �T�                   �=      �=       U�=      >       �U�                  �=      >       S                        �      �       U�      �       S�      �       �U��             S                          �      �       T�      �       V�      �       �T��             T             V                    �      �       q u ��      �       U                   �      �      
 q u s8"��      �       U                                 +       U+      G       SG      K       �U�K      �       S�      �       �U�                                 +       T+      K       �T�K      l       Tl      �       \�      �       �U#                   #      +       u K      s       s                        #      +       r t �K      T       r t �T      l       st �l      s       s| �                  �      �       ��                  �      �       P                  /      B       @�                  /      B       Q                          >      7>       U7>      �>       V�>      �>       �U��>      �>       U�>      ?       V                        >      7>       T7>      �>       �T��>      �>       T�>      ?       \                        >      7>       Q7>      �>       �Q��>      �>       Q�>      ?       �Q�                         >      7>       U7>      �>       V�>      �>       �U��>      �>       U�>      ?       V                    ">      �>       S�>      ?       S                       ">      7>       s��7>      �>       Q�>      �>       s���>      ?       Q                   ">      7>       s�&�>      �>       s�&                      �>      �>       P�>      �>       Q�>      ?       P                  ?      ?       \                  ?      ?       |�                 a>      �>       R                a>      �>       t�                 �>      �>       P                  c>      �>       t�                  c>      �>       R                      �l      �l       U�l      Cm       SCm      Gm       �U�                    �l      �l       T�l      Gm       �T�                    �l      �l       Q�l      Gm       �Q�                      �l      �l       R�l      �l       Z�l      Gm       �R�                    �l      �l       X�l      Gm       �X�                      �l      �l       Y�l      Fm       \Fm      Gm       �U#�                  �l      �l       �                   �l      �l       �                    �l      Dm       VDm      Gm       �U#�                �l      m       Q                �l      m       v�                 m      m       P                  �l      m       v�                  �l      m       Q                            r       Ur      �       S�      �       �U�                        �       V                       \       U                       \       P                          �8      �8       U�8      t9       St9      ~9       �U�~9      �9       S�9      �9       �U�                          �8      �8       T�8      y9       ]y9      ~9       �T�~9      �9       ]�9      �9       �T�                      �8      �8       Q�8      �8       ���8      �9       �Q�                          �8      �8       R�8      {9       ^{9      ~9       �R�~9      �9       ^�9      �9       �R�                          �8      �8       X�8      w9       \w9      ~9       �U#�~9      �9       \�9      �9       �X�                          �8      �8       Y�8      u9       Vu9      ~9       �U#�~9      �9       V�9      �9       �Y�                  �8      �8       �                   �8      �8       �                  �8      �8       �                   �8      9       P~9      �9       P                   �8      �8       t��8      �8       U                    �8      9       P~9      �9       P                    �             T      �       u�                    �      �       Q�      �       �Q�                   �             P      �       u�                                                    T      |       t��      �       t��      �       {��      �       T�      �       t��      �       R�             T             t�      #       t�5      <       t�<      �       [�      �       t�                            �      4       Q4      k       u�k      &       Q&      5       u�5      �       Q�      �       u�                 �      �       U                               F       u�F      k       u�@�k      |       u��      �       u��             X      �       u��      �       u� �                                     1       0�1      k       2�k      |       0��      #       0�#      5       4�5      �       0��      �       2��      �       4�                                             |       0��      �       0��      �       P�      �       0��      �      & t��H$t��@$!t��8$!t��!��      �      & r|��H$r}��@$!r~��8$!r��!��      �       P      Z       0�Z      b       Pb      {       0�{      �       P�      �       0�                      1      k       2�#      5       4��      �       2��      �       4�                        �7      �7       U�7      8       S8      p8       �U�p8      v8       U                      �7      �7       T�7      p8       �T�p8      v8       T                       8      8       0�8      ,8       s�,8      R8       SR8      X8       P                      8      8       P8      W8       ]X8      o8       ]                      �7      �7       Pp8      u8       Pu8      v8       u�	                  18      F8       U                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                    �      �       U�      �       �U�                    �      �       T�      �       �T�                 �      �       u                  �      �       u #�                      �      �       U�      �       S�      �       �U�                 �      �       u                  �      �       u #�                        `      t       Ut      �       T�      �       �U��      �       T                    `      f       Tf      �       �T�                    c      �       Y�      �       Y                    t      �       U�      �       U                     t      x       Px      �       y��      �       y�                      �      �       U�      >       �U�>      D       U                                 �             0�             P             0�      (       X(      1       0�1      4       P4      ;       X;      >       P>      D       0�                               �      �       t �      �       t �#��      
       Q
            ' t �#�U#�t �#�����U#�*( �      (       Q(      /       R/      1       0�4      >       Q>      D       0�                    �      �       T�      �       �T�                 �      �       0�                    s      �       P�      �       u                    s      �       p���      �       u #��                0      ^       1�                0      ^       U                   3      G       PG      ^       u                  :      ^       Q                �             0�                �             U                   �             P             u                  �             Q                      @e      Ye       UYe      e       Ve      �e       �U�                          @e      Ye       TYe      �e       \�e      �e       �T��e      �e       \�e      �e       �T�                         @e      Ye       0�Ye      ce       Pce      ue       0�ue      �e       P�e      �e       0��e      �e       P                              Le      ~e       S~e      �e       | �e      �e       �T�e      �e       S�e      �e       S�e      �e       | �e      �e       P                ke      ue       S                ke      ue       V                  ke      ue       0�ue      ue       P                    `      r       Tr      �       �T�                    `             Q      �       �Q�                 `      �       ��I                   `      �       T                 `      �       U                       `      d       u t "�d      k       Pk      r       u t "�r      �       u �T"�                 `      �       ��I                   `      �       U                    r             0�      �       Y�      �       R                   `      z       q 
���z      �       Q                    �      �       P�      �       r ���                  �      �       X                       0      	0       U	0      !0       �`!0      �2       �U�                     0      2       T2      �2       �T�                     0      2       Q2      �2       �Q�                    0      2       q��2      �2       �Q#��                                              t0      x0       0�x0      �0       P�0      �0       p��0      �0       0��0      �0       P�0      �0       p��0      �0       0��0      �0       P�0      �0       p�1      1       0�1      1       P1      "1       p�s1      w1       0�w1      �1       P�1      �1       p��1      �1       0��1      �1       P�1      �1       p�                            t0      �0       U�0      �0       U�0      �0       U1      j1       Us1      �1       U�1      �2       U                    (2      /2       Q/2      ;2       P;2      ;2       p q '�                          �2      �2       U�2      �3       S�3      �3       �U��3      S4       SS4      U4       �U�                    �2      �3       Q�3      U4       �Q�                 �2      �3       T                 �3      U4       T                        T       P                    �,      �,       U�,      ~-       X                 -      ;-       T                 P-      ~-       T                          0      m       Um      q       �U�q      �       U�             �U�             U                      4      �       P�      �       �U#(�             P                      X      m       Rq      �       0�             R                      �      �       T�      �       T�      �       r  $ &4$p"�                      �      �       U�      �       U�      �      	 pz "@�                   �      �      	 py "1��      �      	 py "1�                      �4      �4       U�4      K5       �U�K5      X5       U                      �4      (5       S)5      W5       SW5      X5       u(                  <5      D5       P                  �      �       P                      �6      �6       U�6      �7       S�7      �7       �U�                    �6      �6       T�6      �7       �T�                      �6      �6       Q�6      57       \57      �7       �Q�                      �6      �6       R�6      57       V57      �7       �R�                    �6      �6       X�6      �7       �X�                  �6      �6       U                 7      57       \                    7      7       P7      57       |�                           �      �       U�      �       �U��             U      �       �U��      �       U                      �      C       PC      I       �U#(I      �       P                      �      �       R�             0��      �       R                            ,       TI      ^       T^      q       r  $ &4$p"�                      $      ,       UI      T       UT      q      	 pz "@�                   $      ,      	 py "1�I      q      	 py "1�                          `4      w4       Uw4      �4       �U��4      �4       U�4      �4       �U��4      �4       U                            e4      �4       S�4      �4       S�4      �4       u(�4      �4       S�4      �4       S�4      �4       u(                  �4      �4       P                          �]      �]       U�]      �]       S�]      �]       �U��]      �]       S�]      �]       �U�                          �]      �]       T�]      �]       V�]      �]       �T��]      �]       V�]      �]       �T�                          �]      �]       Q�]      �]       \�]      �]       �Q��]      �]       \�]      �]       �Q�                    �]      �]       P�]      �]       �\                  �]      �]       1�                    �]      �]       U�]      �]       S                           S       US      �       �U�                           o       To      �       �T�                             o       Qo      �       \�      �       �Q�                           o       Ro      �       �R�                      ,      C       VC      J       u(J      �       V                  k      �       ]                   k      o       Po      �       S                      `5      �5       U�5      ~6       S~6      �6       �U�                    `5      �5       T�5      �6       �T�                      `5      �5       Q�5      �5       ]�5      �6       �Q�                      `5      �5       R�5      �5       V�5      �6       �R�                    `5      �5       X�5      �6       �X�                  �5      �5       U                     $      H$       UH$      I$       �U�                       $      +$       T+$      H$       ZH$      I$       �T�                       $      5$       Q5$      H$       [H$      I$       �Q�                       $      5$       R5$      H$       XH$      I$       �R�                  $      6$       U                                 +      �+       U�+      ,       ^,      ,       �U�,      ",       U",      -,       ^-,      :,       U:,      X,       ^X,      e,       U                     +      ?+       T?+      e,       ��                         +      C+       QC+      ,       \,      ,       �Q�,      e,       \                  +      D+       U                   K+      ,       \,      e,       \                   K+      ,       ��,      e,       ��                           K+      �+       ]�+      �+       T�+      ,       ],      :,       ]:,      F,       TF,      e,       ]                             K+      �+       U�+      ,       ^,      ",       U",      -,       ^-,      :,       U:,      X,       ^X,      e,       U                  D,      F,       S                              P+      �+       0��+      ,       _,      ",       0�",      -,       _-,      :,       0�:,      V,       _V,      X,       	��X,      e,       0�                        \+      �+       P,      ",       P-,      :,       PX,      e,       P                   \+       ,       0�,      e,       0�                     �+      �+       S",      +,       SF,      X,       S                    p,      �,       U�,      �,       �U�                      p,      {,       T{,      �,       Y�,      �,       �T�                 p,      �,       U                          @
      �
       U�
      �
       Z�
      �
       �U��
      �
       U�
             Z      �       U                    @
      R
       TR
      �       [                          @
      Y
       QY
      �
       V�
      �
       �Q��
      �
       V�
             �Q�      �       V                            @
      Y
       RY
      �
       S�
      �
       �R��
      r       Sr             �R�      �       S                       ]
      �
       Y�
      �
       y��
      K       Y]      �       Y�      �       Y                 @
      Z
       U                       |
      |
       V|
      �
       v 1$��
      �
       V�
      K       Q      �       v 1$��      �       Q�      �       Q                   |
      �
       [�
      K       [      �       [�      �       [                          |
      �
       P�
      �
       P�
      �
       u�
      �
       z      �       P�      �       u�      �       u                   |
      �
       �([  �
      K       �([        �       �([  �      �       �([                     |
      �
       Y�
      K       Y      �       Y�      �       Y                            |
      �
       0��
      �
       0��
      �
       V�
      �
       U�
      ,       V,      ;       U      �       0��      �       0�                      |
      �
       0��
      �
       0��
      @       ]@      K       }�      �       0�                          |
      �
       1��
      �
       1��
             P             P      &       1�&      C       P      �       1��      �       1�                        �
      �
       t ���
              t ��              u ���      4       T                     
      1
       U1
      2
       �U�                  
      )
       U                            �)      A*       UA*      �*       _�*      �*       �U��*       +       _ +      +       U+      +       _                            �)      >*       T>*      v*       Sv*      �*       �T��*      +       S+      +       �T�+      +       S                            �)      9*       Q9*      �*       V�*      �*       �Q��*       +       V +      +       Q+      +       V                            �)      4*       R4*      �*       \�*      �*       �R��*       +       \ +      +       R+      +       \                          �)      E*       XE*      �*       �X��*       +       �X� +      +       X+      +       �X�                      q*      v*       ��y�v*      �*       S+      +       S                           �)      *       0�*      �*       P�*      �*       0��*      �*       P�*      +       0�+      +       ��                      d*      �*       ^�*       +       ^+      +       ^                      h*      �*       ]�*       +       ]+      +       ]                    P$      $       U$      �)       ��~                              P$      q$       Tq$      �$       S�$      w(       ��~w(      �(       S�(      �(       ��~�(      )       S)      �)       ��~                    P$      $       Q$      �)       ��~                        P$      $       R$      B%       ]B%      G%       �R�G%      �)       ]                    P$      $       X$      �)       �X�                    �$      �$       ^w(      �(       ^�(      _)       ^_)      l)       ~�                                      �$      �$       1��$      )%       ��~���~�"| �G%      �%       ��~���~�"| ��%      d&       ��~���~�"��~��s&      �&       ��~���~�"| ��&      �&       |  ��~�"��~�"��&      �&       ��~���~�"| ��&      w(       ��~���~�"| �w(      �(       ]�(      �(       ��~���~�"| ��(      l)       1�l)      �)       ��~���~�"| �                                   �$      �$       0��$      )%       \G%      �%       \�%      d&       ��~s&      �&       \�&      w(       \w(      �(       0��(      �(       1��(      �(       \�(      Y)       0�Y)      l)       1�l)      �)       \                 )%      5%       3�                                 �$      �$       R�$      )%       ��~G%      s&       ��~s&      �&       7��&      �(       ��~�(      �(       ��~�(      *)       R*)      P)       ��~P)      l)       8�l)      �)       ��~                  )      l)       \                  )      l)       V                            %      )%       SG%      �%       Ss&      �&       S�&      w(       S�(      �(       S�)      �)       S                       
'      /'       Pr'      �'       P�'      �'       PT(      w(       P                               %      )%       0�G%      �&       0��&      (       0�(      !(       P!(      8(       RE(      w(       0��(      �(       0�l)      �)       0�                    �'      �'       ��~# �'      
(       ��~�(      �(       R                   �'      E(       V�(      �(       V                 s&      �&       S                  �&      �&       P                      u%      y%       Py%      s&       ��~l)      �)       ��~                       u%      }%       0�}%      �%       P�%      q&       Vq&      s&       0�l)      �)       V�)      �)       0�                    �%      �%       Pl)      �)       P                      �%      �%       0��%      &       |�&      N&       \N&      d&       |�                    �%      &       S&      d&       S                    /'      r'       U�(      �(       U�)      �)       U                     5'      r'       Q�(      �(       Q�)      �)       Q                     5'      a'       0��(      �(       0��(      �(       1��)      �)       0�                              �"      &#       U&#      �#       ���#      �#       U�#      �#       ���#      �#       U�#      $       ��$      $       U                        �"      !#       T!#      �#       S�#      �#       �T��#      $       S                              �"      &#       Q&#      �#       ���#      �#       Q�#      �#       ���#      �#       Q�#      $       ��$      $       Q                                �"      &#       R&#      �#       ]�#      �#       �R��#      �#       R�#      �#       ]�#      �#       R�#      $       ]$      $       R                    �"      �"       X�"      $       ��                  $      $       _                                       �"      &#       0�&#      M#       XM#      �#       ^�#      �#       X�#      �#       X�#      �#       0��#      �#       X�#      �#       0��#      $       X$      $       ^$      $       	��$      $       0�                       �"      &#       P�#      �#       P�#      �#       P$      $       P                   �"      �#       0��#      $       0�                     9#      �#       _�#      �#       _$      $       _                             	      H	       UH	      X	       \X	      _	       �U�_	      
       \
      
       �U�
      
       \                             	      D	       TD	      \	       ^\	      _	       �T�_	      
       ^
      
       �T�
      
       ^                       	      H	       QH	      U	       SU	      
       �Q�                             	      H	       RH	      V	       VV	      _	       �R�_	      
       V
      
       �R�
      
       V                      i	      
       ]
      
       �U
      
       ]                        m	      q	       Pq	      	
       w 	
      
       ��
      
       w                      m	      �	       ^�	      �	       S
      
       ^                      u	      
       _
      
       �Q����33$�T"�
      
       _                        P      �       U�      �       S�      �       �U��      	       S                        P      z       Tz      �       V�      �       �T��      	       V                  �      	       Q                       �      �       \�      �       \�      �       T�      	       \                     �      �       1��      �       ]�      �       }��      	       ]                 v             U                 �      �       S                 �      �       S                                  %       U%      4       V4      5       �U�5      J       VJ      K       �U�K      ?       V                         -      3       S3      4       v 4      5       �U5      =       SK      ?       S                                   -             0�      K       PK      �       0��      �       P�      �       0��      �       P�             0�             P      (       0�(      -       3�-      ?       0�                            �             U      �       S�      �       �U��      �       S�              �U�              S                          �             T      �       Z�      �       �T��              Z              T                  �              Q                           �             0�      R       [R      V       {�V      �       [�      �       [�      �       {��      �       [�             0�                                 �      !       0�!      =       P=      l       0�l      �       P�      �       0��      �       P�      �       0��              P              0�                  �      �       Q                    p      }       U}      �       Y                      p      �       T�      �       X�      �       T                  �      �       Q                   w      �       0��      �       P                          �      �       R�      �       Q�      �       R�      ^       Q^      h       R                         �      �       0��      �       Y�      P       YP      T       y�T      ^       Y^      h       0�                     �      �       3��      �       P�      h       3�                        �             0�             R             r�      7       R                         �      �       r �      �       r �             r              q7      ^       r                           K       Pf      r       P                    D      j       Pj      o       p�                      �      �       U�             S             �U�                 �      �       u8                          �             U      #       S#      ,       �U�,      �       S�      �       �U�                 �      �       u8                    �      +       \,      �       \�      �       0�                 ?      w       \                 ?      w       S                  Q      w       T                 Q      w       P                 Q      w       R                                  7       U7      i       Si      o       �U�o      �       S�      �       �U��      �       S                                   T      l       \l      �       �T�                                  4       Q4      j       Vj      o       �Q�o      �       V�      �       �Q��      �       V                                          �      �       U�             X      >       ��>      �       �U��              U       4        �U�4       b        Ub       |        ��|       �        �U��       !       U!      �"       �U��"      �"       ���"      �"       U                                                �      �       T�             ^      >       T>      �       ^�              T               ^       4        �T�4       b        ^b       |        T|       �        ^�       �        T�       >"       ^>"      E"       TE"      �"       ^�"      �"       T�"      �"       ^                                �      �       Q�      >       ]F      �       ]�      �       }��              ]4       T!       ]T!      \!       }�\!      "       ]"      "       }�"      Q"       ]Q"      T"       } p "�T"      �"       ]                                   u �       �        u �       �        ��>"      ["       ��                                                         �             0�      5       P5      >       S�      �       S�      �       R�      �       S�      �       R�              0�4       b        0�b       k        Pk       |        S�       �        S�       �        p ��       !       0��!      �!       S�!      
"       R
"      &"       S&"      >"       Rw"      |"       S�"      �"       S�"      �"       0�                                           �      F       0�F      �       V�      �       V�              0�4       |        0�|       �        V�       T!       0�T!      5"       V<"      t"       Vt"      |"       P|"      �"       V�"      �"       0��"      �"       V�"      �"       0�                                           �      F       1�F      �       \�      �       P�      �       \�              1�4       |        1�|       �        \�       T!       1�T!      �!       \�!      "       \"      �"       \�"      �"       1��"      �"       \�"      �"       1�                           �      �       0��      �       0��             	 p �-)�4       >       	 p �-)�>       b        _�       �        _�"      �"       _                                       �      0       0�0      >       Ye      �       Y�              0�4       n        0�n       |        Y�       �        1��       !       0��!      >"       Y["      s"       Y�"      �"       Y�"      �"       0�                               �      e       0�e      �       T�              0�4       �        0��       �!       0��!      �!       T>"      ["       0�|"      �"       0�                      T!      p!       Q�!      �!       Q|"      �"       Q                    �       �        P>"      ["       P                          �      �       U�      �       \�      �       �U��             \             �U�                    �      �       S�      �       S�             S                    �      �       P�             P                            0       {        Q{       �        [�       �        Q�       �        [�       �        Q�       �       [                          3       ]        X]       �        Y�       �        X�       �        Y�       �        X�       �       Y                           3       �        0��       �        Z�       �        0��       f       Zi      k       Zk      �       0�                         3       Y        0�Y       y       	 s �-)�y       �        x �-)��       �        0��       �        S�       �        0��       �       S                         3       �        0��       �        \�       �        0��       k       \k      �       0�                      ~       �        P�       �        P�       �       P                   �       �        Q�       �       Q                      �              R             XB      k       R                          f      Cf       UCf       g       S g      5g       �U�5g      �i       S�i      j       Uj      xl       S                 f      f       u                     %f      ,g       V5g      xl       V                                   %f      {f       ��{f      �f       \�f       g       \=g      �g       \�g      qh       \qh      |h       ��|h      Oi       \Oi      Ti       7��i      j       ��j      �j       0��j      �j       \                    Df      hf       P�f      �f       P                    %f      {f       0�;i      Ti       ��~�i      j       0�                 �g      h       0�                �g      h       �v                  �g      h       S                 h      qh       A�                      h      .h       z�.h      3h       Z3h      :h       z�                 h      qh       S                      *h      3h       P:h      Lh       Plh      qh       P                  Mh      _h       P                   �f      �f       ��zj      j       0�cl      hl       0�                  �g      �g       P                    �f      �f       Sj      zj       S�j      ik       S                       �f      �f       P�f      �f       ��~j      zj       ��~�j      ik       ��~                    �j      �j       R�j      4k       ��~                  5j      Jj       P                          �f      �f       	��j      (j       	��(j      vj       \vj      zj       |��j      4k       \4k      ik       	��                    j      "j       P4k      Lk       P                  �f      �f       �x  j      j       �x                    �f      �f       Sj      j       S                 4k      Lk       s                     Ti      �i       Sik      cl       Shl      xl       S                       vi      zi       Pzi      �i       ��~ik      cl       ��~hl      xl       ��~                      �k      �k       R�k      <l       ��~hl      xl       ��~                    �i      �i       P�i      �i       P                      vi      �i       	��ik      �k       	���k      7l       \hl      xl       \                    �i      �i       Pik      �k       P                vi      �i       �1z                  vi      �i       S                            �i      �i       P�i      �i       X�k      �k       X�k      <l       ��~<l      bl       Xhl      xl       ��~                      �k      0l       Phl      jl       Pll      xl       P                 ik      �k       s                 i      ;i       �Fv                  i      ;i       S                         )        U                         )        T                         )        R                           %        Q%       )        t �����@$t�����!�                      �      �       U�      �       S�      �       �U�                 �      �       u                       �      �       U�             S             �U�                      �      �       T�             V             �T�                      �      �       Q�             \             �Q�                      �      �       R�             ]             �R�                     �      �       0��      �       P�             Q                      �9      �9       U�9       :       \ :      %:       �U�                      �9      �9       T�9      ":       ]":      %:       �T�                         �9      �9       0��9      �9       p��9      �9       P�9      �9       ^�9      :       P                      �;      �;       U�;      <       ^<      <       �U�<      =       ^                  �;      �;       T�;      =       �T�                      �;      �;       Q�;      <       ]<      <       �Q�<      =       ]                            �;      �;       \�;      �;       U�;      <       \<      J<       \J<      N<       UN<      =       \                     �;      <       V<      <       P<      =       V                                        �;      �;       R�;      
<       �<      -<       R-<      J<       �Y<      y<       Ry<      ~<       �~<      �<       R�<      �<       ��<      �<       R�<      �<       ���<      �<       R�<      �<       ��<      =       R                  �;      �;       sx�<<      J<       sx�                 �<      �<       U                     ;      2;       U2;      �;       T                    D;      t;       Py;      �;       P                    c;      t;       Ry;      �;       R                  ;      2;       U                        �:      �:       U�:      �:       T�:      ;       U;      ;       T                    �:      �:       P;      ;       P                      �:      �:       Q�:      �:       q���;      ;       Q                 �:      �:       U                  d      �       P                    �      �       U�      (       �U�                    �      �       T�      (       �T�                    �      �       Q�      (       �Q�                  �      (       X                  	             U                 	             P                          �      �       U�      �       U�      �       P�      �       u p '��      �       P                  c:      m:       P                 =      �=       U                      4=      I=       QX=      f=       0��=      �=       Q                      =      �=       R�=      �=       R�=      �=       q  $ &4$u"�                      �=      �=       T�=      �=       T�=      �=      	 uz "@�                   �=      �=      	 uy "1��=      �=      	 uy "1�                     ?      B?       UB?      @       [                       ?      E?       TE?      �?       U�?      @       �T�                     ?      I?       XI?      @       �X�                      �?      �?       S���?      �?       S�P��?      �?       �P�                   #?      I?       XI?      W?       �X�                  #?      $?       uȑ                   I?      W?       XW?      W?      
 p x "#���                  I?      W?       x ?&�W?      W?       P                W?      c?       Y                W?      c?       {̑                  W?      c?       Qc?      c?      
 q r "#���                  W?      c?       q ?&�c?      c?       R                �?      �?       r�                    �?      �?       T�?      �?      
 t u "#���                  �?      �?       t ?&��?      �?       U                �?      �?       P                �?      �?       r�                   �?      �?       Q�?      �?      
 q x "#���                  �?      �?       q ?&��?      �?       X                  �?      �?       S�?      �?      
 q s "#���                  �?      �?       s ?&��?      �?       Q                 �?      �?       P                  �?      �?       R�?      �?      
 r t "#���                  �?      �?       r ?&��?      �?       T                  �J      �J       U�                  �J      �J       P                 �J      �J       �k�  �                  �J      �J       ��                  �J      �J       P                  �K      �K       U                  �K      �K       Q                      �K      L       TL      L       �T�L      0L       T                 �K      0L       U                  L      0L       T                  L      0L       U                  L      0L       Q                      0L      IL       TIL      QL       �T�QL      nL       T                 4L      nL       U                  QL      nL       T                  QL      nL       U                  \L      nL       P                        pL      �L       U�L      �L       S�L      �L       �U��L      �L       U                       pL      �L       U�L      �L       S�L      �L       �U��L      �L       U                      zL      �L       U�L      �L       S�L      �L       �U�                  �L      �L       V                              �L       M       U M      LN       VLN      UN       �U�UN      lN       VlN      �N       U�N      �N       V�N      �N       �U�                            �L      _M       T_M      NN       \NN      ]N       �T�]N      �N       T�N      �N       \�N      �N       �T�                              �L      M       QM      N       _N      UN       �Q�UN      lN       _lN      �N       Q�N      �N       _�N      �N       �Q�                              �L      tM       RtM      �M       ���M      FN       ]FN      UN       �R�UN      ]N       ��]N      �N       R�N      �N       ��                            
M      tM       RtM      �M       ���M      FN       ]UN      ]N       ��]N      lN       R�N      �N       ��                          
M      M       QM      FN       _UN      lN       _�N      �N       _�N      �N       �Q�                        
M      FN       \UN      lN       \�N      �N       \�N      �N       �T�                  N      N       0��N      �N       P                       M      5M       S5M      GM      
 s 2%s "#�NM      N       SUN      lN       S�N      �N       S                           M      !M        ~ �!M      tM       YtM      �M       ��UN      ]N       ��]N      lN       Y�N      �N       ��                   hM      N       SUN      ]N       S�N      �N       S                   hM      N       VUN      ]N       V�N      �N       V                      pM      tM       PtM      N       ��UN      ]N       ���N      �N       ��                    pM      �M       ^�M      
N       0�UN      [N       ^�N      �N       ^                 �M      �M       ^                 �M      �M       V                  �M      �M       U                 �M      �M       P                   �M      �M       T�M      �M       v � $ &3$v("�                          �N      �N       Q�N      GO       \GO      NO       �Q�NO      _O       Q_O      ~O       \                          �N      �N       R�N      KO       ^KO      NO       �R�NO      _O       R_O      ~O       ^                      �N      �N       X�N      NO       �X�NO      ~O       X                        �N      �N       Y�N      MO       _MO      NO       �Y�NO      ~O       _                      �N       O       S O      ,O       s~�,O      ;O       S                        �N      �N       S�N      �N       Y�N      IO       ]NO      ~O       Y                      �N      �N       S�N      IO       } 1�NO      ~O       S                   �N      EO       VNO      ~O       V                         �N      �N       Q�N      GO       \GO      NO       �Q�NO      _O       Q_O      ~O       \                         �N      �N       Q�N      GO       \GO      NO       �Q�NO      _O       Q_O      ~O       \                 1O      ;O       \                 cO      ~O       Q                      U      3U       T3U      _U       �T�_U      zU       T                          U      2U       Q2U      ^U       S^U      _U       �Q�_U      nU       QnU      zU       S                     U      4U       0�4U      <U       P_U      zU       0�                   U      ,U       U_U      zU       U                   U      ,U       u��_U      zU       u��                      #U      /U       P_U      gU       PgU      zU       u�#h                AU      YU       w                 AU      YU      	 q  $ &�                        �U      �U       U�U      �U       S�U      �U       �U��U      �U       S                    0]      4]       U4]      W]       �U�                    0]      V]       TV]      W]       �T�                      `]      e]       Ue]      f]       �U�f]      s]       U                      `]      e]       Te]      f]       �T�f]      s]       T                            �]      ^       U^      ^       S^      ^       �U�^      "^       S"^      )^       U)^      *^       �U�                            �]      ^       T^      ^       V^      ^       �T�^      #^       V#^      )^       T)^      *^       �T�                            �]      ^       Q^      ^       \^      ^       �Q�^      %^       \%^      )^       Q)^      *^       �Q�                          �]      ^       \^      ^       �Q�^      %^       \%^      )^       Q)^      *^       �Q�                          �]      ^       V^      ^       �T�^      #^       V#^      )^       T)^      *^       �T�                          �]      ^       S^      ^       �U�^      "^       S"^      )^       U)^      *^       �U�                  ^      )^       P                    0^      V^       TV^      W^       �T�                    `^      v^       Uv^      �^       �U�                    `^      s^       Ts^      �^       �T�                    `^      z^       Qz^      �^       �Q�                   `^      z^       Qz^      �^       �Q�                   `^      s^       Ts^      �^       �T�                   `^      v^       Uv^      �^       �U�                  d^      �^       R                  �^      �^       U                 �^      �^       P                          �^      �^       U�^      1_       S1_      7_       �U�7_      f_       Sf_      �_       U                            �^      �^       T�^      4_       \4_      7_       �T�7_      R_       TR_      f_       \f_      �_       T                            �^      �^       Q�^      6_       ]6_      7_       �Q�7_      G_       QG_      f_       ]f_      �_       Q                     _      ,_       0�E_      G_       0�y_      �_       3�                        �^      �^       U�^      _       S7_      E_       SG_      f_       Sf_      �_       U                      �^      _       V7_      E_       VG_      {_       V{_      �_       u(                  \_      f_       P                 _      ,_       ]                 _      ,_       \                 _      ,_       S                    _      '_       P'_      ,_       �L                 _      ,_       S                 _      _       1�                    �`      �`       U�`      �`       �U�                    �`      �`       T�`      �`       �T�                       a      a       Ua      a       �U�a      a       U                       a      a       Ta      a       �T�a      a       T                       a      6a       U6a      �a       \�a      �a       �U�                       a      .a       T.a      Xa       VXa      �a       �T�                       a      6a       Q6a      _a       S_a      �a       �Q�                  7a      �a       P                  %a      7a       1�                    %a      6a       U6a      7a       \                   ;a      _a       S_a      a       �Q�                   ;a      Xa       VXa      a       �T�                 ;a      a       \                ;a      a       1�                  ;a      _a       S_a      a       �Q�                  ;a      Xa       VXa      a       �T�                ;a      a       \                 Ia      a       T                  ga      xa       U                  ja      xa       R                            �a      �a       U�a      �a       S�a      �a       �U��a      �a       S�a      �a       U�a      �a       �U�                            �a      �a       T�a      �a       V�a      �a       �T��a      �a       V�a      �a       T�a      �a       �T�                            �a      �a       Q�a      �a       \�a      �a       �Q��a      �a       \�a      �a       Q�a      �a       �Q�                          �a      �a       \�a      �a       �Q��a      �a       \�a      �a       Q�a      �a       �Q�                          �a      �a       V�a      �a       �T��a      �a       V�a      �a       T�a      �a       �T�                          �a      �a       S�a      �a       �U��a      �a       S�a      �a       U�a      �a       �U�                  �a      �a       P                        �a       b       U b      "b       �U�"b      9b       U9b      �d       S                        �a       b       T b      "b       �T�"b      ;b       T;b      �d       V                        �a       b       Q b      "b       �Q�"b      +b       Q+b      �d       �Q�                          �a       b       R b      !b       _!b      "b       �R�"b      .b       R.b      �d       _                          �a       b       X b      b       \b      "b       �X�"b      ?b       X?b      �d       \                        �a       b       Y b      "b       �Y�"b      Jb       YJb      �d       �Y�                            bb      c       ]c      Kc      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&�Kc      �c       ]�c      �c      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&��c      ed       ]ed      �d      5 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&�                        �b      �b       Roc      �c       R�c      �c       Rd      d       R                                    nb      �b      	 >u r ��b      �b      + >u O} (  / 0@K$(	 1$#/��O'��b      c      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'�c      Kc       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'�Kc      Uc      	 >u r �Uc      _c      + >r Ov (  / 0@K$(	 1$#/��O'�_c      �c      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'��c      �c       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'��c      ed      M >Ov (  / 0@K$(	 1$#/��O'O} (  / 0@K$(	 1$#/��O'�ed      �d       >Ov (  / 0@K$(	 1$#/��O'O�Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&(  / 0@K$(	 1$#/��O'�                            ;b      �b       TKc      ~c       T~c      �c       p �c      �c       Td      d       Td      :d       �                             ?b      �b       XKc      {c       X{c      �c       p�c      �c       Xd      :d       X:d      �d       ��                         ?b      �b       p�b      �b       � #Kc      �c       p�c      �c       � #d      :d       � #                         ?b      �b       p�b      �b       � #Kc      �c       p�c      �c       � #d      :d       � #                         ?b      �b       p�b      �b       � #Kc      �c       p�c      �c       � #d      :d       � #                         ?b      �b       p�b      �b       � #Kc      �c       p�c      �c       � #d      :d       � #                          Jb      �b       YKc      �c       Y�c      �c       Yd      :d       Y:d      �d       ��                         Jb      �b       p�b      �b       � #Kc      �c       p�c      �c       � #d      :d       � #                     Jb      Qb       QQb      Yb      
 q r "#���Yb      bb       ]                   Jb      Qb       q ?&�Qb      bb       R                    �b      �b       P�b      1c       ��                    �b      c       } p �c      c      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                 Kc      oc       V                 Kc      oc       ]                      Yc      cc       Qcc      kc      
 q r "#���kc      oc       R                     Yc      cc       q ?&�cc      kc       Rkc      oc       q ?&�                    �c      �c       Y�c      �c       w                     �c      �c       } p ��c      �c      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                    6d      :d       R:d      �d       ��                 6d      :d       � #�����                    ;d      ed       } p �ed      yd      8 �Q| " $ &s  $ &�Q| " $ &s  $ &?&"#��@&p �                      �d      �d       U�d      �d       S�d      e       �U�                    �d      �d       T�d      e       �T�                 �d      �d       t ����1$u"�
���                       �d      �d       0��d      �d       s��d      �d       Se      e       s�                      �d      �d       P�d      �d       ^e      e       ^                 �d      �d       U                       e      ,e       U,e      -e       �U�-e      3e       U                       e      ,e       T,e      -e       �T�-e      3e       T                    �e      �e       U�e      f       �U�                    �e      �e       T�e      f       Y                  �e      f       X                         �e      �e       0��e      �e       P�e      �e       0��e      �e       0��e      f       P                        Pm      �m       U�m      �m       X�m      �m       �U��m      �m       U                        Pm      �m       T�m      �m       �T��m      �m       T�m      �m       �T�                      Pm      �m       Q�m      �m       �Q��m      �m       Q                  Pm      om       Q�m      �m       Q                  Pm      om       U�m      �m       U                  �m      �m       Q                  �m      �m       U                  �m      �m       P                    tm      �m       0��m      �m       R                   �m      �m       T�m      �m       T                  tn      �n       ��                  tn      �n       Q                  �n      �n       U                  �n      �n       Q                    �      �       U�      �       �U�                    �      �       T�      �       �T�                  �      �       U                      �       �        U�       y       �U�y      �       U                       �              0�      m       Pt      y       Py      �       0�                          �       �        p��       F       XF      _       0�_      y       Xy      {       p�{      �       t �#�                     �              0�      m       Uy      �       0�                        �              S      9       Y=      B       QB      k       Yy      �       S                        �              Q#      &       R&      Q       Qc      m       Q                      �               Z#      Q       ZQ      c       Qc      t       Z                                 R1      m       R                      @       _        U_       �        �U��       �        U                  D       �        Q                      R       U        q p "�U       �        R�       �        R                  _       �        U                           @       j        0�j       �        X�       �        U�       �        X�       �        U�       �        0�                    j       �        P�       �        P                    �             U      H       ��~                          �      �       T�      7       S7      �       ��~�      �       S�      H       ��~                          �      �       Q�      	       \	      D       �Q�D             \      H       �Q�                    �      �       R�      H       ��~                    �      �       X�      H       ��~                        �      �       Y�      ?       ]?      D       �Y�D      H       ]                        ,      7       0�7      �       SD      �       S�      �       0�                   �      2       V�      H       V                          ,      �       V�      �       vx��      �       VD      �       V�      �       vx��      �       V�      �       vx��      �       V                    �      �       Pt      �       P                      O      [       P[      �       _D      �       _                        [      h       ~�h             ^      �       ~�D      o       ^                       �      �       q��      �       Q�      �       q��      �       Q                                    U       7        �U�                                   U       7        �U�                         7        T                         7        U                                         P       !       	 q ����!       ,        P,       3       	 q ����3       7        t �����                          p      �       U�      �       �U��      �       U�      �       �U��      �       U                   :      @       4�@      n       u r #�                     6      @       0�@      j       Pp      �       P                      :      n       Rn      p       r�p      y       R                     @      n       r n      y       ry      �       X                    H      M       TM      Q       x��Q      �       T                         �      �       6��             T             t�             T$      /       T                       �      �       0��             P      !       P$      /       P                        �             X             x�      !       X$      /       X                     �             x              x$      /       x                       �      �       R�      �       y���      !       R$      /       R                    w      �       U�      �       T                    �      �       0��      �       T                 �      �       T                   �      �       U�      �       �U�                 �      �       0�                 �      �      
 ��G     �                 �      �       T                   �      �       U�      �       �U�                 �      �       0�                 �      �      
 ��G     �                          �      �       U�      l       u�p      t       u�t      y       Uy      �       u��      �       U�      n       u�                            �      l       [p      y       [�      �       R�      �       [�      g       Rg      n       [                              �      l       4�p      y       4��      �       4��      �       z����             z~���             x ��G     "���      0       z���g      n       4�                         �      �       0��      l       Yp      y       Y�      �       Yg      n       Y                           �      �       4��      '       S'      l       R�      �       R�      �       Sg      n       S                                     �      l      
 G     �p      t      
 G     �t      �       Z�      �       z��      �       p��      �       Z�      �      
 G     ��      �       Z�      �       z��      �       z~��      �       P�      g       Qg      n      
 G     �                          �      6       R6      g       Qg      l       R�      �       Qg      n       R                                     �             r 1$ $ &G     "�      6       Z6      X       q 1$ $ &G     "�X      l       Zp      �       Z�      �       P�      �       Z�             z}�             x ��G     "�      :       Z:      I       p ��G     "�I      n       Z                                  '      	 x ��'      ^      F s y "1&1$ $ &G     "�8$
��
��#%!
����G     "���^      g       Pg      l      F s y "1&1$ $ &G     "�8$
��
��#%!
����G     "����      �       Pg      n      	 x ��                  �      0       q ��8$p��!�0      W       q ��8$q��!�                            :       Z:      I       p ��G     "�I      g       Z                    �      �       U�      �       �U�                  �      �       P                            �       �        U�       ^       S^      `       �U�`      r       Sr      t       �U�t      ~       U                        �       �        T�       	       U	      t       �T�t      ~       T                                   P      _       V`      s       V                          0       O        UO       f        �U�f       u        Uu       |        �U�|       �        U                          0       O        TO       f        �T�f       y        Ty       |        �T�|       �        T                              0       O        QO       _        V_       e        Ue       f        �Q�f       r        Qr       |        V|       �        Q                              0       O        RO       Y        SY       e        Qe       f        �R�f       y        Ry       |        S|       �        R                      I       a        \a       e        Rf       |        \                                      U       %        S%       &        �U�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                    �       �        Q�       �        �Q�                    �       �        R�       �        �R�                    �       �        U�       �        �U�                    �       �        T�       �        �T�                      `      �       U�             S             �U�                  �             P                    �      �       �H��      �       Q                                  �      P       UP      C       VC      N       UN      g       �U�g      �       U�      �       V�      �       ���             �U�      �       V                                  �      5       T5      N       SN      g       �T�g      �       S�      9       ��~9             �T�      �       S�      �       �T��      �       S                      �      j       Q�R�n      r       Q�R�C      �       Q�R�                                  �      U       XU      g       �X�g      d       Xd      �       ��~�             �X�      �       X�      �       ��~�      �       �X��      �       X                                  �      U       YU      g       �Y�g      d       Yd      �       ��~�             �Y�      �       Y�      �       ��~�      �       �Y��      �       Y                             8      P       u P      C       v C      N       u g      �       u �      d       v       n       v �      �       v                           �       S�      �       ��~                                         _��      C       _�R��      �       _�R��      �       _���      9       ��~��      �       _���      �       _��                                    y 	����      C       y 	���y	����      d       y 	���y	���      n       y 	���y	����      �       y 	���y	���                       	      U       0�g             0�             ��~      �       0�                           	      U       0�g      �       0��             ��~      �       0��      �       ��~�      �       0�                                 C       _�      �       _�      �        ��~��      9      
 ��~��~�      '       _'      �        ��~��      �        ��~�                        �      C       ^�      �       ^�             ~ ��~�      '       ^'      �       ~ ��~�                             �              u "�              U       C       s�6$���� "��      �        u "��      d       s�6$���� "�      B       s�6$���� "��      �       s�6$���� "�                   �      C       R�      �       R                       �      C       y 	���      �       ]      �       ]�      �       ]                             C       \�      �       \      �       \�      �       \                     	             } z "�      #       Z#      C       p 6$����} "�                 	      C       y	��                   �      �        } -( �      9        } -( �                   �      �       | ~ -( �      9       | ~ -( �                        �      �       Q�             ��~      '       Q'      �       ��~                          �      %       R%      �       ��~      E       RE      �       x�      �       R                   v      �       } 6&��      �       ]                    v      �       | 6&��      �       \            
 ~ ��~6&�                                x      d       x��d      �       ����                    )      0       Q0      z       ��~                         e       0�e      j       ��~                      �      �       Z�             S             T      0       S                    �             [      9       [                  �      9       ]                      J      �       U�      �       w �      �       R                    V      Y       QY      �       ��~                    a      �       Q�      �       ��~                   �      �       w �      �       Z                     �      �       ��~�             R             r|��      �       R                  �      �       V                      �      �       z����             P      D       z���                        r       P                               	 s p ��      r      	 } p ��                       r      	 ~ p ��                       r      	  p ��                          9       Q9      r       �p �                                U      j       r}���                         1       T1      �       r~���                       �       Y                 �      �       Q                              ���                              V                              v                             `      �       U�      �       �U��             U      �       �U��      *       U*      [       �U�                            `      �       T�      	       S	             �T�      �       S�      *       T*      [       S                            `      �       Q�      
       V
             �Q�      �       V�      *       Q*      [       V                                `      �       R�      �       �R��      9       R9             �R�      (       R(      �       �R��      *       R*      [       �R�                     �      �       u �             u              �U                          �      �       \|             \(      �       \�      �       \*      [       \                             �      �       v�      �       X|             X(      �       X�      �       X�      �       X*      [       X                       "      /       0�/      7       Q             Q             r q �      (       P                                      v             p �             q �      %       } �%      N       v��      (       v��                      "      -      	 q �����-      N      	 z �����      (      	 z �����                       �      �       [�      �       {��      �       [�      �       [*      ;       [                       �             \             T      p       t�p      |       T*      ;       \                          �             X             Q      p       qx�p      x       Q�      �       P�      �       p��      �       P*      ;       X                             �      �       q 3%��             P|             q 7�      �       Q�      �       Q*      3       P3      ;       q 3%�                          `       P`      c       U                   �      �       R�      �       R                  �      �       ^                   �      �       ]�      �       }��      �       ]                       �      l       [l      w       {�w      ~       [�      �       [;      K       [                                      \       +       U+      Q       u�Q      \       U;      K       \                                         X       '       Q'      Q       q|�Q      \       Q�      �       Y�      �       y��      �       Y;      K       X                                          p 2%�             Q              p 2%�\      _       p 3�_      e       P�      �       P;      K       Q                    /      >       P>      A       T                   �      �       Q�      �       Q                     �      �       U�      �       u��      �       UK      [       U                         �      �       \�      �       | p "#��      �       | p "��      �       | p "#��      �       | q "�K      [       \                         �      �       X�      �      
 p 1$x "#��      �       p 1$x "��      �      
 p 1$x "#��      �      
 q1$x "#�K      [       X                        �      �       p 1%��      �       QK      S       QS      [       p 1%�                      �      �       r ���      �       q ���      �       | p "���                   <      �       Z�      �       z��      �       Z                     H      W       \W      c      
 t 2$| "#�c      �       t 2$| "��      �      
 t 2$| "#�                     H      W       XW      c       x t "#�c      �       x t "��      �       x t "#�                  K      W       P                 c      �       t 2$| "�                    n      �       U�      �       [                                �      �        r r 
|p p 
�"q q 
m6"@%��      �      4 t 2$| "��t 2$| "��
|p p 
�"q q 
m6"@%��      �      1 t 2$| "��t 2$| "��
|p 
�"q q 
m6"@%��      �      I t 2$| "��t 2$| "��
|p 
�"t 2$| "#��t 2$| "#��
m6"@%��      �      . t 2$| "#��t 2$| "#��
m6p 
�"r "@%��      �      I t 2$| "#��t 2$| "#��
m6t 2$| "#��t 2$| "#��
�"r "@%��      �      * t 2$| "#��t 2$| "#��
�q "r "@%��      �      I t 2$| "#��t 2$| "#��
m6t 2$| "#��t 2$| "#��
�"r "@%�                                            �      "	       U"	      �	       �U��	       
       U 
      �
       V�
      �
       U�
      �
       V�
      a       �U�a      y       Vy      }       U}      �       V�             U             V      ,       U,      Z       VZ      �       �U�                                          �      "	       T"	      �	       �T��	      �
       S�
      �
       T�
      -       S-      a       w a             S      2       �T�2      ?       w ?      g       �T�g      �       S�      �       ���      �       S                            �      �       Q�      !	       �Q�!	      "	       Q"	      �
       �Q��
      �
       Q�
      �       �Q�                            �      �       R�      !	       �R�!	      "	       R"	      �
       �R��
      �
       R�
      �       �R�                            "	      �	       0�!
      /
       P,      6       B�#      2       0�?      Y       0�b      g       0�                      "	      �	       V<      2       VT      Y       V                         "	      /	       Tx	      �	       0��	      �	      	 t q "v ��	      �	       q t "v #��      �       1��      2       T                         "	      F	       XF	      f	       1�f	      �	       U~      �       ~��      2       X                           "	      �	       ��~�#�%      <       s<      ~       ^~      2       ��~�#�G      J       sJ      Y       ^                       "	      �	       w �	      �	       U<      ~       0�~      2       w                                �      	       S	      !	       ��~"	      �
       ��~�
      �
       S�
      �       ��~�      �       P�      �       ��~�      �       ��~                                        �      !	       R"	      �	       ��~�	      �	       R�	      �
       ��~�
      �
       R�
      y       ��~y      �       R�      �       ��~�      �       R�             ��~      #       R%      ,       R,      �       ��~                   �	      �	       ����	      
       Q                     "	      F	       \�      �       u �      2       \                  x	      �	       v t �                                ~
      �
       ��~�
      y       ��~�      �       ��~�             ��~6      #       ��~2      ?       ��~Y      b       ��~g      �       ��~                                ~
      �
       ��~�
      y       ��~�      �       ��~�             ��~6      #       ��~2      ?       ��~Y      b       ��~g      �       ��~                                          ~
      �
       S�
      -       S-      a       w a      y       S�      �       S�             S6             S      #       �T�2      ?       w Y      b       �T�g      �       S�      �       ���      �       S                                      ~
      �
       P�
      �
       ��~�
      y       ��~�      �       P�      �       ��~�      �       P�             ��~6      #       ��~2      ?       ��~Y      b       ��~g      �       ��~                                            �
      �
       _�
             _      a       ^a      y       _�      �       _             _6      �       _�      �       P�      �       ��~2      ?       ^g      �       _�      �       U�      �       ��~�      �       _                                �
             ^t      y       ^�      �       ^             ^6      #       ^Y      \       ^\      b       ~ �g      �       ^                   �
      �
       4�a      y       2��      �       1�             8�                         ~
      �
       \�
             \a      y       \�      �       \�             \6      v       \                            �
      �
       P�
      /       Pa      y       P�      �       P             P6      J       P                                 ~
      �
       0��
      y       0��      �       0��             0�6      Z       0�Z      ^       P^      #       V2      ?       0�Y      b       Vg      �       V                     �
              3$�      a       ~ 3$�2      ?       ~ 3$�                    �
             R             ]                              E       ]E      M       UM      a       ]2      ?       ]                         a       _2      ?       _                           /       R/      a       S2      6       S                         a       \2      ?       \                             /       P/      8       v�8      a       V2      :       V                   >      E       ]E      ^       U                   �      �       ]�      �       ]                         �      �       V�      �       _�      �       U�      �        | "��             _�      �       V                       �      �       s � ����} "��      �       s �p ����} "��      �       s ���~�����} "��      �       s � ����} "�                   s      w       s�      �       ]                         s      w       Uw      �       V�      �       P�      �       S�      �       U�      �       s | "��      �      	 s | " "�                 s      w       s � ����s"�                            @       �        U�       y       �U�y      �       U�      �       �U��             U      Q       �U�                                  @       �        T�       ,       \,      y       �T�y      �       T�      �       �T��      �       T�      �       \�      (       T(      Q       \                                @       �        Q�       5       V5      y       �Q�y      �       Q�      �       �Q��      �       V�             Q      Q       V                      �       �        U�      �       U      ,       U                           �       �        S�       �        s ��       �        t���      �       t���      �       |��      (       t��(      ,       |��                      �       '       ]�      �       ]      Q       ]                        �       x       _y      �       _�      �       _      Q       _                        �       v       ^y      �       ^�      �       ^      Q       ^                     �       �        P�       �        p ��       �        v���      �       v��                    �       �        Q�      �       Q                 �              v                     <      B       PB      K       Vb      f       V                     ,      W       \W      [       T_      r       \                    <      [       Xb      y       X                             1       U1      e       �U�e      v       U                               5       T5      d       Sd      e       �T�e      v       T                   .      1       u 1      9       U                �@     �"@     �"@     #@     #@     8#@     8#@     e#@     f#@     w#@     x#@     �#@     �#@     �$@     �$@     �$@     �$@     �%@     �%@     @&@     @&@     m&@                     W      �      �      �                      \      b      f      h                      �      �      �      �                                                 (      ?      G      K                                    (      ?      G      K                                    (      ?      G      K                      K      O      [      [      [      n                      K      O      [      n                      w      w      w      w            �      �      �                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �                               #      ,      0      @      L      P      V      `      m      �      �                      �      �      �                   0                      �      �      �            8      B                      �      �      �      �                      �	      �	      �	      �	                       
      
      
      
      
      
      #
      *
      1
      9
      A
      E
      I
      L
                       
      
      
      
      
      
      #
      *
      1
      9
      A
      E
                      
      
      
      
      
      
      *
      *
      .
      1
      9
      =
      L
      T
      W
      [
      _
      a
                      
      
      
      
      
      
      *
      *
      .
      1
      9
      =
      L
      T
      W
      [
                      
      
      
      
      =
      @
      E
      I
      g
      v
                      
      
      
      
      =
      @
      E
      I
      g
      s
                      
      #
      *
      .
      I
      I
      T
      W
      [
      _
      v
      �
                      
      #
      *
      .
      I
      I
      T
      W
      [
      _
      v
      �
                                              &      )      4      8      J      M      b      f      t      |      �      �                                              &      )      4      8      J      M      b      f      t      |      �      �                                              &      )      4      8      J      M      b      f      t      |      �      �                            	            "      -      0      8      <      f      i      m      q      �      �      �      �                            	            "      -      0      8      <      f      i      m      q      �      �      �      �                            	            "      -      0      8      <      f      i      m      q      �      �      �      �                                  )      -      <      ?      F      J      U      ]      i      m      q      q                                  )      -      <      ?      F      J      U      ]      i      m      q      q                                  )      -      <      ?      F      J      U      ]      i      m      q      q                                  0      4      C      F      M      Q      ]      b      q      q      �      �      �      �      �      �                                  0      4      C      F      M      Q      ]      b      q      q      �      �      �      �      �      �                                  0      4      C      F      M      Q      ]      b      q      q      �      �      �      �      �      �                      "      &      ?      C      q      q      q      t            �      �      �      �      �      �      �                                  "      &      ?      C      q      q      q      t            �      �      �      �      �      �      �                                  "      &      ?      C      q      q      q      t            �      �      �      �      �      �      �                                  Q      U      �      �      �      �      �      �      �      �      �      �      �      �                      Q      U      �      �      �      �      �      �      �      �      �      �                      q      q      �      �      �      �      �      �      �      �      �      �                                  q      q      �      �      �      �      �      �      �      �      �      �                                  q      q      �      �      �      �      �      �      �      �      �      �                                  �      �      �      �      �      �      �      �      �                                        �      �      �      �      �      �      �                                        `      `      h      r      |            �      �      �      �      �      �      �      �                      `      `      h      r      |            �      �      �      �      �      �                      r      |            �      �      �      �      �      �      �      �      �                      r      |            �      �      �      �      �      �      �                      �      �      P      o             2      �      �                      �            s      �      �      �      9      `                            $      �      �      �      �      x      �      �      �                      '      =      �            `      x      �      �      �                            x      @      H      �                      �      �             @                      �      �      �      �                      �      �      �      �                      �      �      h      �                      �             H      h                      �      �      �      �      �            	                  K                      `      `      i      x      |            �      �                      q      x      |            �      �                      �      �      �                            �      �      �      �                                        ,                      �       �       �       �                       �       �       �       �                       �       �       �       �                       /!      4!      ?!      O!                      K"      N"      U"      _"                      i%      i%      o%      �%      �%      �%      �%      �%      �%      �%                      �%      �%      �%      �%      �%      �%                      A&      F&      M&      ]&                      �&      �&      �&      �&       '      '                      �&      �&      �&      �&       '      '                      �&      �&      �&      �&                      �&      �&      �&       '                      [(      a(      e(      j(                      )      
)      )      )                      �*      �*      �*      +                      �*      �*      +      0+      `+      c+      k+      �+      �+      �+                      �+       ,      @,      �-      �-      �/                      �,      -      �.      �.                      -      /-      �.       /      8/      X/                      w-      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      w-      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      w-      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      z-      }-      �-      �-      �-      �-      �-      �-      �-      �-      �-      �-                      0.      T.      �.      �.                      �/      �/      �/      �/      �/      �/                      I2      _2      g2      k2      o2      r2                      I2      _2      g2      k2                      _2      g2      k2      o2      v2      �2                      _2      g2      k2      o2      v2      �2                      �2      .3      p3      �3                      �2      �2      �3      �3                      �2      3      p3      �3                      �3      �3      �3      �3      4      4      
4      4                      <6      J6      h6      h6                      p7      �7      �7      �7      �7      �7      �7      �7      �7      �7      �7      �7      �7      8                      p7      �7      �7      �7      �7      �7      �7      �7      �7      �7       8      8                      �7      �7      �7      �7                      C8      T8      [8      [8      _8      d8      �8      �8      �8      �8       9      9                      %9      69      :9      J9      K9      k9      p9      �9      �9      �9                      %9      69      :9      ?9      P9      k9      p9      �9      �9      �9                      P9      c9      p9      w9                      �9      �9      �9      �9      �9      �9      �9      �9                      +:      >:      Q:      V:      Z:      _:                      �:      �:      �:      �:      �:      �:      �:      �:                      M;      `;      a;      l;      p;      r;                      ==      _=      `=      f=      i=      p=                      N=      _=      `=      f=      i=      p=                      �=      �=      �=      �=      �=      �=      �=      �=                      �=      �=      �=      �=      �=      �=                      �=      �=      �=       >                      �=      �=      �=       >                      >      >      !>      D>      H>      J>      L>      P>                      2>      D>      H>      J>      L>      P>                      }>      }>      �>      �>      �>      �>      �>      �>                      �>      �>      �>      �>      �>      �>                      9?      U?      `?      p?                      A      >A      HA      HA      JA      MA      YA      �A      �A      �A      �A      �B      �B      �B                      yA      �A      �A      �A      �A      �B      �B      �B                      �A      �A      �A       B                       B      �B      �B      �B                      B      #B      'B      0B      8B      �B      �B      �B                      0B      0B      8B      @B                      GB      �B      �B      �B                      GB      vB      �B      �B                      `B      dB      iB      vB                      �C      �C      �C      ZD      �D      �D                      �D      �D      �D      E                      DF      ^F      mF      �G      �G      ?J      DJ      JJ      QJ      UJ      `J      �J      �J      �J      K      )K                      LG      �G      �G      �G                       H      �H      �J      �J      K      )K                      �H      �H      �H      �H                      I      tI      }I      #J      �J      �J                      5K      zK      �K      �K                      �M      �M      �M      �M      �M      �M                      �N      �N      �N      �N                      �O      �O      �O      �O                      zQ      jS      jS      �S      �S      `T      nT      wT      �T      �T      �T       U                      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R                      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R                      �R      �R      �R      �R      �R      �R      �R      �R      �R      �R                      �R      �R      �R      �R      �R      �R      �R      �R                      qS      zS      �S      �S      �S      �S      �S      �S      �S      �S                      qS      zS      �S      �S      �S      �S      �S      �S      �S      �S                      qS      zS      �S      �S      �S      �S      �S      �S      �S      �S                      zS      }S      �S      �S      �S      �S      �S      �S      �S      �S                      zS      }S      �S      �S      �S      �S      �S      �S      �S      �S                      zS      }S      �S      �S      �S      �S      �S      �S      �S      �S                      �S      �S      �S      T                      �S      �S      �S      T                      �S      �S      �S      T                      8W      `W      �W      �W                      xW      �W      �W      �W                      �X      Y      XY      XY                      RZ      VZ      YZ      pZ      tZ      vZ      �Z      �Z                      �[      �[      �[      �[                      �[      �[      \      \      \      q\      �\      �\      �\      �\       ]      ]                      \      \      \      \      \      )\      �\      �\      �\      �\      �\      �\       ]       ]      ]      ]                      n]      s]      w]      }]                      �_      �_      �_      �_      �b      �b                      �_      �_      �_      �_                      &a      *a      .a      Va      Pb      Zb      ^b      cb                      Za      ja      wa      ~a                      �a      �a      �b      �b                      �a      �a      �b      �b                      b      :b      �b      �b                      �d      �d      �e      �e      �e      �e                      �d      �d      �e      �e      �e      �e                       e      5e      he      e                       e      5e      pe      e                      �f      �f      g      7g      �g      �g      �g       i      6i      �i                       g      7g      i       i      6i      �i                      Gg      Lg      Pg      ^g                      +k      Dk      Ik      Mk      �k      �k      �k      �k                      Mk      jk      �k      �k                      �l      �l      �l      �l                      �m      �m      �m      n                      �n      �n      �n      �n      �n      �n      �n      �n                      /s      @s      `s      fs      hs      xs                      �s      t      	t      t      Dt      It                      t      t      t      "t                      �v      �v      �v      �v                      Ex      �x      y      /y      Py      ty                      y      "y      "y      /y      Py      [y                      �y       z      �z      g{      r{      �{                      P{      T{      ]{      g{                      z      �z      �{      �{                      Zz      �z      �{      �{                      hz      �z      �z      �z                      |      |      |      �|      �|      �|      �|      �|      �|      �|      �|      �|      �|      .}                      �}      ?~      @�      ��                      �}      ~      @�      h�                      ~      ;~      h�      ��                      H~      �~      ��      ��      N�      i�                      Y~      �~      ��      ��      N�      i�                      Y~      ]~      c~      �~      ��      ��                      �~      �~      �~      �~                      �~      �~      �~      �~                      ��      ��      ��      ��                      N�      W�      W�      i�                      �~                        )      @                      �      ��      p�      ��      i�      p�                      �      �      �      �      �      �      i�      p�                      �      �      �      �      i�      p�                      ��      h�      �      N�                      ��      '�      ,�      1�      6�      :�                      �      '�      ,�      1�      6�      :�                      у      ��      ��      ��      ��      ��      �      �      �      �      �      $�                      ��      ��      �      �      �      �      �      $�                      |�      ��      ��      �      �      ��      ��      ��      �      �                      ��      ��       �      �      �      �      X�      c�                      Ç      ч      ��      ��                      ��      ��      ��      ��                      6�      �      0�      5�      ��      ��                      [�      ��      ��      �      ��      ��                      ��      ��      ��      ɋ                      ɋ      ��      ��      �      ��      ��                      ɋ      ��      ��      ��                      ��      �      �      ��                      �      �      0�      5�      ��      ��                      x�      x�      z�      ��                      ��      ��      ��      ��      ��      ��      ��      ͎      ю      �                      ��      ��      ��      ��                      ��      ��      ��      Б      ԑ      ��                      �      �      #�      b�      m�      $�      8�      F�                      {�      $�      8�      F�                      X�      z�      }�      ��                      t�      z�      }�      ��                      h�      ��      �      �      �      �                      �      ��      �      �                      d�      h�      m�      ��      8�      P�                      ��      ��      ��      ��      �      �                      �      )�      ��      ��                      �      )�      ə      ��                      M�      w�      �      �                      U�      w�      �      �                      ��      h�      ��      ��      �      E�      `�      {�      ��      ��      +�      g�                      ��      $�      ��      ��      ��      ��      �      �      �      E�      `�      {�      ��      ��      +�      g�                      ��      �      �      �      ��      ��                      V�      Z�      ^�      ��      ��      ��      �       �      %�      E�                      ��      ̜      ̜      ќ      ؜      ۜ                      )�      D�      ��      ��      �      �      ��      ��                      h�      l�      v�      =�      ��      �      �      ��      E�      `�      {�      ��      ��      +�      g�      ��                      ��      ŝ      �      #�      '�      2�      7�      =�      ��      ��      E�      P�                      @�      c�      ��      Ġ                      z�      ~�      ��      ��                      =�      Y�      �      �      ��      �                      I�      ��      ��      ը                      ��      ��      ģ      ף                      ��      ��      ��       �                      (�      ,�      0�      D�                      Х      L�      d�      ��      ��      �      ��      ӫ                      ��      զ      �      �                      ��      ��      ��      ��                      �      7�      ��      ��      ը      &�      &�      p�      �      b�      t�      ~�                      &�      M�      \�      d�                      M�      \�      d�      y�                      ը      �      �      &�      &�      C�      �      ��      �      b�      t�      ~�                      ��      ��      ũ      �                      &�      &�      &�      4�      9�      C�                      Q�      U�      Y�      c�                      �      ��      ��      ƪ                       �      )�      >�      C�      K�      p�      u�      ��      `�      e�                      p�      p�      u�      ��                      ;�      H�      `�      `�                      ��      ��      ��      ��      ��      í      �      �       �      ��      ��       �       �      �      W�      s�                      8�      b�      f�      j�      ��      ��      ʯ      د                      @�      b�      f�      j�      ��      ��      ʯ      د                      �      �      ��      ʯ                      ��      �      ��      ʯ                      ��      ��      ��      ��                      ˭      ��      �       �      ��      ��       �       �                      ˭      ��      ��      ��                      F�      J�      N�      {�      �      0�                      ��      ð      ʰ      ̰                      �      �      �      h�      ��      Q�                      �      h�      ��      Q�                      "�      $�      ��      Q�                      ��      ��      ��      ۲      
�      �      C�      C�                      ߲      �      �      ��                      b�      g�      ��      �      ��      ô                      ��      �      ��      ô                      ǳ      ɳ      ��      ô                      )�      -�      1�      L�      ��      ��      ��      ��                      P�      Z�      b�      g�                      Դ      ״      ڴ      �      ��      �                      P�      P�      `�      v�      ��      ǵ                      ��      ��      ��      ��                      c       c       g       �                       p      �      �      �                      �      �      �      �                      �      �      �      �                      �      �      (      �      �      �                                                          "      &      *      -      0      4      8      @      H      L                                        "      &      *      -      0      4      8      @      H      O      S                      �      �      �      8                      �      �      �      �      �      �      �      �      �      �                                                           �      �      �      �      �      �      �                                           #                      �!      Z#      b#      p#                      �+      �+      �+      �+                      D.      K.      Y.      `.                      �.      �.      �.      �/                      �.      �.      �.      �.                      A5      A5      H5      N5      T5      f5                      y5      �5      �5      �5                      7      	7      7      �7      �9      �9                      p8      �8      �8      �8      �9      �9                      �9      :      	:      :      :      F:                      �:      �:      �:      �:                      �:      �:      �:      ;                      �@      gB      �B      �B      C      `D      E      #E                      �A      �A      �A      B                      �A      �A      �A      B                      �H      �H      I      I      
I      I      I      )I                      �J      �J      �J      �J                      K      ;K      ?K      FK                      �K      L      L      +L      1L      �L       M      `N                      gN      pN      pN      yN      �N      �N                      O      &O      0O      LO                      �O      �O      �O      HP      `P      lP                      �Q      �Q      �Q      	R                      �Q      �Q       R      	R                      �T      U       U      =U                      �V      W      �W      �W                       W      �W      �W      �W                      SW      SW      YW      \W      _W      bW      eW      iW      mW      pW      sW      wW      {W      �W      �W      �W                      \W      _W      bW      eW      iW      mW      pW      sW      wW      {W      �W      �W      �W      �W                      ~X      <Y      _Y      �Y      �Y      �Y      �Y      �Y                      �X       Y      �Y      �Y      �Y      �Y                      �]      �]      �]      �]      �]      Xa      �a      Mb      �b      �b      +c      �c      td      �d      e      �g                      �]      �]      �]      �]      �]      �]      �e      f      f      �f      �f      �f                      �e      �e      f      f       f      $f      ,f      ?f      Cf      Gf                      $f      ,f      ?f      Cf      Gf      Kf      Nf      af                      �_      �_      �_      `                      �_      �_      �_      �_      �_      �_                      `      �`      e      �e      Vg      �g                      /e      Be      ae      je                      g      �g      �g      �g                      �`      �`      �`      Xa      �f      �f      �f      g                      i      .i      3i      Ji                      �k      �k      �k      
l                      �k      �k      Ql      Xl      \l      `l      il      xl      l      �l                      7l      Ql      Xl      \l                      xl      l      �l      �l      �l      �l                      �m      �o      �q      mr      	t      �|      K}      �}      �}      <~      A~      h�                      �m      �o      �y      �y      z      �|      K}      y}      �}      �}      A~      h�                      �m      �o      �~      �      �      1�      R�      h�                      �m      �n      �n      �n      �n      �n      �n      �n      �n      �n      q      �      R�      h�                      �n      �n      �n      �n      �n      �n      �n      Qo                      z      kz      vz      �|      K}      y}      �}      �}      A~      V~      �      �                      z      \z      �{      �|      K}      y}      �}      �}      �      �                      |      |      #|      '|                      |      #|      '|      +|      .|      A|                      �      �      �      �      �      �      �      �                      �      �      �      �      �      �      �      �                      �q      �q      r      Dr      	t      t                      �t      �x      y}      �}                      �x      y      y       y                      y      y      )y      Gy                      p      �q      ~r      	t      �|      K}      �}      �}                      �p      �q      s      �s      �s      	t      �|      �|      �}      �}                      7q      :q      >q      Uq                      �s      �s      �s      �s                      �|      �|      �|      "}                      �      E�      ��      ,�                      �      �      �      �      "�      9�      <�      @�      ��      ,�                      ��      ��      ��      ��      ��      Á      Ɂ      ́                      ]�      s�      v�      z�      �      ��                      ȃ      �      1�      8�                      Ǆ      ��      �      1�                      g�      ��      �      %�      )�      +�                      ��      ��      ��      ˆ      φ      �      ��      ʇ                      ��      ��      �      0�                      ΍      ��      Ȓ      �                      ��      �      �      O�                      &�      �      ��      �      �      (�      p�      ��      ��      ��                      `�      ��      ږ      �      ��      ��      ��      ��                            K�      \�      `�      ږ       �                      f�      f�      k�      ��                      ��      p�      ��      ݚ      �      5�                      8�      $�      (�      O�      ��      ��                      �      �      2�      <�      <�      H�                       �      �      ,�      m�      q�      v�      0�      H�                      ��      �      $�      0�                      `�      ��      ��      X�      ��      ��       �      �      ܭ      �                      ��      X�      ��      ��       �      �      ܭ      �                      ��      X�      ��      ��       �      �      ܭ      �                      ��      x�       �      �                      ۩      �      �      x�       �      �                      `�      ��      ��      ƫ      Ϋ      Ϋ      Ϋ      ث      �      �      Z�      ��                      ̨      �      &�      E�                      �      :�      ��      ��                      L�      P�      +�      ��      ��      կ                      P�      d�      �      &�                      �      ٬      �      �      ��      ܭ      �      �      ��      ��                      ì      ì      ʮ      J�      `�      ��                      ֱ      ݱ      �      �      �      �      �      K�      R�      |�                      ٲ      e�      i�      x�                      ޲      �      �      �      #�      &�      /�      1�                      ��      "�      #�      )�      *�      .�      0�      2�                      {�      ��      ��      ��      ��      ��                      z�      ��      ��      ��      ö      Ŷ                      �      V�      H�      ��                      Y�      _�      �      �      ��      =�      ù      й      �      #�      ��      л      ��      ̼      �      ��      ��      �      �      �      .�      �      �      ��      ��      ��      ��      ��      ��      	�      �      ;�      @�      y�      ~�      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��      ��                      Y�      _�      ��      q�      ��      ��      ��      �      �      8�      ��      ��                      �      '�      y�      ��                      '�      =�      ��      ��      ��      �      &�      ;�      ��      M�      ��      ��      }�      ��                      ��      M�      }�      ��                      ��      ��      ��      ��      �      �      �      �      �      �      �      �       �      (�      0�      4�                      ��      ��      �      �      �      �      �       �      (�      0�      4�      8�                      �      #�      ;�      ��      Q�      {�                      ��      ̼      8�      ��      M�      ~�                      9�      P�      y�      ��                      P�      `�      ��      ��      ��      p�                      ��      ��      ��      ��                      �      �      �      $�                      ��      ��      V�      y�      ��      �                      ��       �      ��      ��                      �       �      ��      ��                       �      5�      s�      ��                      ��      ��      ��      	�                      ��      ��      -�      ��                      ��      ��      ��      ��                      ��      ��      ��      ��      {�      ��                      ��      ��      �      &�                      ��      �      ~�      ��                      �      ��      ��      ��      ��      ��      ��      ��                      u�      ��      ��      ��                      ��      ��      H�      V�      ��      �      p�      }�                      ��      �      H�      V�                      t�      ��      p�      }�                      ��      ��      ��      ��                      ��      ��      ~�      ��                      '�      �      �      �      ��      ��      �      (�                      �      �      �      ��      ��      ��      �      �                      p�      N�      9�      u�      ��      ��                      ��      ��      V�      ]�      ��      ��                      ��      ��      ]�      u�      ��      ��                      ��      %�      9�      >�      ��      ��                      1�      =�      >�      V�      ��      ��                      ��      ��      �      -�      ��      ��                      ��      ��      ��      ��                      ��      ��      ��      ��                      )�      w�      ��      ��                      �      �      �      �                      q�      ��      '�      1�                      �      ��      ��      �                      ��      �      ��      K�                      �      ��      ��      p�                      ��      N�      @�      y�      p�      ��                      �      ,�      3�      F�                      ]�      '�      ��      ��                      F�      ��      �      H�                      ��      �      K�      ��                      n�      ��      u�      ��                      ��      ��      ��      �      ��      ��                      �      ��      ̼      ޼      �      �      ��      ��                      (�      ��      ̼      ޼      �      �      ��      ��                      m�      ��      �      �                      �      W�      Z�      ��      ��      ��                      }�      :�      @�      ��                      @�      _�      _�      ��      ��      �      ��      ��                      P�      _�      _�      e�      e�      p�      ��      ��      ��      ��                      L�      N�      ��      ��      ��      ��                      ��      ��      ��      ��      ��      �      �      �       �      ��      �      ��      ��      ��                      ��      ��      ��      ��      Q�      ]�      `�      d�      q�      x�      ��      ��      ��      ��      ��      ��                      ��      ��      �      �      )�      ,�      d�      i�      x�      }�      ��      ��      ��      e�      e�      p�      ��      �                      ��      e�      e�      p�                      ��      ��      ��      ��                      W�      �      (�      H�      v�      ��      �       �                      [�      _�      c�      q�      v�      M�      (�      (�      �       �                      ��      ��      
�      �      5�      8�      N�      Z�      d�      l�                      ��      �      �      �      l�      {�      ~�      ��                      �      �      ��      ��                      �      #�      8�      <�      ��      ��                      p�      ��      0�      p�      ��      ��      ��      ��      �      `�      ��      �                      4�      ��      ��      �                      <�      ��      ��      ��                      ��      ��      ��      ��      ��      ��      �      `�                      ��      �      ��      ��                      �      V�      ��      ��                      d�      l�      o�      s�      w�      ��      ��      ��                      l�      o�      s�      w�      ��      ��      ��      ��      ��      ��                      �            0      >                      0      �      0      >                      �      �      �      �                      �      =      P      �                      X      7      �      @      `      u      �      �                      �      �      �      0      �      �                      �      �      �      �                      {      �      �      �                      �      �      �      �                      �      X      �      X                                                               �                  |      �      �                      '!      )!      -!      D!      L!      \!      `!      b!                      �!      �!      �!      ;"      C"      �"      �"      w&                      1"      4"      �#       %      H%      w&                      $       %      H%      t%      w%      w&                      $      )$      /$      D$      D$       %      H%      t%      w%      w&                      �$       %      H%      t%      w%      w&                      �$       %      H%      X%      |%      w&                      �'      �'      �'      �'                      �(      �*      8,      �,                      M)      �*      8,      `,                      �/      ?0      C0      P1      �1      �1                      �/      40      �1      �1                      X4      _4      i4      �4      �4      �4                      5      (5      08      �8                      �:      �:      v>      �>                      ;      P;      R>      v>                      �>      W?      `?      o?                      ?      ?      ?      R?      `?      o?                      �?      6@      `@      �@                      FD      �D      �D      E                      pE      �E      3F      �F                      �E      �E      �E      �E      3F      3F      `F      `F                      �H      �H      �H      5I                      iJ      �J      �K      {M      �M      �M                      �K      sM      �M      �M      �M      �M                      �N      �N      �N      �N      �N      �N      �N      �N                      �N      �N      �N      �N      �N      �N      �N      �N      O      O      O      �O      �P      Q      @Q      `Q      �Q      �Q      �Q      R      hX      �X                      �O      yP      Q      @Q                      1P      AP      MP      yP      Q      @Q                      "R      VU      �W      �W      �W      UX      �Z      }[      �[      �[                      HR      �T      �W      �W      �[      �[                      �W      UX      �Z      }[                      �U      6V      �X      �X                      �W      �W      �X      `Z      }[      �[                      �X      Y      "Y      EY      SY      -Z                      	\      \      \      .\      :\      =\                      �\      �^      X_      �_      �_      `      P`      �`                      	]      `]      �_      �_      p`      �`                       ]      `]      �_      �_      p`      �`                      `^      c^      l^      o^      z^      �^      P`      p`                      �^      B_      `      8`      �`      �`                      �^      B_      `      8`      �`      �`                      b       �       �       �                       �      �      �      �                      �      �      �      �                                                              �             5      I                                        Y                      �      �      �      �      �      �      �      �      �      �                       	      T	      X	      [	      ]	      _	                      �	      �	      �	      �	                      �      #      8      8      <      B      H      J                      p      �      �      �      �      �                                        �      �      �                                  .      J      `      1      1      9      �      �      �      �      �      �                      `      �      �      �      �            �      �                      E      �      �      �      �      �      �      �      �      p                      V      �      �      n      �      p                      �      �      �      �                      �      �      �      �                      �      F      X      ]      `      �                      S      �      �      �                      {      �      �      �                      �      �                                   g      �      �      �      �      �                      �            �                            x      �      �      �                      P      �      �      =      P      ^                      �      �      �      �      �      �                       !!      (!      H!      V!                      "       "      m"       #      #      ##                      5$      B$       *      *                      �$      �$      �$      �$      �(       *      0.      x.      �.      �.                      �(       *      0.      x.      �.      �.                      [%      d%      p%      t%      w%      {%      �%      �%      �%      �%      �%      �%      �%      �&       *      X*      �-      .                      �'      �'      �'      �(                      X*      �-      .      0.                      `+      w+      |+      �+                      w+      |+      �+      �+                      �+      B,      �,      (-                      �,      �,      �,      �,                      `-      �-      �-      �-                      &/      �/      00      �0                      z1      �3      �3      �3                      �1      �1       2      2      2      &2                      2      2      *2      V2      `2      �2                      2      2      *2      22      <2      Q2                      �2      �2      �2      �2                      �2      �2      �2      �2                      �3       4      (4      P4      `4      u4                      �4      �4      �4      �4                      �4      �4      �4      �4                      �4      �4      �4      �4                      �4      �4      �4      5                      �5      �5      
6      x6      �6      �8      �8      �8      �8      �8                      06      x6      �6      �7      �7      8      �8      �8                      �6      �6      7      `7      �7      8      �8      �8                      �9      (:      �:      �:      �:      �:                      �<      �<      �<      �<                      �<      �<      �<      (=      1=      6=                      �=      a?      �?      X@                      �@      �A       B      �B      �B      �C                      �@      "A      LA      �A       B       B      HC      �C                      �@      "A      UA      �A      HC      �C                       B      *B      ,B      gB      mB      �B      C      HC                      �C      �C      �C       D      D      	D                      pD      �D      �D      �D      �D      �D      �D      �D      �D      �D                      �D      �D      E      E      )E      ,E      8E      ;E      VE      �E      �F      �F                      yF      �F      `H      xH                      I      (I      (I      -I      5I      :I                      aI      wI      |I      �I                      �J      �P      Q      �U      +V      pZ      pZ      sZ      �Z      o                      �J      �J      �J      �M      �M      �M      �M      �P      Q      �R      +V      XV      CZ      \Z      G^      �^      �^      o                      �M      �P      �^      �_      Rj      o                      �M      &N      �^      �^      �^      �^      _      �_      Rj      :m      qm      o                      _      �_      Rj      m      qm      o                      �O      �O      �O      fP      :m      qm                      �_      .a      Pa      Rj                      `      `      !`      a      �b      �b      .f      �h      �h      Rj                      �f      ,h      hi      �i                      Pa      Za      ea      �b      �b      �b      �b      �b      �b      .f                      *b      Wb      _b      �b                      �d      �e      f      .f                      �S      �S      �Z      �[                      0T      �T      �T      �U                      jV      �X      �X      �X      �[      :]      W]      G^                      rW      �W      \      6\      W]      2^      ?^      G^                      `]      p]      p]      u]      y]      |]                      |]      2^      ?^      G^                      �]      2^      ?^      G^                      �W      �W      �W      �W                      X       X      "X      %X      -X      2X      5X      uX                      �[      \      \      
\                      �\      1]      1]      :]                      �X      �X      �X      CZ      �Z      �Z      �[      �[      :]      W]                      �Y      CZ      �[      �[      :]      W]                      v      �      �            �      @                      �      �      �      �                                        .      �      �      8      �                      @      �      �                                         �      �                                         D      L      L      �      �                      �	      �      �      �      �      �                      P
      g
      k
      o
                      g
      k
      u
      �
                      �
      �      �      �                                        &                            u      u      �                            K      `      i                            H      �                    &      0      �             �%                            �      �      �      �             �      �      0      �             �%                                  <      H      V      V                            $      +      .      H      Q      V      �      �      �      @      �      �            �      �      �      �      +       5       �       �                       �      �      @      �      +       5                       �      �      @      �      �      �      +       5                             �                  �      �      0      �      �       �       �       	!      $      H$      W$      i$                                  "      �      0      �      �       �       �       	!      $      H$      W$      i$                                  "      0      0      �      0      �      �       �       �       	!      $      H$      W$      i$                      {      �      �       �       �       	!      $      H$      W$      i$                      �      �      �       �       �       	!      $      H$      W$      i$                      �      �      �      �      �      �      �       �       �       	!      $      H$      W$      i$                             �      �       �       �       	!      $      H$      W$      i$                      A      �      �       �       �       	!      $      H$      W$      W$      _$      i$                      �       �       _$      i$                      |      �      �      @             �             +       5       R       �       �       H$      M$                            p             +                       /      �      �      �                      8!      $      M$      W$      i$      %      (%      �%                      �!      $      M$      W$      i$      w$      ,%      v%      �%      �%                      �!      -"      �%      �%                      �"      �"      M$      W$                            �      �      �             H      �             �      �                      `      �             H      �      �                             G       P       U                       {       �       �       �                       �       �       �       U      Y      �      �      �                      /      6      B      n      �      �                      �      �      �      �                      �      �      �      	                            %      (      d                      9	      �	       
      =
                      �      �      �      �                      :      C      P      e      u      y      }      �                      �      �      �      �      `      �      0      M      M      p      �      0      �      9      A      �                      M      M      M      �      u      }                      �      �      �      �                      �      �      �                  p      �      9      A      u      }      �                      �                  p      �      9      A      u      }      �                      #      H      L      Z      �      p                      3      �            9                      �                        A      h      }      }                      �                                        �      �      �      	      	      `      �      0      p      �      0      h      h      k      u      �      9      A      �      �                      �      �      �      �      �      	      	      `      �      �             0      p      �      9      A      �      �                      �      �      {      �      9      A                      	      	      	      h                      �      �      �      �      �      `      �      �             0      p      �                            �      0      h      h      k                      z      �      �      �                      �      �      �      �                      0      7      I      i      p      x                      �                  ?      `      p                      x      {            �                      �      �      �      �      �      �                      �      �      �      �      �      �                      `      `      p      %      �%      �&                      �      �      �      �      �      �      �      �      �      &      (      /      8      G      L      `      �             *%      K%                      !      &      (      +      =      @      L      �      �      `      �      �      *%      K%                      ~      �      �                            &      `      �      �                      p      �             *%      K%      %      �%      �&                      �       Z!      �#      *%                      F"      f#      K%      v%      �%      �&                      �"      �"      �"      �"      �"      f#      K%      v%      �%      &      &      &      &      �&                      �"      f#      K%      v%                      �&      �&      �&      o(                      '      '      '      F(      M(      b(                      (      	(      (      F(      M(      X(                      �(      �(      �(      �(      �(      �(      �(      �(                      &)      �)      �,      �,                      &)      �)      �,      �,                      �)      �)      �)      �+      �+      �,      �,      �,                      a*      f*      l*      �+      �+      �,      �,      �,                      �+      �+      �+      ,                      �,      �,      �,      �,      �,      H/      2      �2      �2      5      *5      �5                      a.      /      2      �2                      n.      �.      �.      /      2      �2                      �3      5      �5      �5                      W4      �4      �4      5      �5      �5                      5      5      *5      �5      �5      �5      �5      �5                      P5      m5      s5      �5                      T/      2      �2      �2      �2      �2                      n/      �/      �2      �2                      �0      �0      �0      �0      1      1      1      01                      H1      �1      �2      �2                      �      �      �      �      �      �                      n      z      �      q      �      �      �      �       	      

      
      "
                      �            
      "
                      �            V      �                      b      �      �      �                      X      �      �      �      0      4      H      @      P      s                            ;      p            V      s                      �      �      �                              v      z      �      �      �                      �      �      �      �      �      �      �      �      �      �                      �                  �      �      �             �              @       �       �$      �$      �%                      �                               #                      @      �      X      �                      �      �      X      �                      �      �      �      J             �      �      �                      h$      �$      �$      9%                      �      �      �       Q!      �!      p"      9%      N%      [%      �%                             �      �      �      �       J!      �!      p"      9%      N%      [%      �%                      5      x      �!      p"      9%      N%      [%      �%                      �!      p"      9%      N%      [%      �%                      �!      �!      �!      p"      9%      N%      [%      �%                      �!      �!      �!      +"      /"      7"      ;"      >"      E"      Z"      9%      N%      [%      �%                      #      h$      �$      �$      N%      [%                      "#      P#      X#      |#      �#      h$                      B      �      �      �      �$      �$                      �      �      �      �      �      %                      	      �      @       �                       �                  @      �      �      �      A                      �                                                     a      h      l      w      �      �      �      �      �      �      �      	      
      �
      �
      �      �      %      5      �                      �      		      
      �
      �
      �      �            5      �                      
      �
      �      �      �      ,                      
      �
      �
      �
      �
      �
      �                                                    �
      �      �      �      ,            5      �                      �      `                  0	      
      �
      �
                      J      R      Z      �      0	      P	                      k      �      �      �                      �      �      �      �                      �      �                                  �      �      �      �                                        !                      �	      �	      �	      
                                        $      @      :      �      �      �      �      �      �      �             &!      /!                      �      T      �      �                      �      A      �      �                      $      *      �      (      @      f      �      �      �                  �      �      �             �                       $      *      �      �            �      �      �             m                             <      @      f      �      �                      �      8      @      f                      �      +      @      f                      �      (      m       �                       ^      �      P      `      �      m      �      �                  �      �                    �       &!                      �      �      �                  m      �       !                      �      .      J      ]      @      P                      ]      #      `      x      �      )      }      }                      /      @      x      �      )      j      �      �      f      }                      �            )      @      x      �                      j      �      �      �      �      �      �       �                       T!      `!      g!      l!                      `!      g!      l!      !      P#      k#                      �!      �"      �"      #                      �"      �"      �"      #                      �"      �"      �"      �"                      0      :      ?      f      p      �                      �      �      �      �      0      @      @      D      H      N                      �      �      �      �                      	      `      p      u      y      {      �      �                      '      P      T      \                             C      �      �                      H      X      b      j      �      �             �      �      )      �       !      0#      @#      (%      =%                      �      �      �      �      �      �      �      �      �      �      �            (      �             �      �       !      0#      @#      (%      =%                      �      �                   (%      =%                      �      �      �      �      �      �      �      �                      U      �       !      #      #      $#      @#      �#      �#      (%      =%      �&                      i      �      �"      �"      H$      P$                      �      �      �       �       !      @!      �!      �"                      �      �      �      �                      �      �      �      �                      M      �      �       �                       x      �      �       �                             �      @!      �!      @#      �#      �#      H$      P$      (%      p&      �&                      w            �      �                      �"      #      #      $#      =%      p&      �&      �&                      �"      �"      �"      �"                      �"      �"      �"      �"                      �"      #      #      $#                      `%      p&      �&      �&                      :&      j&      �&      �&                      �)      �)      �)      \*      �*      �*      +      �+                      �)      *      !*      H*      +      8+      �+      �+      �+      �+      �+      �+                      -      -      *-      �-                      �.      �.      �.      �.                      0      =0      A0      �0      �3      �3      �3      �3      �3      r4                      H0      H0      K0      f0      i0      n0                      g1      i1      m1      |1                      W5      n5      |5      5                      �6      �6      /=      I=      u@      }@                      =      &=      m@      u@                      �>      �?      �?      �?      `@      m@                            :      p      �                      Z      �      �      �                      �      �      �                         *      �                      !      &      ,      /      1      4      6      U      ^                  
                  $      1                      b      o      �      �      �      �      �      �      �      �      (      v      w      {      �      �                      b      o      (      Y      d      v      w      {      �      �                      �      �      �      �      �      �                      �      �      �      �                      |      $	      x	      B
      h
      |
                      V      �      �      �      �      �                      �                              �      H      Q      Y      d      �      �      �            !      :      d      �                            �      �      �      �      �                      �      �      �      �      ~      �                      �            N      �                      �      /      Y      �                      F      L      Q      �      �      �                      �      _      g      �                      �            (      <                      `      �      �      4                       `      o      t      y      |      �      �      �      �      �      �      0                       `      o      t      y      |      �      �      �      �      �      �      �      �      0                       *!      6!      9!      =!      C!       "      ,"      /"      P"      �"                      *!      /!      9!      =!      C!      P!      �!       "      P"      �"      �"      �"                      �!       "      �"      �"                      �!      "      �"      �"                      P"      �"      �"      �"                      X"      �"      �"      �"      �"      �"                      `$      �$      �%      �%                      �$      �%      �%      �%                      �&      �&      �&      �&      �&      �&      �&      �&      �&      �'      �'      0(      @(      v(                      5)      p)      w)      �)      �)      �*                      +      +      +      G+                      �+      ,      	,      s,                      �,      4-      /      �/                      �,      0-      /      �/                      P-      a-      h-      �-      �-      �.      �.      �.      �.      /                      �0      �0      �0      �0                      31      �1      �1      �1                      75      75      A5      p5      �5      �5                      7      s8      w8      �8      �8      �8      �8      �8      �8      �8      �8      o9      �9      �9                      	7      7      7      @7      o8      o8                      P:      T:      Y:      �:      �:      �:                      �B      �B      �D      �D                      �B      �B      �B      �B                      "C      )C      0C      <C      CC      NC                      {I      K      XK      �K                      L      L      L      %L      0L      PL                      nN      `O      �R      �R                      �N      �N      �N      IO                      `O      P      NR      �R                      �O      �O      �O      �O      NR      QR      SR      �R                      dP      vP      vP      �P      �P      �P      �P      �P      �P      (Q      �Q      NR      �R      �S                      Q      (Q      �Q      �Q      �Q      NR      �R      �S                      
R      FR      �R      �R                      �R      tS      ~S      �S                      (Q      wQ      |Q      Q      �Q      �Q                      {U      :W      5Z      LZ                      �W      �W      �W      �X      �X      �X                      �Z      [      �\      h]                       [      �[      \      �\      h]      �]                      {^      B_      �a      �a                      �_      �`      �a      �a                      �`      Ha      `a      �a                      �b      �c      �c      �c       e      Je                      jd      qd      td      �d                      �f      �f      �f      �f      �f      �f                      �g      �g      
h      �i      �i      j                      �g      �g      �h      �i      �i      j                      Ti      �i      �i      j                      >j      Ij      Oj      �j                      m       n       p      p      (p      �r      s      _t      jt      �t      0u      wu      v      Iv                      �m      �m      �m      �m                      n       n       p      p                      hp      �p      �r      �r      �t      �t                      tp      zp      �p      �p      �r      �r                      �p      �p      �p      �p                      �p      �r      0u      @u                       q      �r      0u      @u                      �q      �q      �q      �q      �q      �r                      �n      �n      �n      Ho                      �v      w      	w      ;w                      vw      7x      Ux      �x                      x      7x      Ux      bx      �x      �x                      �y      z      �~                             kz      �}      �}      �}      p~      �~                      �|      �|      �|      P}                      ��      ��      ��      ��      ��      ��      ȁ      ��                      ��      ��      ��      ��      ȁ      ��                      ��      ��      �      ��      ȁ      ��      �      ��                      �      �      0�      h�                      ��      ��      Љ      0�                      ؆      �      ��      ��      Ї      ��      ��      ��      Љ      0�                      t�      ��      Ї      F�       �      0�                      Ї      ه      �      3�      7�      <�                      S�      ��      ��      p�      ��      ��      Љ       �                      ��      �      ��      p�      ��      ��      ��      ��                      4�      4�      5�      L�                      t�      t�      u�      ��                      ��      ڋ      ڋ      �                      ��      �      �      �      �      ��      ��      ��      �      ^�                      ��      q�      O�      W�                      q�      ��      W�      W�      ��      ��                      ��      �      �      �      �      ��      W�      ��      �      ^�                      �      �      �      ~�      ��      ��                      �      �      �      �      Ď      ��                      ��      ��      ��      �                      ��      ��      ��      ʏ                      ��      �      p�      ��                      0�      c�      ��      ��                      ��      ��      ��      ��                      ��      ��      ȓ      �      $�      *�                      �      ��       �      �                      P�      j�      z�      �      З      ��                      �      ��      ��      З      ��      ��      ��      �                      h�      ��      ��      ��      ��      ��                       �      p�      ��      ��                      8�      8�      <�      K�      M�      R�                      ��      Z�      ^�      i�      o�      x�      x�      z�                      ��      ř      ͙      ԙ                      �      �      �      �      0�      ��      �      ��      ��      ��      ��       �      H�      h�      d�      ��      ��      ��      ˧      ˪                      �      �      k�      ��      0�      ��      ��      ��      H�      h�      d�      ��      ˧      ˪                      �      �      ��      ��      ��      �      ��      ��                      �      �      ��      ��      ��      �                      q�      ��      �      �      �      �      �      �      �      �      �      "�      H�      h�                      ��      �      �      ��      �      x�                      Ħ      U�      Z�      ��                      �      �      �      �      ��      �      ��      ��                      �      ��      �      �      ��      ��      8�      H�      h�      @�      ��      ˧                      w�      y�      )�      ]�      ��      ��      ��      ˧                      ī      ��      ��      ��      ��      ��      @�      O�      ��      ��                      ��      @�      X�      ��                      Y�      p�      0�      `�                      ��      `�      c�      p�                      p�      ��      ��      0�      ��      �      h�      p�      ��      �                      δ      ��      ��      0�      ��      �      h�      p�      ��      �                      δ      �      ��      �      �      е      ��      0�      ��      �      h�      p�      ��      �                      ��      ��      `�      ��      #�      W�                      ��      ��      `�      ˹      й      �      �      �      �      ��      @�      ��      #�      W�                      ��      ��      `�      �      @�      ��                      4�      6�      8�      8�      :�      =�      @�      B�      D�      J�      P�      R�      T�      W�      Z�      \�      ^�      d�      z�      |�      ~�      ��      ��      ��                      8�      :�      =�      @�      B�      D�      J�      P�      R�      T�      W�      Z�      \�      ^�      j�      p�      |�      ~�      ��      ��      ��      ��                      d�      j�      p�      z�      ��      ��      ��      ��                      ��      ��      ��      ��      ��      ˹                      �      h�      p�      ��      �      #�                      
                         .      .      1      J                      h      u      �      R                      �      �      �      �      �      �                      �      �      �      �      �      �                      �      �      �      �                      �      �      )      �                      �      �      4      p                      �      �            
                      ?      N      R      c      f      �                      �      �      	      	      	      	      	      "	                      e	      �	      �	      �	                      e	      �	      �	      �	      �	      �	                      �
      �      M      l      {      �                      �
      �
                              "      /      6      9      C      �      {      �                      �      �      �      �      {      �                                                    0                                  >      Q                      M      l      �                                  &      +                   #      (      Q      �      �                            &      �      �            �             #      (      Q                      o      �      �      �      (      Q                      #      8      U      �      �      �                      �      �      V      �                      Q      t      |      %      @      P                                  Q      t      �      �      �      �      (      d      d      �      �      %      @      P            �                      Q      j      o      t      �      �      �      6      h      �             %      @      P      (      �                      Q      j      o      t      �                        &      *             %      @      P      (      �      �      �                      �      �      �                            �      �      �            '      ,      3      \      ^      �                            /       @       s!                      &      "       @       s!                      &      @      �             �       s!                      �      �      i!      s!                      �             !      `!                      �      �      �                             "      (#      H#      U#                      "      "      "      2"      6"      :"                      :"      ="      B"      F"      W"      j"                      F"      H"      K"      O"      x"      z"      z"      �"                      �"      (#      H#      U#                      �"      �"      �"      �"      �"      #                      e$      m$      r$      r$      z$      �$      �$      �$                      �$      �$      �$      !&      �(      �(                      �$      �$      �$      �$      ~%      �%      �%      !&                      j&      �&      �&      �&                      �&      k(      �(      �(                      0'      \(      i(      k(      �(      �(                      H'      �'      �'      0(      i(      k(      �(      �(                      �'      �'      (      (      i(      k(      �(      �(      �(      �(                      m)      �)      h*      �*      �,      R-                      p*      �*      �,      R-                      p*      p*      x*      �*      �*      �*      �*      �*                      -      -      -      -      -      3-                      �)      �)      �)      *                      !*      !*      +*      D*                      (+      �+      �+      O,      �,      �,                      (+      �+      ,      O,      �,      �,                      �+      �+      �+      �+      �+      �+      �+      �+      �+      �+                      �+      �+      �+      �+      �+      �+      �+      �+      �+      �+      ,      ,                      �+      �+      �+      �+      �+      �+      �+      �+      �+      �+                      �.      �.      �.      M/      N/      T/      W/      ]/                      t0      �0       1      51                      w4      �4       6      7                      �4      �4      h6      �6                      �4      �4      z6      �6                      5      @5      x5      �5      �5       6                      �7      �7      �7      �7      �7      U8                      U8      �:      �:      }?                      U8      �:      �:      3;      ?      (?      h?      }?                       9      09      39      �9                      �9      �:      ?      (?      h?      }?                      h:      �:      ?      (?                      h:      q:      z:      �:      ?      (?                      �:      �:      3;      ?      (?      h?                      �:      �:      =      p>                      �:      �:      �:      �:      �=      p>                      �:      �:      �=      
>      >      `>                      �:      �:      �=      �=      �=      >      .>      `>                      �=      �=      P>      `>                      �;      �;      �;      �;                      �;      
=      p>      ?                      �;      �;       <      3<      B<      �<                       <      3<      o<      �<                      �<      �<      �<      �<                      @@      P@      x@      x@      z@      �@                      A       A      �A      �A       B      �B      �B      �C      �C      �C                       B      B       C      @C      �C      �C                      ?D      ?D      CD      eD                      G      G      uG      �I                      
J      J      J      J      !J      +J      TJ      \J                      J      J      +J      8J      =J      HJ      \J      \J                      LJ      TJ      \J      iL      �L      `V                      �J      �J      K      K      S      JS                      K      iL      �L      �L      �L      �L      =O      =O                      �K      L      8L      iL      �L      �L                      �M      =O      �T      �U                      �M      �M      �M      �M      �M      �M      �M      �M                      �M      �M      �M      �M                      �N      �N      �T      �T                      �N      �N      �N      �N      O      
O      
O      O                      U       U      6U      HU                      �O      XR      @V      `V                      �P      �P      �P      �P      �P      Q                      sQ      xQ      �Q      �Q      �Q      �Q      �Q      �Q                      XR      �R       V       V                      pS      |S      �S      �S      �S      �S      �S      �S                      T      �T      �U      �U                      �U       V       V      @V                      iL      iL      qL      �L                      �X      �X      Y      Y                      <Y      @Y      �Y      �Y                      @Y      EY      XY      �Y      �Y      �[                      @Y      EY       Z      X[                      �[      �[      �[      �[                      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\                      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\      �\                      Y]      }]      P_      p_      |_      �_                      �]      y^      �^      �^      @_      P_                      C^      C^      I^      Y^      Y^      a^      d^      h^                      �^      �^      �^      �^      �^      �^                      �^      �^      �^      �^      �^      _                      �_      �_      	`      (a      6a      :a      Pa      �a      �a      ch                      D`      I`      Q`      {`      �`      (a      �a       d      d      d      d      @d      �e      �e      f      �f      �f      hg      pg      ch                      �`      �`      �`      (a      �g      �g                      �`      a      a      "a                      �a      �a      �a      �a      �a      b      !b      �b      �b      �b      �c      �c      f      xf                      �a      �a      �a      b      b      b                      8f      Ff      Of      df      hf      of                      c       c      �f       g      8g      hg      �g      ch                      2c      6c      9c      =c      Ac      Ec      Hc      Lc                      }c      �c      �c       d      pg      �g      �g      �g                      @d      �d      e      `e      �e      f      �f      �f      hg      pg                      Xd      �d      e      `e                      e      e      e      `e                      �e      �e      �e      �e                      �e      �e      �e      �e                      �h      Nk      hk      �k      �k      �k      �k      �v                      �h      �h      �k      �m      �u      �u                      �h      �h      l      �m      �u      �u                      �h      �h      �l      �m                      �h      �h      �l      �m                      �h      �h      6m      �m                      'l      *l      /l      Cl      xl      xl                      i      !i      )i      �j      �m      �m      �m      �n       o      �q       r      @t      `t      �u      av      �v      �v      �v                      pi      `j       o      p      8p      �p      �s       t       u      0u      �v      �v                      �i      `j       o      �o      8p      �p       u      0u                      �o      p      �s       t      �v      �v                      n      on      |n      �n      p      8p      0u      Pu                      n      3n      p       p      0u      >u                      �p      �p      `t      u      �u      �u      av      �v                      �p      �q      8r      �s       t      @t      Pu      �u                      9q      9q      `r      �r      0s      �s      Pu      �u                      �j      k      �q       r      @t      `t      �v      �v                      mk      rk      uk      �k      �n      �n      �n      �n      �n      �n                      �k      �k      �k      �k      �k      �k      �k      �k                      �k      �k      �k      �k      �k      �k                      v      v      v      av                      0v      5v      9v      Pv                       w      Bw      x      Xx      �x      �x                      �w      �w      �w      x      �x      �x                      �x      �x      �x      �x      �x      �x      �x      �x                      �x      �x      �x      Ey      Ey      /{      2{      Z{      o{      �{                      �y      �y      �y      �y                      �y      �z      �{      �{                      -z      5z      8z      @z      �{      �{                      �z      /{      2{      Z{      o{      �{                       |      �}      �}      i�                      @|      z}      �}      :~      �      �      b�      i�                      �|      �|      �|      g}      �}      :~                      �|      ,}      @}      \}      �}      :~                      ŀ      �      �      "�      9�      ;�                      "�      )�      C�      C�      T�      _�      b�      g�                      _�      b�      g�      ł      ł      ��      ��      ڄ      �      @�                      %�      -�      A�      T�                      k�      *�      �      @�                      ��      ��      ��      ��      �      @�                      @�      ��      ��      ڄ      �      �                      ��      �      $�      6�      9�      v�       �      ��      ��      Ր      &�      �                      ܅      �      $�      6�      9�      J�       �      �      1�      ��      ��      Ր      &�      �                      j�      �      �      �       �      {�      ��      �      1�      ��      ��      Ր      &�      �                      ��      ̆      �      Ň                      Ɔ      Ɇ      �      l�      ��      Ň                      Ї      Ї      �       �      '�      {�      ��      ܋      1�      ��      ��      Ր      &�      �                      ��      �      1�      ��      ��      Ր      &�      �                      F�      ��      ��      Ր      &�      �                      Վ      W�      [�      ��      ��      Ր      &�      �                      �      6�      9�      ��      Ր      &�                      �      6�      9�      ��                      0�      6�      9�      k�      s�      ��                      Ր      ��      ��      �                      ��      G�      G�      T�                      ޒ      1�      5�      @�      P�      T�                             "       '       +       .       g       �       �                       >       K       N       Q       V       c                             H      L      \                                        1                      �      �      �      7                      !      >      P      i                      z      z            d      l      �                      �      �      �      �                      �                                                                                          !      %      ?      K                                        !      %      8                      �      �      �      7                      �      �      E      r      u      �                        ,                      �      �      P      P      ]      r      u      y      �      �      �      �                      �      �            ,                      �      �      �      �                      �      	      "	      #	                      P	      S	      a	      �	      �	      -
      1
      4
      H
      �                      �	      �	      H
            p      �                      P
      r
      p      �                      �
      �
      �      �                      �	      -
      1
      4
                      	
      -
      1
      4
                      ~      �      �      �      �      �                      �      s      |      �      �      �                            f      |      �                      x      |      �      �                      @      G      G      e      g      z                      �      �      �      �      �                            �      �      �      �      �                            �      �      �      �                      C      �      �            0      �      �      �                      u      �      �      �      �      �                      �      �      0      �                      �                   %                      �      �            0      0      �      �      �                      �            �      �      �      �      �      P                      �            �      �      �      �      �      P                      �            �      �      �      3      �      P                      �                   @                      p      p      t      �      �      �                      t      w      z      �                      �      �      �      �                            �      �      F                            W      W      ]                      W      W      ]      b      e      �      �      �             %                      e      l      p      �      �      �      �      �                      �      �      �      �      �                  
                                  �      �      �      �      �      �                         +      @      3!      H!      :#                      �      �      �      �                                   �      �      {      �      �      �        "      �"      �"      �"                      �                  �      �!      �!      �"      �"      �"      :#                      �      �      �!      �!                      �      �      �      �      �      �      �      �                                        p      $#      :#                      p      u      y      �                      B#      D#      G#      J#      Y#      \#      a#      n#      r#      #      �#      �#       $      �)       4      @4      g5      o5      �7      8                      \$      d$      s$      %      g5      o5                      �$      �$      �$      %      g5      o5                      %      ('      �7      8                      N%       &      6&      ('      �7      8                      s%      �%       '      ('                      �%      �%      �&      �&      �&      �&      �7      �7      �7      �7                      5'      @'      H'      �'      �7      �7                      �'      0)       4      @4                      �'      �'      �'      0)       4      @4                      �)       4      @4      g5      o5      �7      8      B8                      �)      �)      �)      �)      �)      �)      �)      �)      �)      �)                      y*      ~*      �*      �*      06      �7                      y*      ~*      �*      �*      =6      �7                      %+      y+      �,      h-      �-      �-      05      g5      o5      �5                      2+      @+      �,      h-                      U+      p+      �-      �-      05      g5      o5      �5                      �+      �,      �-      .      �4      5                      `,      `,      d,      g,      p,      �,                      ..      �.      @4      i4      5      05                      ..      N.      [.      �.      @4      i4      5      05                      ..      N.      d.      �.      @4      i4      5      05                      ..      @.      �.      �.      �.      �.                      �.      �0      i4      �4      �5      6      8      78                      y/      �/      �/      �/                      �/      �/      (0      �0      i4      �4      �5      6      8      78                      �0      �0      �5      6      8      78                      i4      i4      k4      �4                      �5      �5      �5      �5                      �0      �1      02      �3      78      B8                      &1      �1      02      �3      78      B8                      &1      81      B2      .3      @3      p3      78      B8                      &1      81      �2      �2      �2      �2                      �2      �2      3      3      @3      P3                      r3      v3      z3      �3                      �8      �8      �8      (:      H:      �:                      �8      �8      �8      %:      H:      �:                      9       :      H:      a:      u:      �:                      49      >9      A9      G9      M9      P9      V9      Z9      f9      i9      �9      �9                      49      >9      A9      G9      M9      P9      V9      Z9      f9      i9      �9      �9                      >9      A9      G9      J9      P9      V9      Z9      f9      i9      l9      r9      u9      �9      �9                      >9      A9      G9      J9      P9      V9      Z9      f9      i9      l9      r9      u9      �9      �9                      J9      M9      l9      r9      u9      �9      �9      �9                      J9      M9      l9      r9      u9      �9      �9      �9                      �:      �:      �:      �:      �:      *;                      �:      �:      �:      �:      �:      �:                      �:      �:      �:      �:                      �:      �:      �:      ;                      G;      G;      \;      �;                      �;      3<      H<      e<                      �;      �;      H<      ]<                      �;      �;      �;      3<                      �<      �<      �<      �<      �<      �<                      �<      �<      �<      �<      �<      �<                      =      =      =      /=      H=      �=                      =      =      =      /=      H=      �=                                  
      U                      3      6      6      ?                      �            �      �                      �      �      �	      �	                      �                  O                      �      �      �                        -      �      0      `      x      @      (      3      B"      P"      �"      �"                      P      �      0      `      x      j             @      B"      P"      �"      �"                      \      _      u      �      0      `      x      �      B"      P"      �"      �"                      \      _      u      �      �      �      0      `      x      �      B"      P"      �"      �"                      �            0      X      �"      �"                      R      U      X      [                      �      '      >      �                                   (      3                      �      �      �                             ^      (      n      B"      P"      X"                      ^      ^      k      t                      }      }      �      �                      �      
      �!      �!                      �      �      �       �       "      "                      &      U      �!      �!      ("      B"                      b      �      �!      �!                      �      �      �       !      �!      "                      �      �      �      �                      +       [       "      ("                      C$      �%       &      J&                      E$      $       &      J&                      �       0      6      W                      �      �      �      �      0      H      M      T      e      o      o      �      �      �                      �      �      �      �      �      �                      �      �      �      �      �      t      �      �                      	      
      �
      �                      (      �      ;      �                      �      �      �      ?                      �      0      3      7      ;      ?                      �	      �	      �	      �	                      `
      d
      h
      v
                      �      �      �      �      �            p      v      �      �                      �      �      �      �      �      0      �                    `       f       \"      f"      �#      �#      E$      E$      �$      �$      B)                      �            �      �      �      �      �                  0             *       f       s       �       �       #"      \"      f"      s"      f#      �#      �#      �#      Y%      �%      �%      �%      �%      �%      2&      �&      �&      �&      �'      �'      �(      �(      ,)      B)                      �      �      �      �      s"      T#      $      2$      J'      �'                      N      a      ~      )      %      "%      &      $&                      �      �      �      �      �      �      �       �       �       �!      �&      '      �'      �(                      �      �      �      �      �      #      �       �       �       �       �       �       !      !      !      �!      �'      �(                      (      1      ;      @      T      T      Y      �      �      �      �      �      �&      �&                      2$      E$      E$      E$      E$      e$      p$      �$      '      1'      �(      !)                      2$      E$      E$      e$      p$      �$      �(      �(                      _)      f)      �)      �)      �)      K*      `*      �*      �*      �*      �*      �*      �*      �*                      _)      f)      �)      �)      �)      8*      `*      �*      �*      �*      �*      �*                      &+      [+      ^+      e+      p+      �+                      0+      [+      ^+      e+      p+      �+                      �+      �+      P,      �,                      K-      �-      �.      �.      /      /                      �-      .      P.      �.      �.      	/      /      �/                      �-      	.      P.      s.      �.      �.                      �.      �.      �.      	/      /      �/                      /      +/      1/      y/                      �       >      �      �                                                    %      )      �      �      �                      `      �      �      �                      �      �      �      $                      �      �      �      �      �      �                      8      k      �      �      	      	      �	      �	      �	      �	                      �      �      �	      �	                      �      	      	      �	                      �	      |
      �
      �                      K
      R
      R
      |
      �      �                      K
      R
      �      �                      �
      �
      �
      �
                      �
      �
      �
      �
                                        �      �      �                                        0                      P      r            �      �      �                      �                   �                      �      �      �      �             ^                      x      {      �      �      �      �                      `	      
      
      
                      �	      �	      �	      �	                      @
      @
      N
      R
      U
      Z
                      |
      �
      �
      �
      �
      K      �      �      �      �                      �
      �
      �
            !      )                      �      �            ,      P      x                      k      p      �      �      �      �                      `      `      d      �                      �      �      �      �                            4      9      |      �      �            &      +      4      8      �                      1      4      9      |      #      &      +      4      �      �                      �      y      �      �                      W      W      [      w                      I      I      �      �      �      �                      �      �      {      e      p      t                                  3      7      9      G      G      O      Q      U                                  #      1                      g      x      i      x                      �      �      �      �                                        \                             
                                    +      P      �      �      �                      /      /      1      B                      �       �       @"      T"                      !      J!      X!      \!      m!      �!      �"      �"                      0#      �#      �#      �#      �#      �#       $      $                       $       $      '$      +$      1$      6$                      �$      0%      P%      �&       '      �(      �(       )      p)      �)                      �$      �$      P%      q&      p)      �)                      �$      �$      �$      �$      &      S&                      0'      h'      m'      r'      �(       )      �)      �)                      �'      @(      �(      �(                       )      :)      J)      P)      _)      p)                       +       +      ;+      D+                      "+      %+      D+      G+      K+      ,      ,      e,                      �+      �+      �+       ,      (,      0,      @,      `,                      p,      p,      w,      �,                      �,      -      -      ;-                      �-      Q.      `.      `.                      q.      t.      �.      �.      �/      �/                      �.      �.      �.      �.      �/      �/                      "/      (/      (/      (/      )/      +/                      N/      T/      U/      o/                      8      $8      ,8      K8      O8      Q8                      �8      �8      �8      �8      �9      �9                      �8      �8      �8      �8                      �:      �:      �:      �:      �:       ;      ;      ;                       ;      #;      &;      2;                      <;      @;      H;      x;      �;      �;                      �;      �;       <      0<      <<      =                      f=      �=      �=      �=                      R>      [>      a>      �>                      #?      #?      $?      '?      *?      1?      E?      I?      M?      P?      S?      W?      W?      _?      c?      f?      n?      r?                      4?      7?      8?      ??      I?      M?      P?      S?      W?      W?      _?      c?      f?      n?      r?      v?                      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?      �?      �?      @      @                      �@      �@      �@      A      ;A      �A      �F      rG      rG      �G      �I      
J      
J      J      J      �J                      �F      �F      �F      �F      �F      �F      �F      �F                      �F      �F      �F      �F      %G      %G                       J      J      
J      J      �J      �J      �J      �J                      �A      �A      �G      �G                      �A      �A      �G      �G                      &B      .B      8B      PB      {B      �B                      �B      C      {C      �C      �C      	E      	E      �E      �E      �F      H       H      �I      �I                      �B      	C      {C      �C      H      H                      �C      �C      �C      �D      �E      �F      �I      �I                      �C      �C      �C      �D       F      iF      pF      �F      �I      �I                      �C      �C      �I      �I                      uD      uD      �I      �I                      E      0E      4E      `E                      C      C       C      2C      6C      GC                      @H      GH      cH      �H                      qH      qH      sH      �H                      �H      �H      �H      �H                      I      I      )I      II      LI      pI                      zL      zL      ~L      �L                      �L      FN      XN      pN      �N      �N                      M      N      XN      pN      �N      �N                      SM      hM      hM      
N      N      N      XN      `N      �N      �N                      �N      �N      �N      �N      �N      �N                      �N      �N       O      ,O                      �O      dP      R      �S      �S      �S      U      U                      .P      2P      6P      9P      <P      @P      DP      LP      TP      XP                      2P      6P      9P      <P      @P      DP      LP      TP      XP      \P                      R      R      2R      6R      :R      =R      @R      DR      HR      PR      XR      \R                      6R      :R      =R      @R      DR      HR      PR      XR      \R      `R                      qR      sR      }R      �R      �R      �R                      �U      �U      �U       V      V      V      �V      �V                      QY      _Y      cY      cY      hY      tY      zY      }Y      �Y      �Y      �Y      �Y                      �[      \      �\      �\                      �]      �]      �]      �]      �]      �]                      �]      ^      ^      !^      %^      *^                      �^      �^      �^      _      @_      E_      P_      p_      t_      y_                      �_      �_      �_      �_      �_      &`                      �_      �_      �_      �_      &`      3`      7`      i`      �`      �`                      .`      3`      7`      ``                      �_      �_      i`      v`      z`      �`                      q`      v`      z`      �`                      %a      %a      )a      .a      2a      7a                      �a      �a      �a      �a      �a      �a                      +b      1b      3b      6b      ?b      Cb      Jb      Yb      ^b      bb                      Pc      Sc      Uc      Yc      \c      oc                      �d      �d      �d      �d      �d      �d      �d      �d                      �d      �d      �d      �d                      �f      �f      8g      �i      j      "j      (j      xl                      �f      �f      �g      �g      Xi      �i      j      "j      (j      �j      �j      xl                      �f      �f      j      "j      (j      zj      �j      ik                      �f      �f      �f      �f      j      j                      >j      zj      �j      4k                      �f      �f      Xi      �i      ik      cl      hl      xl                      \i      qi      vi      �i                      �i      �i      �k      cl      hl      xl                      �i      �i      �k      3l      hl      xl                      �g      �h      �j      �j                      h      qh      qh      �h      �j      �j                       h      qh      qh      �h      �j      �j                      �l      �l      �l      m                      Pm      om      �m      �m                      �m      �m      �m      �m                      n      n      n      'n      Dn      Mn      Sn      Xn                      n      n      n      #n                      �n       o      6o      >o      �o      �o      �p      �q      �q      xr      }r      �r      �r      �r      �r      �r                      �p      �p      �p      q      "q      2q      Rq      Yq      �q      �q                      q      q      2q      :q      cq      jq      �q      �q                      q      q      :q      Bq      nq      uq      �q      �q                      "q      "q      uq      �q                       o      o      "o      )o      Ho      Ho      ns      ps      �s      �s      �s      �s                      Ho      Po      �o      �o      �o      �o                      �o      �o      �o      Ep                      �o      �o      Ep      �p                      �o      �o      �p      �p                      xr      }r      �r      �r      �r      �r      �r      �r                      �r      Cs      Ls      Ps      P�      Y�      _�      d�                      Cs      Ls      Ps      bs      ��      Є                      �s      �s      �t      �t                      �t      �t      �|      �|                      �t      �t      �t      4u      Du      Pu                      4u      Du      Pu      yu      �u      �u                      yu      �u      �u      �u      �u      �u                      �u      �u      �u      v                      �v      �v      Ѕ       �                      �v      �v      Ѕ      �                      �v      �v      �       �                      �v      �v      w      �w                      w      �w      �w      �w                      �v      w      ��      ��      ��      ��      �      0�                      �v      w      ��      ��                      ؀      W�      d�      ��      �      0�                      �w      qx      }x      �x                      �x      �y      �      �      n�      u�                      {      �{      �{      |                      {      ${      ={      L{      [{      f{      r{      �{                      1{      ={      L{      X{      f{      r{      �{      �{                      |      �|      w�      r�      ��      ��      ��      ��                      w�      i�      ��      ��                      |�      ��      ��      ��      ��      ��      ��      ��                      ��      ��      ��      O�      ��      ��                      ��      ��      �      �                      &�      O�      ��      ��                      �|      �|      �      P�      @�      ��      ��      Ѕ      	�      7�      G�      ��      |�      ��      ,�      g�       �      {�      ��      #�                      �|      �|      8�      �      ��      �      �      >�                      O�      O�      �      �                      c�      ��      ��      ѐ                      ~�      ��      ��      ��      ��      ��                      ђ      �      �      ��            �      �      �                      �      ��      �      �                      H�      M�      Q�      c�                      o�      ��      �      �                      E�      E�      T�      `�                      E�      T�      l�      v�      ~�      ��                      �      P�            ��      ؏      ��                      �      �      �      �      �      �      �      ��                      +�      C�      F�      M�      T�      T�      �      �                      @�      b�      ��      Ѕ                      �      2�      G�      R�                      ,�      g�      '�      /�                      H�      g�      '�      /�                      �      �      �      ,�      /�      5�                      <�      ��      �      �                      ܗ      �      '�      [�      `�      ��                      Ù      ˙      ϙ      
�                      ��      ��      ��      ��                      ݛ      ��      T�      ^�                      �      >�      ^�      r�                      ��      ��      ��      ��      ŝ      �                      ,}      ,}      A}      M}                      ,}      1}      5}      A}      Y}      �}                      �}      �}      �}      ~                      H~      �~      8      A                      L~      W~      Z~      \~                      p~      �~      �~      �~      �~      �~                      ��      �      (�      _�      d�      q�      ��      χ      ��      Ӌ                      
�      A�      D�      Q�                      �      �      �      8�                      ��      ��      ��      �      ��      χ      ��      Ӌ                      �      '�      O�      w�                      H�      �      u�      |�      �      O�                      H�      T�      T�      W�                      �       �      7�      G�                      ��      
�      7�      G�                      ;�      ;�      =�      `�                      y�      ��      ��      ��                      ��      ��      ��      ��                      ��      n�      Ӌ      ,�      g�      t�                      ��      ��      �      ,�                      ��      ݈      ��      �                      ݈      ��      �      ��                      ��      �      Ӌ      �                      t�      ��      ��      ��                      ��      ƌ      {�      ��                      w�      �      ��      ��                      }�      ��      ��      ,�      ,�      H�      H�      ��      ��      ҥ      ҥ      ��      ��      ��      Ц      ��      `�      �       �       �       �      ��                      ��      ��      ̞      ڞ      ��      �      ȣ      ��                      ��      �      ��      ��      ��      ��                      �      ,�      ,�      H�      H�      ȣ       �      ��      ��      ҥ      ҥ      ��      ��      ��      Ц      ��      `�       �      X�      ��      ��      �       �       �       �       �      0�      ��                      �      ��      ��      �      �      ,�      ,�      H�      H�      ȣ       �      ��      ��      ҥ      ҥ      �      Ц      ��      `�       �      p�      ��      ��      �       �       �      0�      ��                      ��      ȣ       �      ��      ��      ҥ      ҥ      �      Ц      p�      `�       �      p�      ة      ��      �       �       �      0�      ��                      *�      1�      A�      K�                      ��      ��      ��      ʡ                      ��      �      !�      6�                      T�      a�      a�      ��      ��      ȣ       �      ��      ��      ҥ      ҥ      �      Ц      p�      p�      ة      Ъ      �       �       �                      n�      s�      ��      �                      �      �      �      ��                      Ȥ      -�      Ц      J�      h�      p�                      y�      y�      ��      ��      ��      ��      ��      ��      ��      ǫ                      �      �      �      �                      Ĩ      Ψ      Ԩ       �      ��      ��      ª      Ъ                      ة      �      �      �      �      ��                      �      %�      )�      0�      7�      `�                      W       e       p       }       �       �                       �       �       �       �             Q      R      _      h      t      y      �                      �      g      �      �      g      n                      w      �      �      �      !      $                      �      �      !      #                      �      �      �      �      �      !      $      0                      �            	                            @      j      n      p                      ,      2      H      H                      @      �      H      �                      h      �      H      h      k      o                      �      �      �      �      �      �                      �       �       �      �                      �       j      8      Q                      �      �            s            0      �      �                      �             P      [                      �      �      P      [                      �      �      �             @      P                             s      �             @      P                      �      �      �      �      0      @                      �      �      �      �      0      @                      �      �      �                            �      �      �      �      �      �                      (	      /	      S      ~      �      ?                      �	      �	      �	      
                      e
      l
      p
      r
      v
      y
      ~
      �
      �
      y      �      �      �      �      �      �      �      �      �      �      �            ,      #      Y      b      g      �                      �      �      �                            �      ~      �      �                      �      �      �      9                                        !      *      �                      j      �      �      �                                                    X@                   h@                   @@                   p@                   p@                   p	@                   �	@                   �@                  	 �F                  
  �F                   ��H                    `i                   `i                   `i                   (`i                   xai                   �bi                   �ti                                                                                                                                                                                                                                             ��                     `i                  `i             (     0�H             ;     �@             =     �@             P     @             f     �ti            u     �ti            �     �@             �     �ti     0           ��                �     `i             �     �\I             �     ��F             �    ��                �     i"@     >           �"@               ��                !   ��                0   ��                8   ��                D   ��                Q   ��                Z    �ui            h    �ui            t    �ui            �   ��                �     �B@             �     !C@             �     mC@             �     wC@             �     �C@             �     �C@                ��                   ��                   
 ��F     �       0   ��                n    pF@     1       �y    �F@     H       9     G@            J    G@     k       V    �G@     X       c    �G@     z       x    `H@     /       �    �H@     �       �    @I@            �    `I@     #       �    �I@     �       �   
  �F     �           pJ@     �       $    pK@     \       ;    �K@     7      J    M@     �       p    �M@           �    �N@     �       �    PO@           �    pP@     �       �     Q@     >       �    @Q@     <           �Q@     �       $     R@     (       8    PR@     -       O    �R@     m       h    �b@     #       �    �g@     }       �    pl@           �     �@     \       �   
 �F     �       �    �@     y          `�@     &           ��@     &       :    ��@     �       Q    ��@     D       i    ж@     D       |     �@     �       �    ��@     �       �    0�@     �       �    ��@     �       �    `�@     �            �@     �       7    ��@           A    P�@     >      M    0�@     �      [    ��@           �    ��@     F      �     �@     C	      �   ��                �    P�@     3       �    ��@     �       �    0 A     �       �    � A     �           �A     �      $    `A            :    �A            P    �A            ]    �A            f    �A            p    �A            y    �A     G       �    0A     M       �    �A            �    �A            �    �A     (       �    �A     \      �    0	A     8       �    p	A     8       �    �	A            �    �	A            �    �	A     �          �A     +          �A     �            �A     �       )   
  �F            7    0A     �      @    A     �      K    �A     !       X     A     
       g    A            v     A     �       �    A     9      �    PA     S       �    �A            �    �A     �       �    �A     �      �    �A           �    �A     �       	    @A     �       	    �A     �       ,	    �A            9	    �A     �       Z	    � A     	      h	    �"A     W       s	    0#A     7      �	    p(A     �      �	    P+A     i      �	    �/A     R       �	     0A     	       �	    00A     �      �	     2A     x      �	    �3A     �       
     4A     G       
    P4A     0       3
    �4A     9       F
    �4A     &       ]
    �4A     �      r
    �9A            
    �9A           �
    �:A           �
    =A     y      �
    �DA           �
    �EA     
      �
    �JA     7      �
    �MA     /            NA     |           �NA           (    �OA     f       9    0PA     ]       S    �PA     �       _    `QA     7       m    �QA     <       �    �QA     :       �     RA     7       �    `RA     7       �    �RA     P       �    �RA     U       �    PSA     �       �    �SA     �       �    �TA     �      �    PWA     �           YA     �      5    gA     �      I    �A     �      i    ��A           q    ��A     �       �    ��A     �      �    `�A     ?      �   
  �F     $       �   
  �F             �    ��A     �      �   
 ��F     $       �    ��A     c          �A     �           �A           -     �A           =    0�A     �      [    �A     �      i    ��A     u
      v   
 �F           �   
 `�F     p      �    0�A     7       �    p�A     l      �    �A           �     �A     
       �    �A            �     �A     b          
  �F     p           ��A     ~           �A     R       7    p�A     �       A   
  �F            P    �A     5      _    P�A     ,	      m    ��A     �       {   
 �F     `       �   
 ��F     @       �   
 ��F            �   
 ��F            �   
 @�F            �   ��                C    ��A     )           ��A                ��A     O       *     B            ?      B            U    0 B            l    P B     n       �    � B     �       �    �B     �       �    `B            �    �B            �    �B     �       �    0B            �    @B     x       �    �B                �B     M            B     =      B    `B     Q       Q    �B     !      h    �B     T      x    P	B     �      �     B           �     B     �      �    �B           �    �B     P       �    0B           �     PB     �      �    @B     �      �    0B     Q          � B     p            !B     �      (   
 ��F     �      4     &B     n       A    p&B     &      �     �'B     �      X    @.B     :      d    �1B     �       r    @2B     P      �     �3B     
       �   
  �F     �       �    �3B     �       �    p4B     �	      �     >B     %       *Y    P>B     �       �     ?B           �     @B     �       �    �@B     �           �AB     �          �CB           '    �DB     �      8    PFB     c       J    �FB     1       Z     GB            l    GB     <       �    PGB     C       �    �GB     H       �    �GB     9       �    0HB     �       �    �HB     y      �    `MB     �       �     NB     ~      �    �[B     �         
 `�F               
 p�F            *   
 ��F     (       =   
 ��F            S   
 ��F            f   
  �F     `          ��                �    ``B            �    �`B     	       �    �`B            �    �`B     ;       �    �`B     V            wB                PaB            4    paB            O    �aB     3       _    �aB     
       v    �aB     !       �    bB     A       �    `bB     
       �    pbB     
       �    �bB     
       �    �bB     
       �    �bB     
           �bB     
           �bB     
       )    �bB     
       :    �bB     	       N    �bB     
       a     cB     �       s    �cB            �   
  �F            �    �cB     �       �    �dB     
       �    �dB            �    �dB            �    �dB     x       �    peB                �eB     (           �eB     �       *    pfB     T       8    �fB     �      N    `hB     a       ]    �hB     ~       o    PiB     o           �iB     �      �   
  �F     P       �    �mB     
      �    �nB     �       �    �oB     ;       �    �oB     �      �    �rB           
    �vB     K       #    @wB     �       /    �wB     6      D    0yB            Z    PzB     D       |    �zB     �       �    �{B     �       �    0|B     D      �    �}B     >      �    �~B     Q       �     B     �      �     �B     �           ��B     �          ��B     Z       $    ��B     W       8    P�B     �
      F     �B     V       U    `�B     �      f    �B     �           ��B     �      �    @�B     �       �   
 ��F     P       �    ��B     �       �    ��B     N       �    ЕB     T      �   
  �F     �	      �    0�B     �          ��B     G       #    0�B     /       6    `�B     ^       H    ��B     m       b    0�B     j       y    ��B           �    ��B     E      �    �B     Y       �   
  �F     �       �    p�B     �       �    0�B     �      �    0�B     ?&      �   
 ��F               
  �F     �         
  �F            0   
 ��F     L      C   
  �F     �       \   
 `�F     `       v   
  �F     @       �   
  �F     (       �   
 ��F            �   
 0�F            �   
 ��F            �   
 ��F               
 ��F               
 ��F     (       /   ��                :    p�B     I       Q    ��B            a    ��B            o    ��B     x           `�B            �    p�B            �    ��B     O       �    ��B            �    ��B     .       �     �B            �    0�B     
       
    @�B     M           ��B            '    ��B     �      ;    `�B     �      I    P�B     �      _    ��B     
      n    ��B     
       �   
 ��F     `       �     �B     <       �    @�B     4       �    ��B     Y       �    ��B     9       �     �B     �      �   
 ��F     �	      �   
 ��F               
 ��F     (       $   
 P�F            9   
 @�F            P   ��                V    �B     V       d    p�B            r    ��B     h       �    ��B     �       �    ��B     5       �    ��B     #      �    �B     �       �    ��B     �      �    ��B     �            �B     [           ��B     �      ;    P�B     u       W    ��B     �       i    � C     
       y   
 ��F     0       �    � C     �       �    pC     �       �     C     t       �    �C     �       �    0C     �      �    �C     '      �    �C     �          �C     J         
 ��F     t       -   
 @�F     P       F   
 �F            ^   ��                g    �*C            |     +C     O       �    P+C            �    `+C            �    p+C            �    �+C            �    �+C     t       �     ,C     t            �,C                 �,C     Q       -     -C     6       ;     P-C     �      I     0/C     /       Y     `/C     �       l      0C           |      5C     0      �     P6C     
       �    
 `�F     P       �     `6C     %       �     �6C            �     �6C     
      �     �;C     �      �     p@C     �      !    0CC     6       !    pCC           )!   
 ��F     �      6!   
 ��F            M!   
 ��F            f!   
 ��F     (       z!   ��                �!    �PC             �!    �PC            �!    �PC     /       �!    �PC            �!    QC     L       �!    `QC     q      �!    �SC     l       �!    PTC     
       
"   
  �F     0       "    `TC     �       +"     UC     �       9"   
 ��F     �       N"    �UC     k      \"   
 @�F     P       o"   
  �F            �"   
  �F            �"   
 ��F     4       �"   
 ��F             �"   
 ��F             �"   
 `�F            �"   
 @�F            #    @aC     A       !#   
 0�F            4#   ��                :#    �aC            H#    �aC     	       V#    �aC     c       j#     bC     �       }#    �bC            �#     cC            �#    cC            �#     cC            �#    0cC            �#    @cC     N       �#    �cC     �       �#    �dC     -      $    �gC     �       $    phC     
       .$   
 @�F     @       ;$    �hC     �      P$     jC            ^$    @jC     h       w$    �jC     U       �$    kC     �       �$   
  �F             �$   
  �F             �$   
 ��F            �$    �kC     �      �$   
  �F     4       �$   
 ��F     4       %    �mC     ?      "%   
 `�F            1%   
 @�F            B%   
 ��F            V%   
 ��F            n%   
 ��F            }%   
 `�F            �%    ��C     E      �%   
 ��F     P       �%   
 ��F            �%   
 ��F            �%   ��                �%    �C     �       �%   
  �F             �%   
  �F     �       �%    ��C     �       �%    ��C            &    ІC            &    ��C             #&     �C            1&     �C     {       E&    ��C     �       X&    p�C            k&    ��C     G       {&    ��C     �      �&    ��C     �       �&    �C     6       �&    P�C     �       �&    ��C     
       �&   
 @�F     0       �&    ��C     y       �&    p�C     g       '    ��C     �       '    ��C     @      ''    ��C     �       5'    ��C     G      E'   
 ��F            K'    �C     4       h'    0�C     �       }'    �C           �'   
 ��F     �      �'     �C     �      �'    �C     �      �'   
 ��F     P       �'    �C     �       �'    p�C     I       (    ��C     $      #(    ��C     I      5(   
 ��F             =(   
 ��F            I(   
 p�F            Y(   ��                `(    ��C     �       o(    p�C     "       �(   
 pG            �(    ��C            �(    ��C     �       �(    p�C            �(    ��C            �(    ��C            �(    ��C     3       �(     �C     $       
)    0�C     `       !)    ��C     �       5)    0�C     ]      H)    ��C     $       Z)    ��C     (       h)    ��C     '      {)     �C     W      �)    ��C     �      �)    `�C     P      �)    ��C     :       �)    ��C     $       �)     �C     I       �)    p�C     �       *    @�C     $       *    p�C     e       .*    ��C     �       A*    ��C            S*     �C     3       h*    @�C     �       |*    ��C            �*    �C            �*    0�C     	      �*    @�C     !      �*    p�C            �*    ��C            �*    ��C            �*    ��C     �       +    `�C     	      '+    p�C            <+    ��C            O+    ��C     !       ^+    ��C            s+    ��C     	       �+     �C            �+     �C     �       �+    ��C     �       �+    ��C     �       �+     �C     �       	,    ��C     x       &,    0�C     6       ;,    `YD     ?       M,    p�C            h,    ��C            �,    ��C            �,    ��C     i      �,     �C     �       �,    ��C           �,    ��C     �       �,    ��C     -      -    ��C     �      2-    `�C     
       E-   
 �G     `       S-    p�C     E      e-    ��C     /       w-    ��C     V       �-    P�C           �-    p�C     t       �-    ��C     u       �-    p�C     �      �-     �C     �       �-    ��C     �       .    ��C     X       .    �C     �       5.    ��C     �       P.    ��C     P      h.    ��C           �.    � D     �       �.    �D     B      �.    �D     �      �.    `D     G       �.    �D     G       �.     D           �.    D     
      /     D     �      /     D     )       #/    PD     1       2/    �D     (       G/    �D     �      Y/    �D     =      k/    �D     �       |/    �D     (      �/    �D     K      �/    D     -      �/    @ D     )      �/    p#D     
       0    �#D     �      0    �'D     J       &0   
 �G     D       70    �'D     Z      I0   
 �G            `0   
 �G            x0   
 �G            �0    0+D     J       �0   
 `G     ,       �0    �+D     �       �0   
 @G            �0   
  G     <       �0    p,D     t       1   
 �
G     L       1    �,D           11   
 �G     P       A1     0D     g      P1   
  
G     �       b1    p<D     v      t1    �>D     	      �1     ED     �       �1    �ED     �      �1    �HD     �       �1    `ID     j      �1    �JD     2      �1    LD           �1    0PD     V       2    �PD     U       2    �PD     ?       -2    0QD     ?       A2    pQD     \       S2    �QD     n      c2    @WD     Q      ~2    �XD     &       �2    �XD     �       �2    �YD     r       �2     ZD     �      �2   
 �G            �2   
 �G            3    �]D     B       !3   
 @G     T       43    @^D            F3    P^D            X3    `^D     �       i3   
 �G     �       y3   
 �G            �3   
 `G            �3   
 PG            �3    `_D     K      �3   
 �	G     <       �3   
 �	G            �3    �pD     �       4    pqD           &4    �uD           D4    �vD     1      `4    �wD     G
      q4   
 `G            {4   
 �G     0      �4   
 �G            �4   
 XG            �4   
 �G            �4   
 @G            �4   
 PG            �4   ��                5    @�D     �      5     �D            :5     �D     �      Z5    ��D     �       l5    p�D     w       ~5    p�D     w       �5    ��D     3       �5    0�D            �5    @�D            �5    P�D            �5    p�D     �      6     �D     �       %6    ��D     H       86    @�D            K6    P�D     �      g6   
 �G            y6     �D     m      �6    ��D     �	      �6    ��D     x      �6     �D     �      �6    ��D     �      7    ��D     X       7     �D            .7    �D     5      K7    P�D     U      f7    ��D     <       }7    �D     "      �7     �D     }       �7    ��D     
       �7   
 �)G             �7    ��D     �      �7    ��D     \      �7    �D     Q       8    @�D           68    P�D     I       Q8    ��D     K       f8    �D     �      �8    ��D           �8    ��D     P      �8    0�D     �      �8    ��D     ?      �8    0�D     p      9    ��D     f       (9    �D     �      89    ��D     4      H9    0�D     �      g9    ��D     �      z9    ��D            �9    ��D     =      �9    ��D            �9     �D     �      �9    �E     �       �9    �E     `       :    �E     e       ':    `E            D:    �E     �      `:    PE     O      v:   
 �)G            �:   ��                �:    �E     �       �:    �E     �       �:    PE     �      �:     E            �:    0E            ;    @E            #;    PE     9       1;    �E     9       ?;    �E     �       N;    0E     �      ^;    P)E     Q       r;    @,E     u       �;    (E     V       �;    PNE           �;    `$E     �       �;    p(E     �       �;    �RE     �       �;    `RE     �       �;    �E     m       �;    0E     �       
<    �E     C      .<    E     �      W<    �!E     #      s<    �#E     �       �<    %E     t       �<    �%E     Q       �<    �%E     �      �<    �'E     �       �<    �)E     �      �<    �,E     f      =    0.E     �      +=    �2E     z      :=     9E           Q=    pPE     �       `=     QE     4      {=   
 �eG            �=   ��                �=    �SE     �       �=    pTE     �       �=    UE     �       �=    �UE     d       �=    `VE     �       �=    WE           �=     YE     [       �=    �YE     �      �=    p[E           �=    �]E     �       >    @^E     %       >    p^E     	      *>    �_E     �      >>    @aE            R>    PaE            h>    `aE     p       ~>    �aE     �      �>    �cE            �>    �cE            �>    �cE            �>    �cE     !       �>     dE            �>    @dE            �>    PdE     �      ?     gE           ?     iE     l       ?    �vE     :      0?    �yE     9       =?    zE     ?       Q?    PzE     %      c?    �|E     S       x?   ��                �?    �|E            �?    �|E            �?     }E     g       �?    p}E            �?    �}E            �?    �}E     C      �?    �~E     �       �?    �E     �       @   
 �hG     0       @    �E     �      2@    ��E     �      E@    ЄE            S@    P�E     �      d@    �E     )       q@    @�E     G       ~@    ��E     9       �@    ЉE     ?       �@    �E     j      �@    ��E            �@    ��E            �@    ��E            �@    ��E     �      A    p�E     *       A    ��E     �      7A    ��E     $       EA    ��E     S       YA   ��                bA    �E     �      mA    ��E     �       �A    `�E     R       �A    ��E     ~       �A    @�E     2      �A    ��E     �       �A    0�E            �A    @�E            �A    P�E            �A    p�E            �A    ��E     .      �A    ��E     A      B    �E     �      B    �E     b      &B   
 �lG     D       3B   
  lG     L       :B   
 �}G     x       AB   
 `~G     x       HB   
 �~G     |       OB   
 `G     |       VB   
 �mG            _B   
 �lG            hB    `�E     �      �B     �E     �      �B    ��E     	       �B   ��                �B    ��E     c       �B    P�E     �      �B    ��E     �       �B    ��E     ,      �B    `�E     L       C   ��                C    ��E     )       /C    �E     f      >C   
 ��G     �       LC    ��E     p       �C    ��E     c       ZC    `�E     �       nC    P�E     c       zC    ��E     $      �C    ��E     /      �C     �E     	       �C    0�E     �      �C     �E     �       �C     �E            �C     �E     s      D    ��E     �       D    0�E            %D    P F             8D     �E     E      QD     �E     )       jD    0�E     e      D    ��E     _      �D    @�E     D       �D    ��E     �       �D    p�E     D       �D    ��E     H       �D    �E     �       E    ��E     D       E    @�E     P       E    ��E            *E    ��E             ;E    ��E     1       QE    �E     1       eE    P�E     %       yE    ��E            �E    ��E            �E    ��E     d       �E    0�E            �E    @�E     6       �E    ��E            F    ��E            F    ��E     �      8F    ��E           HF    ��E     �      _F    ��E     �      {F    ��E     f       �F    ��E     �       �F    ��E            �F    ��E     (       �F    ��E     �       �F    ��E     g       �F    ��E     �       �F    � F     �      �F    ��E     �       G    ��E     Y       'G     �E     �       <G    ��E           LG    ��E     ]      \G    p F     �       lG    `F     �       �G    PF     �      �G    �F     �      �G    pF     �      �G    @F            �G    �F     x       �G    @	F     $      �G    @1F            H    `1F     T       H    �1F     J       3H    p
F     8      DH    �4F            UH     5F     d       lH    p5F     J       �H    �F     �       �H    `F           �H    rF     Z      �H    �F     �       �H   
 ��G     P      �H    F     c       I    �F     x       !I     F     h       8I    pF     {      MI    �F     �       mI    �F            �I    �F     	      �I     F     �       �I     F     �
      �I    �F            �I    �F            �I    �F            J    �F            /J    �F     2       AJ    F     5       UJ    PF     `       hJ    �F     `       zJ     F     >       �J    P F     Q       �J    �"F     �       �J    `#F     �      �J    �(F     j       �J    `)F     i       K     +F     �      !K    �)F     �       6K    p*F     �       MK    �,F     F      cK     /F     �      nK    1F     '       �K    2F     '       �K    @2F     <       �K    �2F     �       �K    `3F     F      L    �4F     '       L    �5F     �      <L    �8F     }       [L     9F            rL     9F     U       �L    �9F     b       �L    �9F     h      �L    `@F     �       �L    0AF     �       �L    �AF     x       �L    @BF     X       M    �BF     c/      M   
 ��G            +M   
  �G            >M   
 �G            QM   
  �G            dM   
 ��G     X       tM   ��                ~M    p�F     7       �M    ��F     �       �M    @�F     �       �M    ��F            �M    �F     #       �M    @�F     
       �M   
 ��G             N    P�F     �      /N    ��F           @N     �F     �      QN   
 ��G     (       mN   
  �G     U       �N   
 ��G     (       �N   
 ��G     @       �N   ��                �N    ��F     &       �N    ��F     V       �N    P�F            �N    `�F            �N    p�F            �N   ��                O   ��                     ��                O    (`i             O    xai             .O  
 �G     (       HO   �k@     �       ZO                     bO   ��F            qO  
 �!G            �O  
 �6G            �O   `�@     |       �O                     �O    �1@     �      �O  
 �0G            P  
 ��G     @       P  
  AG     (       2P   0r@     �      EP    �3@     ?      nP                     uP  
 `G     p       �P  
 @�F     P       �P    T@     P       �P  
 @?G     (       �P  
  G            �P   �f@            �P    �ji            �P    ��E           	Q  
 PG            Q  
  �G     h       +Q    �@     +       BQ  
  G             \Q  
 �1G            uQ  
 08G            �Q  
 @G     h       �Q    ?1@     W       �Q    @ui     (       �Q  
 �(G            �Q  
 `eG     H       R  
 �'G            %R  
 �4G            >R   @�@            NR  
 �4G            gR   0\@     �       �R  
 �<G     (       �R  
 @G     h       �R   @�@     �       �R    �E@     �       �R   І@     �       �R    �@     �       �R    @�F     �       S  
 `$G            #S    Pn@            5S   ��@     �       JS    '@     5       ]S                     eS    P�@     q      vS    �@     1       �S    0�@     +       �S   Щ@     �       �S    0�@            �S  
 �AG     (       �S  
 07G            �S  
 pG            T  
 @>G     (       T  
 �G            ,T    P�@     �      :T  
 �PG     �      JT    ��@     �       ]T    �@     g       jT    pn@     �       wT  
 7G            �T  
 `�F     �       �T  
 �wH           �T  
 �&G            �T  
 �%G     (       �T  
 `G            �T  
  <G     (        U  
   G     �       U    ИF     �      *U  
 �6G            CU   ��@     w       NU                     UU  
 04G            nU   ��@            zU   ��@     a       �U  
 P0G            �U    m&@     9       �U  
 @G     h       �U  "  P(@     )       �U  
  G     P       �U  
 �8G            V  
 @EG     (        V    �@     }       1V    ��E     4      CV  
 �DG     (       XV  
  -G     �      jV  
 �0G            �V  
 �GG     (       �V    ��@     S       �V    �/@     j      �V    ��@     F       �V    �e@            W    f@     f       *W  
 3G            CW    28@     �      QW  
  'G            cW    �@     6       sW  
 �G     h       �W  
 �"G            �W  
 �1G            �W  
  CG     (       �W   Pp@     �       �W                     �W  
 �1G            X   `�@     9       X  
 @:G     (       5X   ��E     *       GX  
  >G     (       \X    �@     �      oX  
 �G     h       �X   `�@     �       �X    c@     w       �X  
 @GG     (       �X  
 1G            �X  
 �5G            �X  
 �'G            Y  
 �?G     (       Y   ��@     �      'Y    Px@     �      6Y  
 0G            PY  
 �G            jY    �@     �       �Y  
 6G            �Y    �{@     3       �Y  
 �2G            �Y  
 `G            �Y    �`@     &       Z  
 `gG     x       (Z   P�@     x       7Z  
 �@G     (       LZ  "  �$@     "       iZ                     pZ  
 05G            �Z    ��@     �       �Z  "  �"@     I       �Z   �ti             �Z  
 ��G             �Z  
 �:G     (       �Z    ��@     /       �Z  
 �G            [  
 ��G     ��      [  
 p0G            5[  
 p1G            N[  
  "G            `[    `i             m[  
  BG     (       �[  
 @FG     (       �[   У@     6       �[   ��E     �       �[    pui            �[  
 �G            �[     o@     �       �[   g@            \    0S@     \       \  
 %G            %\  
 �HG     �      8\  
 P3G            Q\  
 �G     h       e\  
 �6G            ~\  
 �=G     (       �\  
 p7G            �\                     �\   ��@            �\    @�@     ;       �\    ��@     �       �\  
 �$G            ]  
 �CG     (       #]  
 ��F     �       4]  
 �!G             M]  
 �EG     (       b]  
  *G     @       �]  
 P6G            �]    `hi     (       �]  
 �;G     (       �]   ��@            �]    ��@     �       �]    �R@            �]  
 �G            ^    ��@     �       ^     �@             ^   �bi             -^  
 �2G            F^  
 8G            _^  
  G            q^  
 �G            �^  
 �G             �^  
 �FG     (       �^   `�@     B       �^   ��@     h       �^     �@     6      �^  
 �G            �^  "  �$@     "       _     D@     �      0_    �&@     3       C_  
  G            U_  
 `)G             m_  "  �$@     �       �_    (@     D       �_  
 #G            �_  
 09G            �_   Pa@     f       �_     �@     c       `  
 �2G            `  
 �/G            4`  
  �F     �       E`   @�@     �      V`   ��@     |       l`  
 `�F     �       }`   `�@            �`  
 `�F     �       �`  
 �G            �`  
 �@G     (       �`    q'@     4       �`  
 �%G     8       �`  
 �"G            a     S@            a  "  �(@            a  
 P2G            4a   `�@     (       Ja  
 �G     h       ]a  
 �G            oa     a@            a  
 ��G             �a    ��@           �a    ��@     g       �a    lui            �a  
 �0G            �a  
 @G             �a                     b    �ji            b  "  x#@     "       .b  
 �$G            Hb  
 @BG     (       ]b     ui            `b    �w@     i       sb  
 �'G            �b    �@     ?       �b    p{@     Q       �b  
 �>G     (       �b   �\@     �      �b   ��F            �b  
 `�G             �>    p	@             �b     �@     ^       �b  
 @G     h       c  
 �G            -c  
 G            ?c    �~@     �       Qc  
 @CG     (       fc    �z@     �       xc  
 �tH           �c    ��@     6       �c                     �c    @�@            �c  
  EG     (       �c  
 �4G            �c    ��@            �c  
 �"G     0       d   @�F     7       d  
 P7G            2d  
 �9G     (       Gd  
 � G           Yd    pv@     �       id    �hi            sd    xui            {d    �ui            �d   �@            �d  
 @G            �d   ��@            �d  
 �5G            �d  
 �7G            �d   ��@     x      	e  
 ��F     �       e  
 `&G            ,e     }@     �       ?e  "  #@     2       Se    )@     8       ne    `�@     f       }e    �@           �e    0�@     p       �e  
 p3G            �e   ��F     �       �e                     �e    �'@     1       �e  
 p8G            f  
 �3G            ,f    C@             Bf    ��F     -       Qf  
 %G            cf    hui            mf   �E     :       �f  
 PG            �f    p�@     �      �f  
 �!G            �f  
 �&G            �f  
 �G             �f   �a@           �f  
 �;G     (       g  
 �3G            +g  
 �5G            Dg   ��@     ^       Sg  
 �9G            lg    a@     #       g  
 �rH            �g    �S@             �g    �)@     �       �g  
 �HG     @       �g  
 �1G            �g  
 0&G            h                     h  
  ?G     (       #h    |@     i       4h    ��@     �      Dh  
  %G     H       ^h     �A     	2      hh  
 @'G     8       �h  
 03G            �h    p�@     F       �h    ��@     �      �h    �ui     (       �h  
  =G     (       �h  
 @DG     (       �h  
 01G            i  
 9G            0i    ��@     6       ?i     �@     g       Ui   ��@     4       li  
 @�F     �       �i   ��F            �i    8C@             �i   ��E     �      �i    �F            �i  
 �CG     (       �i  
  GG     (       �i                     �i  
 �8G            j   @�@     �      j  
 �'G            6j   ��@            Ij  
 P9G            bj    @�@     Q      sj  
 ��F     P       �j  
 �7G            �j   p�@     3       �j  
 p9G            �j  
 �yH     p      �j    `�@     C       k                     k    �9@     k      *k  
 �=G     (       ?k  
 �G            Qk  
  �G     H       fk   �D            {k   ��F            �k    ��@     !       �k    �@            �k    ��@     �       �k  "  #@     2       �k  
 �G            �k  
 P5G            l  
  $G            l     �@            $l  
 00G            =l  
 �2G            Vl   0g@     A       el  
 P1G            ~l    0�A     �       �l    ��@            �'    �@            �l  
 @@G     (       �l                     �l  
 �(G     8       �l    ��@     f       �l  
 p2G            �l    ��@     F       m  
 �'G            m  
  �G            )m  
 �/G            Bm   �@     $      \m   ��@     .       qm  
 �$G            �m  
 �6G            �m  
 �BG     (       �m                     �m  
 P4G            �m  "  �%@     �       �m    ��@     6        n   �d@     !       n  
 �>G     (       (n  
 �4G            An  "  �(@            In    N)@     �       dn   �p@     ^      vn                     ~n     �@     �       �n    P+@     [       �n    p�@            �n  
 @HG     @       �n    @F@     &       �n    b@     �       /Z                     o   P�@     1      ,o    �ui            8o    Pw@     �       Io   �S@     V       \o                     io  
 �&G            �o    :-@     Q       �o  
 P/G            �o    �m@     �       �o  
 �3G            �o                     �o    kui            �o  
  "G     (       p  
 �G            (p    �U@     �      9p   ��@     x       Sp  
 �7G            lp  
 p4G            �p    �@            �p    �-@     J      �p    �@     V       �p    ",@           �p  
 PG            q                     q   @�@     V       q  
 0G            8q   �^@            Nq  
 @�F     P       aq  
 @G     H       sq     �F     V       �q  
  @G     (       �q    �@     �       �q     �@            �q    X>@     �      �q  "  8#@     -       �q                     �q  
 @G     h        r  
 �.G     (       r   0�D     �      0r   �k@            Hr  
 8$G            br  
 @*G     �      sr    ��@     c      �r  
 `G            �r  
  :G     (       �r  
 `�G     P       �r   ��@     �       �r  
  �G            �r  
 pG            s  
  �G     @       "s    ��@     S       <s                     Bs    �ti             Ns    �+@     I       ts    `T@     Q      �s                     �s     v@     p       �s    {6@     �      �s    @     a      �s  
  DG     (       �s   ��E     �       �s                     �s  
 @=G     (       �s  
 �'G            t  
 'G            ,t  
 p6G            Et  
 �EG     (       Zt  
 0G            tt  
 �8G            �t  
 �G           �t  
 @$G            �t    �ni            �t    �+@     .       �t   �X@     !      �t  
 �GG     (       �t  "  �(@            �t  
 ��F     �       u    ��@            #u                     *u    @�@     �      8u  
 @G            Ju    @�@     ;       cu  
 �&G            uu  
  )G     H       �u    P�@            �u  
 �&G             �u                     �u  "  @&@     -       �u  
 �FG     (       �u  "  @&@     -       v   0NE            v  
 �"G            #v    ��@     �       3v  
 02G            Lv     �@     .       [v                     bv    ��@           rv    <'@     5       �v    |C@             �v  
 P$G            �v  
 @�G     P       �v  
 �?G     (       �v   	 �F             �v    ��@     c       �v  
 �eG     x       w                     w  
 �/G            7w   �Y@     g      Gw    д@     /       Uw  
  HG     (       jw    @`@     �       |w    @a@            �w  
 4G            �w  
  G     h       �w  
 �G            �w   �c@     Y       �w  "  f#@            x  
 06G            'x  
 �DG     (       <x    ��@     I       \x  
 2G            ux   ��@     O       �x  
 �#G            �x  
 �G            �x  
  ;G     (       �x  
 0/G            �x  
 �G            �x  
 p#G            y   �g@     d       y    @�@            (y    P�@            8y   ph@     7      Sy  
  (G     �       my  
  &G     0       y  
 �G            �y    ��@     �       �y   �f@     [       �y   и@     Z      �y   �d@     #       �y  
  �F     `           �bi     �      �y  
 p&G            z    @�F     �      (z  
 P8G            Az  "  y(@     )       Gz    ��@     L      Wz    ��@     V       gz    �*@     u       �z    @�@            �z  
 �G             �z  
 0G            �z  
 �pH            �z  
 p5G            �z   ЉF            �z   �@            {    ��@     ,       {    �'@     6       6{    ��@     :       I{   �@           b{    `�@     /      x{   ��@            �{  
 /G            �{  
 �fG     x       �{  
 �G            �{  
 �)G     @       �{  
 �8G            	|  
 x$G            #|    g@            4|   ��@     ;      @|  
 @#G     0       Z|    @z@     �       o|    p@     &       }|   0�@     '       �|    �ti             �|    �|@     u       &    �ui             �|     �F           �|    ��E     �       �|  "  8#@     -       �|    �ji            �|  
 �0G            }    �D            -}  
 �<G     (       B}  
 �G     0       \}    d@     y       m}  
 `"G     8       �}  
 �G     8       �}  
 �BG     (       �}  
 �5G            �}  
 �&G            �}  
 P&G            �}  
  �G     P       ~  
 �:G     (       )~    ��@     �       :~  
 �3G            R~  
 @�G     H       e~  
 p/G            ~~  
 0G            �~    P�@     >       �~  
  G     0       �~  
 �$G            �~  
 P"G            �~    ��@            �~  
 @;G     (           c@               
 @G            :  
 �(G            T  
 �#G     8       n  
 @AG     (       �   `�@     �       �    �@     J      �    �}@     �       �  
 @<G     (       �    �D            �    `�F     f      �  
 `fG     0       �    #3@     �       3�   ��@     '       K�   ��@     6      X�                     _�  
  'G            q�                     y�  
 `hG     0       ��   �@     (       ��   �^@     �       ��  
 �gG     x       ɀ  
  FG     (       ހ  
  G            ��  "  �#@     -      �    �C@     3       0�  
 @&G            B�    `�@     ~       I�   @�@     2       W�    @�@     6       h�   ��F            y�    �&@     .       ��  
  �F     �       ��  
 �/G            ��    �ji            ��  
 ��G     P       ؁    �@     �       �  
 �$G     (       �   ��@            �   �@            "�  
 �#G     @       <�  
 �G     h       O�  
 �AG     (       d�    (ui            k�  
 �G            }�    S@            ��  "  �(@            ��    �B@             ��  
 5G            ��  
 �G            ǂ     f@            ߂  
 �7G            ��    �ui             �    [6@             �     �@     F      !�    �_@     �       5�  
 `G     (       O�   �d@           ^�    ;5@            uU                     ��  
 ��G            ��  
 �'G             crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.5420 dtor_idx.5422 frame_dummy object.5432 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_mouse fb.cpp filesystem.cpp ipc.cpp runtime.cpp graphics.cpp text.cpp _ZL9fontState _ZL7library _ZL8mainFont ../src/gfx/sse2.asm memcpy_sse2.loop memcpy_sse2_unaligned.loop memset32_sse2.loop memset32_sse2.ret memset64_sse2.loop memset64_sse2.ret font.cpp ftinit.c ft_default_modules ftbase.c hash_num_compare hash_bucket destroy_size find_unicode_charmap memory_stream_close ft_recompute_scaled_metrics ft_raccess_sort_ref_by_id hash_str_compare ft_trig_pseudo_rotate.isra.2 ft_trig_arctan_table ft_trig_pseudo_polarize.isra.3 ft_trig_prenorm.isra.4 ft_property_do _ft_face_scale_advances.isra.6.part.7 FT_Match_Size.part.8 FT_Outline_Get_CBox.part.14 FT_Outline_Render.part.15 FT_Vector_Transform.part.16 FT_Outline_Transform.part.17 FT_Vector_Unit.part.19 destroy_charmaps.part.23 FT_List_Add.part.24 FT_List_Remove.part.25 FT_List_Finalize.part.27 FT_GlyphLoader_Done.part.20 ft_glyphslot_done destroy_face find_variant_selector_charmap.isra.10 ft_raccess_guess_table raccess_guess_apple_generic.isra.18 raccess_guess_apple_single raccess_guess_apple_double raccess_make_file_name raccess_guess_linux_cap raccess_guess_vfat raccess_guess_darwin_hfsplus raccess_guess_darwin_newvfs raccess_guess_linux_double_from_file_name raccess_guess_linux_netatalk raccess_guess_linux_double raccess_guess_darwin_ufs_export open_face hash_insert IsMacResource open_face_PS_from_sfnt_stream.isra.28 open_face_from_buffer ft_open_face_internal truetype.c tt_get_kerning tt_get_metrics_incr_overrides TT_Load_Glyph_Header tt_loader_set_pp ft_var_get_value_pointer tt_cvt_ready_iterator TT_MulFix14_long_long Current_Ppem Read_CVT Write_CVT Move_CVT Direct_Move_X Direct_Move_Y Direct_Move_Orig_X Direct_Move_Orig_Y Round_None SetSuperRound Dual_Project Project_x Project_y Compute_Funcs Direct_Move Direct_Move_Orig SkipCode opcode_length Ins_MIRP Ins_DELTAP tt_size_init tt_driver_init tt_driver_done tt_face_get_location tt_size_reset tt_size_select tt_size_reset_iterator ft_var_apply_tuple Compute_Point_Displacement Ins_IP TT_Done_Context tt_glyphzone_done tt_size_done_bytecode tt_size_done ft_var_done_item_variation_store tt_done_blend Update_Max TT_Load_Context tt_size_run_prep TT_Hint_Glyph TT_Access_Glyph_Frame TT_Forget_Glyph_Frame ft_var_readpackedpoints ft_var_readpackeddeltas Current_Ratio Move_CVT_Stretched Write_CVT_Stretched Read_CVT_Stretched Current_Ppem_Stretched TT_Load_Simple_Glyph tt_slot_init tt_face_done ft_var_load_avar tt_face_vary_cvt tt_face_load_cvt ft_var_load_item_variation_store TT_Load_Composite_Glyph tt_property_get TT_Get_VMetrics tt_get_advances tt_get_var_blend Ins_Goto_CodeRange.part.5 Ins_UNKNOWN Round_To_Grid Round_To_Half_Grid Round_Down_To_Grid Round_Up_To_Grid Round_To_Double_Grid Round_Super Round_Super_45 Ins_JMPR Move_Zp2_Point Ins_MDRP.isra.48 tt_delta_interpolate.part.51 TT_Vary_Apply_Glyph_Deltas load_truetype_glyph _iup_worker_interpolate.part.53 Ins_IUP tt_size_request ft_var_to_normalized.isra.55 TT_Get_MM_Var fvar_fields.5740 fvaraxis_fields.5741 tt_set_mm_blend gvar_fields.5612 TT_Set_Var_Design TT_Set_Named_Instance TT_Get_Var_Design TT_Get_MM_Blend ft_var_get_item_delta.isra.57 tt_apply_mvar tt_face_init trick_names.7460 sfnt_id.7489 TT_Set_MM_Blend ft_var_load_hvvar tt_hvadvance_adjust tt_vadvance_adjust tt_hadvance_adjust tt_get_interface tt_services tt_property_set Normalize.isra.64.part.65 Ins_SxVTL Pop_Push_Count tt_loader_init TT_Load_Glyph tt_glyph_load tt_service_gx_multi_masters tt_service_metrics_variations tt_service_truetype_engine tt_service_truetype_glyf tt_service_properties type1.c t1_get_ps_name t1_ps_get_font_info t1_ps_get_font_extra t1_ps_has_glyph_names t1_ps_get_font_private T1_Get_Multi_Master T1_Set_MM_WeightVector T1_Get_MM_WeightVector parse_buildchar parse_private read_binary_data T1_GlyphSlot_Done T1_Driver_Init T1_Driver_Done T1_GlyphSlot_Init T1_Parse_Glyph_And_Get_Char_String T1_Parse_Glyph T1_Compute_Max_Advance T1_Get_Advances t1_allocate_blend parse_weight_vector parse_blend_design_positions parse_blend_design_map T1_Done_Metrics T1_Done_Blend T1_Load_Glyph T1_Face_Done t1_get_name_index parse_dict t1_keywords read_pfb_tag parse_blend_axis_types parse_subrs mm_axis_unmap t1_parse_font_matrix t1_services T1_Get_Track_Kerning t1_ps_get_font_value t1_get_glyph_name mm_weights_unmap T1_Get_MM_Blend T1_Get_Var_Design T1_Get_MM_Var t1_set_mm_blend.isra.2 T1_Set_MM_Design T1_Set_Var_Design T1_Set_MM_Blend T1_Reset_MM_Blend T1_Size_Get_Globals_Funcs.isra.4 T1_Size_Request T1_Size_Init T1_Size_Done t1_get_index T1_Read_Metrics check_type1_format T1_Open_Face T1_Face_Init t1_service_ps_name t1_service_glyph_dict t1_service_ps_info t1_service_properties t1_service_kerning t1_service_multi_masters cff.c cff_cmap_encoding_init cff_cmap_encoding_done cff_cmap_encoding_char_index cff_cmap_encoding_char_next cff_cmap_unicode_init cff_sid_to_glyph_name cff_cmap_unicode_char_index cff_cmap_unicode_char_next cff_get_kerning cff_ps_has_glyph_names cff_get_is_cid cff_get_cid_from_glyph_index cff_set_mm_blend cff_get_mm_blend cff_set_mm_weightvector cff_get_mm_weightvector cff_get_mm_var cff_set_var_design cff_get_var_design cff_set_instance cff_hadvance_adjust cff_metrics_adjust cff_parse_integer cff_get_standard_encoding cff_standard_encoding cff_fd_select_get cff_get_var_blend cff_done_blend cff_slot_done cff_driver_init cff_driver_done cff_cmap_unicode_done cff_vstore_done cff_slot_init cff_make_private_dict cff_index_done cff_get_cmap_info cff_get_ps_name cff_parse_real power_tens cff_get_name_index cff_charset_compute_cids cff_blend_check_vector cff_blend_build_vector cff_index_get_pointers cff_index_get_sid_string cff_get_ros cff_ps_get_font_info cff_ps_get_font_extra cff_size_get_globals_funcs.isra.7 cff_size_select cff_size_done cff_size_request cff_size_init cff_index_read_offset.isra.8 cff_index_access_element cff_index_get_name cff_index_init cff_get_glyph_data cff_free_glyph_data cff_slot_load cff_glyph_load cff_get_advances cff_subfont_done.part.12 cff_face_done do_fixed.isra.13 power_ten_limits cff_parse_font_bbox cff_parse_num.isra.16 cff_parser_run cff_field_handlers cff_load_private_dict cff_parse_vsindex cff_parse_maxstack cff_parse_cid_ros cff_parse_multiple_master cff_parse_private_dict cff_parse_blend cff_parse_font_matrix cff_get_interface cff_services cff_get_glyph_name cff_subfont_load cff_face_init cff_header_fields.6734 cff_isoadobe_charset cff_expert_encoding cff_expert_charset cff_expertsubset_charset cff_service_multi_masters cff_service_metrics_variations cff_service_ps_info cff_service_ps_name cff_service_glyph_dict cff_service_get_cmap_info cff_service_cid_info cff_service_properties cff_service_cff_load type1cid.c parse_expansion_factor parse_font_name cid_slot_done cid_driver_init cid_driver_done cid_get_postscript_name cid_ps_get_font_info cid_ps_get_font_extra cid_get_ros cid_get_is_cid cid_get_cid_from_glyph_index cid_slot_init cid_load_glyph cid_slot_load_glyph cid_face_done cid_parse_font_matrix parse_fd_array cid_get_interface cid_services cid_size_get_globals_funcs.isra.0 cid_size_request cid_size_init cid_size_done cid_face_init cid_field_records cid_service_ps_name cid_service_ps_info cid_service_cid_info cid_service_properties pfr.c pfr_cmap_init pfr_cmap_done pfr_cmap_char_index pfr_cmap_char_next pfr_get_advance pfr_face_get_kerning pfr_extra_item_load_stem_snaps pfr_extra_item_load_bitmap_info pfr_slot_done pfr_slot_init pfr_extra_item_load_kerning_pairs pfr_extra_item_load_font_id pfr_aux_name_load pfr_get_service pfr_services pfr_get_metrics pfr_glyph_close_contour.isra.0 pfr_get_kerning pfr_glyph_line_to.isra.3 pfr_glyph_load_rec pfr_slot_load pfr_face_done pfr_face_init pfr_header_fields pfr_phy_font_extra_items pfr_metrics_service_rec type42.c t42_get_ps_font_name t42_ps_get_font_info t42_ps_get_font_extra t42_ps_has_glyph_names t42_ps_get_font_private T42_Driver_Done T42_Size_Select T42_Size_Request T42_GlyphSlot_Done T42_GlyphSlot_Init T42_Size_Init T42_Face_Done T42_Driver_Init t42_get_name_index t42_parse_sfnts t42_parse_font_matrix T42_Get_Interface t42_services t42_get_glyph_name t42_is_space t42_parse_charstrings t42_parse_encoding T42_GlyphSlot_Load T42_Size_Done T42_Face_Init t42_keywords t42_service_glyph_dict t42_service_ps_font_name t42_service_ps_info winfnt.c fnt_cmap_init fnt_cmap_char_index fnt_cmap_char_next winfnt_get_header FNT_Size_Select FNT_Load_Glyph fnt_font_done winfnt_get_service winfnt_services FNT_Size_Request fnt_font_load winfnt_header_fields FNT_Face_Init fnt_cmap_class_rec winmz_header_fields winne_header_fields winpe32_header_fields winpe32_section_fields winpe_rsrc_dir_fields winpe_rsrc_dir_entry_fields winpe_rsrc_data_entry_fields FNT_Face_Done winfnt_service_rec pcf.c pcf_cmap_init pcf_cmap_done pcf_cmap_char_index pcf_cmap_char_next pcf_get_charset_id pcf_property_set pcf_property_get pcf_driver_init pcf_driver_done PCF_Size_Select PCF_Size_Request PCF_Glyph_Load pcf_seek_to_table_type pcf_driver_requester pcf_services PCF_Face_Done.part.0 PCF_Face_Done pcf_find_property.isra.1 pcf_get_bdf_property pcf_get_metric pcf_metric_header pcf_metric_msb_header pcf_compressed_metric_header pcf_get_accel pcf_accel_header pcf_accel_msb_header pcf_load_font pcf_toc_header pcf_table_header pcf_property_header pcf_property_msb_header pcf_enc_header pcf_enc_msb_header PCF_Face_Init pcf_cmap_class pcf_service_bdf pcf_service_properties bdf.c _bdf_atol ddigits a2i _bdf_atos by_encoding _bdf_parse_end bdf_cmap_init bdf_cmap_done bdf_cmap_char_index bdf_cmap_char_next bdf_get_charset_id BDF_Size_Select BDF_Glyph_Load _bdf_list_ensure _bdf_list_done _bdf_add_comment bdf_driver_requester bdf_services _bdf_atoul.part.0 _bdf_atous.part.1 BDF_Size_Request bdf_free_font.part.3 BDF_Face_Done _bdf_list_split empty bdf_get_font_property.part.5 bdf_get_bdf_property _bdf_add_property.isra.7 _bdf_properties BDF_Face_Init _bdf_parse_start bdf_cmap_class _bdf_list_join.constprop.11 _bdf_list_shift.constprop.12 _bdf_parse_properties _bdf_parse_glyphs hdigits nibble_mask bdf_service_bdf sfnt.c get_sfnt_table sfnt_is_postscript sfnt_ps_map sfnt_is_alphanumeric sfnt_get_name_id compare_offsets tt_cmap_init tt_cmap0_char_index tt_cmap0_char_next tt_cmap0_get_info tt_cmap2_get_subheader tt_cmap2_char_index tt_cmap2_char_next tt_cmap2_get_info tt_cmap4_init tt_cmap4_set_range tt_cmap4_next tt_cmap4_char_map_linear tt_cmap4_char_map_binary tt_cmap4_char_index tt_cmap4_get_info tt_cmap6_char_index tt_cmap6_char_next tt_cmap6_get_info tt_cmap8_char_index tt_cmap8_char_next tt_cmap8_get_info tt_cmap10_char_index tt_cmap10_char_next tt_cmap10_get_info tt_cmap12_init tt_cmap12_next tt_cmap12_char_map_binary tt_cmap12_char_index tt_cmap12_get_info tt_cmap13_init tt_cmap13_next tt_cmap13_char_map_binary tt_cmap13_char_index tt_cmap13_get_info tt_cmap14_init tt_cmap14_char_index tt_cmap14_char_next tt_cmap14_get_info tt_cmap14_char_map_def_binary tt_cmap14_char_map_nondef_binary tt_cmap14_find_variant tt_cmap14_char_var_index tt_cmap14_char_var_isdefault tt_cmap_unicode_init tt_get_glyph_name tt_cmap_unicode_char_index tt_cmap_unicode_char_next tt_get_cmap_info tt_face_get_colr_layer tt_face_palette_set tt_face_get_kerning tt_sbit_decoder_load_metrics tt_sbit_decoder_load_byte_aligned tt_sbit_decoder_load_bit_aligned sfnt_get_interface sfnt_services tt_face_load_kern tt_face_free_sbit tt_face_goto_table tt_face_find_bdf_prop sfnt_get_charset_id tt_face_load_hmtx tt_face_get_metrics tt_name_ascii_from_other tt_name_ascii_from_utf16 tt_cmap14_ensure tt_cmap14_get_def_chars tt_cmap14_get_nondef_chars tt_cmap14_variant_chars tt_cmap14_char_variants tt_cmap14_variants tt_face_load_gasp tt_face_get_name tt_face_free_colr tt_face_free_cpal tt_face_free_ps_names tt_face_free_name sfnt_done_face sfnt_stream_close tt_cmap14_done tt_cmap_unicode_done tt_face_load_colr tt_face_load_cpal tt_face_load_any tt_sbit_decoder_load_image tt_sbit_decoder_load_compound tt_face_colr_blend_layer tt_face_load_strike_metrics tt_face_set_sbit_strike tt_face_load_sbit tt_face_load_pclt pclt_fields.6446 tt_face_load_name name_table_fields.6388 name_record_fields.6389 langTag_record_fields.6390 tt_face_load_post post_fields.6441 tt_face_load_maxp maxp_fields.6374 maxp_fields_extra.6375 tt_face_load_hhea metrics_header_fields.6481 tt_face_build_cmaps tt_cmap_classes sfnt_load_face tt_encodings.4952 tt_cmap2_validate tt_cmap4_validate tt_cmap6_validate tt_cmap8_validate tt_cmap10_validate tt_cmap12_validate tt_cmap13_validate tt_cmap14_validate sfnt_table_info tt_cmap4_char_next tt_cmap12_char_next tt_cmap13_char_next tt_face_load_cmap load_post_names tt_face_get_ps_name.part.8 tt_face_get_ps_name sfnt_get_name_index sfnt_get_glyph_name tt_face_load_font_dir offset_table_fields.6327 table_dir_entry_fields.6310 tt_face_load_generic_header header_fields.6358 tt_face_load_bhed tt_face_load_head tt_face_load_os2 os2_fields.6430 os2_fields_extra1.6431 os2_fields_extra2.6432 os2_fields_extra5.6433 sfnt_init_face woff_header_fields.5096 ttc_header_fields.4966 tt_cmap0_validate tt_face_load_sbit_image get_apple_string.constprop.17 get_win_string.constprop.18 sfnt_get_ps_name hexdigits sfnt_interface sfnt_service_sfnt_table sfnt_service_ps_name sfnt_service_glyph_dict sfnt_service_bdf tt_service_get_cmap_info autofit.c af_sort_and_quantize_widths af_cjk_get_standard_widths af_cjk_hints_compute_blue_edges af_cjk_hints_init af_cjk_snap_width af_latin_snap_width af_dummy_hints_init af_indic_hints_init af_indic_get_standard_widths af_latin_get_standard_widths af_latin_hints_link_segments af_latin_hints_init af_autofitter_init af_autofitter_done af_warper_compute_line_best af_warper_weights af_glyph_hints_reload af_latin_hints_compute_segments af_axis_hints_new_edge af_glyph_hints_align_strong_points af_cjk_metrics_scale_dim af_cjk_metrics_scale af_indic_metrics_scale af_latin_hints_compute_edges af_latin_metrics_scale_dim af_latin_metrics_scale af_glyph_hints_done af_face_globals_free af_get_interface af_services af_cjk_compute_stem_width.isra.0 af_hint_normal_stem af_glyph_hints_save.isra.5 af_latin_compute_stem_width.isra.7 af_latin_align_linked_edge af_dummy_hints_apply af_cjk_hints_detect_features af_iup_interp.part.11 af_glyph_hints_align_weak_points af_loader_compute_darkening.isra.15 af_face_globals_new af_autofitter_load_glyph af_property_get_face_globals af_property_get af_property_set af_warper_compute.constprop.22 af_cjk_hints_apply af_indic_hints_apply af_latin_hints_apply af_cjk_metrics_init_widths af_cjk_metrics_init_blues af_cjk_metrics_check_digits.isra.17 af_cjk_metrics_init af_indic_metrics_init af_latin_metrics_init_widths af_latin_metrics_init_blues af_latin_metrics_init af_service_properties pshinter.c psh_hint_table_record psh_globals_scale_widths psh_globals_set_scale pshinter_get_globals_funcs pshinter_get_t1_funcs pshinter_get_t2_funcs t1_hints_open t2_hints_open ps_hinter_init psh_globals_new psh_globals_destroy ps_hints_close t1_hints_stem ps_hints_t1stem3 ps_hints_t1reset t2_hints_stems ps_hints_t2mask ps_hints_t2counter psh_hint_table_done ps_mask_table_done psh_hint_table_activate_mask.isra.3 psh_hint_table_find_strong_points.isra.4 psh_hint_table_init.isra.12 ps_mask_table_alloc ps_mask_ensure.isra.16 ps_mask_set_bit ps_dimension_add_t1stem ps_hints_stem.part.17 ps_mask_table_merge_all psh_blues_set_zones_0.constprop.26 psh_blues_set_zones psh_hint_align ps_hints_apply.part.21 ps_hinter_done ps_dimension_set_mask_bits pshinter_interface raster.c New_Profile End_Profile Insert_Y_Turn Split_Conic Split_Cubic Bezier_Up Bezier_Down Conic_To Cubic_To Sort Vertical_Sweep_Init Vertical_Sweep_Span Vertical_Sweep_Drop Vertical_Sweep_Step Horizontal_Sweep_Init Horizontal_Sweep_Span Horizontal_Sweep_Drop Horizontal_Sweep_Step ft_black_reset ft_black_set_mode ft_raster1_init ft_raster1_set_mode ft_black_done Line_Up Line_To Render_Single_Pass ft_black_render ft_black_new ft_raster1_get_cbox ft_raster1_render ft_raster1_transform smooth.c gray_raster_reset gray_raster_set_mode ft_smooth_init ft_smooth_set_mode gray_raster_done gray_hline gray_record_cell gray_convert_glyph_inner func_interface gray_convert_glyph gray_raster_render gray_set_cell gray_render_line gray_line_to gray_move_to gray_raster_new ft_smooth_get_cbox ft_smooth_render_generic ft_smooth_render ft_smooth_render_lcd ft_smooth_render_lcd_v gray_render_cubic.isra.0 gray_cubic_to gray_render_conic.isra.1 gray_conic_to ft_smooth_transform ftgzip.c huft_build inflate_blocks_reset inflateReset inflateEnd adler32 ft_gzip_stream_close ft_gzip_free zcfree ft_gzip_alloc zcalloc ft_gzip_check_header inflate_flush inflateInit2_.constprop.4 inflate inflate_mask border cpdext cpdist cplext cplens fixed_tl fixed_td ft_gzip_file_fill_output ft_gzip_file_io ft_gzip_stream_io ftlzw.c ft_lzw_check_header ft_lzwstate_get_code ft_lzwstate_stack_grow ft_lzw_stream_io ft_lzw_stream_close psaux.c afm_compare_kern_pairs PS_Conv_Strtol ft_char_table PS_Conv_ToInt skip_literal_string skip_string skip_procedure ps_parser_skip_PS_token ps_parser_skip_spaces ps_parser_to_token ps_parser_to_token_array ps_parser_to_int ps_parser_to_bytes ps_parser_init ps_parser_done ps_parser_to_fixed ps_parser_to_coord_array ps_parser_to_fixed_array ps_parser_load_field ps_parser_load_field_table t1_builder_done t1_builder_close_contour cff_builder_done cff_builder_add_point cff_builder_close_contour ps_builder_done t1_decrypt cff_random t1_cmap_std_done t1_cmap_standard_init t1_cmap_expert_init t1_cmap_custom_init t1_cmap_custom_done t1_cmap_custom_char_index t1_cmap_custom_char_next psaux_get_glyph_name t1_cmap_unicode_init t1_cmap_unicode_char_index t1_cmap_unicode_char_next t1_decoder_parse_metrics cf2_hintmap_map cf2_hintmap_insertHint cf2_glyphpath_computeOffset ps_table_release t1_decoder_done afm_parser_done t1_cmap_unicode_done ps_table_done afm_parser_init ps_table_new ps_table_add cf2_arrstack_setNumElements cf2_arrstack_push t1_builder_add_point PS_Conv_ToFixed ps_tofixedarray ps_builder_init cf2_getSeacComponent cf2_hint_init t1_make_subfont ps_decoder_init t1_builder_add_contour cff_builder_add_contour t1_builder_init t1_builder_check_points t1_builder_add_point1 t1_builder_start_point cff_builder_init cff_check_points cff_builder_add_point1 cff_builder_start_point t1_lookup_glyph_by_stdcharcode_ps t1_decoder_init cf2_decoder_parse_charstrings afm_tokenize afm_key_table afm_stream_skip_spaces.part.0 afm_stream_read_one afm_stream_read_string afm_parser_read_vals ps_builder_close_contour.isra.1 cf2_builder_moveTo cff_decoder_prepare cf2_glyphpath_hintPoint.isra.35 cf2_hintmap_build cf2_buf_readByte.part.39 cf2_stack_pushInt.part.43 cf2_stack_setReal.part.48 cf2_stack_pushFixed.part.44 cf2_stack_pushInt cf2_stack_pushFixed cf2_stack_popFixed cf2_stack_getReal cf2_stack_pop cf2_free_instance cf2_doStems.isra.54 cf2_glyphpath_pushPrevElem cf2_getT1SeacComponent.isra.58 cf2_glyphpath_closeOpenPath.part.60 cf2_glyphpath_lineTo cf2_glyphpath_moveTo cf2_glyphpath_pushMove cf2_glyphpath_curveTo cf2_doFlex t1_builder_check_points.part.61 ps_builder_check_points.isra.63.part.64 ps_builder_add_point1.part.65 ps_builder_start_point.part.66 cf2_builder_cubeTo cff_check_points.part.67 cf2_computeDarkening.part.71 t1_cmap_std_char_index.part.72 t1_cmap_std_char_index t1_cmap_std_char_next afm_parser_next_key.constprop.76 afm_parser_parse cff_decoder_init cf2_hintmask_read cf2_builder_lineTo cf2_stack_popInt cf2_interpT2CharString readFromStack.7928 readFromStack.7926 readFromStack.7923 readFromStack.7921 psaux_interface psnames.c compare_uni_maps ps_unicodes_char_index ps_unicodes_char_next ps_get_macintosh_name ps_get_standard_strings psnames_get_service pscmaps_services ft_get_adobe_glyph_index.part.0 ps_unicode_value ps_unicodes_init ft_extra_glyph_name_offsets ft_extra_glyph_names ft_extra_glyph_unicodes pscmaps_interface ftsystem.c ft_ansi_stream_close ft_ansi_stream_io ft_alloc ft_free ft_realloc ftdebug.c ftbitmap.c _DYNAMIC _GLOBAL_OFFSET_TABLE_ af_mlym_nonbase_uniranges FT_Done_GlyphSlot longjmp FT_Done_Memory af_khms_nonbase_uniranges af_cyrl_titl_style_class FT_Stream_ReadULong strcpy _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface af_osma_dflt_style_class t1_builder_funcs af_knda_script_class FT_Request_Metrics _Z10surfacecpyP7SurfaceS0_8Vector2i4Rect setjmp af_latp_uniranges cff_cmap_unicode_class_rec FT_DivFix af_mong_script_class af_lisu_nonbase_uniranges ft_validator_init mousePos FT_Stream_OpenGzip af_tibt_uniranges ps_parser_funcs FT_Stream_ReleaseFrame af_limb_nonbase_uniranges af_mymr_dflt_style_class af_copt_dflt_style_class tt_cmap_unicode_class_rec _Z20DrawGradientVertical4Rect10RGBAColourS0_P7Surface renderBuffer af_adlm_uniranges pshinter_module_class af_bamu_uniranges af_grek_sups_style_class FT_Stream_Close af_gujr_dflt_style_class FT_Vector_Transform_Scaled af_sund_script_class tt_cmap6_class_rec FT_Stream_ReadUShortLE FT_Init_FreeType ft_module_get_service FT_Raccess_Guess FT_GlyphSlot_Own_Bitmap af_glag_uniranges FT_Reference_Face FT_Stream_ReadUShort _Z10lemon_readiPvm memmove FT_Get_Sfnt_Name ft_mem_qalloc FT_Set_Debug_Hook FT_Stream_ReadUOffset FT_List_Finalize af_kali_script_class af_cyrl_subs_style_class af_orkh_nonbase_uniranges af_olck_script_class af_nkoo_uniranges FT_Load_Glyph af_blue_strings FT_Vector_Polarize ft_mem_alloc FT_Done_Face af_cyrl_sups_style_class tt_driver_class ft_mac_names af_cher_uniranges af_cyrl_nonbase_uniranges af_osge_uniranges af_tavt_script_class af_latn_nonbase_uniranges FT_Bitmap_Blend af_deva_dflt_style_class ft_mem_dup getenv af_kali_dflt_style_class ft_mem_free FT_Lookup_Renderer af_taml_dflt_style_class _Z12lemon_map_fbP6FBInfo tt_cmap2_class_rec _Znwm af_tibt_nonbase_uniranges af_cakm_dflt_style_class af_copt_script_class FT_Stream_ReadAt FT_Stream_OpenLZW af_cyrl_script_class af_script_classes af_shaw_dflt_style_class af_armn_script_class FT_Face_GetVariantsOfChar _Z12DrawGradientiiii10RGBAColourS_P7Surface FT_New_Memory_Face FT_Library_SetLcdFilterWeights FT_Library_SetLcdGeometry af_latn_sinf_style_class _Z8LoadFontPc af_buhd_uniranges FT_Render_Glyph tt_cmap12_class_rec af_kali_uniranges af_mong_dflt_style_class af_goth_script_class ft_synthesize_vertical_metrics qsort af_mlym_dflt_style_class FT_GlyphLoader_CheckPoints af_sylo_script_class ft_lzwstate_reset af_orkh_script_class _Z13AddNewWindowsv tt_cmap4_class_rec ps_property_get FT_GlyphLoader_Prepare af_avst_script_class af_osge_dflt_style_class af_grek_c2sc_style_class af_armn_uniranges af_lisu_script_class ps_property_set FT_Get_Kerning af_osma_nonbase_uniranges af_hani_nonbase_uniranges _Z19PointInWindowProperP8Window_s8Vector2i af_glag_dflt_style_class FT_Get_Char_Index af_latn_sups_style_class af_taml_uniranges FT_Palette_Set_Foreground_Color ft_smooth_lcd_renderer_class ft_mem_realloc af_latn_script_class _ZN8ListNodeIP8Window_sEC2Ev memcpy af_grek_smcp_style_class FT_Outline_Reverse _ZplRK8Vector2iS1_ __TMC_END__ t1_decoder_funcs af_orya_script_class FT_Outline_Translate af_sinh_uniranges ft_adobe_glyph_list af_sund_dflt_style_class af_none_dflt_style_class af_khms_uniranges __DTOR_END__ af_hebr_script_class af_cakm_script_class FT_Stream_ExitFrame ft_lzwstate_done dragOffset af_nkoo_nonbase_uniranges FT_Done_Size ft_validator_error FT_MulDiv af_dsrt_nonbase_uniranges af_blue_stringsets af_latn_ordn_style_class tt_cmap14_class_rec af_cyrl_dflt_style_class af_osma_script_class af_cyrl_sinf_style_class malloc FT_GlyphLoader_CheckSubGlyphs FT_Face_GetVariantSelectors FT_Set_Charmap af_geok_uniranges af_geok_script_class pcf_driver_class af_lao_nonbase_uniranges af_cari_script_class af_indic_writing_system_class af_geor_dflt_style_class mouseSurface af_telu_script_class FT_Stream_Read FT_Get_SubGlyph_Info FT_RoundFix af_sinh_nonbase_uniranges FT_Get_Advance FT_List_Add __dso_handle af_latn_smcp_style_class af_cprt_dflt_style_class af_saur_uniranges af_shaw_nonbase_uniranges af_thai_nonbase_uniranges af_beng_script_class FT_Stream_Seek FT_Stream_TryRead FT_New_Size af_sund_uniranges _ZN8ListNodeIP8Window_sEC1Ev FT_Set_Default_Properties _Z10lemon_openPKci af_limb_uniranges af_autofitter_interface _ZN4ListIP8Window_sE8add_backES1_ _Z11SendMessagem13ipc_message_t af_hebr_uniranges af_avst_dflt_style_class FT_GlyphLoader_Rewind FT_Get_Sfnt_Table af_latn_titl_style_class af_tfng_dflt_style_class pfr_driver_class FT_New_GlyphSlot FT_Stream_ReadULongLE cff_driver_class ft_property_string_set t1_driver_class af_orkh_uniranges af_lao_script_class _Z10lemon_seekili af_deva_uniranges af_kali_nonbase_uniranges FT_FloorFix _ZdlPv af_latb_dflt_style_class FT_Stream_GetUShortLE tt_cmap8_class_rec af_none_uniranges FT_Error_String ps_table_funcs FT_Outline_Decompose FT_Face_GetCharVariantIndex drag af_sinh_dflt_style_class af_taml_nonbase_uniranges __mlibc_entry backgroundColor _ZN4ListIP8Window_sEixEj af_ethi_nonbase_uniranges af_guru_script_class fb FT_Set_Pixel_Sizes af_beng_uniranges FT_Atan2 FT_Get_Charmap_Index af_none_script_class FT_Vector_NormLen FT_Trace_Get_Name t1_cmap_classes FT_Get_CMap_Format tt_cmap10_class_rec af_mong_nonbase_uniranges af_mlym_uniranges FT_Get_Glyph_Name af_glag_script_class FT_Select_Charmap ft_sid_names FT_Outline_Render strtol FT_Property_Set af_cprt_script_class af_grek_titl_style_class FT_Outline_Transform af_hebr_nonbase_uniranges FT_New_Memory af_cyrl_smcp_style_class af_hani_script_class af_latn_uniranges FT_Request_Size keymap_us lastKey active FT_Stream_GetULongLE af_osma_uniranges FT_Stream_GetULong af_goth_dflt_style_class af_cyrl_ordn_style_class FT_Raccess_Get_DataOffsets bdf_driver_class af_copt_uniranges FT_Face_Properties _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm FT_New_Library _Z22RemoveDestroyedWindowsv FT_Get_Module af_latn_c2sc_style_class FT_Stream_Open strrchr _Z14ReceiveMessageP13ipc_message_t af_cari_dflt_style_class af_knda_dflt_style_class memcpy_sse2_unaligned FT_Bitmap_Init af_dsrt_uniranges mouseData af_shaper_get_elem af_tfng_nonbase_uniranges FT_Remove_Module af_lao_uniranges af_cans_nonbase_uniranges af_latb_uniranges FT_GlyphLoader_Reset af_tfng_script_class af_khms_dflt_style_class af_grek_c2cp_style_class FT_Stream_Skip af_adlm_dflt_style_class FT_Get_Font_Format t1_standard_encoding FT_MulFix _Z16memcpy_optimizedPvS_m af_cjk_writing_system_class af_nkoo_dflt_style_class af_cprt_nonbase_uniranges strcat af_mymr_script_class FT_Get_Next_Char FT_Get_Advances af_deva_nonbase_uniranges TT_RunIns af_beng_nonbase_uniranges af_latn_pcap_style_class FT_List_Up FT_Outline_Get_Orientation closeButtonSurface af_shaw_script_class af_dsrt_script_class af_orkh_dflt_style_class af_bamu_dflt_style_class FT_Attach_File FT_Outline_Get_Bitmap FT_Stream_ExtractFrame winfnt_driver_class FT_Trace_Get_Count memset32_sse2 ft_lzwstate_io FT_Bitmap_New af_geor_script_class af_bamu_script_class fseek af_cans_dflt_style_class FT_Stream_ReadFields af_avst_nonbase_uniranges ft_hash_str_insert af_armn_dflt_style_class FT_Vector_Rotate cff_cmap_encoding_class_rec af_cyrl_c2sc_style_class FT_GlyphLoader_New af_arab_dflt_style_class ft_standard_glyph_names FT_Get_TrueType_Engine_Type memchr _Z8DrawCharciihhhP7Surface af_osge_script_class af_telu_uniranges psnames_module_class af_shaper_buf_create ft_debug_init FT_Vector_From_Polar FT_Stream_ReadChar FT_Load_Sfnt_Table _ZN10win_info_tC1Ev af_sylo_uniranges af_grek_sinf_style_class af_grek_uniranges FT_Vector_Unit af_tavt_dflt_style_class af_latn_subs_style_class FT_Stream_Free af_olck_dflt_style_class TT_New_Context FT_Outline_Embolden af_latb_script_class strstr af_arab_uniranges FT_Outline_Check af_latn_dflt_style_class FT_Load_Char af_avst_uniranges ps_builder_funcs af_vaii_dflt_style_class FT_Raccess_Get_HeaderInfo FT_Stream_GetUOffset af_geor_uniranges af_dsrt_dflt_style_class af_gujr_script_class strncmp af_hebr_dflt_style_class _ZN4ListIP8Window_sE6get_atEj FT_Get_Renderer ft_hash_str_lookup af_nkoo_script_class af_grek_dflt_style_class _ZdlPvm _Z18memset64_optimizedPvmm FT_Select_Metrics strncpy FT_Sfnt_Table_Info _Z11PointInRect4Rect8Vector2i FT_Vector_Transform af_dummy_writing_system_class FT_Done_FreeType _Z13PointInWindowP8Window_s8Vector2i FT_Stream_EnterFrame windowCount FT_Set_Char_Size FT_MulDiv_No_Round __cxa_atexit af_cari_nonbase_uniranges _Z8DrawRectiiii10RGBAColourP7Surface af_sylo_dflt_style_class FT_Set_Transform af_latn_c2cp_style_class memcmp mouseDown af_khmr_nonbase_uniranges af_orya_uniranges FT_Matrix_Invert ft_glyphslot_alloc_bitmap af_cyrl_c2cp_style_class af_guru_dflt_style_class FT_Get_Sfnt_Name_Count _Z15DrawBitmapImageiiiiPhP7Surface ft_hash_num_init _Z8DrawRectiiiihhhP7Surface af_osge_nonbase_uniranges isalpha ft_hash_str_init af_telu_dflt_style_class ft_corner_orientation pfr_cmap_class_rec sfnt_module_class FT_Bitmap_Done af_latp_script_class FT_Outline_Copy FT_Cos _Z10DrawStringPcjjhhhP7Surface _ZN4ListIP8Window_sEC1Ev fread tt_cmap13_class_rec af_writing_system_classes af_shaper_get_cluster ft_glyphslot_set_bitmap af_goth_nonbase_uniranges af_style_classes FT_Get_Sfnt_LangTag af_tfng_uniranges af_tibt_script_class t1_cmap_standard_class_rec FT_GlyphLoader_CreateExtra cff_decoder_funcs af_sund_nonbase_uniranges cff_builder_funcs FT_Face_GetCharsOfVariant fopen __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface FT_Matrix_Multiply memset FT_Select_Size _Z15InitializeFontsv main af_ethi_script_class ft_lzwstate_init ftell af_saur_script_class af_bamu_nonbase_uniranges af_buhd_nonbase_uniranges af_ethi_dflt_style_class af_cher_script_class af_vaii_nonbase_uniranges af_beng_dflt_style_class af_hani_uniranges af_goth_uniranges font_default _Z5floord FT_Matrix_Multiply_Scaled af_arab_script_class _ZdaPv t42_driver_class FT_Outline_Get_CBox fclose FT_Add_Module af_vaii_uniranges FT_Get_Color_Glyph_Layer af_cari_uniranges autofit_module_class FT_List_Remove af_cakm_nonbase_uniranges isprint _ZN4ListIP8Window_sED2Ev af_buhd_script_class _ZN4ListIP8Window_sED1Ev ps_hints_apply af_knda_uniranges FT_Outline_Done af_latp_dflt_style_class FT_List_Insert strcmp FT_Set_Renderer _Z11lemon_writeiPKvm memset64_sse2 af_glag_nonbase_uniranges t1_cmap_unicode_class_rec af_mlym_script_class _fini FT_Get_CMap_Language_ID ft_raster1_renderer_class sprintf af_thai_dflt_style_class FT_Matrix_Check FT_Angle_Diff af_adlm_script_class FT_Palette_Select FT_Get_X11_Font_Format af_khmr_dflt_style_class af_mymr_nonbase_uniranges af_thai_uniranges FT_GlyphLoader_Add _ZN4ListIP8Window_sE10get_lengthEv af_geok_dflt_style_class af_deva_script_class FT_Face_GetCharVariantIsDefault af_lisu_dflt_style_class ft_mem_strcpyn af_gujr_uniranges af_olck_uniranges af_vaii_script_class af_tibt_dflt_style_class af_none_nonbase_uniranges af_guru_uniranges ft_glyphslot_free_bitmap FT_Open_Face FT_Property_Get ft_glyphslot_preset_bitmap af_arab_nonbase_uniranges af_cyrl_uniranges af_latb_nonbase_uniranges FT_Attach_Stream ft_service_list_lookup FT_Stream_New ft_hash_num_lookup tt_default_graphics_state af_cher_nonbase_uniranges FT_Bitmap_Convert af_cher_dflt_style_class _Znam FT_Done_Library FT_List_Iterate _Z24CreateFramebufferSurface6FBInfoPv FT_Sin af_mymr_uniranges af_tavt_uniranges t1_expert_encoding af_grek_pcap_style_class FT_Trace_Enable FT_Stream_GetChar FT_List_Find _Z13lemon_readdirimP12lemon_dirent FT_Library_Version FT_Render_Glyph_Internal FT_Outline_EmboldenXY FT_Hypot af_hani_dflt_style_class ft_smooth_lcdv_renderer_class af_olck_nonbase_uniranges af_latin_writing_system_class af_buhd_dflt_style_class af_geok_nonbase_uniranges ft_validator_run FT_CMap_New af_guru_nonbase_uniranges FT_Get_Track_Kerning FT_Match_Size FT_Stream_GetUShort _edata FT_Get_First_Char FT_Bitmap_Copy FT_Gzip_Uncompress _ZN4ListIP8Window_sEC2Ev redrawWindowDecorations af_saur_dflt_style_class af_shaper_get_coverage af_sinh_script_class af_telu_nonbase_uniranges ft_hash_str_free af_knda_nonbase_uniranges af_orya_nonbase_uniranges af_grek_script_class af_grek_ordn_style_class af_cans_uniranges af_copt_nonbase_uniranges t1_cmap_expert_class_rec af_limb_script_class FT_Vector_Length af_lao_dflt_style_class psaux_module_class af_orya_dflt_style_class af_lisu_uniranges FT_New_Face af_tavt_nonbase_uniranges af_geor_nonbase_uniranges af_khmr_uniranges FT_Reference_Library af_thai_script_class FT_GlyphLoader_Done af_latp_nonbase_uniranges af_adlm_nonbase_uniranges af_gujr_nonbase_uniranges af_khms_script_class ft_mem_qrealloc _Z10DrawWindowP8Window_s FT_Get_Name_Index af_taml_script_class af_shaper_buf_destroy FT_Bitmap_Embolden ft_standard_raster _Z10surfacecpyP7SurfaceS0_8Vector2i FT_Get_Module_Interface FT_CMap_Done strlen af_cakm_uniranges toupper ft_grays_raster FT_Stream_OpenMemory ft_corner_is_flat ft_smooth_renderer_class af_cans_script_class af_saur_nonbase_uniranges _ZN4ListIP8Window_sE9remove_atEj FT_Add_Default_Modules af_cprt_uniranges FT_Tan ft_mem_strdup FT_Activate_Size FT_Trace_Disable _Z11lemon_closei t1cid_driver_class af_limb_dflt_style_class font_old t1_cmap_custom_class_rec FT_Get_Postscript_Name af_ethi_uniranges ft_hash_num_insert FT_Stream_Pos af_grek_nonbase_uniranges tt_cmap0_class_rec af_khmr_script_class fbInfo af_shaw_uniranges FT_CeilFix _ZdaPvm memcpy_sse2 af_grek_subs_style_class af_mong_uniranges FT_Library_SetLcdFilter af_cyrl_pcap_style_class windows _Z12RefreshFontsv FT_Outline_New FT_Palette_Data_Get af_sylo_nonbase_uniranges ft_lcd_padding _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i afm_parser_funcs af_armn_nonbase_uniranges  .symtab .strtab .shstrtab .interp .hash .dynsym .dynstr .rela.plt .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .dynamic .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_str .debug_loc .debug_ranges                                                                                 X@     X                                    #             h@     h      �                            )             @@     @      0                          1             p@     p                                    9      B       p@     p                                 C             p	@     p	                                    >             �	@     �	                                  I             �@     �      q�                            O             �F     �                                   U              �F      �     ��                             ]             ��H     ��     ��                             g              `i      `	                                  s             `i     `	                                   z             `i     `	                                   �             (`i     (`	     P                           �             xai     xa	                                 �             �bi     �b	                                    �             �ti     �t	     (                              �      0               �t	     +                             �                      �t	     �                             �                      {{	                                   �                      �{	                                 �                      ��     �                             �                      �.     U�                            �                      �                                   �      0               �     �~                                                �`      ~D                                                 0�2     ��                                                  �`4     ��         G                	                      �5     ��                                                   X�5                                  