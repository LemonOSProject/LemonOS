ELF              ��4   �6      4    (           � ��'  �'           �'  ķķ�   �        �W  �  �                 �    UU���  VW�����_^�Y  �    �i���f�f�f�f�f��L�=L�t$�    ��tU���hL��Ѓ��Í�&    f�Í�&    ��&    ��L�-L����������t(�    ��tU���PhL��҃��Í�&    �t& �Í�&    ��&    ��=`� ugU�d���V�̷S�з��̷����9�s�v ���d����d�9�r��'����    ��t��h���Q~�����`��e�[^]�Í�&    ��&    ��    ��t'U���hh�h���~������	�����&    f�������L$����q�U��Q��  f���/ �E� ����P�  ����h����  ������P��  ���E�<
tơ@�Pjj�E�P��   ��������tك�ht��  ����f�f�f�f�f�f�f��S�  ��.5  ��h   �7  ����t�T$�@   �P��   �P��[Ít& S��  ���4  ��j �t$�V  ����1���x���t$R��������[Í�    S�  �î4  ���D$�p�E  ��1�[Í�&    ��&    S�U  ��~4  ���D$�D$P�t$�D$(�p�7  ��[�f�S�%  ��N4  ���T$��t���D$�D$PR�D$(�p�?  ����[Í�&    S��   ��4  ���t$�t$�D$�p�M  ��[Í�&    �S�   ���3  ��jj �D$�p�!  ��[Í�&    �t& �1�Í�&    ��    1�Í�&    ��    S�e   �Î3  ���t$jj�D$P������[Í�&    �v WVS�|$�/   ��X3  ��W�
  �t$$j��PW������� 9�[^��_����Ë$ÐU��01�WVS�������3  ��(��   �����9�   C�   P���8  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p���1���   �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � �����T  ��X   �g�����&    �t& ��  �1  ǀ`      ���ǀ\      �    �B    ���ǀ      �    �B    �� �ǀ       �    �B    ǀT      ǀX      ǀL      ǀP      ǀD      ǀH      Í�&    �UWVS�������0  ���|$0� ��&    ���T  �   ��X   ��  �w ��  ��t܋�`  �t$�|$0����  �|$0��\  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s��\  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ���`  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$��������B1ҋD$~Q��@�����   ��   �E���  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,����E$���~�� �Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ�������������`  ���K�����  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~�� ��N,����ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��t  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS��������,  ���D$ ����   �P���)փ� C���  �N�A=����~   �y���1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o��\  ����   ��t�J+J�ʋO)�9�|W�  ��[^_]Í�&    �v ��L  ��P   ����� ���� t
f=��t<�u���D  ��H   뱍�&    ���\  롍�&    ���T  ��X   ��[^_]Í�&    �v �G9�`  tU9�ta���t�B�G��t�����G1�)Q���wW�  ���4�����&    �t& �o�������&    ���`  룍�&    �ǃ\      듍t& WVS�t$������H+  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS�2�����[*  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��A  �G�P�������   �P9���   �T$�+  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ�L  ��P   %��� =�� tDf����t=���t8�s
  1���[��^_]Í�&    �p���V
  ����[^_]Í�&    �t& ���D  ��H   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ������$�f���T$1��: t�t& ����< u�Í�    Í�&    ��&    �UWV1�S�P�����y(  ���|$ �l$$�f��D5 �7����U�����7��9��� ����[^_]Ít& �UWVS�t$�\$�L$��t}�A�S9���9���	ЍV�����tm��	Ȩue���ȉڃ��ύ�&    �v �(�����j�9�u����9�t'���B9�v�D�D�B9�v	�D�D�� [^_]Í�&    �ȉٍ<0��&    f�������Q�9�u��͍�&    ��&    VS�4�����]'  ���t$V����ZY�t$�P��������[^ËD$�L$��t& �����t	�8�u�Ð1�Í�&    ��    �D$�8 t��&    ���8 u�Í�&    U1�WVS�������&  ���t$ �|$$���u�'��&    �t& ���.��t��PW�k�������u����[^_]Í�&    �v U1�WVS�P�����y&  ���t$ �|$$���u�'��&    �t& ���.��t��PW��������t����[^_]Í�&    �v WVS�t$�������&  �|$��tV��d  ��WV�����XZWV�k��������d  9�t<1Ҁ8 u��d  ��[^_Í�&    f��  �P�㍴&    ���d  ��u�1���f�ǃd      1���f�VS�\$�t$��8�u"��t(�   ������t��8�t���)�[^Ít& �1�[^)�Í�&    f�UWVS�D$�\$�l$�0���8�u`��t@�<(��u�[��&    ��t,9�t8�����0���8�t�����[)�^_]Í�&    f�1�1�[)�^_]Ít& ���[��)�^_]�����������ōt& �UWVS�����ë$  ���t$ �|$$��t& ��t)�������P�  ����$�}  ��9��t����[^)�_]Í�    UWVS�"�����K$  ���l$0�D$8�t$4�D$���&    �v ��t1;l$t+�����E ��P�  ����$�  ��9��E t����[^)�_]Í�&    ��&    WVS�t$�������#  ��V�������$������4$�����������Pj W�!  XZVW������[^_ÐS�U�����~#  �� j j j �D$ P�t$8j�k  �D$,��8[�f�S�%�����N#  ��j j j j �t$(j�>  ��([Í�&    f�S�������#  �� j �D$P�t$8�t$8�t$8j�  �D$,��8[Í�&    ��&    S�������"  �� j �D$P�t$8�t$8�t$8j��  �D$,��8[Í�&    ��&    S�u����Þ"  �� j �D$P�t$8�t$8�t$8j�  �D$,��8[Í�&    ��&    S�5�����^"  �� j �D$P�t$4�t$<�t$8j�G  �D$,��8[Í�&    ��&    S�������"  ���t$�t$�t$�������[Í�&    �t& S��������!  ���t$�t$�t$�������[Í�&    �t& S�����þ!  ���t$�t$�t$� �����[Í�&    �t& S�e����Î!  ���t$�t$�������[Í�&    ��&    �S�5�����^!  ���t$�������1�[ÐS������>!  ��j �t$�������   ��u
����[Ív ��P������1҃���[�f�f�f�f�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��S�����þ   ����D��0�t$������[Í�&    �t& S�e����Î   ����D��0�t$������[�f�f�f�f�f���T$�   �JЃ�	v���1���A����ËD$��߃�A������Í�&    �t& �1��|$z��Ít& �1��|$@��Ít& ��D$��0��	����Í�&    ��&    ��T$�   �JЃ�	v���1���A�����Í�&    ��&    ��D$��!��]����Í�&    ��&    ��T$�� ����	��	���Í�&    �v Í�&    ��&    �1�Í�&    ��    VS�$�����M  ���t$V��������u��[^Í�&    f���V��������������[^Í�    �D$��_Í�&    ��D$�� �f�f�f�f�1�Í�&    ��    �����  ��`��  1�Í�&    �v S�����î  �� j j j �D$ P�t$8j�����D$,��8[�f�1��f�f�f�f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f��ķ���t6U��S�ķ����&    �v �Ѓ�����u��[]Í�&    ��&    �������  
Lemon:  > test1234

         zR |�         e����    D Gu Cu|   $   @   ����<    A�NE H^A�  4   h   ����:    A�NBD HKDA HCA�       �   ����"    A�NG HC� (   �   ���.    A�NJDG HA�   ,   �   ���9    A�NKJAG HCA� (      ���(    A�NDDG HA�   (   L   ���$    A�NBBG HA�      x  $���          �   ���       (   �  ���&    A�NDBBE HA�@   �   ���;    A�A�A�RA I$B(C,A0HC�A�D�        ���       D   $  ����   A�F�A�A�N<Z@J0�
A�A�A�A�M      l  P����       T   �  �����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `   �  t����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   <  �����    A�A�A�WA H��A�A�  �   t  x����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0     ����            ����!       @   ,  ����K    A�A�A�C�N Z,A0K JC�A�A�A�8   p  �����    A�A�A�A��
�A�A�A�H   4   �  @���0    A�A�NE FADC HC�A�   �  8���#          �  T���       D     `���V    A�C�A�A�N j(A,A0H GC�A�A�A� D   T  x���V    A�C�A�A�N j(A,A0H GC�A�A�A� D   �  �����    A�A�A�`AA HAAA H\
�A�A�J ,   �  ����G    A�A�w
�A�FC�A�  \     �����    A�A�A�A�M
�C�A�A�JE
�C�A�A�FD
�E�A�A�A @   t  (���Z    A�A�A�A�N ^,A0U MA�A�C�A�@   �  D���r    A�A�A�A�N0u<A@U0NA�A�C�A�L   �  ����O    A�A�A�RA ]DBA FAAA HA�A�A�   0   L  ����.    A�N(B,B0B4E8D<B@LA�  0   �  |���'    A�NBB B$B(D,B0HA�  0   �  x���2    A�N(B,E0D4D8D<B@LA�  0   �  ����2    A�N(B,E0D4D8D<B@LA�  0     ����2    A�N(B,E0D4D8D<B@LA�  0   P  ����2    A�N(B,E0D4D8D<B@LA�  (   �  ����%    A�NDDD HA�   (   �  ����%    A�NDDD HA�   (   �  ����%    A�NDDD HA�   $   	  ����!    A�NDD HA�      0	  ����    A�ND HC� 8   T	  ����E    A�NBD HL
C�DCA HEC�(   �	  ����!    A�A�A�[�A�A�$   �	  ����%    A�NHD HA�  $   �	  ����%    A�NHD HA�     
  ����            
  ����          4
  ����          H
  ����          \
  ����          p
  ����           �
  ���          �
  ���          �
  ���          �
  ���          �
  ���       D   �
  ���J    A�A�NE HG
A�A�JCA HHD�A�     0  ���          D  ���          X  ���          l  ���       0   �  ���.    A�N(B,B0B4E8D<B@LA�     �  ���       <   �  ���   A�A�A�A�C �
C�A�A�A�A 8     �����    A�A�A�A��
�A�A�A�P       ����    ����                    i�r�                                                                                @� � �GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o                      t�          ��          a�          i�          ��          ķ          ̷          Է          �     	     `�     
                           ��   ķ         ̷      (   ��      ;   ��      =    �      P   P�      f   `�    
 u   d�    
 �   Ё      �   h�    
             ���   ȷ      �   ��      �    �      �            ��  ��                  ��           ���           ��  ���    1  �    	 <  �    	 H  (�    
 W  4�    
 a  0�    
 k   �    
 x  �    
 �           ���  8�    
 �           ���           ���           ���           ���           ���           ���           ��             ���  Է      �  �%       �    
   P�K     �  D�    	    �    
 "  ��!     *  @��     8   �     (  `�    
 H  ��2     S  `�     [  ���    
 l   �     	 t  p��     {  �    
 �  L�    	 �  з     �  @�%     �  P�.     �  ��     �  ��     �  0�     �  ���    �  �     �  �    	 �  ��J     �  @�     �  @�     
 �   �       �%     
  ��r       �      2  t�        �     -  А     5  ���     O  ��%     <  p�0     C  ��(     I  �2     �  @�    	 �  ��&     U  �    	 N  ��%     g  ��     o  ���     w   �.     �  ���     �   �Z     �  p��    �  ���     �  ��     �  ��<     �  ��     �  P�.     �   �O     �  ��:     �  L�     
 �  `�    �  ��     �  ��$     �   �     	    �"        �       p�        p�     %  �    	 2  @�G     9  a�      ?  P�V     m  H�    	 G  P�     U  @�&     [  З     c  ��9     j  ��E     q  L�     	 x  d�     
 }  0�2     �  �     �  �V     �   �!     �  @�!     �  И     �  ��'     �  ��#     �  p�;     �  p�2     �  p�     P  Њ�     crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp fileio.c allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns string.c p.1056 filesystem.c syscall.c stdstreams.c stdout.c ctype.c _liballoc.c memory.c _GLOBAL_OFFSET_TABLE_ putchar l_allocated strcpy l_max_inuse syscall liballoc_init liballoc_unlock lemon_read isblank currentDirectory _stderr memcpy l_inuse __TMC_END__ __DTOR_END__ lemon_open islower tolower feof malloc __x86.get_pc_thunk.ax __dso_handle ispunct isspace _stdin fflush lseek strncasecmp isxdigit liballoc_lock strrchr calloc strcat fseek lemon_write promptStringStart isupper strncmp liballoc_alloc strncpy strcasecmp realloc strtok __x86.get_pc_thunk.bx fdopen isalpha fread strdup fopen __bss_start memset main ftell _stdout fclose isgraph isalnum isprint promptString strcmp _fini strcspn liballoc_free fputc isdigit fwrite access _edata _end lemon_seek iscntrl strspn strlen toupper lemon_close strchr fputs lemon_readdir  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .ctors .dtors .got.plt .data .bss .comment                                                   t�t                     !         ���   �                 '         a�a                    -         i�i                    5         ���  D                 ?         ķ�'                    F         ̷�'                    M         Է�'                   V         ��'  l                   \         `�L(                    a      0       L(  +                               x(  �     3         	              H1  �                               6  j                  