ELF          >    x @     @       0          @ 8  @                   @       @     �       �               UH��S�� @ �   H���i��Test ELF         zR x�        ����    A�CA�GCC: (GNU) 8.2.0                                  x @                   � @                   � @                                       ��                     x @                 � `                  � `                  � `              main.c __bss_start _edata _end  .symtab .strtab .shstrtab .text .rodata .eh_frame .comment                                                                                  x @     x                                     !             � @     �       	                              )             � @     �       4                              3      0               �                                                          �       �                           	                      �                                                           �      <                              