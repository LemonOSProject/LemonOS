ELF              ��4   B      4    (  
         � ��.  �.            0   � �`  �                    �=  ��U��8�i�mN�A90  �8��8���%�  ]�U��S���l��0�9�sy�U��E��j j j RPj��  �� �E���    �`��d�)�Ӊȉ�i��  �M��h�)щ�¡l�Уl��E��    �`��d��E�h��x����l�    ��]���U��WVS����j�  ���ǃ�W�  ���=t��t��E�   �E�   ���u��u�P�  ���t��	   �   ��VSP�  ����e�[^_]�U��WVS��  fǅ���� fǅ���� fǅ����@ fǅ����  ǅ����    ��j��  ���Ã�S��  ���t��t��   �   ��WVP�  ���t�ǅH���	   ǅL���   ����L�����H���P��  ���E�    �}�.�E�    �}��E����E�����  �E��߃E��̃�������P�  ���E����������|���P�  ��������tw��������u��p���t�p� �P���������=  t)=  w	=
  t�=  t=  t��E�    ��E�   ��E�   ��E�   ��n����p�����  �E�    �}�.�E�    �}��E����E�����  �E��߃E��̡<��@������� �E�    �t���P�%  ��9E�����t[�t��EЍ������PQR�
  ��������t��EЍ������PQR��  ��������������� �E���E�    �}���   �E�    �}���   �Eč��   �E����E����� ����"����E����E����� ����!��؋E����E����� ���� ��ЋE������E���WVSRjjQP�=  �� �E��[����E��A����}���   �}��}� t�  �}��W  �}���  �  �t��t���P�  �����������RSP�  ���t��t��������j RP�  ���������P����t���$�����j RP�Z  ����(�������T�������T�����P���S�}  ����  �t��t���P�  ������,�����RSP�`  ���t��t���4�����j RP��  ����4�������X����t���<�����j RP�  ����@�����\�������\�����X���S��  ���D  �t��t���P�g  ������D�����RSP�  ���t��t���L�����j RP�9  ����L�������`����t���T�����j RP�  ����X�����d�������d�����`���S�5  ���   �t��t���P��  ������\�����RSP�  ���t��t���d�����j RP�  ����d�����h����t���l�����j RP�n  ����p�������l�������l�����h���S�  ����t���t�����j RP�+  ����t����t���|�����j RP�
  ���U��������� <t~�t��E���j RP��  ���E���x_�t��E���j RP�  ���E���x@�t��E���j RP�  ���E��� �t��E���j RP�~  ���E���~�   ��    ��t]�p��E��   ��Ph�   h�   h�   j j h���  �� �E��   �Eċ@��j j j RPj�  �� �  �t��E���j RP��  ���]��t��E���j RP��  ���U��������� <������   �t��E���j RP�  ���]��t��E���j RP�  ���U���������  �����������������<��@��t�ǅp���    ǅt���    ����t�����p���P�h   ���E��   �Eċ@��j j j RPj�  �� ����������U��E�     �E�@    �]ÐU��E�     �E�@    �]ÐU���(��j�s  ���E��E�    �E�    �E�    �E�    ���E�P�������E�U��U�P�U�P�U��P�M�E�U�A�Q�E� ��u
�E�U���E�@�U��E�P�E�P�E�U�P�E�@�P�E�P��ÐU��E�@]ÐU����E�@9Er�    �M�P� ��Q�6�E� �E��E�    �E�;Es�E�� �E��E���M�E��P�@��Q�E�� U����E�@9Er�    �M�P� ��Q�   �E� �E��E�    �E�;Es�E� �E�E���E�P�@�E�U�E� ��t�E� �U�R�P�E�@��t�E�@�U���} u
�E��E��E�@�P��E�P�E�@9E����t�E�P�E�P���u���	  ���M�E�U��Q�E�� U���(��j�m  ���E��E�    �E�    �E�    �E�    ���E�P�������E�U��U�P�U�P�U��P�M�E�U�A�Q�E�@��u�E�U�P��E� �U�P�E��E��E�U��E�@�P�E�P���U����'  #  �E�    ��U�E�ЋU��E��E�;Er�E��U�����  �"  �E�E�E�E���U��B�E��E�H�M���m�}w��E�E��E��E���U��B�E��E��H�M����m�} uߋE��U��WVS���  ��W"  �E���E�E���D   �E�    ��Ѕ�u��D   �E�    ���E����D   �E�    �����E䋃H   9E�s	��H   �E���u��A  ���E��}� u%���  ���  ���� ���  ���  �    �l�E��     �E��@    �E��U�P��D   �E�E��P�E��@   �E��@    �E��@�ƿ    �����P� ��������Q�E��e�[^_]�U��WVS��L�Y  ��1!  �E�    �E�    �E�    �E�    �E�E��E� �,  �}� u5���  ���  ���� ���  ���  �  ��j�������  ���  ��u-���u��K��������  ���  ��u��
  �    �{  ���  �E��E�    ���  ���C  ���  �P���  �@)ЉE��E�    �E����    ;E؉�E��
  ���  �E��E�   ��  �EЋP�EЋ@)ЉE��E��    �M�9E��s�EЉ��  �E��E��E�    �E���9E�sk�EЋ@��t�EЋ@�E��  �}�u���  �E��E�    �|  ���u��9������EЉP�EЋ@���d  �EЋ@�UЉ�EЋ@�EЋEЋ@���  �EЃ��EЉP�EЋ@�@����EЋ@�     �EЋ@�@    �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eȃ}� t�   +EȉEȋUԋE�ЉEԋEȍP�Eԃ���  �E��@  �EЋ@�E��E�)E��m��E���9E��"  �EЍP�EЋ@��EЋ@� �UЋR�P�EЋ@��EЉP�EЋ@�@����EЋ@�     �EЋ@�UЉP�EЋ@�U��P�EЋ@�U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�EЋ@���EԋEԃ��EԋEԃ��Eă}� t�   +EĉEċUԋE�ЉEԋEčP�Eԃ���W  �E���  �EЋ@�E��t  �E̋@���>  �EЋP�E�ЉE��E�)E��m��E̋@)E��E���9E��  �E̋P�E�Ѓ��ẺP�E̋@�Ủ�E̋@�E̋E��@    �E��@����E̋UЉP�E̋U��P�E̋U�P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�����0�x�����P� 9Ɖ��s�Ɖ������0�x�Ẽ��EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��  �E̋@���  �E̋@�E��E�)E��m��E̋@)E��E���9E���   �E̋P�E�Ѓ��E��E��@����E̋P�E��P�E��Ủ�E��U��P�E��U�P�E��UЉP�E̋@�U���E̋U��P�EЋP�E�ЍP�EЉP�u��    �����P� ��������Q�E����EԋEԃ��EԋEԃ��E��}� t�   +E��E��UԋE�ЉEԋE��P�Eԃ����  �E��   �E̋@�Ẽ}� ������EЋ@��uC�}�u���  �E��E�    �4���u���������EЉP�EЋ@��t#�EЋ@�UЉ�EЋ@�EЃ}� ���������X  �    �e�[^_]�U��WVS��,�%  ���  �} u#���  ���  ���� ���  ���  �9  �E��� ���E�}�w	�E+E�E��  �E���E��E��@=���tx���  ���  ���� ���  ���  �E��@%��� =�� t �E��@��=��  t�E��@��=�   u���  ���  ���� ���  ���  �b  �  �E��@�E������P� �M��I�ο    )��������Q�E܋P�E��@)ЍP�E܉P�E��@�ޭދE��@��t�E��@�U����E�� ��t�E�� �U��R�P�E�� ��u�E��P�E܉P�E܋@����   ���  9E�u�E܋@���  ���  9E�u
ǃ�      �E܋ ��t�E܋ �U܋R�P�E܋@��t�E܋@�U܋������P� �M܋I�ο    )��������Q�E܋@��P�u��y  ���G���  ��t=���  �P���  �@)ЉE؋E܋P�E܋@)ЉEԋE�;E�~	�E܉��  ��  �e�[^_]�U��S���  �  �U�U�U�U��R���%������E��E��Pj �u��?������E��]���U��S���^  ��6  �} u���u�������    �1  �} u���u��������  �E�E�E��� ���E��}�w	�E�+E��E���   �E���E�E�@=���tz���  ���  ���� ���  ���  �E�@%��� =�� t �E�@��=��  t�E�@��=�   u���  ���  ���� ���  ���  �   �    �_�E�@�E�E�;Er�E�U�P�a   �E�;�W   ���u��������E���u��u�u����������u��������E�]��Ë$Ë$�U��������  �    ]�U��������  �����  �    ]�U��S�������  �M�U��j j j QRj���   �� �E�]���U������e  �    ]�U��WVS�r���N  �E�]�M�U�u�}�i�[^_]�U��S���G���#  �M�U��j j j QRj�������� �E�]���U��S�������  �U�U�U�U���j j �u��u��uj���j����� ��]���U���������  �E�������E����	��E����	��E��	ЉE�E�@�E��E�    �E9E�}G�E�    �E9E�}2�U�E�E�@�M�U��Ѝ�    �E�E��E��ƃE�뱐��U��S���0���  �U��j j j j Rj �������� ��E�]��� U���������  �M�U�E �M�U�E�} y�EE�E    �} y�EE�E    �E������E���	��E�	ЉE�E$�@�E��E�    �E�;E}k�U��EE$�@9�}Y�E�    �E�;E}D�U�E�E$�@9�}2�U��EE$�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��������  �} y�EE�E    �} y�EE�E    �E�������E����	��E��	ЉE�E�@�E��E�    �E�;E}k�U��EE�@9�}Y�E�    �E�;E}D�U�E�E�@9�}2�U��EE�@�M��U�Ѝ�    �E�E��E�봃E�덐��U��� �1���  �E�E�E�E��E��}��E��f�E��m��]��m��E��E�������v�E�����E���U��S��4�7  ���  �U���������P��H����E��Eԃ��d$��$���l��������E��E�    �E�   �E�    �E�;E��   �E�    �E�;E��   �U�E�E�@�������U�E���E�ȉE��U���ЉE�E��E�P�E�����U���ЉE�ЍP�E��E�@�U�������U���ЉE�ЍP�E��E�@�U�������E��F����E�E�E��$�����]��Ë$�U��WVS��<������r  �u�M�U�}���EԈMЈỦ��E��E�    �}���   �U���`���E��� ���E��E�    �}�]�E�   �����#E܉E������Ѕ�t7�}��u��MЋE� �EE�EċE�E��u WVQjjRP������� �E�띃E��f�����e�[^_]�U��WVS��,�����  �EȋM�U�E�MԈUЈE��E�    �E� ��tC�}��u��]ԋM�U�EЉE� �����u WVSQRP�]������� �E��E볐�e�[^_]�U��S���9���  ���u����������]���U��S�������  ���u���������]���U��S��������  ���u����������]���U��S��������  ���u����������]���U��S������{  ���u���^�������]���U��S���x���T  ���u����������]���U��S���Q���-  �M�U��j j j QRj�������� �E�]���U��S�������  �U��j j j j Rj!�������� ��]���U��S��������  �M�U��j j j QRj���M����� ��]���U��WVS��,�����Ï  ���u�E������E��h�   �J������Ɖ��    �*   ����V�  ���u��E��U�P�E��U���ֺ   �ǉ��E�@���EЋE�@���EԋUЋE�������P�������E܋E��Uȉ��   �Ủ��   �UЉ��   �Uԉ��   �U؉��   �U܉��   �E��e�[^_]�U��VS������å  �E�@��P�������u��t��V�?  ����h�   V��������e�[^]�U��S���}�����U  �E���   �E�@�ЋE�@����Q�M���   RPj j �"����� �E�    �E��P�L  ��9E�����t0�U�E��RP�E  �����M���   ��QP�҃��E�뷋E���   �E�@��RP���������]���U��S��$������Ù  �E�    �E��P��  ��9E�������   �U�E��RP�  ���P�U�P�U�P�U�@�E��U�E9�}Y�U�E9�}O�U�E�E9�~@�U�E�E9�~1�U�E��RP�`  ��������P�҃��E�U􉐤   �	�E��L�����]���U��S��������
  �U���   �ыU��QR���  ��������P�҃���]���U��S�������
  �U��R���Y   ���Eƀ�   ��Eƀ�   ��Eƀ�   ��Eƀ�   ���]���U��S���V���2
  �U��R���-   ����]���U���2���
  �E�     �E�@    �]ÐU��S���������	  �E� �E�E� ��t���u��������琋]��ÐU��������	  �E�@]ÐU��������	  �E�@9Er	�    � �+�E� �E��E�    �E�;Es�E�� �E��E���E��@�� Game Over, Press ENTER to Reset        zR |�        ����'    A�Bc�      <   �����    A�BD���� (   `   ���u    A�BF���h�A�A�A�   �   b���G   A�BI���   �   ����    A�BU�     �   ����    A�BU�     �   ~����    A�B��      ���    A�BG�     ,  ����b    A�B\�    L  <����    A�B��    l  ����    A�B��    �  ����7    A�Bs�     �  ����r    A�Bn� ,   �  ����&   A�BF����A�A�A�   ,   �  ����4   A�BF���'�A�A�A�   ,   ,  ����~   A�BF���q�A�A�A�       \  C���K    A�BD�C��     �  j���f   A�BD�^��   �  ����          �  ����          �  ����    A�BP�     �  ����    A�BY�        }���6    A�BD�n��     0  ����    A�BP�  (   P  ����*    A�BC���`�A�A�A�     |  ����6    A�BD�n��      �  ����?    A�BD�w��     �  �����    A�B��     �  0���7    A�BD�m��       C����    A�B��    (  ����    A�B��    H  ����Q    A�BM�     h  ����C   A�BD�;��   �  ���       (   �  ����    A�BF�����A�A�A�(   �  �����    A�BF���x�A�A�A�    �  ���&    A�BD�^��        ���&    A�BD�^��      @  ���'    A�BD�_��      d  ���'    A�BD�_��      �  ���'    A�BD�_��      �   ���'    A�BD�_��      �  #���6    A�BD�n��      �  5���2    A�BD�j��        C���4    A�BD�l��      <  b���P    A�BD�H�� (   `  /����    A�BF�����A�A�A�    �  b���(    A�BD�`��  $   �  ����N    A�BB��F�A�A�    �  �����    A�BD����     �  �����    A�BD����        :���D    A�BD�|��     D  ����#    A�B_�      d  ����9    A�BD�q��     �  ����    A�BQ�     �  ����Q    A�BM�                                                                                                                                                                                                                                                                                                                                                                                                             `�`�@@@�@@@�@@@�d   �                                                                                                                                                                                                                                                                                                            <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;              GCC: (GNU) 8.2.0                        ��          ��          Ц           �           �          `�                                ���  ��                   ���            ��   ��        ��     (   D�     3   H�     ?   ��     N   ��     [   ��     n   �7     ~   )�r     �   ��&    �   ��4    �            ���            ���            ���            ���            ���            ��             ���    �        |�       ��     )  �7     ;  t�     A  ǡ6     `  D��   "  �  $�   "  �  ��     �  ��2     �  ��*     �  �9   "  �  @�     �  њ6     �  ��     �  ߠ&       �9   "    ��     "  �?     .  ���     F  ��4    M  >��   "  n  $�     �  l�     �  ¥(   "  �  +�'     �  ���     �  [��     �  ¥(   "  �  ,�     �  0�     �  $�   "    �#   "  2  s�K     9  r�P   "  H  p�     Q  r�P   "  `  4�     o  
�   "  �  ���       ��      �  <�     �  ]�6     �  R�'     �  ��f    �  ��     �  (�       ��       c��     1  9�C    T  ��     p  Q�N     �  8�     �  ^�Q   "  �  Z��     �  \��   "  �  M�u     �  `�       `�        F��     8  h�     H  `�     U  �Q     _  y�'     f  
�   "  ~  /�4     �  ��'     �  ��     �  G    �  �&     �   �     �  ��b   "  �  `�      �  ��      �  .�D       �   "  3  �#   "  J  ��'     R  H�   "  �  ��~     snake.asm main.cpp l_memRoot l_bestBet l_pageSize l_pageCount l_warningCount l_errorCount l_possibleOverruns liballoc_memset liballoc_memcpy allocate_new_page malloc.localalias.0 _liballoc.c syscall.c ipc.c graphics.cpp text.cpp window.cpp _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx l_allocated _Z12GetVideoModev snake _Z13_CreateWindowP10win_info_t _ZN4ListI8Vector2iE9add_frontES0_ _ZN8ListNodeI8Vector2iEC1Ev l_max_inuse _Z14_DestroyWindowPv syscall _ZN4ListIP6WidgetED2Ev liballoc_unlock ReceiveMessage _Znwm _ZN4ListIP6WidgetED1Ev l_inuse SendMessage _Z11PaintWindowP6Window malloc _ZN4ListI8Vector2iE8add_backES0_ __x86.get_pc_thunk.ax tickCounter _ZN6WindowD1Ev _ZdlPv _Z4Waitv _Z15HandleMouseDownP6Window8Vector2i _ZN6WindowD2Ev liballoc_lock frameWaitTime _ZN8ListNodeI8Vector2iEC2Ev _ZN4ListIP6WidgetEC1Ev calloc _ZN6WindowC1Ev gameOver _ZN6WindowC2Ev timerFrequency _ZN4ListI8Vector2iEC2Ev _Z8DrawCharciihhhP7Surface applePos liballoc_alloc _ZdlPvm realloc _Z8DrawRectiiii10RGBAColourP7Surface __x86.get_pc_thunk.bx snakeMapCells _Z12CreateWindowP10win_info_t _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window rand_next _ZN4ListIP6WidgetEixEj _Z10DrawStringPcjjhhhP7Surface _ZN4ListI8Vector2iE9remove_atEj _Z5Resetv lastUptimeSeconds __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface lastUptimeTicks font_default _Z5floord _ZdaPv _ZN4ListI8Vector2iEC1Ev _Z12_PaintWindowPvP7Surface _Z4randv liballoc_free pmain _Znam snakeCellColours _ZN4ListI8Vector2iE6get_atEj _edata _end _Z13HandleMouseUpP6Window _ZN4ListI8Vector2iE10get_lengthEv _ZN4ListIP6WidgetEC2Ev _ZdaPvm _ZN4ListIP6WidgetE10get_lengthEv  .symtab .strtab .shstrtab .text .rodata .eh_frame .got.plt .data .bss .comment                                                   ���   /&                 !         ���&                     )         Ц�&  �                 3          � 0                   <          � 0  @                  B         `�`4  \                  G      0       `4                                 t4  �  	            	              T;  s                               �A  P                  