ELF              ��4   P�      4    (           � �^  ^            `   � ��
  �        �W  �@  �                 �    UU���R+  VW�����_^�g  �    �i���f�f�f�f�f����=��t$�    ��tU���h���Ѓ��Í�&    f�Í�&    ��&    ����-�����������t(�    ��tU���Ph���҃��Í�&    �t& �Í�&    ��&    ��=�� ugU�����V��S���������9�s�v ����������9�r��'����    ��t��h���Q~��������e�[^]�Í�&    ��&    ��    ��t'U���h��h���~������	�����&    f������U��S��   ������L���Pj R�:  ���E��E�    �E�    �E�    �}� ��  �E����EԋE���E��E�`   �E�H   ��hp  �V  ���Ã��u��u��u��uԍ�L�����PS�\  �� �]�E�ƀ�   /�E�ƀ�    �E��   ����L�����RP�5  ���E��   ��P�3  ���P��E����   <fuy�E��   ��P�3  ���P��E����   <euS�E��   ��P�]3  ���P��E����   <lu-�E��   ��P�73  ���P��E����   <.u�   ��    ��t�E��@a�E�ǀ�      �EЃ�u�E�ǀ�      ����P�u��#  ���E��E���у���L���RPQ�9  ���E�E�d�E��Pc�$���9��F����E�L�E�    �6�����]��ÍL$����q�U��VSQ��<�ȋ �E�f�$��f�&��f� �2 f�"�2 �(�    �,�File�0� Man�4�ager�8� ��h ��c  ������j h\��7  ������h^�h`���#  ���E���u���$  ���E����u���'  ��� �� ��u�j�u�P�$  �����u���#  ����h^�hj��r#  ���E���u��q$  ���E����u��`'  �������u�j�u�P�#  �����u��g#  ����h^�hw��#  ���E���u��$  ���E����u�� '  �������u�j�u�P�E#  �����u��#  ���4������E�P�s8  ����������   �EЃ�u��y�EЃ�u����P��   ��뾋EЃ�u2�E���f�EދE�f�E��Eމ��E܉ơ���VSP�  ��넋EЃ��x�������P�  ���q8  ���[�������P�  ����D���U����}u�}��  u��h ��!   �����U�����h��  j��������ÐU��Ef�   �Ef�@  �Ef�@  �Ef�@  �]ÐU����E���u�u�u�u�uP�  �� ����E��Eǀ�       ���U����E�@ �E�@a��t�E�   ��j j j j Pj�E7  �� �E���   ��uP����P�f4  ����    �E�   ��j P�4  ��������t����P��  ����ÐU��VS�E�@���r  �E�@��������X��E�@�H��E�@�P�E�@���uh�   h�   h�   SQRP�4  �� �E�@��������X��E�@�H��E�P�E�@�������E�@���uh�   h�   h�   SQRP��  �� �E�@�H��E�@�U�R���uj`j`j`jQPR�  �� �E�@�H��E�P�E�@ЍP��E�@���uj`j`j`jQRP�t  �� �E�@�H��E�@�P�E�@�uj`j`j`QjRP�F  �� �E�@�H��E�@�P�E�X�E�@؃��uj`j`j`QjRP�  �� �E���   ��u@� ��E�P�E�X�E�@�������؃����uQj0j0RP�u  �� �   �E���   ��u=���E�P�E�X�E�@�������؃����uQj0j0RP�'  �� �I�E���   ��u;���E�P�E�X�E�@�������؃����uQj0j0RP��  �� �E�P�E�@Ѓ��ËE�P�E�@�������E�@X��)ЉE�����uj j j SRP�v  �� ��e�[^]ÐU����E� �E�E� ��t�E� �E����u���%  ���E��E��ًE�     �E�@    �E�@    ���f�f��UWVS��  �ÓU  ���|$$�D$ �l$(	��t��UW�t$,�*  �������)�����RW�t$,�  ����u
��[^_]�f����VW�t$,�V�}*  ����[^_]�f��T$�D$�Í�    �T$�Í�&    �v S�3  ���T  ��h�  ��������� [��Í�&    �t& �VS�  ���T  ���t$��&    �t& �������t�������Vh�  �t�����[^Í�&    ��&    VS�
  ��uT  ���t$�> t-��&    �[�����t����F���Ph�  �"������> uڃ�[^Ít& UWVS�`
  ��#T  ���t$ �|$$�T$(��   t*�B���t�v ���>�����u��[^_]Í�&    �t& ������R��WV�-  ����tӉ>��t̉~��tĉ~��[^_]Í�&    �t& ���1��|$�D$�D$��f�D$�l$�T$�l$�D$�D$�D$������)�Ð�	  WS  UWVS��,�T$H�|$@�D$�t$T�D$P�l$D�L$L�T$��y�1��T$��y�1���Ё�   ���	ډ�% �  ����	�	ËF�\$�D$��~v;n}q�D$�t$T����D$�D)��l$T�D$���&    ���9u~C�]��)�;\$OD$��P�t$�E�L$ ����������P�\$�N�����;t$u���,[^_]Í�&    ��    VS�  ��UR  ���t$j j j j Vj �\0  ��$��[^� f��`  'R  UWVS��,�|$@�t$D�D$�L$L�D$P�\$T�T$X�l$\��y|$H1���y�1�����������	�	E�T$�D$��~\;u}W�D$H��D$�D��D$�
f���9u~9�]������)�;\$OT$H��R��t$�L$ ��P�\$�H�����;t$u���,[^_]Í�&    �  WQ  UWVS��,�t$@�l$D�D$�L$L�D$P�|$T��yt$H1���y�1��؉������� �  ��	�	G�T$�D$��~i;o}d�D$H��D$�D��D$��t& ���9o~C�G�_������)����;\$OT$H��R�t$�L$ ���P�\$�n�����;l$u���,[^_]Í�&    ��    UWVS�  ��sP  ��<�D$`�l$\�|$T�t$d�@
�D$ �D$X�@���B>��H����T$�D$�$�������D$,�E�������   ;~��   D$D$P�D$�D/��T$H�D$�D$@�D��D$��&    �v �D$H����   �N9L$@��   �T$@�D$�T$�U��&    f��n�T$�L� �n�ύ��\ �^�P�T�^�P�T�L$9L$t7�D$�N���T$9�~$���u��xu��xu��L$9L$uύ�    9|$t�T$��)T$9~�F�����,[^_]Í�&    ��&    UWVS�@  ��O  ��L�l$p�t$`�|$x���������yt$h1��L$d��y�L$dL$l�D$d    �L$h���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$hf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��P�t$|j�t$|W�,����� 9t$h�_�����L[^_]Í�&    UWVS�p  ��3M  ��L�l$p�L$`�t$d�|$x���������y�L$`L$h�D$`    ��yt$l1��L$l���k  ;w�b  �L$t�|$x����f�L$���D$��f�L$�D$�T$�T$t���D$lf�������\$�D$f�T$�����\$�D$f�T$�D$�D$�D$t�����\$�D$f�D$�����\$ �D$f�D$�D$�������1��l$x�D$�����\$(�D$�\$0���&    �t& ��9}��   �t$�D$��U�D$�|$B���D$�D$B��f�D$@�l$@�\$>�l$B�D$>��P�D$ ���D$(�l$D�\$B�l$F�D$B��P�L$4�D$<�l$H�\$F�l$J�D$F��Pj�t$|W�t$|�\����� 9t$l�_�����L[^_]Í�&    UWVS�  ��cK  ���l$4�|$0�L$8�T$<�E��~v�G)Ѕ�~m��    ��1��T$�D$�|$4��t& ��E+D$9�~D�G����    ��Q�O���MP�T$�E���2����D$EP�9�����9w���[^_]Í�&    f�UWVS���D$,�l$(�t$4�|$0�@�t$�D$�E�D$�D$,�X����   �E)�����   �D$,�t$�$    �H��&    f���~i�U��)���~^1����&    ��    �U��)�9�~;�$�t$��Ë��������   u�T$�ʋL$���T$,�J��9�|��D$,�X�$�$9�}�E�D$+D$;$�s�����[^_]Ë$Ë$�f��S�   ������ñI  ���D$��D�P�  ��[Í�&    �S������ÆI  ���t$�  ��[Ív S������fI  ���t$�H  ��[Ív S������FI  ���t$�������[Ív S�c�����&I  ���t$�  ��[Ív S�C�����I  ���t$��  ��[�f��UWVS� ������H  ���D$<�|$8�t$0�D$�G�D$�D$D�������D$�D$@�D$�j��&    f���@   ��   ��    ��   ��   ��   ��   �  ��   �)  ��   �P  ���w  ��9|$��  �.���y��t$H�t$�t$�L$QjjW�t$P������� ��@   �s����t$H�t$�t$�L$QjjW�D$P�HQ������ ��    �L����t$H�t$�t$�L$QjjW�D$P�HQ������ ��   �%����t$H�t$�t$�L$QjjW�D$P�HQ�M����� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������� ��   ������t$H�t$�t$�L$QjjW�D$P�HQ������ ��������t$H���t$�t$�D$PjjW�D$P����P�~����� 9|$�b�����[^_]Í�&    f�UWVS������ÃF  ���D$@�t$0�|$4�l$D�D$��D$<�D$��t3��&    ������t$LU�t$�t$�t$LW��Q�?������ ��uՃ�[^_]�f�f�f�f�f�f��Ð��&    ��&    Ð��&    ��&    �D$�@Ð��    �D$�@Ð��    �D$�@ Ð��    UW1�V1�S������ïE  ���l$0�t$4h�   h�   h�   �u�u�u�u�R����E�D$,�� �l$0���|$0�D$    ��t& �|7
t^�����t$�J  ��9�~S���t$8��  P��  P��  P�D$GP�G��P�D7P�����G�� ��9���D$1��f��|$0��l$0�O�t$4j j j jj�t$ Q������ �t$4h�   h�   h�   �ujj �E��P�r����� �t$4h�   h�   h�   jjj�E��P�J����� �t$4h�   h�   h�   jj�E��P�E��P������<[^_]Ð�t& U1�WV1�S�l�����/D  ���|$0�D$    �G���&    f��<0
tN����P��  ��9�~G���t$8j j j �D$ GP�G��P�G�0P������G�� ��9�G��D$1�멍v ��[^_]Í�&    �UWVS������ÓC  ���t$ �l$$�F ��~J1���&    ��    �F����    ��R�V(��P�F�U��EF����P�  ��9~ Ń�[^_]Ð��&    �t& ���  ��C  �D$ǀ     ���(�����T$�P�T$�P�T$�P�T$�PÐ��&    ��&    WVS�|$��������B  ��W�  �T$ ���r=   $��h   j V��  XZWV�  ��[^_Ít& ��W�w  YZPV��  ���Ő��&    �WVS�t$������PB  �|$����<����W�6  �FXX�FZWP�W  �D$(�F�D$,�F�D$0�F�D$4���F[^_Ít& WVS�t$�-������A  �|$�F�N�P��F���|$ ��   Wh�   h�   h�   jRQP������ Wh�   h�   h�   j�F��P�FF��P�F��P�T����� Wh�   h�   h�   �F��Pj�F��P�v�)����� Wh�   h�   h�   �F��Pj�F��P�FF��P������� [^_�Wj`j`j`jRQP������� Wj`j`j`j�F��P�FF��P�F��P������ Wj`j`j`�F��Pj�F��P�v������ Wj`j`j`�o�����t& UWVS������ã@  ���t$0�|$4�F�n�N�P��F���l$���~ ��   ���n\�L$�N�L$����  ����  ����  ��Wh����h�����t$RP�t$ �������j WV������Wj j j �V�������F��P�V����ЋVX��F��)�P�t$(�P����� ��[^_]Ít& ���W��h�   �h�   ��h�   ��QRP�t$ �x����V�� W��h�   ��h�   �h�   ���P�R�N�Q�RFP�F��P�>����� Wj`j`j`j�F��P�v�F��P������ Wj`j`j`j�F��P�FF��P�F��P������� Wj`j`j`�F��Pj�F��P�v������� Wj`j`j`�F��Pj�F��P�FF��P������ ��[^_]Í�&    ��    ��Wh--��h22���t$RP�t$ �c�����jWV������Wh�   h�   h�   �k�����&    ��&    ���Wh��-�hȠ2�뮃�Wh�77�h�<<��VS������E>  ���t$�T$,�V��P�����D$ �F�D$$�F�D$(�F����P�
  �V�F(�F�V�F ��[^Ít& WVS�t$�������=  �|$����d����W��  �F�$��	  �FZYWP��  �D$(�F�D$,�F�D$0�F�D$4���F[^_Í�&    �t& ��G   ��w=  �D$�@    �@    �@    ��x�����T$�P�T$�P�T$�P�T$�PË$�S�c�����&=  �� j j j �t$4�D$$Pj�+  �D$,��8[�f�S�3������<  ��j j j j �t$(j!��  ��([Í�&    f�S�������<  ��j j j �t$(�t$(j��  ��([Í�&    UWVS������Ó<  ��(�l$<U�T����$�   �D$�����+   �T$����1����FjtUPǆ�   ����ǆ�   �����V�  �}�m����    ���� ��f��� vf��� wd���   ������P�  �����   ���   ���   ��ǆ�       ǆ�       Ɔ�    Ɔ�    ��[^_]Í�&    ��&    �ȃ���P�  ��롍�&    ��    S������Æ;  ���D$�p�u�����[��7�����g;  UWVS���l$0�T$�Eu(�����   S�����   �EP�EPj j ������� �E���   ��~?1����   �v 9�v\�M ��t1��v ���	9�u��A�������WP��E��9�̋��   ��t	��S�Ѓ���S�u�\$�������,[^_]Ð�    ��&    f�UWVS���D$0�l$4�|$8�p��~G� 1ۉD$��&    ��&    9�t<�D$��t1�f���� 9�u��@�P�H9�~9�|&��9�uσ�[^_]Í�&    �    ��&    f�H9�~�P9�~̅�t�T$1���&    ����9�u��T$�D$���@�P�R�D$@�����   ��[^_]Í�&    ��&    S���\$���   ��xn;CsY���t1Ґ���	9�u��A���P�R���   ��;Ss-���t1��t& ����	9�u��A��[Í�&    ��&    ��    ��&    f�ǃ�   ������1�[Í�&    ��&    �VS�R�����9  ���t$ j�E����T$ ���     �P��@    ��t�V��P�F�F��[^Ív ��F�F��[^ÐU��E�]�Mfof ��������]�U��E�]�M��~4fn�fo@�f��fs�f��fs�f��fs�f��f ������]Ð������                S�s�����68  ��h   �7  ����t�T$�@   �P��   �P��[Ít& S�3������7  ��j �t$�  ����1���x���t$R��������[Í�    S������ö7  ���D$�p�  ��1�[Í�&    ��&    S������Æ7  ���D$�D$P�t$�D$(�p��  ��[�f�S������V7  ���T$��t���D$�D$PR�D$(�p��  ����[Í�&    S�S�����7  ���t$�t$�D$�p�  ��[Í�&    �S�#������6  ��jj �D$�p��  ��[Í�&    �t& �1�Í�&    ��    1�Í�&    ��    S������Ö6  ���t$jj�D$P������[Í�&    �v WVS�|$������`6  ��W�U  �t$$j��PW������� 9�[^��_�����f�f��U��01�WVS�[�����6  ��(��8
  �����9�4
  C�4
  P���8  �����ڃ��  �  ����   �@ ����   �@ �   �D$   �   �)��    ���A    ���A    �A    �A    ��ux�A    ����   �p�¨�1���8
  �     �@    2z�p�@   �@    ��[^_]Í�&    �t& ��   �D$   �`�����&    ��&    �L$�D8 ��t��D8 ���s����D8 �i�����&    �v 1��D$   ������D$   �   � �����4  ��8   �g�����&    �t& ������4  ǀ@      �¨�ǀ<      �    �B    � �ǀ8
     �    �B    ��ǀ4
      �    �B    ǀ4      ǀ8      ǀ,      ǀ0      ǀ$      ǀ(      Í�&    �UWVS� ������3  ���|$0� ��&    ���4  �   ��8   ��  �w ��  ��t܋�@  �t$�|$0����  �|$0��<  ��8���a  �V�N�D$    �D$   ��)͉,$9���   �H�P�D$    �Ɖȉщl$)�1�9$�s��<  �$�T$9�s&�F����   �P�H�Ƌl$)�1�9$�r�9�rڋV����  ��)���9��  �J�j��t��)Ѓ�)�9���   �ʋJ�j��u�F���)�)�9���   �F��u��|$t-�D$�d����F����  �0�g���f��ȉщ��/����t& ���@  ����  �D$    �:����t& ��|$tًD$�����F���T  �0���,�����&    �t& �ՉM�L$�E�U�M(�L$0�u �M,�J�E$���������B1ҋD$~Q��@�����   ��   �E���  ����[^_]Í�&    �v ՋL$0�E�B�U�T$�E    �u �ЉU(1҉M,�����E$���~�Ƙ�Q�>�4$�v�9ǉQ���B�B�$��@��8�p���l����   )�Ń����`�����&    �t& ��H�P���$    �D$    ���D$    �щ�������������@  ���K�����  1���[��^_]ÍF��V�F�F$����F    �L$0�T$�v ~�ǘ��N,�����ЉV(�/1҉<$�Q�9ŉQ���B�B��$��@��(�x��u4���   �F��t  �����F�F$����F�F    �F    �x����   )�ƃ����Í�&    ��&    �UWVS�@�����0  ���D$ ����   �P���)փ� C���  �N�A=����~   �y�Š�1ҋA)E �GU+A�i���V�G�A�ޭޅ�t�U ����   �j�o��<  ����   ��t�J+J�ʋO)�9�|W�  ��[^_]Í�&    �v ��,  ��0   ����� ���� t
f=��t<�u���$  ��(   뱍�&    ���<  롍�&    ���4  ��8   ��[^_]Í�&    �v �G9�@  tU9�ta���t�B�G��t������G1�)Q���wW�  ���4�����&    �t& �o�������&    ���@  룍�&    �ǃ<      듍t& WVS�t$������P.  �t$��V�P���������   �¿   �^��ڃ��J��B�9˹    r\��t$�  �   ��t�@ �   ��u	�@ �   ��)�����Ӎ�&    ��&    ��    ��9�u������9�t@�Q� 9�v5�Q�D 9�v)�Q�D 9�v�Q�D 9�v�Q�D 9�v�D [^_Ít& UWVS������c-  ���t$4�l$0���>  ���V  �U���)Ѓ� Cŉ��A  �G�P�������   �P9���   �T$�+  ��V�������T$�ǃ��   �J�������   �D$�L ����&    �9�u��t$�ǃ�ƅ�t����t�A�F��t�Q�V��U����������[^_]Í�&    f��Ѓ�,  ��0   %��� =�� tDf����t=���t8�s  1���[��^_]Í�&    �p���V  ����[^_]Í�&    �t& ���$  ��(   븃�1�U��������j�����&    ��    ��V����������J�����&    ��    �Ɖ�����f�f�f��UWVS���\$(�l$ �T$$����   ��   �K��T$�؃��p��B�9���   �,$��t.�M�U �$�K���t�}�U�K��<$��u�U�M�$�K�)����\$1ۊ\$����������	��<$	ދ\$���Í�&    ��&    �0��9�u��t$�������)�9�t)���t#�P��t�P��t�P��t�P��t�P����[^_]É��ɍ�&    ��    UWVS�t$�D$�|$����   �V������,�   �(�v �1�y�����r��z�9�u�|$�t$����v��������S���t#�7��3��t�T7��T3���t�W�S[^_]Í�&    ��&    ����f�f�f�f�f�f��T$1��: t�t& ����< u�Í�    Í�&    ��&    �UWV1�S��������)  ���|$ �l$$�f��D5 �7����U�����7��9��� ����[^_]Ít& �UWVS�t$�\$�L$��t}�A�S9���9���	ЍV�����tm��	Ȩue���ȉڃ��ύ�&    �v �(�����j�9�u����9�t'���B9�v�D�D�B9�v	�D�D�� [^_]Í�&    �ȉٍ<0��&    f�������Q�9�u��͍�&    ��&    VS������å(  ���t$V����ZY�t$�P��������[^ËD$�L$��t& �����t	�8�u�Ð1�Í�&    ��    �D$�8 t��&    ���8 u�Í�&    U1�WVS�^�����!(  ���t$ �|$$���u�'��&    �t& ���.��t��PW�k�������u����[^_]Í�&    �v U1�WVS��������'  ���t$ �|$$���u�'��&    �t& ���.��t��PW��������t����[^_]Í�&    �v WVS�t$������`'  �|$��tV��D  ��WV�����XZWV�k��������D  9�t<1Ҁ8 u��D  ��[^_Í�&    f��  �P�㍴&    ���D  ��u�1���f�ǃD      1���f�VS�\$�t$��8�u"��t(�   ������t��8�t���)�[^Ít& �1�[^)�Í�&    f�UWVS�D$�\$�l$�0���8�u`��t@�<(��u�[��&    ��t,9�t8�����0���8�t�����[)�^_]Í�&    f�1�1�[)�^_]Ít& ���[��)�^_]�����������ōt& �UWVS�0������%  ���t$ �|$$��t& ��t)�������P��  ����$�  ��9��t����[^)�_]Í�    UWVS������Ó%  ���l$0�D$8�t$4�D$���&    �v ��t1;l$t+�����E ��P�S  ����$�F  ��9��E t����[^)�_]Í�&    ��&    WVS�t$�M�����%  ��V�������$�
����4$�����������Pj W�!���XZVW������[^_ÐS�������$  �� j j j �D$ P�t$8j��  �D$,��8[�f�S������Ö$  ��j j j j �t$(j�  ��([Í�&    f�S������f$  �� j �D$P�t$8�t$8�t$8j�g  �D$,��8[Í�&    ��&    S�c�����&$  �� j �D$P�t$8�t$8�t$8j�'  �D$,��8[Í�&    ��&    S�#������#  �� j �D$P�t$8�t$8�t$8j��  �D$,��8[Í�&    ��&    S������æ#  �� j �D$P�t$4�t$<�t$8j�  �D$,��8[Í�&    ��&    S������f#  ���t$�t$�t$�������[Í�&    �t& S�s�����6#  ���t$�t$�t$�������[Í�&    �t& S�C�����#  ���t$�t$�t$� �����[Í�&    �t& S�������"  ���t$�t$�������[Í�&    ��&    �S������æ"  ���t$�������1�[ÐS������Æ"  ��j �t$�������   ��u
����[Ív ��P������1҃���[�f�f�f�f�f��S�s�����6"  �� j j j �D$ P�t$8j�;   �D$,��8[�f�S�C�����"  ��j �t$0�t$0�t$0�t$(j�   ��([�f��WVS�D$�L$�T$�\$�t$ �|$$�i[^_�f�f�f�f�f�f�f��S������æ!  ��j j j j j j������ ��&    ��    ���f�f�f�f�f�f���T$�   �JЃ�	v���1���A����ËD$��߃�A������Í�&    �t& �1��|$z��Ít& �1��|$@��Ít& ��D$��0��	����Í�&    ��&    ��T$�   �JЃ�	v���1���A�����Í�&    ��&    ��D$��!��]����Í�&    ��&    ��T$�� ����	��	���Í�&    �v Í�&    ��&    �1�Í�&    ��    VS������U   ���t$V��������u��[^Í�&    f���V��������������[^Í�    �D$��_Í�&    ��D$�� �f�f�f�f�1�Í�&    ��    �����  �����  1�Í�&    �v S������ö  �� j j j �D$ P�t$8j�����D$,��8[�f�1��f�f�f�f�f�f�������t6U��S������&    �v �Ѓ�����u��[]Í�&    ��&    �������     / r /file.bmp /binfile.bmp /folder.bmp          Ї��8�       zR |�        ���)    A�Be�     <   "���>    A�Bz�     \   @����    A�B�� (   |   �����   A�BB����A�A�       �   ����   A�BG���(   �   ����z   D Gu Eutu|ux    �   ���U    A�BQ�      ����(    A�Bd�     8  ����    A�BV�  |   X  ����~    A�A�A�A�N U$A(A,D0H E$K(A,D0H G
A�A�A�A�CC$C(A,G0H CA�A�A�A�     �  ����
          �  ����              ����$    A�NE HD� 0   $   ���B    A�A�N^DE HA�A�  4   X  ���L    A�A�NcAE HHA�A�   \   �  4����    A�A�A�A�N n
A�A�A�A�LC$F(D,A0H YA�A�A�A�   �  d���?    Cy H     �����    K�A�A�A�C@�DAHDLYPL@IA�A�A�A� 8   T  @���.    A�A�NFB B$B(A,B0HC�A� H   �  4����    K�A�A�A�C@�DAHFLHPL@IA�A�A�A� H   �  �����    K�A�A�A�C@�DAHDLJPL@IA�A�A�A� <   (  L���b   A�A�A�A�NPL@�A�A�A�A�X   h  |����   A�A�A�A�N`&dph_l]pDtBxD|A�H`MA�A�A�A�   X   �  �����   A�A�A�A�N`&dph_l]pBtDxA|D�H`MA�A�A�A�   H      d����    A�A�A�A�N0O4K8J<\@H0HA�A�A�A� 8   l  �����    A�A�A�A�C(�A�A�A�A�   �  ����          �  q���           �  d���(    A�SJ HA�     �  p���    A�ND HA�       l���    A�ND HA�     <  h���    A�ND HA�     `  d���    A�ND HA�     �  `���    A�ND HA�   �  \���W   A�A�A�A�N0�4D8D<F@BDBHALDPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0P4D8D<F@BDBHALHPH0M4G8D<F@BDBHALKPH0MA�A�A�A�T   �  ����s    A�A�A�A�N0q4G8A<D@DDDHALDPK0GA�A�A�A�       ����          (  ����          <  ����	          P  ����	          d  ����	       �   x  ����{   A�A�C�C�N0H4E8E<E@CDCHCLCPO0e<D@H0G4D8H<H@HDHHILFPK0c4B8B<B@BDBHDLAPH0D4E8E<E@CDBHBLGPH0D4E8E<E@BDBHBLGPH0D4E8E<E@BDBHGLGPHA�A�A�A� \   \	  X����    A�C�A�C�N0f<A@H0G4D8B<B@BDHHILHPK0YA�A�A�A� H   �	  ����s    A�A�A�A�N d$K(G,V0H HA�A�A�A�     
  ����A       d   
  ���g    A�A�A�RA LMEBA FAAA HA
�A�A�ECA FAAA H@   �
  ���\    A�A�A�VL IDAA aD�A�A�   �   �
  ,���K   A�A�A�nEEE B$A(A,A0HAEEE B$G(J,G0HAEEE G$B(G,C0HAEEE G$B(G,J0HA
�A�A�AABBB B$A(A,A0HABBB B$G(J,G0HABBB G$B(G,C0HABBB �  �  ����`   A�A�A�A�N0Z4A8E<E@DDAHALDPH4B8A<A@H4A8B<B@BDSHXLDPH0C
A�A�A�A�FC4H8G<G@DDAHALDPK0A4G8H<G@FDGHDLGPH0A4B8B<B@BDGHCLGPH0A4B8B<B@BDGHJLGPH0A4B8B<B@GDBHGLCPH0A4B8B<B@GDBHGLJPH0C
A�A�A�A�NC4A8E<E@DDAHALDPH4B8A<A@H4A8E<E@EDT0C
4A8E<E@BC4A8E<E@ (   H  \���\    A�A�Nr WA�A�@   t  ����d    A�A�A�VL TAAA aD�A�A�      �  ����L          �  ����       0   �  ����.    A�N(B,B0B4D8E<B@LA�  0     ����'    A�NBB B$B(D,B0HA�  0   H  ����)    A�NBB B$D(D,B0HA�  `   |  ����   A�A�A�A�N<E@a4M8A<A@g0g<G@H0y
A�A�A�A�OE<D@H0      �  ����     A�NG HA� x     �����    L�A�A�A�C0Q8G<H@EDEHBLBPH0w8H<A@H0Q<A@E0C8A<C@LA�A�A�A�B0����X   �  �����    A�A�A�A�C0]
A�A�A�A�HD<F@J0IA�A�A�A�0   �  X����    A�CkC La
A�P]C� <     ����_    A�A�NF Lh
A�A�DLA�A�   $   P  d���<    A�NE H^A�  4   x  |���:    A�NBD HKDA HCA�       �  ����"    A�NG HC� (   �  ����.    A�NJDG HA�   ,      ����9    A�NKJAG HCA� (   0  ����(    A�NDDG HA�   (   \  ����$    A�NBBG HA�      �  ����          �  ����       (   �  ����&    A�NDBBE HA�@   �  ����;    A�A�A�RA I$B(C,A0HC�A�D�   D      �����   A�F�A�A�N<Z@J0�
A�A�A�A�M      h  �����       T   |  �����   A�A�A�A�N0
C�A�A�A�K�
A�C�A�A�A `   �  ����   A�A�A�A�N �
A�A�A�A�Ka
A�A�A�A�Kt(C,A0H   4   8  \����    A�A�A�WA H��A�A�  �   p  ����   A�A�A�A�N0V<A@H0c<A@H0C
C�A�A�A�Jr
A�C�A�A�HM
C�A�A�A�MS<C@H0U<A@H0<      4���   A�A�A�A�C �
C�A�A�A�A 8   @  ����    A�A�A�A��
�A�A�A�P      |  x���!       @   �  ����K    A�A�A�C�N Z,A0K JC�A�A�A�8   �  �����    A�A�A�A��
�A�A�A�H   4     4���0    A�A�NE FADC HC�A�   H  ,���#          \  H���       D   p  T���V    A�C�A�A�N j(A,A0H GC�A�A�A� D   �  l���V    A�C�A�A�N j(A,A0H GC�A�A�A� D      �����    A�A�A�`AA HAAA H\
�A�A�J ,   H  ����G    A�A�w
�A�FC�A�  \   x  �����    A�A�A�A�M
�C�A�A�JE
�C�A�A�FD
�E�A�A�A @   �  ���Z    A�A�A�A�N ^,A0U MA�A�C�A�@     8���r    A�A�A�A�N0u<A@U0NA�A�C�A�L   `  t���O    A�A�A�RA ]DBA FAAA HA�A�A�   0   �  t���.    A�N(B,B0B4E8D<B@LA�  0   �  p���'    A�NBB B$B(D,B0HA�  0     l���2    A�N(B,E0D4D8D<B@LA�  0   L  x���2    A�N(B,E0D4D8D<B@LA�  0   �  ����2    A�N(B,E0D4D8D<B@LA�  0   �  ����2    A�N(B,E0D4D8D<B@LA�  (   �  ����%    A�NDDD HA�   (     ����%    A�NDDD HA�   (   @  ����%    A�NDDD HA�   $   l  ����!    A�NDD HA�      �  ����    A�ND HC� 8   �  ����E    A�NBD HL
C�DCA HEC�0   �  ����.    A�N(B,B0B4E8D<B@LA�  0   (  ����-    A�NBD D$D(D,B0HA�  (   \  ����!    A�A�A�[�A�A�,   �  ����3    A�NBB B$B(B,B0H     �  ����           �  ����          �  ����          �  ����            ����            ����           0  ����          D  ����          X  ����          l  ���          �  ���       D   �   ���J    A�A�NE HG
A�A�JCA HHD�A�     �  ���          �  ���             ���            ����       0   ,  ���.    A�N(B,B0B4E8D<B@LA�     `  ���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               ������    ����            ������        К����        ������        �����        P�����        ������                                                                                                                                                                                                                                                                                                                           <<  66      66666 >0  c3fc 6n;3n         f<�<f   ?          ?          `0 >cs{og> ? 303? 3003 8<630x ?003 33 ?30 3333 33>0           ?  ?  0 30  >c{{{ 33?33 ?ff>ff? <ff< 6fff6 FF F <fsf| 333?333  x00033 gf66fg Ff cwkcc cgo{scc 6ccc6 ?ff> 333;8 ?ff>6fg 383 ?- 333333? 33333 ccckwc cc66c 333 c1Lf  0`@  6c           �       0>3n >ff;   33 800>33n   3? 6   n33>06nffg   0 00033f66g    3kc   3333   333   ;ff>  n33>0x  ;nf   >0 >,   3333n   333   ck6   c66c   333>0  ?&? 88   8 n;                                               $                                                         `                           `                                   8$$ T                                              @8 0                                                             8$$A$8    <<|B~<~<>    $8<|<|~~<B|B@BB<|<|>~BBDBD~@(  @   @@p                                                 8H$*�$ (   B0BB@@BB @BDBBBB@@BBD@fbBBBB@BBDBD D   @    @  @                                                 8 �(d  (   NPBB@@BB  ~0�BB@B@@@BX@~ZBBBB@BBD$D    >|<>< >|8F<<<<<^>|BBDBB~                                   8 $H$   | ~ R|B|\<B  0 �B|@B||@~`@ZFBBBB<BBT(   BBBBB|BBXZBBBB`@ BBD$B 2                                   $P      b>BB>  @ �~B@B@@BB`@ZBB|B|BBT$    BB@BB BB`ZBBBB@< BBTBL                                   �
"J       B BB0~�BB@B@@BBX@BBB@BHBB|B@   BB@B| BB`ZBBBB@ BBT$B                                      $
EJ        B@BB 0�BBBB@@FBBD@BBB@FDB$lB@   BBBB@ BBXBBBBB@ B$TBB@                                     $*�F     @<~~||<<|   @ @B|<|~@:B|>B~BB<@<B|<DB~   ><<>> >BFBB<|>@|><B>~                                    $<      @                8                         8               @                                                  @                                                         |  |     @       |  `        GNU C crti.s GCC: (GNU) 8.2.0 GNU C crtn.o              Ч�                           >        ЧP�    src/gfx/sse2.asm NASM 2.14.02 �Ч     %  . @   _    '   �       src/gfx/sse2.asm      Ч!0==?LL==0/!#!0==>=0K�KYKYKYMK>1/""u�                                            t�          ��          Q�          \�          ��           �          �          �          �     	     ��     
     ��          ��                                                                                                                                  ��   �         �      (   ��      ;   ��      =    �      P   P�      f   ��     u   ��     �   Ё      �   ��                 ���   �      �   �      �   �      �            ��  ��                  ��  ��(     F  ��     d           ��q           ��}           ���           ���           ���           ���           ���  ܧ       �  ,�       �  5�       �  @�     �           ���           ���  `��      ��       ��     #  ��     2  ��     <  ��     F  ��     S  ��     f           ��o           ��x  ��                ���           ���           ���           ���           ���           ��             ���  ��     
 �  ��     �  ��K     �  0�.     �  P��    &  ��     K  ��     W  `�.     v  Ї�  "  �  ��`    �  ��     �  ��'     �  ��!     �  ��     �  ��     �  P�.     !  ��       Ж(   "     �2       �        ���    L  ��B     ^  p�A     r  ��     y  0�\     �  ��     �  ��     �  ��-     �  �     �  ��.     �  `�     �  ��     �  �     �   ��     �  ���    �   �t       Ŗ       ��     (  0�J     0  К{    L  �     T  Щ     [  ��K    �  <�   ! 	 �  ��%     �  �     �   �   "  �  (�   ! 	 �  �r     �  \�     �  ��     �  ��U   "    ��      �  t�        ��     &  ��>   "  @  ��	     Z  І)   "  n  `��     �  @�     �  0�\     �  0��       P�%     �  �     �  ��~     �  P��     �  �0     �  �      p�(       `�2       ��W    8  І)   "  L  ��     f  �     4	  ��&     j  �     w  x�   ! 	    �%     �  p�A     �  p�     �   ��     �  p�_     �  ��.     �  �s     �  @�   "     ��       ��Z        ��      p�
     )  0��     N   ��     U  ɖ     k  �    �  P�<     �  �b    �  `��     �   �      �  @�     �  �   ! 	 �   �s     	   �.     "	  p�O     )	  ��:     /	  ��      ;	  0��     a	  д    h	  �z    m	  ��$     s	  ��     �	  ��?     �	  P�   ! 	 U   �     �	  `�   "  �	  �L     �	  Ш"     �	  п     �	  ��$     �	   �      �	   �     �	  ��G     �	  @�\     

  ��   !  
  Q�      !
  ��g     9
  ��V     A
  ��)     ]
  ��     x
   �     �
  @�\     �
  �&     �
   �   "  �
  8��   "  �
  ��     �
  ��     �
  �L     �
  0�9     �
   �E       ��        ��        ��d     !  Ц�     ;  ��2     F  �3     K  ��	     b  ��     j   ��     �  `�V     �  ��!     �  ��!     �  ��     �  �'     �  ��d     �  �#     �   �;     �  ��     �  d�   ! 	 �  ��	        �        ��   "    �2     "  Ч      �  �     .  ��>   "  H  Е�     �
  ���    w  �L      crtstuff.c __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ deregister_tm_clones __do_global_dtors_aux completed.4231 dtor_idx.4233 frame_dummy object.4243 __CTOR_END__ __FRAME_END__ __do_global_ctors_aux /home/computerfido/Desktop/Lemon/FakeSysroot/usr/lib/crt0.o hang main.cpp _Z41__static_initialization_and_destruction_0ii _GLOBAL__sub_I_fileIconBuffer graphics.cpp runtime.cpp text.cpp widgets.cpp window.cpp font.cpp src/gfx/sse2.asm memcpy_sse2.loop memset_sse2.loop memset_sse2.ret bigzero fileio.c allocate_new_page l_pageSize l_pageCount l_warningCount l_memRoot l_bestBet l_errorCount l_possibleOverruns memory.c string.c p.1056 filesystem.c ipc.c syscall.c exit.c ctype.c _liballoc.c _GLOBAL_OFFSET_TABLE_ l_allocated strcpy _Z12GetVideoModev _Z20DrawGradientVerticaliiii10RGBAColourS_P7Surface _ZN15ScrollContainer5PaintEP7Surface _Z7inportbt _Z13_CreateWindowP10win_info_t _ZN10FileButton5PaintEP7Surface _ZN6Button5PaintEP7Surface l_max_inuse _Z14_DestroyWindowPv syscall liballoc_init liballoc_unlock ReceiveMessage _Znwm lemon_read isblank _Z12DrawGradientiiii10RGBAColourS_P7Surface _Z12write_serialc _ZN7TextBoxC2E4Rect memcpy _ZN6ButtonC1EPc4Rect l_inuse __TMC_END__ SendMessage __DTOR_END__ lemon_open islower tolower feof _Z11PaintWindowP6Window malloc windowInfo __x86.get_pc_thunk.ax __dso_handle ispunct _ZN7TextBox5PaintEP7Surface isspace fflush _ZN6Button17DrawButtonBordersEP7Surfaceb _ZTV6Button lseek fd _ZdlPv _ZTV7TextBox strncasecmp __x86.get_pc_thunk.dx _Z15HandleMouseDownP6Window8Vector2i _ZN4ListIP6WidgetE5clearEv isxdigit liballoc_lock _ZN10FileButtonC2EPc4Rect _ZN6Button11OnMouseDownEv _ZN10win_info_tC2Ev _Z18memset32_optimizedPvjm strrchr _ZN6ButtonC2EPc4Rect calloc folderIconBuffer _Z16memcpy_optimizedPvS_m _ZN5Label5PaintEP7Surface strcat _Z12RefreshFilesv fseek lemon_write _Z8DrawCharciihhhP7Surface _ZN10win_info_tC1Ev _ZN6Widget11OnMouseDownEv win exIconBuffer _ZTV15ScrollContainer _ZN7TextBoxC1E4Rect isupper strncmp _Z9AddWidgetP6WidgetP6Window liballoc_alloc _ZN6Bitmap5PaintEP7Surface _ZdlPvm strncpy strcasecmp realloc _Z8outportbth _Z8DrawRectiiii10RGBAColourP7Surface strtok __x86.get_pc_thunk.bx _Z12CreateWindowP10win_info_t fdopen _Z15DrawBitmapImageiiiiPhP7Surface _Z8DrawRectiiiihhhP7Surface _Z13DestroyWindowP6Window isalpha _ZTV6Widget _Z10DrawStringPcjjhhhP7Surface fread strdup fopen __bss_start _Z8DrawRect4Rect10RGBAColourP7Surface memset main ftell font_default _Z5floord _ZTV6Bitmap _ZdaPv _ZN15ScrollContainerC2E4Rect fclose isgraph _Z17is_transmit_emptyv isalnum isprint strcmp _ZN6BitmapC1E4Rect _ZTV10FileButton _fini _ZN7TextBox8LoadTextEPc strcspn _Z12_PaintWindowPvP7Surface _ZN6Widget5PaintEP7Surface liballoc_free _ZN6BitmapC2E4Rect fputc _Znam _ZN10FileButton9OnMouseUpEv _ZN6Widget9OnMouseUpEv isdigit _Z12write_serialPc fwrite access _edata _end _ZN5LabelC2EPc4Rect _Z13HandleMouseUpP6Window lemon_seek exit _ZN6Button9OnMouseUpEv iscntrl _Z10surfacecpyP7SurfaceS0_8Vector2i strspn strlen toupper lemon_close _ZN5LabelC1EPc4Rect strchr fputs font_old _ZTV5Label _ZN7TextBox11OnMouseDownEv memset_sse2 _ZdaPvm lemon_readdir memcpy_sse2 _ZN10FileButtonC1EPc4Rect _Z21surfacecpyTransparentP7SurfaceS0_8Vector2i _ZN15ScrollContainerC1E4Rect  .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .init_array .ctors .dtors .data.rel.ro .got.plt .data .bss .comment .debug_aranges .debug_pubnames .debug_info .debug_abbrev .debug_line .debug_frame .debug_loc                                                  t�t                     !         ���   �@                 '         Q�QA                    -         \�\A  <                  5         ���A  t                 ?          � `                   K         �`                    R         �`                    Y         �`  x                  f         ���`                   o         ���`  (
                  u         ���j  �                   z      0       �j  +                 �              �j                     �              k                    �              %k  B                  �              gk                    �              �k  c                  �              �k                    �              �k                                  �k  �     I         	              �z  �                               p�  �                  